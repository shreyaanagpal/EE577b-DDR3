
module FIFO_DEPTH_P25_WIDTH16 ( clk, reset, data_in, put, get, data_out, 
        empty_bar, full_bar, fillcount );
  input [15:0] data_in;
  output [15:0] data_out;
  output [5:0] fillcount;
  input clk, reset, put, get;
  output empty_bar, full_bar;
  wire   n12, n13, n14, n15, n16, n2314, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
         n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
         n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
         n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
         n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
         n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
         n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
         n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
         n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
         n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
         n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877,
         n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887,
         n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897,
         n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946;
  wire   [4:0] wr_ptr;
  wire   [511:0] mem;
  assign full_bar = 1'b1;

  DFFPOSX1 wr_ptr_reg_0_ ( .D(n1413), .CLK(clk), .Q(wr_ptr[0]) );
  DFFPOSX1 rd_ptr_reg_4_ ( .D(n2316), .CLK(clk), .Q(n16) );
  DFFPOSX1 rd_ptr_reg_0_ ( .D(n1411), .CLK(clk), .Q(n12) );
  DFFPOSX1 rd_ptr_reg_1_ ( .D(n1410), .CLK(clk), .Q(n13) );
  DFFPOSX1 rd_ptr_reg_2_ ( .D(n1409), .CLK(clk), .Q(n14) );
  DFFPOSX1 rd_ptr_reg_3_ ( .D(n1408), .CLK(clk), .Q(n15) );
  DFFPOSX1 wr_ptr_reg_4_ ( .D(n1407), .CLK(clk), .Q(wr_ptr[4]) );
  DFFPOSX1 wr_ptr_reg_1_ ( .D(n1406), .CLK(clk), .Q(wr_ptr[1]) );
  DFFPOSX1 wr_ptr_reg_2_ ( .D(n1405), .CLK(clk), .Q(wr_ptr[2]) );
  DFFPOSX1 wr_ptr_reg_3_ ( .D(n1404), .CLK(clk), .Q(wr_ptr[3]) );
  DFFPOSX1 data_out_reg_15_ ( .D(n2332), .CLK(clk), .Q(data_out[15]) );
  DFFPOSX1 data_out_reg_14_ ( .D(n2331), .CLK(clk), .Q(data_out[14]) );
  DFFPOSX1 data_out_reg_13_ ( .D(n2330), .CLK(clk), .Q(data_out[13]) );
  DFFPOSX1 data_out_reg_12_ ( .D(n2329), .CLK(clk), .Q(data_out[12]) );
  DFFPOSX1 data_out_reg_11_ ( .D(n2328), .CLK(clk), .Q(data_out[11]) );
  DFFPOSX1 data_out_reg_10_ ( .D(n2327), .CLK(clk), .Q(data_out[10]) );
  DFFPOSX1 data_out_reg_9_ ( .D(n2326), .CLK(clk), .Q(data_out[9]) );
  DFFPOSX1 data_out_reg_8_ ( .D(n2325), .CLK(clk), .Q(data_out[8]) );
  DFFPOSX1 data_out_reg_7_ ( .D(n2324), .CLK(clk), .Q(data_out[7]) );
  DFFPOSX1 data_out_reg_6_ ( .D(n2323), .CLK(clk), .Q(data_out[6]) );
  DFFPOSX1 data_out_reg_5_ ( .D(n2322), .CLK(clk), .Q(data_out[5]) );
  DFFPOSX1 data_out_reg_4_ ( .D(n2321), .CLK(clk), .Q(data_out[4]) );
  DFFPOSX1 data_out_reg_3_ ( .D(n2320), .CLK(clk), .Q(data_out[3]) );
  DFFPOSX1 data_out_reg_2_ ( .D(n2319), .CLK(clk), .Q(data_out[2]) );
  DFFPOSX1 data_out_reg_1_ ( .D(n2318), .CLK(clk), .Q(data_out[1]) );
  DFFPOSX1 data_out_reg_0_ ( .D(n2317), .CLK(clk), .Q(data_out[0]) );
  DFFPOSX1 mem_reg_31__15_ ( .D(n1403), .CLK(clk), .Q(mem[511]) );
  DFFPOSX1 mem_reg_31__14_ ( .D(n1402), .CLK(clk), .Q(mem[510]) );
  DFFPOSX1 mem_reg_31__13_ ( .D(n1401), .CLK(clk), .Q(mem[509]) );
  DFFPOSX1 mem_reg_31__12_ ( .D(n1400), .CLK(clk), .Q(mem[508]) );
  DFFPOSX1 mem_reg_31__11_ ( .D(n1399), .CLK(clk), .Q(mem[507]) );
  DFFPOSX1 mem_reg_31__10_ ( .D(n1398), .CLK(clk), .Q(mem[506]) );
  DFFPOSX1 mem_reg_31__9_ ( .D(n1397), .CLK(clk), .Q(mem[505]) );
  DFFPOSX1 mem_reg_31__8_ ( .D(n1396), .CLK(clk), .Q(mem[504]) );
  DFFPOSX1 mem_reg_31__7_ ( .D(n1395), .CLK(clk), .Q(mem[503]) );
  DFFPOSX1 mem_reg_31__6_ ( .D(n1394), .CLK(clk), .Q(mem[502]) );
  DFFPOSX1 mem_reg_31__5_ ( .D(n1393), .CLK(clk), .Q(mem[501]) );
  DFFPOSX1 mem_reg_31__4_ ( .D(n1392), .CLK(clk), .Q(mem[500]) );
  DFFPOSX1 mem_reg_31__3_ ( .D(n1391), .CLK(clk), .Q(mem[499]) );
  DFFPOSX1 mem_reg_31__2_ ( .D(n1390), .CLK(clk), .Q(mem[498]) );
  DFFPOSX1 mem_reg_31__1_ ( .D(n1389), .CLK(clk), .Q(mem[497]) );
  DFFPOSX1 mem_reg_31__0_ ( .D(n1388), .CLK(clk), .Q(mem[496]) );
  DFFPOSX1 mem_reg_30__15_ ( .D(n1387), .CLK(clk), .Q(mem[495]) );
  DFFPOSX1 mem_reg_30__14_ ( .D(n1386), .CLK(clk), .Q(mem[494]) );
  DFFPOSX1 mem_reg_30__13_ ( .D(n1385), .CLK(clk), .Q(mem[493]) );
  DFFPOSX1 mem_reg_30__12_ ( .D(n1384), .CLK(clk), .Q(mem[492]) );
  DFFPOSX1 mem_reg_30__11_ ( .D(n1383), .CLK(clk), .Q(mem[491]) );
  DFFPOSX1 mem_reg_30__10_ ( .D(n1382), .CLK(clk), .Q(mem[490]) );
  DFFPOSX1 mem_reg_30__9_ ( .D(n1381), .CLK(clk), .Q(mem[489]) );
  DFFPOSX1 mem_reg_30__8_ ( .D(n1380), .CLK(clk), .Q(mem[488]) );
  DFFPOSX1 mem_reg_30__7_ ( .D(n1379), .CLK(clk), .Q(mem[487]) );
  DFFPOSX1 mem_reg_30__6_ ( .D(n1378), .CLK(clk), .Q(mem[486]) );
  DFFPOSX1 mem_reg_30__5_ ( .D(n1377), .CLK(clk), .Q(mem[485]) );
  DFFPOSX1 mem_reg_30__4_ ( .D(n1376), .CLK(clk), .Q(mem[484]) );
  DFFPOSX1 mem_reg_30__3_ ( .D(n1375), .CLK(clk), .Q(mem[483]) );
  DFFPOSX1 mem_reg_30__2_ ( .D(n1374), .CLK(clk), .Q(mem[482]) );
  DFFPOSX1 mem_reg_30__1_ ( .D(n1373), .CLK(clk), .Q(mem[481]) );
  DFFPOSX1 mem_reg_30__0_ ( .D(n1372), .CLK(clk), .Q(mem[480]) );
  DFFPOSX1 mem_reg_29__15_ ( .D(n1371), .CLK(clk), .Q(mem[479]) );
  DFFPOSX1 mem_reg_29__14_ ( .D(n1370), .CLK(clk), .Q(mem[478]) );
  DFFPOSX1 mem_reg_29__13_ ( .D(n1369), .CLK(clk), .Q(mem[477]) );
  DFFPOSX1 mem_reg_29__12_ ( .D(n1368), .CLK(clk), .Q(mem[476]) );
  DFFPOSX1 mem_reg_29__11_ ( .D(n1367), .CLK(clk), .Q(mem[475]) );
  DFFPOSX1 mem_reg_29__10_ ( .D(n1366), .CLK(clk), .Q(mem[474]) );
  DFFPOSX1 mem_reg_29__9_ ( .D(n1365), .CLK(clk), .Q(mem[473]) );
  DFFPOSX1 mem_reg_29__8_ ( .D(n1364), .CLK(clk), .Q(mem[472]) );
  DFFPOSX1 mem_reg_29__7_ ( .D(n1363), .CLK(clk), .Q(mem[471]) );
  DFFPOSX1 mem_reg_29__6_ ( .D(n1362), .CLK(clk), .Q(mem[470]) );
  DFFPOSX1 mem_reg_29__5_ ( .D(n1361), .CLK(clk), .Q(mem[469]) );
  DFFPOSX1 mem_reg_29__4_ ( .D(n1360), .CLK(clk), .Q(mem[468]) );
  DFFPOSX1 mem_reg_29__3_ ( .D(n1359), .CLK(clk), .Q(mem[467]) );
  DFFPOSX1 mem_reg_29__2_ ( .D(n1358), .CLK(clk), .Q(mem[466]) );
  DFFPOSX1 mem_reg_29__1_ ( .D(n1357), .CLK(clk), .Q(mem[465]) );
  DFFPOSX1 mem_reg_29__0_ ( .D(n1356), .CLK(clk), .Q(mem[464]) );
  DFFPOSX1 mem_reg_28__15_ ( .D(n1355), .CLK(clk), .Q(mem[463]) );
  DFFPOSX1 mem_reg_28__14_ ( .D(n1354), .CLK(clk), .Q(mem[462]) );
  DFFPOSX1 mem_reg_28__13_ ( .D(n1353), .CLK(clk), .Q(mem[461]) );
  DFFPOSX1 mem_reg_28__12_ ( .D(n1352), .CLK(clk), .Q(mem[460]) );
  DFFPOSX1 mem_reg_28__11_ ( .D(n1351), .CLK(clk), .Q(mem[459]) );
  DFFPOSX1 mem_reg_28__10_ ( .D(n1350), .CLK(clk), .Q(mem[458]) );
  DFFPOSX1 mem_reg_28__9_ ( .D(n1349), .CLK(clk), .Q(mem[457]) );
  DFFPOSX1 mem_reg_28__8_ ( .D(n1348), .CLK(clk), .Q(mem[456]) );
  DFFPOSX1 mem_reg_28__7_ ( .D(n1347), .CLK(clk), .Q(mem[455]) );
  DFFPOSX1 mem_reg_28__6_ ( .D(n1346), .CLK(clk), .Q(mem[454]) );
  DFFPOSX1 mem_reg_28__5_ ( .D(n1345), .CLK(clk), .Q(mem[453]) );
  DFFPOSX1 mem_reg_28__4_ ( .D(n1344), .CLK(clk), .Q(mem[452]) );
  DFFPOSX1 mem_reg_28__3_ ( .D(n1343), .CLK(clk), .Q(mem[451]) );
  DFFPOSX1 mem_reg_28__2_ ( .D(n1342), .CLK(clk), .Q(mem[450]) );
  DFFPOSX1 mem_reg_28__1_ ( .D(n1341), .CLK(clk), .Q(mem[449]) );
  DFFPOSX1 mem_reg_28__0_ ( .D(n1340), .CLK(clk), .Q(mem[448]) );
  DFFPOSX1 mem_reg_27__15_ ( .D(n1339), .CLK(clk), .Q(mem[447]) );
  DFFPOSX1 mem_reg_27__14_ ( .D(n1338), .CLK(clk), .Q(mem[446]) );
  DFFPOSX1 mem_reg_27__13_ ( .D(n1337), .CLK(clk), .Q(mem[445]) );
  DFFPOSX1 mem_reg_27__12_ ( .D(n1336), .CLK(clk), .Q(mem[444]) );
  DFFPOSX1 mem_reg_27__11_ ( .D(n1335), .CLK(clk), .Q(mem[443]) );
  DFFPOSX1 mem_reg_27__10_ ( .D(n1334), .CLK(clk), .Q(mem[442]) );
  DFFPOSX1 mem_reg_27__9_ ( .D(n1333), .CLK(clk), .Q(mem[441]) );
  DFFPOSX1 mem_reg_27__8_ ( .D(n1332), .CLK(clk), .Q(mem[440]) );
  DFFPOSX1 mem_reg_27__7_ ( .D(n1331), .CLK(clk), .Q(mem[439]) );
  DFFPOSX1 mem_reg_27__6_ ( .D(n1330), .CLK(clk), .Q(mem[438]) );
  DFFPOSX1 mem_reg_27__5_ ( .D(n1329), .CLK(clk), .Q(mem[437]) );
  DFFPOSX1 mem_reg_27__4_ ( .D(n1328), .CLK(clk), .Q(mem[436]) );
  DFFPOSX1 mem_reg_27__3_ ( .D(n1327), .CLK(clk), .Q(mem[435]) );
  DFFPOSX1 mem_reg_27__2_ ( .D(n1326), .CLK(clk), .Q(mem[434]) );
  DFFPOSX1 mem_reg_27__1_ ( .D(n1325), .CLK(clk), .Q(mem[433]) );
  DFFPOSX1 mem_reg_27__0_ ( .D(n1324), .CLK(clk), .Q(mem[432]) );
  DFFPOSX1 mem_reg_26__15_ ( .D(n1323), .CLK(clk), .Q(mem[431]) );
  DFFPOSX1 mem_reg_26__14_ ( .D(n1322), .CLK(clk), .Q(mem[430]) );
  DFFPOSX1 mem_reg_26__13_ ( .D(n1321), .CLK(clk), .Q(mem[429]) );
  DFFPOSX1 mem_reg_26__12_ ( .D(n1320), .CLK(clk), .Q(mem[428]) );
  DFFPOSX1 mem_reg_26__11_ ( .D(n1319), .CLK(clk), .Q(mem[427]) );
  DFFPOSX1 mem_reg_26__10_ ( .D(n1318), .CLK(clk), .Q(mem[426]) );
  DFFPOSX1 mem_reg_26__9_ ( .D(n1317), .CLK(clk), .Q(mem[425]) );
  DFFPOSX1 mem_reg_26__8_ ( .D(n1316), .CLK(clk), .Q(mem[424]) );
  DFFPOSX1 mem_reg_26__7_ ( .D(n1315), .CLK(clk), .Q(mem[423]) );
  DFFPOSX1 mem_reg_26__6_ ( .D(n1314), .CLK(clk), .Q(mem[422]) );
  DFFPOSX1 mem_reg_26__5_ ( .D(n1313), .CLK(clk), .Q(mem[421]) );
  DFFPOSX1 mem_reg_26__4_ ( .D(n1312), .CLK(clk), .Q(mem[420]) );
  DFFPOSX1 mem_reg_26__3_ ( .D(n1311), .CLK(clk), .Q(mem[419]) );
  DFFPOSX1 mem_reg_26__2_ ( .D(n1310), .CLK(clk), .Q(mem[418]) );
  DFFPOSX1 mem_reg_26__1_ ( .D(n1309), .CLK(clk), .Q(mem[417]) );
  DFFPOSX1 mem_reg_26__0_ ( .D(n1308), .CLK(clk), .Q(mem[416]) );
  DFFPOSX1 mem_reg_25__15_ ( .D(n1307), .CLK(clk), .Q(mem[415]) );
  DFFPOSX1 mem_reg_25__14_ ( .D(n1306), .CLK(clk), .Q(mem[414]) );
  DFFPOSX1 mem_reg_25__13_ ( .D(n1305), .CLK(clk), .Q(mem[413]) );
  DFFPOSX1 mem_reg_25__12_ ( .D(n1304), .CLK(clk), .Q(mem[412]) );
  DFFPOSX1 mem_reg_25__11_ ( .D(n1303), .CLK(clk), .Q(mem[411]) );
  DFFPOSX1 mem_reg_25__10_ ( .D(n1302), .CLK(clk), .Q(mem[410]) );
  DFFPOSX1 mem_reg_25__9_ ( .D(n1301), .CLK(clk), .Q(mem[409]) );
  DFFPOSX1 mem_reg_25__8_ ( .D(n1300), .CLK(clk), .Q(mem[408]) );
  DFFPOSX1 mem_reg_25__7_ ( .D(n1299), .CLK(clk), .Q(mem[407]) );
  DFFPOSX1 mem_reg_25__6_ ( .D(n1298), .CLK(clk), .Q(mem[406]) );
  DFFPOSX1 mem_reg_25__5_ ( .D(n1297), .CLK(clk), .Q(mem[405]) );
  DFFPOSX1 mem_reg_25__4_ ( .D(n1296), .CLK(clk), .Q(mem[404]) );
  DFFPOSX1 mem_reg_25__3_ ( .D(n1295), .CLK(clk), .Q(mem[403]) );
  DFFPOSX1 mem_reg_25__2_ ( .D(n1294), .CLK(clk), .Q(mem[402]) );
  DFFPOSX1 mem_reg_25__1_ ( .D(n1293), .CLK(clk), .Q(mem[401]) );
  DFFPOSX1 mem_reg_25__0_ ( .D(n1292), .CLK(clk), .Q(mem[400]) );
  DFFPOSX1 mem_reg_24__15_ ( .D(n1291), .CLK(clk), .Q(mem[399]) );
  DFFPOSX1 mem_reg_24__14_ ( .D(n1290), .CLK(clk), .Q(mem[398]) );
  DFFPOSX1 mem_reg_24__13_ ( .D(n1289), .CLK(clk), .Q(mem[397]) );
  DFFPOSX1 mem_reg_24__12_ ( .D(n1288), .CLK(clk), .Q(mem[396]) );
  DFFPOSX1 mem_reg_24__11_ ( .D(n1287), .CLK(clk), .Q(mem[395]) );
  DFFPOSX1 mem_reg_24__10_ ( .D(n1286), .CLK(clk), .Q(mem[394]) );
  DFFPOSX1 mem_reg_24__9_ ( .D(n1285), .CLK(clk), .Q(mem[393]) );
  DFFPOSX1 mem_reg_24__8_ ( .D(n1284), .CLK(clk), .Q(mem[392]) );
  DFFPOSX1 mem_reg_24__7_ ( .D(n1283), .CLK(clk), .Q(mem[391]) );
  DFFPOSX1 mem_reg_24__6_ ( .D(n1282), .CLK(clk), .Q(mem[390]) );
  DFFPOSX1 mem_reg_24__5_ ( .D(n1281), .CLK(clk), .Q(mem[389]) );
  DFFPOSX1 mem_reg_24__4_ ( .D(n1280), .CLK(clk), .Q(mem[388]) );
  DFFPOSX1 mem_reg_24__3_ ( .D(n1279), .CLK(clk), .Q(mem[387]) );
  DFFPOSX1 mem_reg_24__2_ ( .D(n1278), .CLK(clk), .Q(mem[386]) );
  DFFPOSX1 mem_reg_24__1_ ( .D(n1277), .CLK(clk), .Q(mem[385]) );
  DFFPOSX1 mem_reg_24__0_ ( .D(n1276), .CLK(clk), .Q(mem[384]) );
  DFFPOSX1 mem_reg_23__15_ ( .D(n1275), .CLK(clk), .Q(mem[383]) );
  DFFPOSX1 mem_reg_23__14_ ( .D(n1274), .CLK(clk), .Q(mem[382]) );
  DFFPOSX1 mem_reg_23__13_ ( .D(n1273), .CLK(clk), .Q(mem[381]) );
  DFFPOSX1 mem_reg_23__12_ ( .D(n1272), .CLK(clk), .Q(mem[380]) );
  DFFPOSX1 mem_reg_23__11_ ( .D(n1271), .CLK(clk), .Q(mem[379]) );
  DFFPOSX1 mem_reg_23__10_ ( .D(n1270), .CLK(clk), .Q(mem[378]) );
  DFFPOSX1 mem_reg_23__9_ ( .D(n1269), .CLK(clk), .Q(mem[377]) );
  DFFPOSX1 mem_reg_23__8_ ( .D(n1268), .CLK(clk), .Q(mem[376]) );
  DFFPOSX1 mem_reg_23__7_ ( .D(n1267), .CLK(clk), .Q(mem[375]) );
  DFFPOSX1 mem_reg_23__6_ ( .D(n1266), .CLK(clk), .Q(mem[374]) );
  DFFPOSX1 mem_reg_23__5_ ( .D(n1265), .CLK(clk), .Q(mem[373]) );
  DFFPOSX1 mem_reg_23__4_ ( .D(n1264), .CLK(clk), .Q(mem[372]) );
  DFFPOSX1 mem_reg_23__3_ ( .D(n1263), .CLK(clk), .Q(mem[371]) );
  DFFPOSX1 mem_reg_23__2_ ( .D(n1262), .CLK(clk), .Q(mem[370]) );
  DFFPOSX1 mem_reg_23__1_ ( .D(n1261), .CLK(clk), .Q(mem[369]) );
  DFFPOSX1 mem_reg_23__0_ ( .D(n1260), .CLK(clk), .Q(mem[368]) );
  DFFPOSX1 mem_reg_22__15_ ( .D(n1259), .CLK(clk), .Q(mem[367]) );
  DFFPOSX1 mem_reg_22__14_ ( .D(n1258), .CLK(clk), .Q(mem[366]) );
  DFFPOSX1 mem_reg_22__13_ ( .D(n1257), .CLK(clk), .Q(mem[365]) );
  DFFPOSX1 mem_reg_22__12_ ( .D(n1256), .CLK(clk), .Q(mem[364]) );
  DFFPOSX1 mem_reg_22__11_ ( .D(n1255), .CLK(clk), .Q(mem[363]) );
  DFFPOSX1 mem_reg_22__10_ ( .D(n1254), .CLK(clk), .Q(mem[362]) );
  DFFPOSX1 mem_reg_22__9_ ( .D(n1253), .CLK(clk), .Q(mem[361]) );
  DFFPOSX1 mem_reg_22__8_ ( .D(n1252), .CLK(clk), .Q(mem[360]) );
  DFFPOSX1 mem_reg_22__7_ ( .D(n1251), .CLK(clk), .Q(mem[359]) );
  DFFPOSX1 mem_reg_22__6_ ( .D(n1250), .CLK(clk), .Q(mem[358]) );
  DFFPOSX1 mem_reg_22__5_ ( .D(n1249), .CLK(clk), .Q(mem[357]) );
  DFFPOSX1 mem_reg_22__4_ ( .D(n1248), .CLK(clk), .Q(mem[356]) );
  DFFPOSX1 mem_reg_22__3_ ( .D(n1247), .CLK(clk), .Q(mem[355]) );
  DFFPOSX1 mem_reg_22__2_ ( .D(n1246), .CLK(clk), .Q(mem[354]) );
  DFFPOSX1 mem_reg_22__1_ ( .D(n1245), .CLK(clk), .Q(mem[353]) );
  DFFPOSX1 mem_reg_22__0_ ( .D(n1244), .CLK(clk), .Q(mem[352]) );
  DFFPOSX1 mem_reg_21__15_ ( .D(n1243), .CLK(clk), .Q(mem[351]) );
  DFFPOSX1 mem_reg_21__14_ ( .D(n1242), .CLK(clk), .Q(mem[350]) );
  DFFPOSX1 mem_reg_21__13_ ( .D(n1241), .CLK(clk), .Q(mem[349]) );
  DFFPOSX1 mem_reg_21__12_ ( .D(n1240), .CLK(clk), .Q(mem[348]) );
  DFFPOSX1 mem_reg_21__11_ ( .D(n1239), .CLK(clk), .Q(mem[347]) );
  DFFPOSX1 mem_reg_21__10_ ( .D(n1238), .CLK(clk), .Q(mem[346]) );
  DFFPOSX1 mem_reg_21__9_ ( .D(n1237), .CLK(clk), .Q(mem[345]) );
  DFFPOSX1 mem_reg_21__8_ ( .D(n1236), .CLK(clk), .Q(mem[344]) );
  DFFPOSX1 mem_reg_21__7_ ( .D(n1235), .CLK(clk), .Q(mem[343]) );
  DFFPOSX1 mem_reg_21__6_ ( .D(n1234), .CLK(clk), .Q(mem[342]) );
  DFFPOSX1 mem_reg_21__5_ ( .D(n1233), .CLK(clk), .Q(mem[341]) );
  DFFPOSX1 mem_reg_21__4_ ( .D(n1232), .CLK(clk), .Q(mem[340]) );
  DFFPOSX1 mem_reg_21__3_ ( .D(n1231), .CLK(clk), .Q(mem[339]) );
  DFFPOSX1 mem_reg_21__2_ ( .D(n1230), .CLK(clk), .Q(mem[338]) );
  DFFPOSX1 mem_reg_21__1_ ( .D(n1229), .CLK(clk), .Q(mem[337]) );
  DFFPOSX1 mem_reg_21__0_ ( .D(n1228), .CLK(clk), .Q(mem[336]) );
  DFFPOSX1 mem_reg_20__15_ ( .D(n1227), .CLK(clk), .Q(mem[335]) );
  DFFPOSX1 mem_reg_20__14_ ( .D(n1226), .CLK(clk), .Q(mem[334]) );
  DFFPOSX1 mem_reg_20__13_ ( .D(n1225), .CLK(clk), .Q(mem[333]) );
  DFFPOSX1 mem_reg_20__12_ ( .D(n1224), .CLK(clk), .Q(mem[332]) );
  DFFPOSX1 mem_reg_20__11_ ( .D(n1223), .CLK(clk), .Q(mem[331]) );
  DFFPOSX1 mem_reg_20__10_ ( .D(n1222), .CLK(clk), .Q(mem[330]) );
  DFFPOSX1 mem_reg_20__9_ ( .D(n1221), .CLK(clk), .Q(mem[329]) );
  DFFPOSX1 mem_reg_20__8_ ( .D(n1220), .CLK(clk), .Q(mem[328]) );
  DFFPOSX1 mem_reg_20__7_ ( .D(n1219), .CLK(clk), .Q(mem[327]) );
  DFFPOSX1 mem_reg_20__6_ ( .D(n1218), .CLK(clk), .Q(mem[326]) );
  DFFPOSX1 mem_reg_20__5_ ( .D(n1217), .CLK(clk), .Q(mem[325]) );
  DFFPOSX1 mem_reg_20__4_ ( .D(n1216), .CLK(clk), .Q(mem[324]) );
  DFFPOSX1 mem_reg_20__3_ ( .D(n1215), .CLK(clk), .Q(mem[323]) );
  DFFPOSX1 mem_reg_20__2_ ( .D(n1214), .CLK(clk), .Q(mem[322]) );
  DFFPOSX1 mem_reg_20__1_ ( .D(n1213), .CLK(clk), .Q(mem[321]) );
  DFFPOSX1 mem_reg_20__0_ ( .D(n1212), .CLK(clk), .Q(mem[320]) );
  DFFPOSX1 mem_reg_19__15_ ( .D(n1211), .CLK(clk), .Q(mem[319]) );
  DFFPOSX1 mem_reg_19__14_ ( .D(n1210), .CLK(clk), .Q(mem[318]) );
  DFFPOSX1 mem_reg_19__13_ ( .D(n1209), .CLK(clk), .Q(mem[317]) );
  DFFPOSX1 mem_reg_19__12_ ( .D(n1208), .CLK(clk), .Q(mem[316]) );
  DFFPOSX1 mem_reg_19__11_ ( .D(n1207), .CLK(clk), .Q(mem[315]) );
  DFFPOSX1 mem_reg_19__10_ ( .D(n1206), .CLK(clk), .Q(mem[314]) );
  DFFPOSX1 mem_reg_19__9_ ( .D(n1205), .CLK(clk), .Q(mem[313]) );
  DFFPOSX1 mem_reg_19__8_ ( .D(n1204), .CLK(clk), .Q(mem[312]) );
  DFFPOSX1 mem_reg_19__7_ ( .D(n1203), .CLK(clk), .Q(mem[311]) );
  DFFPOSX1 mem_reg_19__6_ ( .D(n1202), .CLK(clk), .Q(mem[310]) );
  DFFPOSX1 mem_reg_19__5_ ( .D(n1201), .CLK(clk), .Q(mem[309]) );
  DFFPOSX1 mem_reg_19__4_ ( .D(n1200), .CLK(clk), .Q(mem[308]) );
  DFFPOSX1 mem_reg_19__3_ ( .D(n1199), .CLK(clk), .Q(mem[307]) );
  DFFPOSX1 mem_reg_19__2_ ( .D(n1198), .CLK(clk), .Q(mem[306]) );
  DFFPOSX1 mem_reg_19__1_ ( .D(n1197), .CLK(clk), .Q(mem[305]) );
  DFFPOSX1 mem_reg_19__0_ ( .D(n1196), .CLK(clk), .Q(mem[304]) );
  DFFPOSX1 mem_reg_18__15_ ( .D(n1195), .CLK(clk), .Q(mem[303]) );
  DFFPOSX1 mem_reg_18__14_ ( .D(n1194), .CLK(clk), .Q(mem[302]) );
  DFFPOSX1 mem_reg_18__13_ ( .D(n1193), .CLK(clk), .Q(mem[301]) );
  DFFPOSX1 mem_reg_18__12_ ( .D(n1192), .CLK(clk), .Q(mem[300]) );
  DFFPOSX1 mem_reg_18__11_ ( .D(n1191), .CLK(clk), .Q(mem[299]) );
  DFFPOSX1 mem_reg_18__10_ ( .D(n1190), .CLK(clk), .Q(mem[298]) );
  DFFPOSX1 mem_reg_18__9_ ( .D(n1189), .CLK(clk), .Q(mem[297]) );
  DFFPOSX1 mem_reg_18__8_ ( .D(n1188), .CLK(clk), .Q(mem[296]) );
  DFFPOSX1 mem_reg_18__7_ ( .D(n1187), .CLK(clk), .Q(mem[295]) );
  DFFPOSX1 mem_reg_18__6_ ( .D(n1186), .CLK(clk), .Q(mem[294]) );
  DFFPOSX1 mem_reg_18__5_ ( .D(n1185), .CLK(clk), .Q(mem[293]) );
  DFFPOSX1 mem_reg_18__4_ ( .D(n1184), .CLK(clk), .Q(mem[292]) );
  DFFPOSX1 mem_reg_18__3_ ( .D(n1183), .CLK(clk), .Q(mem[291]) );
  DFFPOSX1 mem_reg_18__2_ ( .D(n1182), .CLK(clk), .Q(mem[290]) );
  DFFPOSX1 mem_reg_18__1_ ( .D(n1181), .CLK(clk), .Q(mem[289]) );
  DFFPOSX1 mem_reg_18__0_ ( .D(n1180), .CLK(clk), .Q(mem[288]) );
  DFFPOSX1 mem_reg_17__15_ ( .D(n1179), .CLK(clk), .Q(mem[287]) );
  DFFPOSX1 mem_reg_17__14_ ( .D(n1178), .CLK(clk), .Q(mem[286]) );
  DFFPOSX1 mem_reg_17__13_ ( .D(n1177), .CLK(clk), .Q(mem[285]) );
  DFFPOSX1 mem_reg_17__12_ ( .D(n1176), .CLK(clk), .Q(mem[284]) );
  DFFPOSX1 mem_reg_17__11_ ( .D(n1175), .CLK(clk), .Q(mem[283]) );
  DFFPOSX1 mem_reg_17__10_ ( .D(n1174), .CLK(clk), .Q(mem[282]) );
  DFFPOSX1 mem_reg_17__9_ ( .D(n1173), .CLK(clk), .Q(mem[281]) );
  DFFPOSX1 mem_reg_17__8_ ( .D(n1172), .CLK(clk), .Q(mem[280]) );
  DFFPOSX1 mem_reg_17__7_ ( .D(n1171), .CLK(clk), .Q(mem[279]) );
  DFFPOSX1 mem_reg_17__6_ ( .D(n1170), .CLK(clk), .Q(mem[278]) );
  DFFPOSX1 mem_reg_17__5_ ( .D(n1169), .CLK(clk), .Q(mem[277]) );
  DFFPOSX1 mem_reg_17__4_ ( .D(n1168), .CLK(clk), .Q(mem[276]) );
  DFFPOSX1 mem_reg_17__3_ ( .D(n1167), .CLK(clk), .Q(mem[275]) );
  DFFPOSX1 mem_reg_17__2_ ( .D(n1166), .CLK(clk), .Q(mem[274]) );
  DFFPOSX1 mem_reg_17__1_ ( .D(n1165), .CLK(clk), .Q(mem[273]) );
  DFFPOSX1 mem_reg_17__0_ ( .D(n1164), .CLK(clk), .Q(mem[272]) );
  DFFPOSX1 mem_reg_16__15_ ( .D(n1163), .CLK(clk), .Q(mem[271]) );
  DFFPOSX1 mem_reg_16__14_ ( .D(n1162), .CLK(clk), .Q(mem[270]) );
  DFFPOSX1 mem_reg_16__13_ ( .D(n1161), .CLK(clk), .Q(mem[269]) );
  DFFPOSX1 mem_reg_16__12_ ( .D(n1160), .CLK(clk), .Q(mem[268]) );
  DFFPOSX1 mem_reg_16__11_ ( .D(n1159), .CLK(clk), .Q(mem[267]) );
  DFFPOSX1 mem_reg_16__10_ ( .D(n1158), .CLK(clk), .Q(mem[266]) );
  DFFPOSX1 mem_reg_16__9_ ( .D(n1157), .CLK(clk), .Q(mem[265]) );
  DFFPOSX1 mem_reg_16__8_ ( .D(n1156), .CLK(clk), .Q(mem[264]) );
  DFFPOSX1 mem_reg_16__7_ ( .D(n1155), .CLK(clk), .Q(mem[263]) );
  DFFPOSX1 mem_reg_16__6_ ( .D(n1154), .CLK(clk), .Q(mem[262]) );
  DFFPOSX1 mem_reg_16__5_ ( .D(n1153), .CLK(clk), .Q(mem[261]) );
  DFFPOSX1 mem_reg_16__4_ ( .D(n1152), .CLK(clk), .Q(mem[260]) );
  DFFPOSX1 mem_reg_16__3_ ( .D(n1151), .CLK(clk), .Q(mem[259]) );
  DFFPOSX1 mem_reg_16__2_ ( .D(n1150), .CLK(clk), .Q(mem[258]) );
  DFFPOSX1 mem_reg_16__1_ ( .D(n1149), .CLK(clk), .Q(mem[257]) );
  DFFPOSX1 mem_reg_16__0_ ( .D(n1148), .CLK(clk), .Q(mem[256]) );
  DFFPOSX1 mem_reg_15__15_ ( .D(n1147), .CLK(clk), .Q(mem[255]) );
  DFFPOSX1 mem_reg_15__14_ ( .D(n1146), .CLK(clk), .Q(mem[254]) );
  DFFPOSX1 mem_reg_15__13_ ( .D(n1145), .CLK(clk), .Q(mem[253]) );
  DFFPOSX1 mem_reg_15__12_ ( .D(n1144), .CLK(clk), .Q(mem[252]) );
  DFFPOSX1 mem_reg_15__11_ ( .D(n1143), .CLK(clk), .Q(mem[251]) );
  DFFPOSX1 mem_reg_15__10_ ( .D(n1142), .CLK(clk), .Q(mem[250]) );
  DFFPOSX1 mem_reg_15__9_ ( .D(n1141), .CLK(clk), .Q(mem[249]) );
  DFFPOSX1 mem_reg_15__8_ ( .D(n1140), .CLK(clk), .Q(mem[248]) );
  DFFPOSX1 mem_reg_15__7_ ( .D(n1139), .CLK(clk), .Q(mem[247]) );
  DFFPOSX1 mem_reg_15__6_ ( .D(n1138), .CLK(clk), .Q(mem[246]) );
  DFFPOSX1 mem_reg_15__5_ ( .D(n1137), .CLK(clk), .Q(mem[245]) );
  DFFPOSX1 mem_reg_15__4_ ( .D(n1136), .CLK(clk), .Q(mem[244]) );
  DFFPOSX1 mem_reg_15__3_ ( .D(n1135), .CLK(clk), .Q(mem[243]) );
  DFFPOSX1 mem_reg_15__2_ ( .D(n1134), .CLK(clk), .Q(mem[242]) );
  DFFPOSX1 mem_reg_15__1_ ( .D(n1133), .CLK(clk), .Q(mem[241]) );
  DFFPOSX1 mem_reg_15__0_ ( .D(n1132), .CLK(clk), .Q(mem[240]) );
  DFFPOSX1 mem_reg_14__15_ ( .D(n1131), .CLK(clk), .Q(mem[239]) );
  DFFPOSX1 mem_reg_14__14_ ( .D(n1130), .CLK(clk), .Q(mem[238]) );
  DFFPOSX1 mem_reg_14__13_ ( .D(n1129), .CLK(clk), .Q(mem[237]) );
  DFFPOSX1 mem_reg_14__12_ ( .D(n1128), .CLK(clk), .Q(mem[236]) );
  DFFPOSX1 mem_reg_14__11_ ( .D(n1127), .CLK(clk), .Q(mem[235]) );
  DFFPOSX1 mem_reg_14__10_ ( .D(n1126), .CLK(clk), .Q(mem[234]) );
  DFFPOSX1 mem_reg_14__9_ ( .D(n1125), .CLK(clk), .Q(mem[233]) );
  DFFPOSX1 mem_reg_14__8_ ( .D(n1124), .CLK(clk), .Q(mem[232]) );
  DFFPOSX1 mem_reg_14__7_ ( .D(n1123), .CLK(clk), .Q(mem[231]) );
  DFFPOSX1 mem_reg_14__6_ ( .D(n1122), .CLK(clk), .Q(mem[230]) );
  DFFPOSX1 mem_reg_14__5_ ( .D(n1121), .CLK(clk), .Q(mem[229]) );
  DFFPOSX1 mem_reg_14__4_ ( .D(n1120), .CLK(clk), .Q(mem[228]) );
  DFFPOSX1 mem_reg_14__3_ ( .D(n1119), .CLK(clk), .Q(mem[227]) );
  DFFPOSX1 mem_reg_14__2_ ( .D(n1118), .CLK(clk), .Q(mem[226]) );
  DFFPOSX1 mem_reg_14__1_ ( .D(n1117), .CLK(clk), .Q(mem[225]) );
  DFFPOSX1 mem_reg_14__0_ ( .D(n1116), .CLK(clk), .Q(mem[224]) );
  DFFPOSX1 mem_reg_13__15_ ( .D(n1115), .CLK(clk), .Q(mem[223]) );
  DFFPOSX1 mem_reg_13__14_ ( .D(n1114), .CLK(clk), .Q(mem[222]) );
  DFFPOSX1 mem_reg_13__13_ ( .D(n1113), .CLK(clk), .Q(mem[221]) );
  DFFPOSX1 mem_reg_13__12_ ( .D(n1112), .CLK(clk), .Q(mem[220]) );
  DFFPOSX1 mem_reg_13__11_ ( .D(n1111), .CLK(clk), .Q(mem[219]) );
  DFFPOSX1 mem_reg_13__10_ ( .D(n1110), .CLK(clk), .Q(mem[218]) );
  DFFPOSX1 mem_reg_13__9_ ( .D(n1109), .CLK(clk), .Q(mem[217]) );
  DFFPOSX1 mem_reg_13__8_ ( .D(n1108), .CLK(clk), .Q(mem[216]) );
  DFFPOSX1 mem_reg_13__7_ ( .D(n1107), .CLK(clk), .Q(mem[215]) );
  DFFPOSX1 mem_reg_13__6_ ( .D(n1106), .CLK(clk), .Q(mem[214]) );
  DFFPOSX1 mem_reg_13__5_ ( .D(n1105), .CLK(clk), .Q(mem[213]) );
  DFFPOSX1 mem_reg_13__4_ ( .D(n1104), .CLK(clk), .Q(mem[212]) );
  DFFPOSX1 mem_reg_13__3_ ( .D(n1103), .CLK(clk), .Q(mem[211]) );
  DFFPOSX1 mem_reg_13__2_ ( .D(n1102), .CLK(clk), .Q(mem[210]) );
  DFFPOSX1 mem_reg_13__1_ ( .D(n1101), .CLK(clk), .Q(mem[209]) );
  DFFPOSX1 mem_reg_13__0_ ( .D(n1100), .CLK(clk), .Q(mem[208]) );
  DFFPOSX1 mem_reg_12__15_ ( .D(n1099), .CLK(clk), .Q(mem[207]) );
  DFFPOSX1 mem_reg_12__14_ ( .D(n1098), .CLK(clk), .Q(mem[206]) );
  DFFPOSX1 mem_reg_12__13_ ( .D(n1097), .CLK(clk), .Q(mem[205]) );
  DFFPOSX1 mem_reg_12__12_ ( .D(n1096), .CLK(clk), .Q(mem[204]) );
  DFFPOSX1 mem_reg_12__11_ ( .D(n1095), .CLK(clk), .Q(mem[203]) );
  DFFPOSX1 mem_reg_12__10_ ( .D(n1094), .CLK(clk), .Q(mem[202]) );
  DFFPOSX1 mem_reg_12__9_ ( .D(n1093), .CLK(clk), .Q(mem[201]) );
  DFFPOSX1 mem_reg_12__8_ ( .D(n1092), .CLK(clk), .Q(mem[200]) );
  DFFPOSX1 mem_reg_12__7_ ( .D(n1091), .CLK(clk), .Q(mem[199]) );
  DFFPOSX1 mem_reg_12__6_ ( .D(n1090), .CLK(clk), .Q(mem[198]) );
  DFFPOSX1 mem_reg_12__5_ ( .D(n1089), .CLK(clk), .Q(mem[197]) );
  DFFPOSX1 mem_reg_12__4_ ( .D(n1088), .CLK(clk), .Q(mem[196]) );
  DFFPOSX1 mem_reg_12__3_ ( .D(n1087), .CLK(clk), .Q(mem[195]) );
  DFFPOSX1 mem_reg_12__2_ ( .D(n1086), .CLK(clk), .Q(mem[194]) );
  DFFPOSX1 mem_reg_12__1_ ( .D(n1085), .CLK(clk), .Q(mem[193]) );
  DFFPOSX1 mem_reg_12__0_ ( .D(n1084), .CLK(clk), .Q(mem[192]) );
  DFFPOSX1 mem_reg_11__15_ ( .D(n1083), .CLK(clk), .Q(mem[191]) );
  DFFPOSX1 mem_reg_11__14_ ( .D(n1082), .CLK(clk), .Q(mem[190]) );
  DFFPOSX1 mem_reg_11__13_ ( .D(n1081), .CLK(clk), .Q(mem[189]) );
  DFFPOSX1 mem_reg_11__12_ ( .D(n1080), .CLK(clk), .Q(mem[188]) );
  DFFPOSX1 mem_reg_11__11_ ( .D(n1079), .CLK(clk), .Q(mem[187]) );
  DFFPOSX1 mem_reg_11__10_ ( .D(n1078), .CLK(clk), .Q(mem[186]) );
  DFFPOSX1 mem_reg_11__9_ ( .D(n1077), .CLK(clk), .Q(mem[185]) );
  DFFPOSX1 mem_reg_11__8_ ( .D(n1076), .CLK(clk), .Q(mem[184]) );
  DFFPOSX1 mem_reg_11__7_ ( .D(n1075), .CLK(clk), .Q(mem[183]) );
  DFFPOSX1 mem_reg_11__6_ ( .D(n1074), .CLK(clk), .Q(mem[182]) );
  DFFPOSX1 mem_reg_11__5_ ( .D(n1073), .CLK(clk), .Q(mem[181]) );
  DFFPOSX1 mem_reg_11__4_ ( .D(n1072), .CLK(clk), .Q(mem[180]) );
  DFFPOSX1 mem_reg_11__3_ ( .D(n1071), .CLK(clk), .Q(mem[179]) );
  DFFPOSX1 mem_reg_11__2_ ( .D(n1070), .CLK(clk), .Q(mem[178]) );
  DFFPOSX1 mem_reg_11__1_ ( .D(n1069), .CLK(clk), .Q(mem[177]) );
  DFFPOSX1 mem_reg_11__0_ ( .D(n1068), .CLK(clk), .Q(mem[176]) );
  DFFPOSX1 mem_reg_10__15_ ( .D(n1067), .CLK(clk), .Q(mem[175]) );
  DFFPOSX1 mem_reg_10__14_ ( .D(n1066), .CLK(clk), .Q(mem[174]) );
  DFFPOSX1 mem_reg_10__13_ ( .D(n1065), .CLK(clk), .Q(mem[173]) );
  DFFPOSX1 mem_reg_10__12_ ( .D(n1064), .CLK(clk), .Q(mem[172]) );
  DFFPOSX1 mem_reg_10__11_ ( .D(n1063), .CLK(clk), .Q(mem[171]) );
  DFFPOSX1 mem_reg_10__10_ ( .D(n1062), .CLK(clk), .Q(mem[170]) );
  DFFPOSX1 mem_reg_10__9_ ( .D(n1061), .CLK(clk), .Q(mem[169]) );
  DFFPOSX1 mem_reg_10__8_ ( .D(n1060), .CLK(clk), .Q(mem[168]) );
  DFFPOSX1 mem_reg_10__7_ ( .D(n1059), .CLK(clk), .Q(mem[167]) );
  DFFPOSX1 mem_reg_10__6_ ( .D(n1058), .CLK(clk), .Q(mem[166]) );
  DFFPOSX1 mem_reg_10__5_ ( .D(n1057), .CLK(clk), .Q(mem[165]) );
  DFFPOSX1 mem_reg_10__4_ ( .D(n1056), .CLK(clk), .Q(mem[164]) );
  DFFPOSX1 mem_reg_10__3_ ( .D(n1055), .CLK(clk), .Q(mem[163]) );
  DFFPOSX1 mem_reg_10__2_ ( .D(n1054), .CLK(clk), .Q(mem[162]) );
  DFFPOSX1 mem_reg_10__1_ ( .D(n1053), .CLK(clk), .Q(mem[161]) );
  DFFPOSX1 mem_reg_10__0_ ( .D(n1052), .CLK(clk), .Q(mem[160]) );
  DFFPOSX1 mem_reg_9__15_ ( .D(n1051), .CLK(clk), .Q(mem[159]) );
  DFFPOSX1 mem_reg_9__14_ ( .D(n1050), .CLK(clk), .Q(mem[158]) );
  DFFPOSX1 mem_reg_9__13_ ( .D(n1049), .CLK(clk), .Q(mem[157]) );
  DFFPOSX1 mem_reg_9__12_ ( .D(n1048), .CLK(clk), .Q(mem[156]) );
  DFFPOSX1 mem_reg_9__11_ ( .D(n1047), .CLK(clk), .Q(mem[155]) );
  DFFPOSX1 mem_reg_9__10_ ( .D(n1046), .CLK(clk), .Q(mem[154]) );
  DFFPOSX1 mem_reg_9__9_ ( .D(n1045), .CLK(clk), .Q(mem[153]) );
  DFFPOSX1 mem_reg_9__8_ ( .D(n1044), .CLK(clk), .Q(mem[152]) );
  DFFPOSX1 mem_reg_9__7_ ( .D(n1043), .CLK(clk), .Q(mem[151]) );
  DFFPOSX1 mem_reg_9__6_ ( .D(n1042), .CLK(clk), .Q(mem[150]) );
  DFFPOSX1 mem_reg_9__5_ ( .D(n1041), .CLK(clk), .Q(mem[149]) );
  DFFPOSX1 mem_reg_9__4_ ( .D(n1040), .CLK(clk), .Q(mem[148]) );
  DFFPOSX1 mem_reg_9__3_ ( .D(n1039), .CLK(clk), .Q(mem[147]) );
  DFFPOSX1 mem_reg_9__2_ ( .D(n1038), .CLK(clk), .Q(mem[146]) );
  DFFPOSX1 mem_reg_9__1_ ( .D(n1037), .CLK(clk), .Q(mem[145]) );
  DFFPOSX1 mem_reg_9__0_ ( .D(n1036), .CLK(clk), .Q(mem[144]) );
  DFFPOSX1 mem_reg_8__15_ ( .D(n1035), .CLK(clk), .Q(mem[143]) );
  DFFPOSX1 mem_reg_8__14_ ( .D(n1034), .CLK(clk), .Q(mem[142]) );
  DFFPOSX1 mem_reg_8__13_ ( .D(n1033), .CLK(clk), .Q(mem[141]) );
  DFFPOSX1 mem_reg_8__12_ ( .D(n1032), .CLK(clk), .Q(mem[140]) );
  DFFPOSX1 mem_reg_8__11_ ( .D(n1031), .CLK(clk), .Q(mem[139]) );
  DFFPOSX1 mem_reg_8__10_ ( .D(n1030), .CLK(clk), .Q(mem[138]) );
  DFFPOSX1 mem_reg_8__9_ ( .D(n1029), .CLK(clk), .Q(mem[137]) );
  DFFPOSX1 mem_reg_8__8_ ( .D(n1028), .CLK(clk), .Q(mem[136]) );
  DFFPOSX1 mem_reg_8__7_ ( .D(n1027), .CLK(clk), .Q(mem[135]) );
  DFFPOSX1 mem_reg_8__6_ ( .D(n1026), .CLK(clk), .Q(mem[134]) );
  DFFPOSX1 mem_reg_8__5_ ( .D(n1025), .CLK(clk), .Q(mem[133]) );
  DFFPOSX1 mem_reg_8__4_ ( .D(n1024), .CLK(clk), .Q(mem[132]) );
  DFFPOSX1 mem_reg_8__3_ ( .D(n1023), .CLK(clk), .Q(mem[131]) );
  DFFPOSX1 mem_reg_8__2_ ( .D(n1022), .CLK(clk), .Q(mem[130]) );
  DFFPOSX1 mem_reg_8__1_ ( .D(n1021), .CLK(clk), .Q(mem[129]) );
  DFFPOSX1 mem_reg_8__0_ ( .D(n1020), .CLK(clk), .Q(mem[128]) );
  DFFPOSX1 mem_reg_7__15_ ( .D(n1019), .CLK(clk), .Q(mem[127]) );
  DFFPOSX1 mem_reg_7__14_ ( .D(n1018), .CLK(clk), .Q(mem[126]) );
  DFFPOSX1 mem_reg_7__13_ ( .D(n1017), .CLK(clk), .Q(mem[125]) );
  DFFPOSX1 mem_reg_7__12_ ( .D(n1016), .CLK(clk), .Q(mem[124]) );
  DFFPOSX1 mem_reg_7__11_ ( .D(n1015), .CLK(clk), .Q(mem[123]) );
  DFFPOSX1 mem_reg_7__10_ ( .D(n1014), .CLK(clk), .Q(mem[122]) );
  DFFPOSX1 mem_reg_7__9_ ( .D(n1013), .CLK(clk), .Q(mem[121]) );
  DFFPOSX1 mem_reg_7__8_ ( .D(n1012), .CLK(clk), .Q(mem[120]) );
  DFFPOSX1 mem_reg_7__7_ ( .D(n1011), .CLK(clk), .Q(mem[119]) );
  DFFPOSX1 mem_reg_7__6_ ( .D(n1010), .CLK(clk), .Q(mem[118]) );
  DFFPOSX1 mem_reg_7__5_ ( .D(n1009), .CLK(clk), .Q(mem[117]) );
  DFFPOSX1 mem_reg_7__4_ ( .D(n1008), .CLK(clk), .Q(mem[116]) );
  DFFPOSX1 mem_reg_7__3_ ( .D(n1007), .CLK(clk), .Q(mem[115]) );
  DFFPOSX1 mem_reg_7__2_ ( .D(n1006), .CLK(clk), .Q(mem[114]) );
  DFFPOSX1 mem_reg_7__1_ ( .D(n1005), .CLK(clk), .Q(mem[113]) );
  DFFPOSX1 mem_reg_7__0_ ( .D(n1004), .CLK(clk), .Q(mem[112]) );
  DFFPOSX1 mem_reg_6__15_ ( .D(n1003), .CLK(clk), .Q(mem[111]) );
  DFFPOSX1 mem_reg_6__14_ ( .D(n1002), .CLK(clk), .Q(mem[110]) );
  DFFPOSX1 mem_reg_6__13_ ( .D(n1001), .CLK(clk), .Q(mem[109]) );
  DFFPOSX1 mem_reg_6__12_ ( .D(n1000), .CLK(clk), .Q(mem[108]) );
  DFFPOSX1 mem_reg_6__11_ ( .D(n999), .CLK(clk), .Q(mem[107]) );
  DFFPOSX1 mem_reg_6__10_ ( .D(n998), .CLK(clk), .Q(mem[106]) );
  DFFPOSX1 mem_reg_6__9_ ( .D(n997), .CLK(clk), .Q(mem[105]) );
  DFFPOSX1 mem_reg_6__8_ ( .D(n996), .CLK(clk), .Q(mem[104]) );
  DFFPOSX1 mem_reg_6__7_ ( .D(n995), .CLK(clk), .Q(mem[103]) );
  DFFPOSX1 mem_reg_6__6_ ( .D(n994), .CLK(clk), .Q(mem[102]) );
  DFFPOSX1 mem_reg_6__5_ ( .D(n993), .CLK(clk), .Q(mem[101]) );
  DFFPOSX1 mem_reg_6__4_ ( .D(n992), .CLK(clk), .Q(mem[100]) );
  DFFPOSX1 mem_reg_6__3_ ( .D(n991), .CLK(clk), .Q(mem[99]) );
  DFFPOSX1 mem_reg_6__2_ ( .D(n990), .CLK(clk), .Q(mem[98]) );
  DFFPOSX1 mem_reg_6__1_ ( .D(n989), .CLK(clk), .Q(mem[97]) );
  DFFPOSX1 mem_reg_6__0_ ( .D(n988), .CLK(clk), .Q(mem[96]) );
  DFFPOSX1 mem_reg_5__15_ ( .D(n987), .CLK(clk), .Q(mem[95]) );
  DFFPOSX1 mem_reg_5__14_ ( .D(n986), .CLK(clk), .Q(mem[94]) );
  DFFPOSX1 mem_reg_5__13_ ( .D(n985), .CLK(clk), .Q(mem[93]) );
  DFFPOSX1 mem_reg_5__12_ ( .D(n984), .CLK(clk), .Q(mem[92]) );
  DFFPOSX1 mem_reg_5__11_ ( .D(n983), .CLK(clk), .Q(mem[91]) );
  DFFPOSX1 mem_reg_5__10_ ( .D(n982), .CLK(clk), .Q(mem[90]) );
  DFFPOSX1 mem_reg_5__9_ ( .D(n981), .CLK(clk), .Q(mem[89]) );
  DFFPOSX1 mem_reg_5__8_ ( .D(n980), .CLK(clk), .Q(mem[88]) );
  DFFPOSX1 mem_reg_5__7_ ( .D(n979), .CLK(clk), .Q(mem[87]) );
  DFFPOSX1 mem_reg_5__6_ ( .D(n978), .CLK(clk), .Q(mem[86]) );
  DFFPOSX1 mem_reg_5__5_ ( .D(n977), .CLK(clk), .Q(mem[85]) );
  DFFPOSX1 mem_reg_5__4_ ( .D(n976), .CLK(clk), .Q(mem[84]) );
  DFFPOSX1 mem_reg_5__3_ ( .D(n975), .CLK(clk), .Q(mem[83]) );
  DFFPOSX1 mem_reg_5__2_ ( .D(n974), .CLK(clk), .Q(mem[82]) );
  DFFPOSX1 mem_reg_5__1_ ( .D(n973), .CLK(clk), .Q(mem[81]) );
  DFFPOSX1 mem_reg_5__0_ ( .D(n972), .CLK(clk), .Q(mem[80]) );
  DFFPOSX1 mem_reg_4__15_ ( .D(n971), .CLK(clk), .Q(mem[79]) );
  DFFPOSX1 mem_reg_4__14_ ( .D(n970), .CLK(clk), .Q(mem[78]) );
  DFFPOSX1 mem_reg_4__13_ ( .D(n969), .CLK(clk), .Q(mem[77]) );
  DFFPOSX1 mem_reg_4__12_ ( .D(n968), .CLK(clk), .Q(mem[76]) );
  DFFPOSX1 mem_reg_4__11_ ( .D(n967), .CLK(clk), .Q(mem[75]) );
  DFFPOSX1 mem_reg_4__10_ ( .D(n966), .CLK(clk), .Q(mem[74]) );
  DFFPOSX1 mem_reg_4__9_ ( .D(n965), .CLK(clk), .Q(mem[73]) );
  DFFPOSX1 mem_reg_4__8_ ( .D(n964), .CLK(clk), .Q(mem[72]) );
  DFFPOSX1 mem_reg_4__7_ ( .D(n963), .CLK(clk), .Q(mem[71]) );
  DFFPOSX1 mem_reg_4__6_ ( .D(n962), .CLK(clk), .Q(mem[70]) );
  DFFPOSX1 mem_reg_4__5_ ( .D(n961), .CLK(clk), .Q(mem[69]) );
  DFFPOSX1 mem_reg_4__4_ ( .D(n960), .CLK(clk), .Q(mem[68]) );
  DFFPOSX1 mem_reg_4__3_ ( .D(n959), .CLK(clk), .Q(mem[67]) );
  DFFPOSX1 mem_reg_4__2_ ( .D(n958), .CLK(clk), .Q(mem[66]) );
  DFFPOSX1 mem_reg_4__1_ ( .D(n957), .CLK(clk), .Q(mem[65]) );
  DFFPOSX1 mem_reg_4__0_ ( .D(n956), .CLK(clk), .Q(mem[64]) );
  DFFPOSX1 mem_reg_3__15_ ( .D(n955), .CLK(clk), .Q(mem[63]) );
  DFFPOSX1 mem_reg_3__14_ ( .D(n954), .CLK(clk), .Q(mem[62]) );
  DFFPOSX1 mem_reg_3__13_ ( .D(n953), .CLK(clk), .Q(mem[61]) );
  DFFPOSX1 mem_reg_3__12_ ( .D(n952), .CLK(clk), .Q(mem[60]) );
  DFFPOSX1 mem_reg_3__11_ ( .D(n951), .CLK(clk), .Q(mem[59]) );
  DFFPOSX1 mem_reg_3__10_ ( .D(n950), .CLK(clk), .Q(mem[58]) );
  DFFPOSX1 mem_reg_3__9_ ( .D(n949), .CLK(clk), .Q(mem[57]) );
  DFFPOSX1 mem_reg_3__8_ ( .D(n948), .CLK(clk), .Q(mem[56]) );
  DFFPOSX1 mem_reg_3__7_ ( .D(n947), .CLK(clk), .Q(mem[55]) );
  DFFPOSX1 mem_reg_3__6_ ( .D(n946), .CLK(clk), .Q(mem[54]) );
  DFFPOSX1 mem_reg_3__5_ ( .D(n945), .CLK(clk), .Q(mem[53]) );
  DFFPOSX1 mem_reg_3__4_ ( .D(n944), .CLK(clk), .Q(mem[52]) );
  DFFPOSX1 mem_reg_3__3_ ( .D(n943), .CLK(clk), .Q(mem[51]) );
  DFFPOSX1 mem_reg_3__2_ ( .D(n942), .CLK(clk), .Q(mem[50]) );
  DFFPOSX1 mem_reg_3__1_ ( .D(n941), .CLK(clk), .Q(mem[49]) );
  DFFPOSX1 mem_reg_3__0_ ( .D(n940), .CLK(clk), .Q(mem[48]) );
  DFFPOSX1 mem_reg_2__15_ ( .D(n939), .CLK(clk), .Q(mem[47]) );
  DFFPOSX1 mem_reg_2__14_ ( .D(n938), .CLK(clk), .Q(mem[46]) );
  DFFPOSX1 mem_reg_2__13_ ( .D(n937), .CLK(clk), .Q(mem[45]) );
  DFFPOSX1 mem_reg_2__12_ ( .D(n936), .CLK(clk), .Q(mem[44]) );
  DFFPOSX1 mem_reg_2__11_ ( .D(n935), .CLK(clk), .Q(mem[43]) );
  DFFPOSX1 mem_reg_2__10_ ( .D(n934), .CLK(clk), .Q(mem[42]) );
  DFFPOSX1 mem_reg_2__9_ ( .D(n933), .CLK(clk), .Q(mem[41]) );
  DFFPOSX1 mem_reg_2__8_ ( .D(n932), .CLK(clk), .Q(mem[40]) );
  DFFPOSX1 mem_reg_2__7_ ( .D(n931), .CLK(clk), .Q(mem[39]) );
  DFFPOSX1 mem_reg_2__6_ ( .D(n930), .CLK(clk), .Q(mem[38]) );
  DFFPOSX1 mem_reg_2__5_ ( .D(n929), .CLK(clk), .Q(mem[37]) );
  DFFPOSX1 mem_reg_2__4_ ( .D(n928), .CLK(clk), .Q(mem[36]) );
  DFFPOSX1 mem_reg_2__3_ ( .D(n927), .CLK(clk), .Q(mem[35]) );
  DFFPOSX1 mem_reg_2__2_ ( .D(n926), .CLK(clk), .Q(mem[34]) );
  DFFPOSX1 mem_reg_2__1_ ( .D(n925), .CLK(clk), .Q(mem[33]) );
  DFFPOSX1 mem_reg_2__0_ ( .D(n924), .CLK(clk), .Q(mem[32]) );
  DFFPOSX1 mem_reg_1__15_ ( .D(n923), .CLK(clk), .Q(mem[31]) );
  DFFPOSX1 mem_reg_1__14_ ( .D(n922), .CLK(clk), .Q(mem[30]) );
  DFFPOSX1 mem_reg_1__13_ ( .D(n921), .CLK(clk), .Q(mem[29]) );
  DFFPOSX1 mem_reg_1__12_ ( .D(n920), .CLK(clk), .Q(mem[28]) );
  DFFPOSX1 mem_reg_1__11_ ( .D(n919), .CLK(clk), .Q(mem[27]) );
  DFFPOSX1 mem_reg_1__10_ ( .D(n918), .CLK(clk), .Q(mem[26]) );
  DFFPOSX1 mem_reg_1__9_ ( .D(n917), .CLK(clk), .Q(mem[25]) );
  DFFPOSX1 mem_reg_1__8_ ( .D(n916), .CLK(clk), .Q(mem[24]) );
  DFFPOSX1 mem_reg_1__7_ ( .D(n915), .CLK(clk), .Q(mem[23]) );
  DFFPOSX1 mem_reg_1__6_ ( .D(n914), .CLK(clk), .Q(mem[22]) );
  DFFPOSX1 mem_reg_1__5_ ( .D(n913), .CLK(clk), .Q(mem[21]) );
  DFFPOSX1 mem_reg_1__4_ ( .D(n912), .CLK(clk), .Q(mem[20]) );
  DFFPOSX1 mem_reg_1__3_ ( .D(n911), .CLK(clk), .Q(mem[19]) );
  DFFPOSX1 mem_reg_1__2_ ( .D(n910), .CLK(clk), .Q(mem[18]) );
  DFFPOSX1 mem_reg_1__1_ ( .D(n909), .CLK(clk), .Q(mem[17]) );
  DFFPOSX1 mem_reg_1__0_ ( .D(n908), .CLK(clk), .Q(mem[16]) );
  DFFPOSX1 mem_reg_0__15_ ( .D(n907), .CLK(clk), .Q(mem[15]) );
  DFFPOSX1 mem_reg_0__14_ ( .D(n906), .CLK(clk), .Q(mem[14]) );
  DFFPOSX1 mem_reg_0__13_ ( .D(n905), .CLK(clk), .Q(mem[13]) );
  DFFPOSX1 mem_reg_0__12_ ( .D(n904), .CLK(clk), .Q(mem[12]) );
  DFFPOSX1 mem_reg_0__11_ ( .D(n903), .CLK(clk), .Q(mem[11]) );
  DFFPOSX1 mem_reg_0__10_ ( .D(n902), .CLK(clk), .Q(mem[10]) );
  DFFPOSX1 mem_reg_0__9_ ( .D(n901), .CLK(clk), .Q(mem[9]) );
  DFFPOSX1 mem_reg_0__8_ ( .D(n900), .CLK(clk), .Q(mem[8]) );
  DFFPOSX1 mem_reg_0__7_ ( .D(n899), .CLK(clk), .Q(mem[7]) );
  DFFPOSX1 mem_reg_0__6_ ( .D(n898), .CLK(clk), .Q(mem[6]) );
  DFFPOSX1 mem_reg_0__5_ ( .D(n897), .CLK(clk), .Q(mem[5]) );
  DFFPOSX1 mem_reg_0__4_ ( .D(n896), .CLK(clk), .Q(mem[4]) );
  DFFPOSX1 mem_reg_0__3_ ( .D(n895), .CLK(clk), .Q(mem[3]) );
  DFFPOSX1 mem_reg_0__2_ ( .D(n894), .CLK(clk), .Q(mem[2]) );
  DFFPOSX1 mem_reg_0__1_ ( .D(n893), .CLK(clk), .Q(mem[1]) );
  DFFPOSX1 mem_reg_0__0_ ( .D(n892), .CLK(clk), .Q(mem[0]) );
  NAND3X1 U583 ( .A(n2544), .B(n543), .C(n544), .Y(n2233) );
  NOR3X1 U584 ( .A(n2818), .B(n2834), .C(n2850), .Y(n544) );
  NAND3X1 U586 ( .A(n1594), .B(n2673), .C(n2802), .Y(n549) );
  AOI22X1 U587 ( .A(n552), .B(n3626), .C(n553), .D(n3578), .Y(n551) );
  NAND3X1 U589 ( .A(n2527), .B(n2672), .C(n2801), .Y(n548) );
  AOI22X1 U590 ( .A(n557), .B(n3658), .C(n558), .D(n3594), .Y(n556) );
  AOI22X1 U592 ( .A(n560), .B(n3674), .C(n561), .D(n3642), .Y(n554) );
  NAND3X1 U594 ( .A(n564), .B(n2671), .C(n2800), .Y(n563) );
  AOI22X1 U595 ( .A(n552), .B(n3498), .C(n3411), .D(n3450), .Y(n566) );
  NAND3X1 U597 ( .A(n2526), .B(n2670), .C(n2799), .Y(n562) );
  AOI22X1 U598 ( .A(n557), .B(n3530), .C(n558), .D(n3466), .Y(n569) );
  AOI22X1 U600 ( .A(n560), .B(n3546), .C(n561), .D(n3514), .Y(n567) );
  NAND3X1 U602 ( .A(n3398), .B(n2669), .C(n2798), .Y(n571) );
  AOI22X1 U603 ( .A(n552), .B(n3882), .C(n3411), .D(n3834), .Y(n574) );
  NAND3X1 U605 ( .A(n2525), .B(n2668), .C(n2797), .Y(n570) );
  AOI22X1 U606 ( .A(n557), .B(n3914), .C(n558), .D(n3850), .Y(n577) );
  AOI22X1 U608 ( .A(n560), .B(n3930), .C(n561), .D(n3898), .Y(n575) );
  NAND3X1 U609 ( .A(n3396), .B(n2667), .C(n2796), .Y(n579) );
  AOI22X1 U610 ( .A(n552), .B(n3754), .C(n553), .D(n3706), .Y(n582) );
  NAND3X1 U612 ( .A(n2524), .B(n2666), .C(n2795), .Y(n578) );
  AOI22X1 U613 ( .A(n557), .B(n3786), .C(n558), .D(n3722), .Y(n585) );
  AOI22X1 U615 ( .A(n560), .B(n3802), .C(n561), .D(n3770), .Y(n583) );
  NAND3X1 U617 ( .A(n2543), .B(n587), .C(n588), .Y(n2234) );
  NOR3X1 U618 ( .A(n2817), .B(n2833), .C(n2849), .Y(n588) );
  NAND3X1 U620 ( .A(n1594), .B(n2665), .C(n2794), .Y(n593) );
  AOI22X1 U621 ( .A(n552), .B(n3627), .C(n553), .D(n3579), .Y(n595) );
  NAND3X1 U623 ( .A(n2523), .B(n2664), .C(n2793), .Y(n592) );
  AOI22X1 U624 ( .A(n557), .B(n3659), .C(n558), .D(n3595), .Y(n598) );
  AOI22X1 U626 ( .A(n560), .B(n3675), .C(n561), .D(n3643), .Y(n596) );
  NAND3X1 U628 ( .A(n564), .B(n2663), .C(n2792), .Y(n600) );
  AOI22X1 U629 ( .A(n552), .B(n3499), .C(n553), .D(n3451), .Y(n602) );
  NAND3X1 U631 ( .A(n2522), .B(n2662), .C(n2791), .Y(n599) );
  AOI22X1 U632 ( .A(n557), .B(n3531), .C(n558), .D(n3467), .Y(n605) );
  AOI22X1 U634 ( .A(n560), .B(n3547), .C(n561), .D(n3515), .Y(n603) );
  NAND3X1 U636 ( .A(n3398), .B(n2661), .C(n2790), .Y(n607) );
  AOI22X1 U637 ( .A(n552), .B(n3883), .C(n553), .D(n3835), .Y(n609) );
  NAND3X1 U639 ( .A(n2521), .B(n2660), .C(n2789), .Y(n606) );
  AOI22X1 U640 ( .A(n557), .B(n3915), .C(n558), .D(n3851), .Y(n612) );
  AOI22X1 U642 ( .A(n560), .B(n3931), .C(n561), .D(n3899), .Y(n610) );
  NAND3X1 U643 ( .A(n3396), .B(n2659), .C(n2788), .Y(n614) );
  AOI22X1 U644 ( .A(n552), .B(n3755), .C(n553), .D(n3707), .Y(n616) );
  NAND3X1 U646 ( .A(n2520), .B(n2658), .C(n2787), .Y(n613) );
  AOI22X1 U647 ( .A(n557), .B(n3787), .C(n558), .D(n3723), .Y(n619) );
  AOI22X1 U649 ( .A(n560), .B(n3803), .C(n561), .D(n3771), .Y(n617) );
  NAND3X1 U651 ( .A(n2542), .B(n621), .C(n622), .Y(n2235) );
  NOR3X1 U652 ( .A(n2816), .B(n2832), .C(n2848), .Y(n622) );
  NAND3X1 U654 ( .A(n1594), .B(n2657), .C(n2786), .Y(n627) );
  AOI22X1 U655 ( .A(n552), .B(n3628), .C(n553), .D(n3580), .Y(n629) );
  NAND3X1 U657 ( .A(n2519), .B(n2656), .C(n2785), .Y(n626) );
  AOI22X1 U658 ( .A(n557), .B(n3660), .C(n558), .D(n3596), .Y(n632) );
  AOI22X1 U660 ( .A(n560), .B(n3676), .C(n561), .D(n3644), .Y(n630) );
  NAND3X1 U662 ( .A(n564), .B(n2655), .C(n2784), .Y(n634) );
  AOI22X1 U663 ( .A(n552), .B(n3500), .C(n553), .D(n3452), .Y(n636) );
  NAND3X1 U665 ( .A(n2518), .B(n2654), .C(n2783), .Y(n633) );
  AOI22X1 U666 ( .A(n557), .B(n3532), .C(n558), .D(n3468), .Y(n639) );
  AOI22X1 U668 ( .A(n3403), .B(n3548), .C(n561), .D(n3516), .Y(n637) );
  NAND3X1 U670 ( .A(n3398), .B(n2653), .C(n2782), .Y(n641) );
  AOI22X1 U671 ( .A(n552), .B(n3884), .C(n3411), .D(n3836), .Y(n643) );
  NAND3X1 U673 ( .A(n2517), .B(n2652), .C(n2781), .Y(n640) );
  AOI22X1 U674 ( .A(n557), .B(n3916), .C(n558), .D(n3852), .Y(n646) );
  AOI22X1 U676 ( .A(n560), .B(n3932), .C(n561), .D(n3900), .Y(n644) );
  NAND3X1 U677 ( .A(n3396), .B(n2651), .C(n2780), .Y(n648) );
  AOI22X1 U678 ( .A(n552), .B(n3756), .C(n553), .D(n3708), .Y(n650) );
  NAND3X1 U680 ( .A(n2516), .B(n2650), .C(n2779), .Y(n647) );
  AOI22X1 U681 ( .A(n557), .B(n3788), .C(n558), .D(n3724), .Y(n653) );
  AOI22X1 U683 ( .A(n560), .B(n3804), .C(n561), .D(n3772), .Y(n651) );
  NAND3X1 U685 ( .A(n2541), .B(n655), .C(n656), .Y(n2236) );
  NOR3X1 U686 ( .A(n2815), .B(n2831), .C(n2847), .Y(n656) );
  NAND3X1 U688 ( .A(n1594), .B(n2649), .C(n2778), .Y(n661) );
  AOI22X1 U689 ( .A(n552), .B(n3629), .C(n553), .D(n3581), .Y(n663) );
  NAND3X1 U691 ( .A(n2515), .B(n2648), .C(n2777), .Y(n660) );
  AOI22X1 U692 ( .A(n557), .B(n3661), .C(n558), .D(n3597), .Y(n666) );
  AOI22X1 U694 ( .A(n560), .B(n3677), .C(n561), .D(n3645), .Y(n664) );
  NAND3X1 U696 ( .A(n564), .B(n2647), .C(n2776), .Y(n668) );
  AOI22X1 U697 ( .A(n552), .B(n3501), .C(n553), .D(n3453), .Y(n670) );
  NAND3X1 U699 ( .A(n2514), .B(n2646), .C(n2775), .Y(n667) );
  AOI22X1 U700 ( .A(n557), .B(n3533), .C(n558), .D(n3469), .Y(n673) );
  AOI22X1 U702 ( .A(n560), .B(n3549), .C(n561), .D(n3517), .Y(n671) );
  NAND3X1 U704 ( .A(n3398), .B(n2645), .C(n2774), .Y(n675) );
  AOI22X1 U705 ( .A(n552), .B(n3885), .C(n3411), .D(n3837), .Y(n677) );
  NAND3X1 U707 ( .A(n2513), .B(n2644), .C(n2773), .Y(n674) );
  AOI22X1 U708 ( .A(n557), .B(n3917), .C(n558), .D(n3853), .Y(n680) );
  AOI22X1 U710 ( .A(n560), .B(n3933), .C(n561), .D(n3901), .Y(n678) );
  NAND3X1 U711 ( .A(n3396), .B(n2643), .C(n2772), .Y(n682) );
  AOI22X1 U712 ( .A(n3413), .B(n3757), .C(n553), .D(n3709), .Y(n684) );
  NAND3X1 U714 ( .A(n2512), .B(n2642), .C(n2771), .Y(n681) );
  AOI22X1 U715 ( .A(n557), .B(n3789), .C(n558), .D(n3725), .Y(n687) );
  AOI22X1 U717 ( .A(n560), .B(n3805), .C(n561), .D(n3773), .Y(n685) );
  NAND3X1 U719 ( .A(n2540), .B(n689), .C(n690), .Y(n2237) );
  NOR3X1 U720 ( .A(n2814), .B(n2830), .C(n2846), .Y(n690) );
  NAND3X1 U722 ( .A(n1594), .B(n2641), .C(n2770), .Y(n695) );
  AOI22X1 U723 ( .A(n3413), .B(n3630), .C(n3411), .D(n3582), .Y(n697) );
  NAND3X1 U725 ( .A(n2511), .B(n2640), .C(n2769), .Y(n694) );
  AOI22X1 U726 ( .A(n557), .B(n3662), .C(n558), .D(n3598), .Y(n700) );
  AOI22X1 U728 ( .A(n560), .B(n3678), .C(n561), .D(n3646), .Y(n698) );
  NAND3X1 U730 ( .A(n564), .B(n2639), .C(n2768), .Y(n702) );
  AOI22X1 U731 ( .A(n552), .B(n3502), .C(n3411), .D(n3454), .Y(n704) );
  NAND3X1 U733 ( .A(n2510), .B(n2638), .C(n2767), .Y(n701) );
  AOI22X1 U734 ( .A(n557), .B(n3534), .C(n558), .D(n3470), .Y(n707) );
  AOI22X1 U736 ( .A(n560), .B(n3550), .C(n561), .D(n3518), .Y(n705) );
  NAND3X1 U738 ( .A(n3398), .B(n2637), .C(n2766), .Y(n709) );
  AOI22X1 U739 ( .A(n552), .B(n3886), .C(n3411), .D(n3838), .Y(n711) );
  NAND3X1 U741 ( .A(n2509), .B(n2636), .C(n2765), .Y(n708) );
  AOI22X1 U742 ( .A(n557), .B(n3918), .C(n558), .D(n3854), .Y(n714) );
  AOI22X1 U744 ( .A(n560), .B(n3934), .C(n561), .D(n3902), .Y(n712) );
  NAND3X1 U745 ( .A(n3396), .B(n2635), .C(n2764), .Y(n716) );
  AOI22X1 U746 ( .A(n3413), .B(n3758), .C(n3411), .D(n3710), .Y(n718) );
  NAND3X1 U748 ( .A(n2508), .B(n2634), .C(n2763), .Y(n715) );
  AOI22X1 U749 ( .A(n557), .B(n3790), .C(n558), .D(n3726), .Y(n721) );
  AOI22X1 U751 ( .A(n560), .B(n3806), .C(n561), .D(n3774), .Y(n719) );
  NAND3X1 U753 ( .A(n2539), .B(n723), .C(n724), .Y(n2238) );
  NOR3X1 U754 ( .A(n2813), .B(n2829), .C(n2845), .Y(n724) );
  NAND3X1 U756 ( .A(n1594), .B(n2633), .C(n2762), .Y(n729) );
  AOI22X1 U757 ( .A(n552), .B(n3631), .C(n3411), .D(n3583), .Y(n731) );
  NAND3X1 U759 ( .A(n2507), .B(n2632), .C(n2761), .Y(n728) );
  AOI22X1 U760 ( .A(n557), .B(n3663), .C(n558), .D(n3599), .Y(n734) );
  AOI22X1 U762 ( .A(n560), .B(n3679), .C(n561), .D(n3647), .Y(n732) );
  NAND3X1 U764 ( .A(n564), .B(n2631), .C(n2760), .Y(n736) );
  AOI22X1 U765 ( .A(n552), .B(n3503), .C(n3411), .D(n3455), .Y(n738) );
  NAND3X1 U767 ( .A(n2506), .B(n2630), .C(n2759), .Y(n735) );
  AOI22X1 U768 ( .A(n557), .B(n3535), .C(n558), .D(n3471), .Y(n741) );
  AOI22X1 U770 ( .A(n560), .B(n3551), .C(n561), .D(n3519), .Y(n739) );
  NAND3X1 U772 ( .A(n3398), .B(n2629), .C(n2758), .Y(n743) );
  AOI22X1 U773 ( .A(n552), .B(n3887), .C(n3411), .D(n3839), .Y(n745) );
  NAND3X1 U775 ( .A(n2505), .B(n2628), .C(n2757), .Y(n742) );
  AOI22X1 U776 ( .A(n557), .B(n3919), .C(n3407), .D(n3855), .Y(n748) );
  AOI22X1 U778 ( .A(n560), .B(n3935), .C(n561), .D(n3903), .Y(n746) );
  NAND3X1 U779 ( .A(n3396), .B(n2627), .C(n2756), .Y(n750) );
  AOI22X1 U780 ( .A(n3413), .B(n3759), .C(n3411), .D(n3711), .Y(n752) );
  NAND3X1 U782 ( .A(n2504), .B(n2626), .C(n2755), .Y(n749) );
  AOI22X1 U783 ( .A(n557), .B(n3791), .C(n558), .D(n3727), .Y(n755) );
  AOI22X1 U785 ( .A(n560), .B(n3807), .C(n561), .D(n3775), .Y(n753) );
  NAND3X1 U787 ( .A(n2538), .B(n757), .C(n758), .Y(n2239) );
  NOR3X1 U788 ( .A(n2812), .B(n2828), .C(n2844), .Y(n758) );
  NAND3X1 U790 ( .A(n1594), .B(n2625), .C(n2754), .Y(n763) );
  AOI22X1 U791 ( .A(n552), .B(n3632), .C(n3411), .D(n3584), .Y(n765) );
  NAND3X1 U793 ( .A(n2503), .B(n2624), .C(n2753), .Y(n762) );
  AOI22X1 U794 ( .A(n557), .B(n3664), .C(n3407), .D(n3600), .Y(n768) );
  AOI22X1 U796 ( .A(n560), .B(n3680), .C(n561), .D(n3648), .Y(n766) );
  NAND3X1 U798 ( .A(n564), .B(n2623), .C(n2752), .Y(n770) );
  AOI22X1 U799 ( .A(n552), .B(n3504), .C(n3411), .D(n3456), .Y(n772) );
  NAND3X1 U801 ( .A(n2502), .B(n2622), .C(n2751), .Y(n769) );
  AOI22X1 U802 ( .A(n557), .B(n3536), .C(n3407), .D(n3472), .Y(n775) );
  AOI22X1 U804 ( .A(n560), .B(n3552), .C(n561), .D(n3520), .Y(n773) );
  NAND3X1 U806 ( .A(n3398), .B(n2621), .C(n2750), .Y(n777) );
  AOI22X1 U807 ( .A(n3413), .B(n3888), .C(n3411), .D(n3840), .Y(n779) );
  NAND3X1 U809 ( .A(n2501), .B(n2620), .C(n2749), .Y(n776) );
  AOI22X1 U810 ( .A(n557), .B(n3920), .C(n3407), .D(n3856), .Y(n782) );
  AOI22X1 U812 ( .A(n560), .B(n3936), .C(n561), .D(n3904), .Y(n780) );
  NAND3X1 U813 ( .A(n3396), .B(n2619), .C(n2748), .Y(n784) );
  AOI22X1 U814 ( .A(n3413), .B(n3760), .C(n3411), .D(n3712), .Y(n786) );
  NAND3X1 U816 ( .A(n2500), .B(n2618), .C(n2747), .Y(n783) );
  AOI22X1 U817 ( .A(n3409), .B(n3792), .C(n3407), .D(n3728), .Y(n789) );
  AOI22X1 U819 ( .A(n560), .B(n3808), .C(n561), .D(n3776), .Y(n787) );
  NAND3X1 U821 ( .A(n2537), .B(n791), .C(n792), .Y(n2240) );
  NOR3X1 U822 ( .A(n2811), .B(n2827), .C(n2843), .Y(n792) );
  NAND3X1 U824 ( .A(n1594), .B(n2617), .C(n2746), .Y(n797) );
  AOI22X1 U825 ( .A(n3413), .B(n3633), .C(n553), .D(n3585), .Y(n799) );
  NAND3X1 U827 ( .A(n2499), .B(n2616), .C(n2745), .Y(n796) );
  AOI22X1 U828 ( .A(n557), .B(n3665), .C(n3407), .D(n3601), .Y(n802) );
  AOI22X1 U830 ( .A(n560), .B(n3681), .C(n561), .D(n3649), .Y(n800) );
  NAND3X1 U832 ( .A(n564), .B(n2615), .C(n2744), .Y(n804) );
  AOI22X1 U833 ( .A(n3413), .B(n3505), .C(n3411), .D(n3457), .Y(n806) );
  NAND3X1 U835 ( .A(n2498), .B(n2614), .C(n2743), .Y(n803) );
  AOI22X1 U836 ( .A(n557), .B(n3537), .C(n3407), .D(n3473), .Y(n809) );
  AOI22X1 U838 ( .A(n560), .B(n3553), .C(n561), .D(n3521), .Y(n807) );
  NAND3X1 U840 ( .A(n3398), .B(n2613), .C(n2742), .Y(n811) );
  AOI22X1 U841 ( .A(n3413), .B(n3889), .C(n553), .D(n3841), .Y(n813) );
  NAND3X1 U843 ( .A(n2497), .B(n2612), .C(n2741), .Y(n810) );
  AOI22X1 U844 ( .A(n557), .B(n3921), .C(n3407), .D(n3857), .Y(n816) );
  AOI22X1 U846 ( .A(n560), .B(n3937), .C(n561), .D(n3905), .Y(n814) );
  NAND3X1 U847 ( .A(n3396), .B(n2611), .C(n2740), .Y(n818) );
  AOI22X1 U848 ( .A(n3413), .B(n3761), .C(n553), .D(n3713), .Y(n820) );
  NAND3X1 U850 ( .A(n2496), .B(n2610), .C(n2739), .Y(n817) );
  AOI22X1 U851 ( .A(n3409), .B(n3793), .C(n3407), .D(n3729), .Y(n823) );
  AOI22X1 U853 ( .A(n560), .B(n3809), .C(n561), .D(n3777), .Y(n821) );
  NAND3X1 U855 ( .A(n2536), .B(n825), .C(n826), .Y(n2241) );
  NOR3X1 U856 ( .A(n2810), .B(n2826), .C(n2842), .Y(n826) );
  NAND3X1 U858 ( .A(n1594), .B(n2609), .C(n2738), .Y(n831) );
  AOI22X1 U859 ( .A(n3413), .B(n3634), .C(n553), .D(n3586), .Y(n833) );
  NAND3X1 U861 ( .A(n2495), .B(n2608), .C(n2737), .Y(n830) );
  AOI22X1 U862 ( .A(n557), .B(n3666), .C(n3407), .D(n3602), .Y(n836) );
  AOI22X1 U864 ( .A(n560), .B(n3682), .C(n561), .D(n3650), .Y(n834) );
  NAND3X1 U866 ( .A(n564), .B(n2607), .C(n2736), .Y(n838) );
  AOI22X1 U867 ( .A(n3413), .B(n3506), .C(n553), .D(n3458), .Y(n840) );
  NAND3X1 U869 ( .A(n2494), .B(n2606), .C(n2735), .Y(n837) );
  AOI22X1 U870 ( .A(n557), .B(n3538), .C(n3407), .D(n3474), .Y(n843) );
  AOI22X1 U872 ( .A(n560), .B(n3554), .C(n561), .D(n3522), .Y(n841) );
  NAND3X1 U874 ( .A(n3397), .B(n2605), .C(n2734), .Y(n845) );
  AOI22X1 U875 ( .A(n3413), .B(n3890), .C(n553), .D(n3842), .Y(n847) );
  NAND3X1 U877 ( .A(n2493), .B(n2604), .C(n2733), .Y(n844) );
  AOI22X1 U878 ( .A(n557), .B(n3922), .C(n3407), .D(n3858), .Y(n850) );
  AOI22X1 U880 ( .A(n560), .B(n3938), .C(n561), .D(n3906), .Y(n848) );
  NAND3X1 U881 ( .A(n3395), .B(n2603), .C(n2732), .Y(n852) );
  AOI22X1 U882 ( .A(n3413), .B(n3762), .C(n553), .D(n3714), .Y(n854) );
  NAND3X1 U884 ( .A(n2492), .B(n2602), .C(n2731), .Y(n851) );
  AOI22X1 U885 ( .A(n3409), .B(n3794), .C(n3407), .D(n3730), .Y(n857) );
  AOI22X1 U887 ( .A(n560), .B(n3810), .C(n561), .D(n3778), .Y(n855) );
  NAND3X1 U889 ( .A(n2535), .B(n859), .C(n860), .Y(n2242) );
  NOR3X1 U890 ( .A(n2809), .B(n2825), .C(n2841), .Y(n860) );
  NAND3X1 U892 ( .A(n1594), .B(n2601), .C(n2730), .Y(n865) );
  AOI22X1 U893 ( .A(n3413), .B(n3635), .C(n553), .D(n3587), .Y(n867) );
  NAND3X1 U895 ( .A(n2491), .B(n2600), .C(n2729), .Y(n864) );
  AOI22X1 U896 ( .A(n557), .B(n3667), .C(n558), .D(n3603), .Y(n870) );
  AOI22X1 U898 ( .A(n560), .B(n3683), .C(n3401), .D(n3651), .Y(n868) );
  NAND3X1 U900 ( .A(n564), .B(n2599), .C(n2728), .Y(n872) );
  AOI22X1 U901 ( .A(n3413), .B(n3507), .C(n3411), .D(n3459), .Y(n874) );
  NAND3X1 U903 ( .A(n2490), .B(n2598), .C(n2727), .Y(n871) );
  AOI22X1 U904 ( .A(n557), .B(n3539), .C(n558), .D(n3475), .Y(n877) );
  AOI22X1 U906 ( .A(n560), .B(n3555), .C(n561), .D(n3523), .Y(n875) );
  NAND3X1 U908 ( .A(n3397), .B(n2597), .C(n2726), .Y(n879) );
  AOI22X1 U909 ( .A(n3413), .B(n3891), .C(n553), .D(n3843), .Y(n881) );
  NAND3X1 U911 ( .A(n2489), .B(n2596), .C(n2725), .Y(n878) );
  AOI22X1 U912 ( .A(n557), .B(n3923), .C(n558), .D(n3859), .Y(n884) );
  AOI22X1 U914 ( .A(n560), .B(n3939), .C(n561), .D(n3907), .Y(n882) );
  NAND3X1 U915 ( .A(n3395), .B(n2595), .C(n2724), .Y(n886) );
  AOI22X1 U916 ( .A(n552), .B(n3763), .C(n553), .D(n3715), .Y(n888) );
  NAND3X1 U918 ( .A(n2488), .B(n2594), .C(n2723), .Y(n885) );
  AOI22X1 U919 ( .A(n3409), .B(n3795), .C(n558), .D(n3731), .Y(n891) );
  AOI22X1 U921 ( .A(n3403), .B(n3811), .C(n3401), .D(n3779), .Y(n889) );
  NAND3X1 U923 ( .A(n2534), .B(n1415), .C(n1416), .Y(n2243) );
  NOR3X1 U924 ( .A(n2808), .B(n2824), .C(n2840), .Y(n1416) );
  NAND3X1 U926 ( .A(n1594), .B(n2593), .C(n2722), .Y(n1421) );
  AOI22X1 U927 ( .A(n552), .B(n3636), .C(n553), .D(n3588), .Y(n1423) );
  NAND3X1 U929 ( .A(n2487), .B(n2592), .C(n2721), .Y(n1420) );
  AOI22X1 U930 ( .A(n3409), .B(n3668), .C(n558), .D(n3604), .Y(n1426) );
  AOI22X1 U932 ( .A(n560), .B(n3684), .C(n3401), .D(n3652), .Y(n1424) );
  NAND3X1 U934 ( .A(n564), .B(n2591), .C(n2720), .Y(n1428) );
  AOI22X1 U935 ( .A(n552), .B(n3508), .C(n553), .D(n3460), .Y(n1430) );
  NAND3X1 U937 ( .A(n2486), .B(n2590), .C(n2719), .Y(n1427) );
  AOI22X1 U938 ( .A(n3409), .B(n3540), .C(n558), .D(n3476), .Y(n1433) );
  AOI22X1 U940 ( .A(n560), .B(n3556), .C(n561), .D(n3524), .Y(n1431) );
  NAND3X1 U942 ( .A(n3397), .B(n2589), .C(n2718), .Y(n1435) );
  AOI22X1 U943 ( .A(n552), .B(n3892), .C(n3411), .D(n3844), .Y(n1437) );
  NAND3X1 U945 ( .A(n2485), .B(n2588), .C(n2717), .Y(n1434) );
  AOI22X1 U946 ( .A(n3409), .B(n3924), .C(n558), .D(n3860), .Y(n1440) );
  AOI22X1 U948 ( .A(n560), .B(n3940), .C(n561), .D(n3908), .Y(n1438) );
  NAND3X1 U949 ( .A(n3395), .B(n2587), .C(n2716), .Y(n1442) );
  AOI22X1 U950 ( .A(n552), .B(n3764), .C(n553), .D(n3716), .Y(n1444) );
  NAND3X1 U952 ( .A(n2484), .B(n2586), .C(n2715), .Y(n1441) );
  AOI22X1 U953 ( .A(n3409), .B(n3796), .C(n558), .D(n3732), .Y(n1447) );
  AOI22X1 U955 ( .A(n3403), .B(n3812), .C(n3401), .D(n3780), .Y(n1445) );
  NAND3X1 U957 ( .A(n2533), .B(n1449), .C(n1450), .Y(n2244) );
  NOR3X1 U958 ( .A(n2807), .B(n2823), .C(n2839), .Y(n1450) );
  NAND3X1 U960 ( .A(n1594), .B(n2585), .C(n2714), .Y(n1455) );
  AOI22X1 U961 ( .A(n552), .B(n3637), .C(n553), .D(n3589), .Y(n1457) );
  NAND3X1 U963 ( .A(n2483), .B(n2584), .C(n2713), .Y(n1454) );
  AOI22X1 U964 ( .A(n3409), .B(n3669), .C(n558), .D(n3605), .Y(n1460) );
  AOI22X1 U966 ( .A(n560), .B(n3685), .C(n561), .D(n3653), .Y(n1458) );
  NAND3X1 U968 ( .A(n564), .B(n2583), .C(n2712), .Y(n1462) );
  AOI22X1 U969 ( .A(n552), .B(n3509), .C(n553), .D(n3461), .Y(n1464) );
  NAND3X1 U971 ( .A(n2482), .B(n2582), .C(n2711), .Y(n1461) );
  AOI22X1 U972 ( .A(n3409), .B(n3541), .C(n558), .D(n3477), .Y(n1467) );
  AOI22X1 U974 ( .A(n560), .B(n3557), .C(n561), .D(n3525), .Y(n1465) );
  NAND3X1 U976 ( .A(n3397), .B(n2581), .C(n2710), .Y(n1469) );
  AOI22X1 U977 ( .A(n552), .B(n3893), .C(n553), .D(n3845), .Y(n1471) );
  NAND3X1 U979 ( .A(n2481), .B(n2580), .C(n2709), .Y(n1468) );
  AOI22X1 U980 ( .A(n3409), .B(n3925), .C(n558), .D(n3861), .Y(n1474) );
  AOI22X1 U982 ( .A(n560), .B(n3941), .C(n561), .D(n3909), .Y(n1472) );
  NAND3X1 U983 ( .A(n3395), .B(n2579), .C(n2708), .Y(n1476) );
  AOI22X1 U984 ( .A(n552), .B(n3765), .C(n553), .D(n3717), .Y(n1478) );
  NAND3X1 U986 ( .A(n2480), .B(n2578), .C(n2707), .Y(n1475) );
  AOI22X1 U987 ( .A(n3409), .B(n3797), .C(n558), .D(n3733), .Y(n1481) );
  AOI22X1 U989 ( .A(n3403), .B(n3813), .C(n3401), .D(n3781), .Y(n1479) );
  NAND3X1 U991 ( .A(n2532), .B(n1483), .C(n1484), .Y(n2245) );
  NOR3X1 U992 ( .A(n2806), .B(n2822), .C(n2838), .Y(n1484) );
  NAND3X1 U994 ( .A(n1594), .B(n2577), .C(n2706), .Y(n1489) );
  AOI22X1 U995 ( .A(n552), .B(n3638), .C(n553), .D(n3590), .Y(n1491) );
  NAND3X1 U997 ( .A(n2479), .B(n2576), .C(n2705), .Y(n1488) );
  AOI22X1 U998 ( .A(n3409), .B(n3670), .C(n3407), .D(n3606), .Y(n1494) );
  AOI22X1 U1000 ( .A(n560), .B(n3686), .C(n3401), .D(n3654), .Y(n1492) );
  NAND3X1 U1002 ( .A(n564), .B(n2575), .C(n2704), .Y(n1496) );
  AOI22X1 U1003 ( .A(n552), .B(n3510), .C(n553), .D(n3462), .Y(n1498) );
  NAND3X1 U1005 ( .A(n2478), .B(n2574), .C(n2703), .Y(n1495) );
  AOI22X1 U1006 ( .A(n3409), .B(n3542), .C(n558), .D(n3478), .Y(n1501) );
  AOI22X1 U1008 ( .A(n560), .B(n3558), .C(n3401), .D(n3526), .Y(n1499) );
  NAND3X1 U1010 ( .A(n3397), .B(n2573), .C(n2702), .Y(n1503) );
  AOI22X1 U1011 ( .A(n552), .B(n3894), .C(n553), .D(n3846), .Y(n1505) );
  NAND3X1 U1013 ( .A(n2477), .B(n2572), .C(n2701), .Y(n1502) );
  AOI22X1 U1014 ( .A(n3409), .B(n3926), .C(n558), .D(n3862), .Y(n1508) );
  AOI22X1 U1016 ( .A(n560), .B(n3942), .C(n3401), .D(n3910), .Y(n1506) );
  NAND3X1 U1017 ( .A(n3395), .B(n2571), .C(n2700), .Y(n1510) );
  AOI22X1 U1018 ( .A(n552), .B(n3766), .C(n553), .D(n3718), .Y(n1512) );
  NAND3X1 U1020 ( .A(n2476), .B(n2570), .C(n2699), .Y(n1509) );
  AOI22X1 U1021 ( .A(n3409), .B(n3798), .C(n3407), .D(n3734), .Y(n1515) );
  AOI22X1 U1023 ( .A(n560), .B(n3814), .C(n3401), .D(n3782), .Y(n1513) );
  NAND3X1 U1025 ( .A(n2531), .B(n1517), .C(n1518), .Y(n2246) );
  NOR3X1 U1026 ( .A(n2805), .B(n2821), .C(n2837), .Y(n1518) );
  NAND3X1 U1028 ( .A(n1594), .B(n2569), .C(n2698), .Y(n1523) );
  AOI22X1 U1029 ( .A(n552), .B(n3639), .C(n3411), .D(n3591), .Y(n1525) );
  NAND3X1 U1031 ( .A(n2475), .B(n2568), .C(n2697), .Y(n1522) );
  AOI22X1 U1032 ( .A(n557), .B(n3671), .C(n558), .D(n3607), .Y(n1528) );
  AOI22X1 U1034 ( .A(n3403), .B(n3687), .C(n3401), .D(n3655), .Y(n1526) );
  NAND3X1 U1036 ( .A(n564), .B(n2567), .C(n2696), .Y(n1530) );
  AOI22X1 U1037 ( .A(n552), .B(n3511), .C(n3411), .D(n3463), .Y(n1532) );
  NAND3X1 U1039 ( .A(n2474), .B(n2566), .C(n2695), .Y(n1529) );
  AOI22X1 U1040 ( .A(n557), .B(n3543), .C(n558), .D(n3479), .Y(n1535) );
  AOI22X1 U1042 ( .A(n3403), .B(n3559), .C(n3401), .D(n3527), .Y(n1533) );
  NAND3X1 U1044 ( .A(n3397), .B(n2565), .C(n2694), .Y(n1537) );
  AOI22X1 U1045 ( .A(n552), .B(n3895), .C(n3411), .D(n3847), .Y(n1539) );
  NAND3X1 U1047 ( .A(n2473), .B(n2564), .C(n2693), .Y(n1536) );
  AOI22X1 U1048 ( .A(n557), .B(n3927), .C(n558), .D(n3863), .Y(n1542) );
  AOI22X1 U1050 ( .A(n3403), .B(n3943), .C(n3401), .D(n3911), .Y(n1540) );
  NAND3X1 U1051 ( .A(n3395), .B(n2563), .C(n2692), .Y(n1544) );
  AOI22X1 U1052 ( .A(n552), .B(n3767), .C(n3411), .D(n3719), .Y(n1546) );
  NAND3X1 U1054 ( .A(n2472), .B(n2562), .C(n2691), .Y(n1543) );
  AOI22X1 U1055 ( .A(n557), .B(n3799), .C(n3407), .D(n3735), .Y(n1549) );
  AOI22X1 U1057 ( .A(n3403), .B(n3815), .C(n3401), .D(n3783), .Y(n1547) );
  NAND3X1 U1059 ( .A(n2530), .B(n1551), .C(n1552), .Y(n2247) );
  NOR3X1 U1060 ( .A(n2804), .B(n2820), .C(n2836), .Y(n1552) );
  NAND3X1 U1062 ( .A(n1594), .B(n2561), .C(n2690), .Y(n1557) );
  AOI22X1 U1063 ( .A(n552), .B(n3640), .C(n3411), .D(n3592), .Y(n1559) );
  NAND3X1 U1065 ( .A(n2471), .B(n2560), .C(n2689), .Y(n1556) );
  AOI22X1 U1066 ( .A(n557), .B(n3672), .C(n558), .D(n3608), .Y(n1562) );
  AOI22X1 U1068 ( .A(n3403), .B(n3688), .C(n3401), .D(n3656), .Y(n1560) );
  NAND3X1 U1070 ( .A(n564), .B(n2559), .C(n2688), .Y(n1564) );
  AOI22X1 U1071 ( .A(n552), .B(n3512), .C(n3411), .D(n3464), .Y(n1566) );
  NAND3X1 U1073 ( .A(n2470), .B(n2558), .C(n2687), .Y(n1563) );
  AOI22X1 U1074 ( .A(n557), .B(n3544), .C(n558), .D(n3480), .Y(n1569) );
  AOI22X1 U1076 ( .A(n3403), .B(n3560), .C(n3401), .D(n3528), .Y(n1567) );
  NAND3X1 U1078 ( .A(n3397), .B(n2557), .C(n2686), .Y(n1571) );
  AOI22X1 U1079 ( .A(n552), .B(n3896), .C(n3411), .D(n3848), .Y(n1573) );
  NAND3X1 U1081 ( .A(n2469), .B(n2556), .C(n2685), .Y(n1570) );
  AOI22X1 U1082 ( .A(n557), .B(n3928), .C(n558), .D(n3864), .Y(n1576) );
  AOI22X1 U1084 ( .A(n3403), .B(n3944), .C(n3401), .D(n3912), .Y(n1574) );
  NAND3X1 U1085 ( .A(n3395), .B(n2555), .C(n2684), .Y(n1578) );
  AOI22X1 U1086 ( .A(n552), .B(n3768), .C(n3411), .D(n3720), .Y(n1580) );
  NAND3X1 U1088 ( .A(n2468), .B(n2554), .C(n2683), .Y(n1577) );
  AOI22X1 U1089 ( .A(n557), .B(n3800), .C(n3407), .D(n3736), .Y(n1583) );
  AOI22X1 U1091 ( .A(n3403), .B(n3816), .C(n3401), .D(n3784), .Y(n1581) );
  NAND3X1 U1093 ( .A(n2529), .B(n1585), .C(n1586), .Y(n2248) );
  NOR3X1 U1094 ( .A(n2803), .B(n2819), .C(n2835), .Y(n1586) );
  NAND3X1 U1096 ( .A(n1594), .B(n2553), .C(n2682), .Y(n1591) );
  AOI22X1 U1097 ( .A(n552), .B(n3641), .C(n3411), .D(n3593), .Y(n1593) );
  NAND3X1 U1099 ( .A(n2467), .B(n2552), .C(n2681), .Y(n1590) );
  AOI22X1 U1100 ( .A(n557), .B(n3673), .C(n558), .D(n3609), .Y(n1597) );
  AOI22X1 U1102 ( .A(n3403), .B(n3689), .C(n561), .D(n3657), .Y(n1595) );
  NAND3X1 U1104 ( .A(n564), .B(n2551), .C(n2680), .Y(n1599) );
  AOI22X1 U1105 ( .A(n552), .B(n3513), .C(n3411), .D(n3465), .Y(n1601) );
  NAND3X1 U1107 ( .A(n2466), .B(n2550), .C(n2679), .Y(n1598) );
  AOI22X1 U1108 ( .A(n557), .B(n3545), .C(n558), .D(n3481), .Y(n1605) );
  AOI22X1 U1110 ( .A(n3403), .B(n3561), .C(n561), .D(n3529), .Y(n1603) );
  NAND3X1 U1112 ( .A(n3397), .B(n2549), .C(n2678), .Y(n1607) );
  AOI22X1 U1113 ( .A(n552), .B(n3897), .C(n3411), .D(n3849), .Y(n1609) );
  NOR3X1 U1115 ( .A(n15), .B(n16), .C(n3344), .Y(n572) );
  NAND3X1 U1116 ( .A(n2465), .B(n2548), .C(n2677), .Y(n1606) );
  AOI22X1 U1117 ( .A(n557), .B(n3929), .C(n558), .D(n3865), .Y(n1613) );
  AOI22X1 U1119 ( .A(n3403), .B(n3945), .C(n561), .D(n3913), .Y(n1611) );
  NAND3X1 U1120 ( .A(n3395), .B(n2547), .C(n2676), .Y(n1615) );
  AOI22X1 U1121 ( .A(n552), .B(n3769), .C(n3411), .D(n3721), .Y(n1617) );
  NOR3X1 U1122 ( .A(n3428), .B(n3399), .C(n3427), .Y(n553) );
  NAND3X1 U1124 ( .A(n2464), .B(n2546), .C(n2675), .Y(n1614) );
  AOI22X1 U1125 ( .A(n557), .B(n3801), .C(n558), .D(n3737), .Y(n1620) );
  AOI22X1 U1127 ( .A(n3403), .B(n3817), .C(n561), .D(n3785), .Y(n1618) );
  AOI21X1 U1129 ( .A(n16), .B(n3296), .C(n3419), .Y(n1624) );
  OAI21X1 U1130 ( .A(n3296), .B(n16), .C(n3430), .Y(n1626) );
  OAI21X1 U1131 ( .A(n1627), .B(n3838), .C(n3014), .Y(n999) );
  OAI21X1 U1133 ( .A(n1627), .B(n3839), .C(n3036), .Y(n998) );
  OAI21X1 U1135 ( .A(n1627), .B(n3840), .C(n3144), .Y(n997) );
  OAI21X1 U1137 ( .A(n1627), .B(n3841), .C(n3186), .Y(n996) );
  OAI21X1 U1139 ( .A(n1627), .B(n3842), .C(n3334), .Y(n995) );
  OAI21X1 U1141 ( .A(n1627), .B(n3843), .C(n3381), .Y(n994) );
  OAI21X1 U1143 ( .A(n1627), .B(n3844), .C(n3238), .Y(n993) );
  OAI21X1 U1145 ( .A(n1627), .B(n3845), .C(n3285), .Y(n992) );
  OAI21X1 U1147 ( .A(n1627), .B(n3846), .C(n3145), .Y(n991) );
  OAI21X1 U1149 ( .A(n1627), .B(n3847), .C(n3187), .Y(n990) );
  OAI21X1 U1151 ( .A(n1627), .B(n3848), .C(n3067), .Y(n989) );
  OAI21X1 U1153 ( .A(n1627), .B(n3849), .C(n3104), .Y(n988) );
  OAI21X1 U1155 ( .A(n1652), .B(n3850), .C(n2901), .Y(n987) );
  OAI21X1 U1157 ( .A(n1652), .B(n3851), .C(n2875), .Y(n986) );
  OAI21X1 U1159 ( .A(n1652), .B(n3852), .C(n3286), .Y(n985) );
  OAI21X1 U1161 ( .A(n1652), .B(n3853), .C(n3239), .Y(n984) );
  OAI21X1 U1163 ( .A(n1652), .B(n3854), .C(n3382), .Y(n983) );
  OAI21X1 U1165 ( .A(n1652), .B(n3855), .C(n3335), .Y(n982) );
  OAI21X1 U1167 ( .A(n1652), .B(n3856), .C(n2953), .Y(n981) );
  OAI21X1 U1169 ( .A(n1652), .B(n3857), .C(n2927), .Y(n980) );
  OAI21X1 U1171 ( .A(n1652), .B(n3858), .C(n3287), .Y(n979) );
  OAI21X1 U1173 ( .A(n1652), .B(n3859), .C(n3240), .Y(n978) );
  OAI21X1 U1175 ( .A(n1652), .B(n3860), .C(n3383), .Y(n977) );
  OAI21X1 U1177 ( .A(n1652), .B(n3861), .C(n3336), .Y(n976) );
  OAI21X1 U1179 ( .A(n1652), .B(n3862), .C(n3105), .Y(n975) );
  OAI21X1 U1181 ( .A(n1652), .B(n3863), .C(n3068), .Y(n974) );
  OAI21X1 U1183 ( .A(n1652), .B(n3864), .C(n3188), .Y(n973) );
  OAI21X1 U1185 ( .A(n1652), .B(n3865), .C(n3146), .Y(n972) );
  OAI21X1 U1187 ( .A(n3345), .B(n3157), .C(n3415), .Y(n1652) );
  OAI21X1 U1188 ( .A(n1675), .B(n3866), .C(n2876), .Y(n971) );
  OAI21X1 U1190 ( .A(n1675), .B(n3867), .C(n2902), .Y(n970) );
  OAI21X1 U1192 ( .A(n1675), .B(n3868), .C(n3241), .Y(n969) );
  OAI21X1 U1194 ( .A(n1675), .B(n3869), .C(n3288), .Y(n968) );
  OAI21X1 U1196 ( .A(n1675), .B(n3870), .C(n3337), .Y(n967) );
  OAI21X1 U1198 ( .A(n1675), .B(n3871), .C(n3384), .Y(n966) );
  OAI21X1 U1200 ( .A(n1675), .B(n3872), .C(n2928), .Y(n965) );
  OAI21X1 U1202 ( .A(n1675), .B(n3873), .C(n2954), .Y(n964) );
  OAI21X1 U1204 ( .A(n1675), .B(n3874), .C(n3242), .Y(n963) );
  OAI21X1 U1206 ( .A(n1675), .B(n3875), .C(n3289), .Y(n962) );
  OAI21X1 U1208 ( .A(n1675), .B(n3876), .C(n3338), .Y(n961) );
  OAI21X1 U1210 ( .A(n1675), .B(n3877), .C(n3385), .Y(n960) );
  OAI21X1 U1212 ( .A(n1675), .B(n3878), .C(n3069), .Y(n959) );
  OAI21X1 U1214 ( .A(n1675), .B(n3879), .C(n3106), .Y(n958) );
  OAI21X1 U1216 ( .A(n1675), .B(n3880), .C(n3147), .Y(n957) );
  OAI21X1 U1218 ( .A(n1675), .B(n3881), .C(n3189), .Y(n956) );
  OAI21X1 U1220 ( .A(n3345), .B(n3299), .C(n3415), .Y(n1675) );
  OAI21X1 U1221 ( .A(n1693), .B(n3882), .C(n3037), .Y(n955) );
  OAI21X1 U1223 ( .A(n1693), .B(n3883), .C(n3015), .Y(n954) );
  OAI21X1 U1225 ( .A(n1693), .B(n3884), .C(n3190), .Y(n953) );
  OAI21X1 U1227 ( .A(n1693), .B(n3885), .C(n3148), .Y(n952) );
  OAI21X1 U1229 ( .A(n1693), .B(n3886), .C(n3107), .Y(n951) );
  OAI21X1 U1231 ( .A(n1693), .B(n3887), .C(n3070), .Y(n950) );
  OAI21X1 U1233 ( .A(n1693), .B(n3888), .C(n2993), .Y(n949) );
  OAI21X1 U1235 ( .A(n1693), .B(n3889), .C(n2972), .Y(n948) );
  OAI21X1 U1237 ( .A(n1693), .B(n3890), .C(n3191), .Y(n947) );
  OAI21X1 U1239 ( .A(n1693), .B(n3891), .C(n3149), .Y(n946) );
  OAI21X1 U1241 ( .A(n1693), .B(n3892), .C(n3108), .Y(n945) );
  OAI21X1 U1243 ( .A(n1693), .B(n3893), .C(n3071), .Y(n944) );
  OAI21X1 U1245 ( .A(n1693), .B(n3894), .C(n3386), .Y(n943) );
  OAI21X1 U1247 ( .A(n1693), .B(n3895), .C(n3339), .Y(n942) );
  OAI21X1 U1249 ( .A(n1693), .B(n3896), .C(n3290), .Y(n941) );
  OAI21X1 U1251 ( .A(n1693), .B(n3897), .C(n3243), .Y(n940) );
  OAI21X1 U1253 ( .A(n3345), .B(n3300), .C(n3415), .Y(n1693) );
  OAI21X1 U1254 ( .A(n1711), .B(n3898), .C(n3016), .Y(n939) );
  OAI21X1 U1256 ( .A(n1711), .B(n3899), .C(n3038), .Y(n938) );
  OAI21X1 U1258 ( .A(n1711), .B(n3900), .C(n3150), .Y(n937) );
  OAI21X1 U1260 ( .A(n1711), .B(n3901), .C(n3192), .Y(n936) );
  OAI21X1 U1262 ( .A(n1711), .B(n3902), .C(n3072), .Y(n935) );
  OAI21X1 U1264 ( .A(n1711), .B(n3903), .C(n3109), .Y(n934) );
  OAI21X1 U1266 ( .A(n1711), .B(n3904), .C(n2973), .Y(n933) );
  OAI21X1 U1268 ( .A(n1711), .B(n3905), .C(n2994), .Y(n932) );
  OAI21X1 U1270 ( .A(n1711), .B(n3906), .C(n3151), .Y(n931) );
  OAI21X1 U1272 ( .A(n1711), .B(n3907), .C(n3193), .Y(n930) );
  OAI21X1 U1274 ( .A(n1711), .B(n3908), .C(n3073), .Y(n929) );
  OAI21X1 U1276 ( .A(n1711), .B(n3909), .C(n3110), .Y(n928) );
  OAI21X1 U1278 ( .A(n1711), .B(n3910), .C(n3340), .Y(n927) );
  OAI21X1 U1280 ( .A(n1711), .B(n3911), .C(n3387), .Y(n926) );
  OAI21X1 U1282 ( .A(n1711), .B(n3912), .C(n3244), .Y(n925) );
  OAI21X1 U1284 ( .A(n1711), .B(n3913), .C(n3291), .Y(n924) );
  OAI21X1 U1286 ( .A(n3345), .B(n3158), .C(n3415), .Y(n1711) );
  OAI21X1 U1287 ( .A(n1729), .B(n3914), .C(n2995), .Y(n923) );
  OAI21X1 U1289 ( .A(n1729), .B(n3915), .C(n2974), .Y(n922) );
  OAI21X1 U1291 ( .A(n1729), .B(n3916), .C(n3111), .Y(n921) );
  OAI21X1 U1293 ( .A(n1729), .B(n3917), .C(n3074), .Y(n920) );
  OAI21X1 U1295 ( .A(n1729), .B(n3918), .C(n3194), .Y(n919) );
  OAI21X1 U1297 ( .A(n1729), .B(n3919), .C(n3152), .Y(n918) );
  OAI21X1 U1299 ( .A(n1729), .B(n3920), .C(n3039), .Y(n917) );
  OAI21X1 U1301 ( .A(n1729), .B(n3921), .C(n3017), .Y(n916) );
  OAI21X1 U1303 ( .A(n1729), .B(n3922), .C(n3112), .Y(n915) );
  OAI21X1 U1305 ( .A(n1729), .B(n3923), .C(n3075), .Y(n914) );
  OAI21X1 U1307 ( .A(n1729), .B(n3924), .C(n3195), .Y(n913) );
  OAI21X1 U1309 ( .A(n1729), .B(n3925), .C(n3153), .Y(n912) );
  OAI21X1 U1311 ( .A(n1729), .B(n3926), .C(n3292), .Y(n911) );
  OAI21X1 U1313 ( .A(n1729), .B(n3927), .C(n3245), .Y(n910) );
  OAI21X1 U1315 ( .A(n1729), .B(n3928), .C(n3388), .Y(n909) );
  OAI21X1 U1317 ( .A(n1729), .B(n3929), .C(n3341), .Y(n908) );
  OAI21X1 U1319 ( .A(n3345), .B(n3203), .C(n3415), .Y(n1729) );
  OAI21X1 U1320 ( .A(n1747), .B(n3930), .C(n2975), .Y(n907) );
  OAI21X1 U1322 ( .A(n1747), .B(n3931), .C(n2996), .Y(n906) );
  OAI21X1 U1324 ( .A(n1747), .B(n3932), .C(n3076), .Y(n905) );
  OAI21X1 U1326 ( .A(n1747), .B(n3933), .C(n3113), .Y(n904) );
  OAI21X1 U1328 ( .A(n1747), .B(n3934), .C(n3154), .Y(n903) );
  OAI21X1 U1330 ( .A(n1747), .B(n3935), .C(n3196), .Y(n902) );
  OAI21X1 U1332 ( .A(n1747), .B(n3936), .C(n3018), .Y(n901) );
  OAI21X1 U1334 ( .A(n1747), .B(n3937), .C(n3040), .Y(n900) );
  OAI21X1 U1336 ( .A(n1747), .B(n3938), .C(n3077), .Y(n899) );
  OAI21X1 U1338 ( .A(n1747), .B(n3939), .C(n3114), .Y(n898) );
  OAI21X1 U1340 ( .A(n1747), .B(n3940), .C(n3155), .Y(n897) );
  OAI21X1 U1342 ( .A(n1747), .B(n3941), .C(n3197), .Y(n896) );
  OAI21X1 U1344 ( .A(n1747), .B(n3942), .C(n3246), .Y(n895) );
  OAI21X1 U1346 ( .A(n1747), .B(n3943), .C(n3293), .Y(n894) );
  OAI21X1 U1348 ( .A(n1747), .B(n3944), .C(n3342), .Y(n893) );
  OAI21X1 U1350 ( .A(n1747), .B(n3945), .C(n3389), .Y(n892) );
  OAI21X1 U1352 ( .A(n3345), .B(n3249), .C(n3415), .Y(n1747) );
  OAI21X1 U1354 ( .A(wr_ptr[0]), .B(n3392), .C(n1766), .Y(n1413) );
  NAND3X1 U1355 ( .A(n2528), .B(n3390), .C(n2674), .Y(n1412) );
  AOI22X1 U1356 ( .A(n1602), .B(n3343), .C(n1777), .D(n16), .Y(n1769) );
  NOR3X1 U1359 ( .A(n3429), .B(n16), .C(n3344), .Y(n580) );
  OAI21X1 U1360 ( .A(n12), .B(n3344), .C(n3198), .Y(n1411) );
  OAI21X1 U1362 ( .A(n3295), .B(n3427), .C(n2334), .Y(n1410) );
  NAND3X1 U1363 ( .A(n3399), .B(n3427), .C(n1610), .Y(n1773) );
  OAI21X1 U1364 ( .A(n3295), .B(n3428), .C(n1774), .Y(n1409) );
  OAI21X1 U1365 ( .A(n552), .B(n1621), .C(n1610), .Y(n1774) );
  AOI21X1 U1366 ( .A(n3426), .B(n1610), .C(n1777), .Y(n1772) );
  OAI21X1 U1367 ( .A(n2545), .B(n3429), .C(n2333), .Y(n1408) );
  NAND3X1 U1368 ( .A(n1610), .B(n3429), .C(n3400), .Y(n1776) );
  AOI21X1 U1369 ( .A(n1610), .B(n3343), .C(n1777), .Y(n1775) );
  NAND3X1 U1370 ( .A(n14), .B(n3399), .C(n13), .Y(n1770) );
  NAND3X1 U1374 ( .A(n1779), .B(n1780), .C(n1781), .Y(n2314) );
  NOR3X1 U1375 ( .A(n1782), .B(fillcount[0]), .C(n1783), .Y(n1781) );
  OAI21X1 U1376 ( .A(n3200), .B(n3430), .C(n3199), .Y(n1407) );
  NAND3X1 U1377 ( .A(n3425), .B(n1765), .C(n3201), .Y(n1785) );
  AOI21X1 U1379 ( .A(n1765), .B(n3433), .C(n1787), .Y(n1784) );
  OAI21X1 U1380 ( .A(n3423), .B(n3431), .C(n3041), .Y(n1406) );
  NAND3X1 U1381 ( .A(wr_ptr[0]), .B(n3431), .C(n1765), .Y(n1788) );
  OAI21X1 U1382 ( .A(n3078), .B(n3432), .C(n1791), .Y(n1405) );
  AOI21X1 U1383 ( .A(n1765), .B(n3431), .C(n1789), .Y(n1790) );
  OAI21X1 U1384 ( .A(wr_ptr[0]), .B(n3392), .C(n3298), .Y(n1789) );
  OAI21X1 U1385 ( .A(n3424), .B(n3433), .C(n3156), .Y(n1404) );
  NAND3X1 U1386 ( .A(n1765), .B(n3433), .C(n3425), .Y(n1792) );
  OAI21X1 U1387 ( .A(n3425), .B(n3392), .C(n3298), .Y(n1787) );
  OAI21X1 U1390 ( .A(n1794), .B(n3434), .C(n3347), .Y(n1403) );
  OAI21X1 U1392 ( .A(n1794), .B(n3435), .C(n3301), .Y(n1402) );
  OAI21X1 U1394 ( .A(n1794), .B(n3436), .C(n2929), .Y(n1401) );
  OAI21X1 U1396 ( .A(n1794), .B(n3437), .C(n2903), .Y(n1400) );
  OAI21X1 U1398 ( .A(n1794), .B(n3438), .C(n2851), .Y(n1399) );
  OAI21X1 U1400 ( .A(n1794), .B(n3439), .C(n2877), .Y(n1398) );
  OAI21X1 U1402 ( .A(n1794), .B(n3440), .C(n3251), .Y(n1397) );
  OAI21X1 U1404 ( .A(n1794), .B(n3441), .C(n3204), .Y(n1396) );
  OAI21X1 U1406 ( .A(n1794), .B(n3442), .C(n2930), .Y(n1395) );
  OAI21X1 U1408 ( .A(n1794), .B(n3443), .C(n2904), .Y(n1394) );
  OAI21X1 U1410 ( .A(n1794), .B(n3444), .C(n2878), .Y(n1393) );
  OAI21X1 U1412 ( .A(n1794), .B(n3445), .C(n2852), .Y(n1392) );
  OAI21X1 U1414 ( .A(n1794), .B(n3446), .C(n3019), .Y(n1391) );
  OAI21X1 U1416 ( .A(n1794), .B(n3447), .C(n2997), .Y(n1390) );
  OAI21X1 U1418 ( .A(n1794), .B(n3448), .C(n2976), .Y(n1389) );
  OAI21X1 U1420 ( .A(n1794), .B(n3449), .C(n2955), .Y(n1388) );
  OAI21X1 U1422 ( .A(n3250), .B(n3346), .C(n3415), .Y(n1794) );
  OAI21X1 U1423 ( .A(n1812), .B(n3450), .C(n3302), .Y(n1387) );
  OAI21X1 U1425 ( .A(n1812), .B(n3451), .C(n3348), .Y(n1386) );
  OAI21X1 U1427 ( .A(n1812), .B(n3452), .C(n2879), .Y(n1385) );
  OAI21X1 U1429 ( .A(n1812), .B(n3453), .C(n2853), .Y(n1384) );
  OAI21X1 U1431 ( .A(n1812), .B(n3454), .C(n2931), .Y(n1383) );
  OAI21X1 U1433 ( .A(n1812), .B(n3455), .C(n2905), .Y(n1382) );
  OAI21X1 U1435 ( .A(n1812), .B(n3456), .C(n3205), .Y(n1381) );
  OAI21X1 U1437 ( .A(n1812), .B(n3457), .C(n3252), .Y(n1380) );
  OAI21X1 U1439 ( .A(n1812), .B(n3458), .C(n2906), .Y(n1379) );
  OAI21X1 U1441 ( .A(n1812), .B(n3459), .C(n2932), .Y(n1378) );
  OAI21X1 U1443 ( .A(n1812), .B(n3460), .C(n2854), .Y(n1377) );
  OAI21X1 U1445 ( .A(n1812), .B(n3461), .C(n2880), .Y(n1376) );
  OAI21X1 U1447 ( .A(n1812), .B(n3462), .C(n2998), .Y(n1375) );
  OAI21X1 U1449 ( .A(n1812), .B(n3463), .C(n3020), .Y(n1374) );
  OAI21X1 U1451 ( .A(n1812), .B(n3464), .C(n2956), .Y(n1373) );
  OAI21X1 U1453 ( .A(n1812), .B(n3465), .C(n2977), .Y(n1372) );
  OAI21X1 U1455 ( .A(n3202), .B(n3346), .C(n3415), .Y(n1812) );
  OAI21X1 U1456 ( .A(n1830), .B(n3466), .C(n3206), .Y(n1371) );
  OAI21X1 U1458 ( .A(n1830), .B(n3467), .C(n3253), .Y(n1370) );
  OAI21X1 U1460 ( .A(n1830), .B(n3468), .C(n2855), .Y(n1369) );
  OAI21X1 U1462 ( .A(n1830), .B(n3469), .C(n2881), .Y(n1368) );
  OAI21X1 U1464 ( .A(n1830), .B(n3470), .C(n2907), .Y(n1367) );
  OAI21X1 U1466 ( .A(n1830), .B(n3471), .C(n2933), .Y(n1366) );
  OAI21X1 U1468 ( .A(n1830), .B(n3472), .C(n3349), .Y(n1365) );
  OAI21X1 U1470 ( .A(n1830), .B(n3473), .C(n3303), .Y(n1364) );
  OAI21X1 U1472 ( .A(n1830), .B(n3474), .C(n2882), .Y(n1363) );
  OAI21X1 U1474 ( .A(n1830), .B(n3475), .C(n2856), .Y(n1362) );
  OAI21X1 U1476 ( .A(n1830), .B(n3476), .C(n2934), .Y(n1361) );
  OAI21X1 U1478 ( .A(n1830), .B(n3477), .C(n2908), .Y(n1360) );
  OAI21X1 U1480 ( .A(n1830), .B(n3478), .C(n2978), .Y(n1359) );
  OAI21X1 U1482 ( .A(n1830), .B(n3479), .C(n2957), .Y(n1358) );
  OAI21X1 U1484 ( .A(n1830), .B(n3480), .C(n3021), .Y(n1357) );
  OAI21X1 U1486 ( .A(n1830), .B(n3481), .C(n2999), .Y(n1356) );
  OAI21X1 U1488 ( .A(n3157), .B(n3346), .C(n3415), .Y(n1830) );
  OAI21X1 U1489 ( .A(n1847), .B(n3482), .C(n3159), .Y(n1355) );
  OAI21X1 U1491 ( .A(n1847), .B(n3483), .C(n3117), .Y(n1354) );
  OAI21X1 U1493 ( .A(n1847), .B(n3484), .C(n2909), .Y(n1353) );
  OAI21X1 U1495 ( .A(n1847), .B(n3485), .C(n2935), .Y(n1352) );
  OAI21X1 U1497 ( .A(n1847), .B(n3486), .C(n3254), .Y(n1351) );
  OAI21X1 U1499 ( .A(n1847), .B(n3487), .C(n3207), .Y(n1350) );
  OAI21X1 U1501 ( .A(n1847), .B(n3488), .C(n3304), .Y(n1349) );
  OAI21X1 U1503 ( .A(n1847), .B(n3489), .C(n3350), .Y(n1348) );
  OAI21X1 U1505 ( .A(n1847), .B(n3490), .C(n2857), .Y(n1347) );
  OAI21X1 U1507 ( .A(n1847), .B(n3491), .C(n2883), .Y(n1346) );
  OAI21X1 U1509 ( .A(n1847), .B(n3492), .C(n2910), .Y(n1345) );
  OAI21X1 U1511 ( .A(n1847), .B(n3493), .C(n2936), .Y(n1344) );
  OAI21X1 U1513 ( .A(n1847), .B(n3494), .C(n2958), .Y(n1343) );
  OAI21X1 U1515 ( .A(n1847), .B(n3495), .C(n2979), .Y(n1342) );
  OAI21X1 U1517 ( .A(n1847), .B(n3496), .C(n3000), .Y(n1341) );
  OAI21X1 U1519 ( .A(n1847), .B(n3497), .C(n3022), .Y(n1340) );
  OAI21X1 U1521 ( .A(n3299), .B(n3346), .C(n3415), .Y(n1847) );
  OAI21X1 U1522 ( .A(n1864), .B(n3498), .C(n2911), .Y(n1339) );
  OAI21X1 U1524 ( .A(n1864), .B(n3499), .C(n2937), .Y(n1338) );
  OAI21X1 U1526 ( .A(n1864), .B(n3500), .C(n3351), .Y(n1337) );
  OAI21X1 U1528 ( .A(n1864), .B(n3501), .C(n3305), .Y(n1336) );
  OAI21X1 U1530 ( .A(n1864), .B(n3502), .C(n3208), .Y(n1335) );
  OAI21X1 U1532 ( .A(n1864), .B(n3503), .C(n3255), .Y(n1334) );
  OAI21X1 U1534 ( .A(n1864), .B(n3504), .C(n2858), .Y(n1333) );
  OAI21X1 U1536 ( .A(n1864), .B(n3505), .C(n2884), .Y(n1332) );
  OAI21X1 U1538 ( .A(n1864), .B(n3506), .C(n3352), .Y(n1331) );
  OAI21X1 U1540 ( .A(n1864), .B(n3507), .C(n3306), .Y(n1330) );
  OAI21X1 U1542 ( .A(n1864), .B(n3508), .C(n3256), .Y(n1329) );
  OAI21X1 U1544 ( .A(n1864), .B(n3509), .C(n3209), .Y(n1328) );
  OAI21X1 U1546 ( .A(n1864), .B(n3510), .C(n3160), .Y(n1327) );
  OAI21X1 U1548 ( .A(n1864), .B(n3511), .C(n3118), .Y(n1326) );
  OAI21X1 U1550 ( .A(n1864), .B(n3512), .C(n3079), .Y(n1325) );
  OAI21X1 U1552 ( .A(n1864), .B(n3513), .C(n3042), .Y(n1324) );
  OAI21X1 U1554 ( .A(n3300), .B(n3346), .C(n3415), .Y(n1864) );
  OAI21X1 U1555 ( .A(n1881), .B(n3514), .C(n3119), .Y(n1323) );
  OAI21X1 U1557 ( .A(n1881), .B(n3515), .C(n3161), .Y(n1322) );
  OAI21X1 U1559 ( .A(n1881), .B(n3516), .C(n3307), .Y(n1321) );
  OAI21X1 U1561 ( .A(n1881), .B(n3517), .C(n3353), .Y(n1320) );
  OAI21X1 U1563 ( .A(n1881), .B(n3518), .C(n2885), .Y(n1319) );
  OAI21X1 U1565 ( .A(n1881), .B(n3519), .C(n2859), .Y(n1318) );
  OAI21X1 U1567 ( .A(n1881), .B(n3520), .C(n3257), .Y(n1317) );
  OAI21X1 U1569 ( .A(n1881), .B(n3521), .C(n3210), .Y(n1316) );
  OAI21X1 U1571 ( .A(n1881), .B(n3522), .C(n2938), .Y(n1315) );
  OAI21X1 U1573 ( .A(n1881), .B(n3523), .C(n2912), .Y(n1314) );
  OAI21X1 U1575 ( .A(n1881), .B(n3524), .C(n2886), .Y(n1313) );
  OAI21X1 U1577 ( .A(n1881), .B(n3525), .C(n2860), .Y(n1312) );
  OAI21X1 U1579 ( .A(n1881), .B(n3526), .C(n3023), .Y(n1311) );
  OAI21X1 U1581 ( .A(n1881), .B(n3527), .C(n3001), .Y(n1310) );
  OAI21X1 U1583 ( .A(n1881), .B(n3528), .C(n2980), .Y(n1309) );
  OAI21X1 U1585 ( .A(n1881), .B(n3529), .C(n2959), .Y(n1308) );
  OAI21X1 U1587 ( .A(n3158), .B(n3346), .C(n3415), .Y(n1881) );
  OAI21X1 U1588 ( .A(n1898), .B(n3530), .C(n3354), .Y(n1307) );
  OAI21X1 U1590 ( .A(n1898), .B(n3531), .C(n3308), .Y(n1306) );
  OAI21X1 U1592 ( .A(n1898), .B(n3532), .C(n2913), .Y(n1305) );
  OAI21X1 U1594 ( .A(n1898), .B(n3533), .C(n2939), .Y(n1304) );
  OAI21X1 U1596 ( .A(n1898), .B(n3534), .C(n2861), .Y(n1303) );
  OAI21X1 U1598 ( .A(n1898), .B(n3535), .C(n2887), .Y(n1302) );
  OAI21X1 U1600 ( .A(n1898), .B(n3536), .C(n3211), .Y(n1301) );
  OAI21X1 U1602 ( .A(n1898), .B(n3537), .C(n3258), .Y(n1300) );
  OAI21X1 U1604 ( .A(n1898), .B(n3538), .C(n2914), .Y(n1299) );
  OAI21X1 U1606 ( .A(n1898), .B(n3539), .C(n2940), .Y(n1298) );
  OAI21X1 U1608 ( .A(n1898), .B(n3540), .C(n2862), .Y(n1297) );
  OAI21X1 U1610 ( .A(n1898), .B(n3541), .C(n2888), .Y(n1296) );
  OAI21X1 U1612 ( .A(n1898), .B(n3542), .C(n3002), .Y(n1295) );
  OAI21X1 U1614 ( .A(n1898), .B(n3543), .C(n3024), .Y(n1294) );
  OAI21X1 U1616 ( .A(n1898), .B(n3544), .C(n2960), .Y(n1293) );
  OAI21X1 U1618 ( .A(n1898), .B(n3545), .C(n2981), .Y(n1292) );
  OAI21X1 U1620 ( .A(n3203), .B(n3346), .C(n3415), .Y(n1898) );
  OAI21X1 U1621 ( .A(n1915), .B(n3546), .C(n3259), .Y(n1291) );
  OAI21X1 U1623 ( .A(n1915), .B(n3547), .C(n3212), .Y(n1290) );
  OAI21X1 U1625 ( .A(n1915), .B(n3548), .C(n2889), .Y(n1289) );
  OAI21X1 U1627 ( .A(n1915), .B(n3549), .C(n2863), .Y(n1288) );
  OAI21X1 U1629 ( .A(n1915), .B(n3550), .C(n2941), .Y(n1287) );
  OAI21X1 U1631 ( .A(n1915), .B(n3551), .C(n2915), .Y(n1286) );
  OAI21X1 U1633 ( .A(n1915), .B(n3552), .C(n3355), .Y(n1285) );
  OAI21X1 U1635 ( .A(n1915), .B(n3553), .C(n3309), .Y(n1284) );
  OAI21X1 U1637 ( .A(n1915), .B(n3554), .C(n2890), .Y(n1283) );
  OAI21X1 U1639 ( .A(n1915), .B(n3555), .C(n2864), .Y(n1282) );
  OAI21X1 U1641 ( .A(n1915), .B(n3556), .C(n2942), .Y(n1281) );
  OAI21X1 U1643 ( .A(n1915), .B(n3557), .C(n2916), .Y(n1280) );
  OAI21X1 U1645 ( .A(n1915), .B(n3558), .C(n2982), .Y(n1279) );
  OAI21X1 U1647 ( .A(n1915), .B(n3559), .C(n2961), .Y(n1278) );
  OAI21X1 U1649 ( .A(n1915), .B(n3560), .C(n3025), .Y(n1277) );
  OAI21X1 U1651 ( .A(n1915), .B(n3561), .C(n3003), .Y(n1276) );
  OAI21X1 U1653 ( .A(n3249), .B(n3346), .C(n3415), .Y(n1915) );
  NAND3X1 U1654 ( .A(wr_ptr[4]), .B(wr_ptr[3]), .C(put), .Y(n1811) );
  OAI21X1 U1655 ( .A(n1932), .B(n3562), .C(n3213), .Y(n1275) );
  OAI21X1 U1657 ( .A(n1932), .B(n3563), .C(n3260), .Y(n1274) );
  OAI21X1 U1659 ( .A(n1932), .B(n3564), .C(n2865), .Y(n1273) );
  OAI21X1 U1661 ( .A(n1932), .B(n3565), .C(n2891), .Y(n1272) );
  OAI21X1 U1663 ( .A(n1932), .B(n3566), .C(n2917), .Y(n1271) );
  OAI21X1 U1665 ( .A(n1932), .B(n3567), .C(n2943), .Y(n1270) );
  OAI21X1 U1667 ( .A(n1932), .B(n3568), .C(n3310), .Y(n1269) );
  OAI21X1 U1669 ( .A(n1932), .B(n3569), .C(n3356), .Y(n1268) );
  OAI21X1 U1671 ( .A(n1932), .B(n3570), .C(n2866), .Y(n1267) );
  OAI21X1 U1673 ( .A(n1932), .B(n3571), .C(n2892), .Y(n1266) );
  OAI21X1 U1675 ( .A(n1932), .B(n3572), .C(n2918), .Y(n1265) );
  OAI21X1 U1677 ( .A(n1932), .B(n3573), .C(n2944), .Y(n1264) );
  OAI21X1 U1679 ( .A(n1932), .B(n3574), .C(n2962), .Y(n1263) );
  OAI21X1 U1681 ( .A(n1932), .B(n3575), .C(n2983), .Y(n1262) );
  OAI21X1 U1683 ( .A(n1932), .B(n3576), .C(n3004), .Y(n1261) );
  OAI21X1 U1685 ( .A(n1932), .B(n3577), .C(n3026), .Y(n1260) );
  OAI21X1 U1687 ( .A(n3250), .B(n3393), .C(n3415), .Y(n1932) );
  OAI21X1 U1688 ( .A(n1950), .B(n3578), .C(n2335), .Y(n1259) );
  OAI21X1 U1690 ( .A(n1950), .B(n3579), .C(n3357), .Y(n1258) );
  OAI21X1 U1692 ( .A(n1950), .B(n3580), .C(n3005), .Y(n1257) );
  OAI21X1 U1694 ( .A(n1950), .B(n3581), .C(n3027), .Y(n1256) );
  OAI21X1 U1696 ( .A(n1950), .B(n3582), .C(n3261), .Y(n1255) );
  OAI21X1 U1698 ( .A(n1950), .B(n3583), .C(n3214), .Y(n1254) );
  OAI21X1 U1700 ( .A(n1950), .B(n3584), .C(n2893), .Y(n1253) );
  OAI21X1 U1702 ( .A(n1950), .B(n3585), .C(n2867), .Y(n1252) );
  OAI21X1 U1704 ( .A(n1950), .B(n3586), .C(n3358), .Y(n1251) );
  OAI21X1 U1706 ( .A(n1950), .B(n3587), .C(n3311), .Y(n1250) );
  OAI21X1 U1708 ( .A(n1950), .B(n3588), .C(n3262), .Y(n1249) );
  OAI21X1 U1710 ( .A(n1950), .B(n3589), .C(n3215), .Y(n1248) );
  OAI21X1 U1712 ( .A(n1950), .B(n3590), .C(n3162), .Y(n1247) );
  OAI21X1 U1714 ( .A(n1950), .B(n3591), .C(n3120), .Y(n1246) );
  OAI21X1 U1716 ( .A(n1950), .B(n3592), .C(n3080), .Y(n1245) );
  OAI21X1 U1718 ( .A(n1950), .B(n3593), .C(n3043), .Y(n1244) );
  OAI21X1 U1720 ( .A(n3202), .B(n3393), .C(n3415), .Y(n1950) );
  OAI21X1 U1721 ( .A(n1967), .B(n3594), .C(n2945), .Y(n1243) );
  OAI21X1 U1723 ( .A(n1967), .B(n3595), .C(n2919), .Y(n1242) );
  OAI21X1 U1725 ( .A(n1967), .B(n3596), .C(n3359), .Y(n1241) );
  OAI21X1 U1727 ( .A(n1967), .B(n3597), .C(n3312), .Y(n1240) );
  OAI21X1 U1729 ( .A(n1967), .B(n3598), .C(n3216), .Y(n1239) );
  OAI21X1 U1731 ( .A(n1967), .B(n3599), .C(n3263), .Y(n1238) );
  OAI21X1 U1733 ( .A(n1967), .B(n3600), .C(n2868), .Y(n1237) );
  OAI21X1 U1735 ( .A(n1967), .B(n3601), .C(n2894), .Y(n1236) );
  OAI21X1 U1737 ( .A(n1967), .B(n3602), .C(n3313), .Y(n1235) );
  OAI21X1 U1739 ( .A(n1967), .B(n3603), .C(n3360), .Y(n1234) );
  OAI21X1 U1741 ( .A(n1967), .B(n3604), .C(n3217), .Y(n1233) );
  OAI21X1 U1743 ( .A(n1967), .B(n3605), .C(n3264), .Y(n1232) );
  OAI21X1 U1745 ( .A(n1967), .B(n3606), .C(n3121), .Y(n1231) );
  OAI21X1 U1747 ( .A(n1967), .B(n3607), .C(n3163), .Y(n1230) );
  OAI21X1 U1749 ( .A(n1967), .B(n3608), .C(n3044), .Y(n1229) );
  OAI21X1 U1751 ( .A(n1967), .B(n3609), .C(n3081), .Y(n1228) );
  OAI21X1 U1753 ( .A(n3157), .B(n3393), .C(n3415), .Y(n1967) );
  OAI21X1 U1754 ( .A(n1984), .B(n3610), .C(n2895), .Y(n1227) );
  OAI21X1 U1756 ( .A(n1984), .B(n3611), .C(n2869), .Y(n1226) );
  OAI21X1 U1758 ( .A(n1984), .B(n3612), .C(n3265), .Y(n1225) );
  OAI21X1 U1760 ( .A(n1984), .B(n3613), .C(n3218), .Y(n1224) );
  OAI21X1 U1762 ( .A(n1984), .B(n3614), .C(n3361), .Y(n1223) );
  OAI21X1 U1764 ( .A(n1984), .B(n3615), .C(n3314), .Y(n1222) );
  OAI21X1 U1766 ( .A(n1984), .B(n3616), .C(n2946), .Y(n1221) );
  OAI21X1 U1768 ( .A(n1984), .B(n3617), .C(n2920), .Y(n1220) );
  OAI21X1 U1770 ( .A(n1984), .B(n3618), .C(n3266), .Y(n1219) );
  OAI21X1 U1772 ( .A(n1984), .B(n3619), .C(n3219), .Y(n1218) );
  OAI21X1 U1774 ( .A(n1984), .B(n3620), .C(n3362), .Y(n1217) );
  OAI21X1 U1776 ( .A(n1984), .B(n3621), .C(n3315), .Y(n1216) );
  OAI21X1 U1778 ( .A(n1984), .B(n3622), .C(n3082), .Y(n1215) );
  OAI21X1 U1780 ( .A(n1984), .B(n3623), .C(n3045), .Y(n1214) );
  OAI21X1 U1782 ( .A(n1984), .B(n3624), .C(n3164), .Y(n1213) );
  OAI21X1 U1784 ( .A(n1984), .B(n3625), .C(n3122), .Y(n1212) );
  OAI21X1 U1786 ( .A(n3299), .B(n3393), .C(n3415), .Y(n1984) );
  OAI21X1 U1787 ( .A(n2001), .B(n3626), .C(n2870), .Y(n1211) );
  OAI21X1 U1789 ( .A(n2001), .B(n3627), .C(n2896), .Y(n1210) );
  OAI21X1 U1791 ( .A(n2001), .B(n3628), .C(n3220), .Y(n1209) );
  OAI21X1 U1793 ( .A(n2001), .B(n3629), .C(n3267), .Y(n1208) );
  OAI21X1 U1795 ( .A(n2001), .B(n3630), .C(n3316), .Y(n1207) );
  OAI21X1 U1797 ( .A(n2001), .B(n3631), .C(n3363), .Y(n1206) );
  OAI21X1 U1799 ( .A(n2001), .B(n3632), .C(n2921), .Y(n1205) );
  OAI21X1 U1801 ( .A(n2001), .B(n3633), .C(n2947), .Y(n1204) );
  OAI21X1 U1803 ( .A(n2001), .B(n3634), .C(n3221), .Y(n1203) );
  OAI21X1 U1805 ( .A(n2001), .B(n3635), .C(n3268), .Y(n1202) );
  OAI21X1 U1807 ( .A(n2001), .B(n3636), .C(n3317), .Y(n1201) );
  OAI21X1 U1809 ( .A(n2001), .B(n3637), .C(n3364), .Y(n1200) );
  OAI21X1 U1811 ( .A(n2001), .B(n3638), .C(n3046), .Y(n1199) );
  OAI21X1 U1813 ( .A(n2001), .B(n3639), .C(n3083), .Y(n1198) );
  OAI21X1 U1815 ( .A(n2001), .B(n3640), .C(n3123), .Y(n1197) );
  OAI21X1 U1817 ( .A(n2001), .B(n3641), .C(n3165), .Y(n1196) );
  OAI21X1 U1819 ( .A(n3300), .B(n3393), .C(n3415), .Y(n2001) );
  OAI21X1 U1820 ( .A(n2018), .B(n3642), .C(n2922), .Y(n1195) );
  OAI21X1 U1822 ( .A(n2018), .B(n3643), .C(n2948), .Y(n1194) );
  OAI21X1 U1824 ( .A(n2018), .B(n3644), .C(n3166), .Y(n1193) );
  OAI21X1 U1826 ( .A(n2018), .B(n3645), .C(n3124), .Y(n1192) );
  OAI21X1 U1828 ( .A(n2018), .B(n3646), .C(n3084), .Y(n1191) );
  OAI21X1 U1830 ( .A(n2018), .B(n3647), .C(n3047), .Y(n1190) );
  OAI21X1 U1832 ( .A(n2018), .B(n3648), .C(n2984), .Y(n1189) );
  OAI21X1 U1834 ( .A(n2018), .B(n3649), .C(n2963), .Y(n1188) );
  OAI21X1 U1836 ( .A(n2018), .B(n3650), .C(n3167), .Y(n1187) );
  OAI21X1 U1838 ( .A(n2018), .B(n3651), .C(n3125), .Y(n1186) );
  OAI21X1 U1840 ( .A(n2018), .B(n3652), .C(n3085), .Y(n1185) );
  OAI21X1 U1842 ( .A(n2018), .B(n3653), .C(n3048), .Y(n1184) );
  OAI21X1 U1844 ( .A(n2018), .B(n3654), .C(n3365), .Y(n1183) );
  OAI21X1 U1846 ( .A(n2018), .B(n3655), .C(n3318), .Y(n1182) );
  OAI21X1 U1848 ( .A(n2018), .B(n3656), .C(n3269), .Y(n1181) );
  OAI21X1 U1850 ( .A(n2018), .B(n3657), .C(n3222), .Y(n1180) );
  OAI21X1 U1852 ( .A(n3158), .B(n3393), .C(n3415), .Y(n2018) );
  OAI21X1 U1853 ( .A(n2035), .B(n3658), .C(n3028), .Y(n1179) );
  OAI21X1 U1855 ( .A(n2035), .B(n3659), .C(n3006), .Y(n1178) );
  OAI21X1 U1857 ( .A(n2035), .B(n3660), .C(n3126), .Y(n1177) );
  OAI21X1 U1859 ( .A(n2035), .B(n3661), .C(n3168), .Y(n1176) );
  OAI21X1 U1861 ( .A(n2035), .B(n3662), .C(n3049), .Y(n1175) );
  OAI21X1 U1863 ( .A(n2035), .B(n3663), .C(n3086), .Y(n1174) );
  OAI21X1 U1865 ( .A(n2035), .B(n3664), .C(n2964), .Y(n1173) );
  OAI21X1 U1867 ( .A(n2035), .B(n3665), .C(n2985), .Y(n1172) );
  OAI21X1 U1869 ( .A(n2035), .B(n3666), .C(n3127), .Y(n1171) );
  OAI21X1 U1871 ( .A(n2035), .B(n3667), .C(n3169), .Y(n1170) );
  OAI21X1 U1873 ( .A(n2035), .B(n3668), .C(n3050), .Y(n1169) );
  OAI21X1 U1875 ( .A(n2035), .B(n3669), .C(n3087), .Y(n1168) );
  OAI21X1 U1877 ( .A(n2035), .B(n3670), .C(n3319), .Y(n1167) );
  OAI21X1 U1879 ( .A(n2035), .B(n3671), .C(n3366), .Y(n1166) );
  OAI21X1 U1881 ( .A(n2035), .B(n3672), .C(n3223), .Y(n1165) );
  OAI21X1 U1883 ( .A(n2035), .B(n3673), .C(n3270), .Y(n1164) );
  OAI21X1 U1885 ( .A(n3203), .B(n3393), .C(n3415), .Y(n2035) );
  OAI21X1 U1886 ( .A(n2052), .B(n3674), .C(n2986), .Y(n1163) );
  OAI21X1 U1888 ( .A(n2052), .B(n3675), .C(n2965), .Y(n1162) );
  OAI21X1 U1890 ( .A(n2052), .B(n3676), .C(n3088), .Y(n1161) );
  OAI21X1 U1892 ( .A(n2052), .B(n3677), .C(n3051), .Y(n1160) );
  OAI21X1 U1894 ( .A(n2052), .B(n3678), .C(n3170), .Y(n1159) );
  OAI21X1 U1896 ( .A(n2052), .B(n3679), .C(n3128), .Y(n1158) );
  OAI21X1 U1898 ( .A(n2052), .B(n3680), .C(n3029), .Y(n1157) );
  OAI21X1 U1900 ( .A(n2052), .B(n3681), .C(n3007), .Y(n1156) );
  OAI21X1 U1902 ( .A(n2052), .B(n3682), .C(n3089), .Y(n1155) );
  OAI21X1 U1904 ( .A(n2052), .B(n3683), .C(n3052), .Y(n1154) );
  OAI21X1 U1906 ( .A(n2052), .B(n3684), .C(n3171), .Y(n1153) );
  OAI21X1 U1908 ( .A(n2052), .B(n3685), .C(n3129), .Y(n1152) );
  OAI21X1 U1910 ( .A(n2052), .B(n3686), .C(n3271), .Y(n1151) );
  OAI21X1 U1912 ( .A(n2052), .B(n3687), .C(n3224), .Y(n1150) );
  OAI21X1 U1914 ( .A(n2052), .B(n3688), .C(n3367), .Y(n1149) );
  OAI21X1 U1916 ( .A(n2052), .B(n3689), .C(n3320), .Y(n1148) );
  OAI21X1 U1918 ( .A(n3249), .B(n3393), .C(n3416), .Y(n2052) );
  NAND3X1 U1919 ( .A(wr_ptr[4]), .B(n3433), .C(put), .Y(n1949) );
  OAI21X1 U1920 ( .A(n2069), .B(n3690), .C(n2966), .Y(n1147) );
  OAI21X1 U1922 ( .A(n2069), .B(n3691), .C(n2987), .Y(n1146) );
  OAI21X1 U1924 ( .A(n2069), .B(n3692), .C(n3053), .Y(n1145) );
  OAI21X1 U1926 ( .A(n2069), .B(n3693), .C(n3090), .Y(n1144) );
  OAI21X1 U1928 ( .A(n2069), .B(n3694), .C(n3130), .Y(n1143) );
  OAI21X1 U1930 ( .A(n2069), .B(n3695), .C(n3172), .Y(n1142) );
  OAI21X1 U1932 ( .A(n2069), .B(n3696), .C(n3008), .Y(n1141) );
  OAI21X1 U1934 ( .A(n2069), .B(n3697), .C(n3030), .Y(n1140) );
  OAI21X1 U1936 ( .A(n2069), .B(n3698), .C(n3054), .Y(n1139) );
  OAI21X1 U1938 ( .A(n2069), .B(n3699), .C(n3091), .Y(n1138) );
  OAI21X1 U1940 ( .A(n2069), .B(n3700), .C(n3131), .Y(n1137) );
  OAI21X1 U1942 ( .A(n2069), .B(n3701), .C(n3173), .Y(n1136) );
  OAI21X1 U1944 ( .A(n2069), .B(n3702), .C(n3225), .Y(n1135) );
  OAI21X1 U1946 ( .A(n2069), .B(n3703), .C(n3272), .Y(n1134) );
  OAI21X1 U1948 ( .A(n2069), .B(n3704), .C(n3321), .Y(n1133) );
  OAI21X1 U1950 ( .A(n2069), .B(n3705), .C(n3368), .Y(n1132) );
  OAI21X1 U1952 ( .A(n3250), .B(n3394), .C(n3416), .Y(n2069) );
  OAI21X1 U1953 ( .A(n2087), .B(n3706), .C(n3009), .Y(n1131) );
  OAI21X1 U1955 ( .A(n2087), .B(n3707), .C(n3031), .Y(n1130) );
  OAI21X1 U1957 ( .A(n2087), .B(n3708), .C(n3322), .Y(n1129) );
  OAI21X1 U1959 ( .A(n2087), .B(n3709), .C(n3369), .Y(n1128) );
  OAI21X1 U1961 ( .A(n2087), .B(n3710), .C(n3273), .Y(n1127) );
  OAI21X1 U1963 ( .A(n2087), .B(n3711), .C(n3226), .Y(n1126) );
  OAI21X1 U1965 ( .A(n2087), .B(n3712), .C(n2897), .Y(n1125) );
  OAI21X1 U1967 ( .A(n2087), .B(n3713), .C(n2871), .Y(n1124) );
  OAI21X1 U1969 ( .A(n2087), .B(n3714), .C(n3370), .Y(n1123) );
  OAI21X1 U1971 ( .A(n2087), .B(n3715), .C(n3323), .Y(n1122) );
  OAI21X1 U1973 ( .A(n2087), .B(n3716), .C(n3274), .Y(n1121) );
  OAI21X1 U1975 ( .A(n2087), .B(n3717), .C(n3227), .Y(n1120) );
  OAI21X1 U1977 ( .A(n2087), .B(n3718), .C(n3174), .Y(n1119) );
  OAI21X1 U1979 ( .A(n2087), .B(n3719), .C(n3132), .Y(n1118) );
  OAI21X1 U1981 ( .A(n2087), .B(n3720), .C(n3092), .Y(n1117) );
  OAI21X1 U1983 ( .A(n2087), .B(n3721), .C(n3055), .Y(n1116) );
  OAI21X1 U1985 ( .A(n3202), .B(n3394), .C(n3416), .Y(n2087) );
  OAI21X1 U1986 ( .A(n2104), .B(n3722), .C(n2949), .Y(n1115) );
  OAI21X1 U1988 ( .A(n2104), .B(n3723), .C(n2923), .Y(n1114) );
  OAI21X1 U1990 ( .A(n2104), .B(n3724), .C(n3324), .Y(n1113) );
  OAI21X1 U1992 ( .A(n2104), .B(n3725), .C(n3371), .Y(n1112) );
  OAI21X1 U1994 ( .A(n2104), .B(n3726), .C(n3228), .Y(n1111) );
  OAI21X1 U1996 ( .A(n2104), .B(n3727), .C(n3275), .Y(n1110) );
  OAI21X1 U1998 ( .A(n2104), .B(n3728), .C(n2872), .Y(n1109) );
  OAI21X1 U2000 ( .A(n2104), .B(n3729), .C(n2898), .Y(n1108) );
  OAI21X1 U2002 ( .A(n2104), .B(n3730), .C(n3325), .Y(n1107) );
  OAI21X1 U2004 ( .A(n2104), .B(n3731), .C(n3372), .Y(n1106) );
  OAI21X1 U2006 ( .A(n2104), .B(n3732), .C(n3229), .Y(n1105) );
  OAI21X1 U2008 ( .A(n2104), .B(n3733), .C(n3276), .Y(n1104) );
  OAI21X1 U2010 ( .A(n2104), .B(n3734), .C(n3133), .Y(n1103) );
  OAI21X1 U2012 ( .A(n2104), .B(n3735), .C(n3175), .Y(n1102) );
  OAI21X1 U2014 ( .A(n2104), .B(n3736), .C(n3056), .Y(n1101) );
  OAI21X1 U2016 ( .A(n2104), .B(n3737), .C(n3093), .Y(n1100) );
  OAI21X1 U2018 ( .A(n3157), .B(n3394), .C(n3416), .Y(n2104) );
  NAND3X1 U2019 ( .A(wr_ptr[0]), .B(n3431), .C(wr_ptr[2]), .Y(n1674) );
  OAI21X1 U2020 ( .A(n2121), .B(n3738), .C(n2899), .Y(n1099) );
  OAI21X1 U2022 ( .A(n2121), .B(n3739), .C(n2873), .Y(n1098) );
  OAI21X1 U2024 ( .A(n2121), .B(n3740), .C(n3277), .Y(n1097) );
  OAI21X1 U2026 ( .A(n2121), .B(n3741), .C(n3230), .Y(n1096) );
  OAI21X1 U2028 ( .A(n2121), .B(n3742), .C(n3373), .Y(n1095) );
  OAI21X1 U2030 ( .A(n2121), .B(n3743), .C(n3326), .Y(n1094) );
  OAI21X1 U2032 ( .A(n2121), .B(n3744), .C(n2950), .Y(n1093) );
  OAI21X1 U2034 ( .A(n2121), .B(n3745), .C(n2924), .Y(n1092) );
  OAI21X1 U2036 ( .A(n2121), .B(n3746), .C(n3278), .Y(n1091) );
  OAI21X1 U2038 ( .A(n2121), .B(n3747), .C(n3231), .Y(n1090) );
  OAI21X1 U2040 ( .A(n2121), .B(n3748), .C(n3374), .Y(n1089) );
  OAI21X1 U2042 ( .A(n2121), .B(n3749), .C(n3327), .Y(n1088) );
  OAI21X1 U2044 ( .A(n2121), .B(n3750), .C(n3094), .Y(n1087) );
  OAI21X1 U2046 ( .A(n2121), .B(n3751), .C(n3057), .Y(n1086) );
  OAI21X1 U2048 ( .A(n2121), .B(n3752), .C(n3176), .Y(n1085) );
  OAI21X1 U2050 ( .A(n2121), .B(n3753), .C(n3134), .Y(n1084) );
  OAI21X1 U2052 ( .A(n3299), .B(n3394), .C(n3416), .Y(n2121) );
  NAND3X1 U2053 ( .A(n3422), .B(n3431), .C(wr_ptr[2]), .Y(n1692) );
  OAI21X1 U2054 ( .A(n2138), .B(n3754), .C(n2874), .Y(n1083) );
  OAI21X1 U2056 ( .A(n2138), .B(n3755), .C(n2900), .Y(n1082) );
  OAI21X1 U2058 ( .A(n2138), .B(n3756), .C(n3232), .Y(n1081) );
  OAI21X1 U2060 ( .A(n2138), .B(n3757), .C(n3279), .Y(n1080) );
  OAI21X1 U2062 ( .A(n2138), .B(n3758), .C(n3328), .Y(n1079) );
  OAI21X1 U2064 ( .A(n2138), .B(n3759), .C(n3375), .Y(n1078) );
  OAI21X1 U2066 ( .A(n2138), .B(n3760), .C(n2925), .Y(n1077) );
  OAI21X1 U2068 ( .A(n2138), .B(n3761), .C(n2951), .Y(n1076) );
  OAI21X1 U2070 ( .A(n2138), .B(n3762), .C(n3233), .Y(n1075) );
  OAI21X1 U2072 ( .A(n2138), .B(n3763), .C(n3280), .Y(n1074) );
  OAI21X1 U2074 ( .A(n2138), .B(n3764), .C(n3329), .Y(n1073) );
  OAI21X1 U2076 ( .A(n2138), .B(n3765), .C(n3376), .Y(n1072) );
  OAI21X1 U2078 ( .A(n2138), .B(n3766), .C(n3058), .Y(n1071) );
  OAI21X1 U2080 ( .A(n2138), .B(n3767), .C(n3095), .Y(n1070) );
  OAI21X1 U2082 ( .A(n2138), .B(n3768), .C(n3135), .Y(n1069) );
  OAI21X1 U2084 ( .A(n2138), .B(n3769), .C(n3177), .Y(n1068) );
  OAI21X1 U2086 ( .A(n3300), .B(n3394), .C(n3416), .Y(n2138) );
  NAND3X1 U2087 ( .A(wr_ptr[0]), .B(n3432), .C(wr_ptr[1]), .Y(n1710) );
  OAI21X1 U2088 ( .A(n2155), .B(n3770), .C(n3032), .Y(n1067) );
  OAI21X1 U2090 ( .A(n2155), .B(n3771), .C(n3010), .Y(n1066) );
  OAI21X1 U2092 ( .A(n2155), .B(n3772), .C(n3178), .Y(n1065) );
  OAI21X1 U2094 ( .A(n2155), .B(n3773), .C(n3136), .Y(n1064) );
  OAI21X1 U2096 ( .A(n2155), .B(n3774), .C(n3096), .Y(n1063) );
  OAI21X1 U2098 ( .A(n2155), .B(n3775), .C(n3059), .Y(n1062) );
  OAI21X1 U2100 ( .A(n2155), .B(n3776), .C(n2988), .Y(n1061) );
  OAI21X1 U2102 ( .A(n2155), .B(n3777), .C(n2967), .Y(n1060) );
  OAI21X1 U2104 ( .A(n2155), .B(n3778), .C(n3179), .Y(n1059) );
  OAI21X1 U2106 ( .A(n2155), .B(n3779), .C(n3137), .Y(n1058) );
  OAI21X1 U2108 ( .A(n2155), .B(n3780), .C(n3097), .Y(n1057) );
  OAI21X1 U2110 ( .A(n2155), .B(n3781), .C(n3060), .Y(n1056) );
  OAI21X1 U2112 ( .A(n2155), .B(n3782), .C(n3377), .Y(n1055) );
  OAI21X1 U2114 ( .A(n2155), .B(n3783), .C(n3330), .Y(n1054) );
  OAI21X1 U2116 ( .A(n2155), .B(n3784), .C(n3281), .Y(n1053) );
  OAI21X1 U2118 ( .A(n2155), .B(n3785), .C(n3234), .Y(n1052) );
  OAI21X1 U2120 ( .A(n3158), .B(n3394), .C(n3416), .Y(n2155) );
  NAND3X1 U2121 ( .A(n3422), .B(n3432), .C(wr_ptr[1]), .Y(n1728) );
  OAI21X1 U2122 ( .A(n2172), .B(n3786), .C(n3011), .Y(n1051) );
  OAI21X1 U2124 ( .A(n2172), .B(n3787), .C(n3033), .Y(n1050) );
  OAI21X1 U2126 ( .A(n2172), .B(n3788), .C(n3138), .Y(n1049) );
  OAI21X1 U2128 ( .A(n2172), .B(n3789), .C(n3180), .Y(n1048) );
  OAI21X1 U2130 ( .A(n2172), .B(n3790), .C(n3061), .Y(n1047) );
  OAI21X1 U2132 ( .A(n2172), .B(n3791), .C(n3098), .Y(n1046) );
  OAI21X1 U2134 ( .A(n2172), .B(n3792), .C(n2968), .Y(n1045) );
  OAI21X1 U2136 ( .A(n2172), .B(n3793), .C(n2989), .Y(n1044) );
  OAI21X1 U2138 ( .A(n2172), .B(n3794), .C(n3139), .Y(n1043) );
  OAI21X1 U2140 ( .A(n2172), .B(n3795), .C(n3181), .Y(n1042) );
  OAI21X1 U2142 ( .A(n2172), .B(n3796), .C(n3062), .Y(n1041) );
  OAI21X1 U2144 ( .A(n2172), .B(n3797), .C(n3099), .Y(n1040) );
  OAI21X1 U2146 ( .A(n2172), .B(n3798), .C(n3331), .Y(n1039) );
  OAI21X1 U2148 ( .A(n2172), .B(n3799), .C(n3378), .Y(n1038) );
  OAI21X1 U2150 ( .A(n2172), .B(n3800), .C(n3235), .Y(n1037) );
  OAI21X1 U2152 ( .A(n2172), .B(n3801), .C(n3282), .Y(n1036) );
  OAI21X1 U2154 ( .A(n3203), .B(n3394), .C(n3416), .Y(n2172) );
  NAND3X1 U2155 ( .A(n3431), .B(n3432), .C(wr_ptr[0]), .Y(n1746) );
  OAI21X1 U2156 ( .A(n2189), .B(n3802), .C(n2990), .Y(n1035) );
  OAI21X1 U2158 ( .A(n2189), .B(n3803), .C(n2969), .Y(n1034) );
  OAI21X1 U2160 ( .A(n2189), .B(n3804), .C(n3100), .Y(n1033) );
  OAI21X1 U2162 ( .A(n2189), .B(n3805), .C(n3063), .Y(n1032) );
  OAI21X1 U2164 ( .A(n2189), .B(n3806), .C(n3182), .Y(n1031) );
  OAI21X1 U2166 ( .A(n2189), .B(n3807), .C(n3140), .Y(n1030) );
  OAI21X1 U2168 ( .A(n2189), .B(n3808), .C(n3034), .Y(n1029) );
  OAI21X1 U2170 ( .A(n2189), .B(n3809), .C(n3012), .Y(n1028) );
  OAI21X1 U2172 ( .A(n2189), .B(n3810), .C(n3101), .Y(n1027) );
  OAI21X1 U2174 ( .A(n2189), .B(n3811), .C(n3064), .Y(n1026) );
  OAI21X1 U2176 ( .A(n2189), .B(n3812), .C(n3183), .Y(n1025) );
  OAI21X1 U2178 ( .A(n2189), .B(n3813), .C(n3141), .Y(n1024) );
  OAI21X1 U2180 ( .A(n2189), .B(n3814), .C(n3283), .Y(n1023) );
  OAI21X1 U2182 ( .A(n2189), .B(n3815), .C(n3236), .Y(n1022) );
  OAI21X1 U2184 ( .A(n2189), .B(n3816), .C(n3379), .Y(n1021) );
  OAI21X1 U2186 ( .A(n2189), .B(n3817), .C(n3332), .Y(n1020) );
  OAI21X1 U2188 ( .A(n3249), .B(n3394), .C(n3416), .Y(n2189) );
  NAND3X1 U2189 ( .A(wr_ptr[3]), .B(n3430), .C(put), .Y(n2086) );
  NAND3X1 U2190 ( .A(n3431), .B(n3432), .C(n3422), .Y(n1764) );
  OAI21X1 U2191 ( .A(n2206), .B(n3818), .C(n2970), .Y(n1019) );
  OAI21X1 U2193 ( .A(n2206), .B(n3819), .C(n2991), .Y(n1018) );
  OAI21X1 U2195 ( .A(n2206), .B(n3820), .C(n3065), .Y(n1017) );
  OAI21X1 U2197 ( .A(n2206), .B(n3821), .C(n3102), .Y(n1016) );
  OAI21X1 U2199 ( .A(n2206), .B(n3822), .C(n3142), .Y(n1015) );
  OAI21X1 U2201 ( .A(n2206), .B(n3823), .C(n3184), .Y(n1014) );
  OAI21X1 U2203 ( .A(n2206), .B(n3824), .C(n3013), .Y(n1013) );
  OAI21X1 U2205 ( .A(n2206), .B(n3825), .C(n3035), .Y(n1012) );
  OAI21X1 U2207 ( .A(n2206), .B(n3826), .C(n3066), .Y(n1011) );
  OAI21X1 U2209 ( .A(n2206), .B(n3827), .C(n3103), .Y(n1010) );
  OAI21X1 U2211 ( .A(n2206), .B(n3828), .C(n3143), .Y(n1009) );
  OAI21X1 U2213 ( .A(n2206), .B(n3829), .C(n3185), .Y(n1008) );
  OAI21X1 U2215 ( .A(n2206), .B(n3830), .C(n3237), .Y(n1007) );
  OAI21X1 U2217 ( .A(n2206), .B(n3831), .C(n3284), .Y(n1006) );
  OAI21X1 U2219 ( .A(n2206), .B(n3832), .C(n3333), .Y(n1005) );
  OAI21X1 U2221 ( .A(n2206), .B(n3833), .C(n3380), .Y(n1004) );
  OAI21X1 U2223 ( .A(n3345), .B(n3250), .C(n3416), .Y(n2206) );
  NAND3X1 U2224 ( .A(wr_ptr[2]), .B(wr_ptr[0]), .C(wr_ptr[1]), .Y(n1793) );
  OAI21X1 U2225 ( .A(n1627), .B(n3834), .C(n2926), .Y(n1003) );
  OAI21X1 U2227 ( .A(n1627), .B(n3835), .C(n2952), .Y(n1002) );
  OAI21X1 U2229 ( .A(n1627), .B(n3836), .C(n2971), .Y(n1001) );
  OAI21X1 U2231 ( .A(n1627), .B(n3837), .C(n2992), .Y(n1000) );
  OAI21X1 U2233 ( .A(n3202), .B(n3345), .C(n3415), .Y(n1627) );
  NAND3X1 U2234 ( .A(n3433), .B(n3430), .C(put), .Y(n1673) );
  NAND3X1 U2235 ( .A(wr_ptr[2]), .B(n3422), .C(wr_ptr[1]), .Y(n1829) );
  XOR2X1 U2236 ( .A(n3296), .B(n1783), .Y(fillcount[4]) );
  XNOR2X1 U2237 ( .A(n16), .B(n3430), .Y(n1783) );
  AOI21X1 U2238 ( .A(n3429), .B(n2227), .C(n3297), .Y(n1625) );
  AOI21X1 U2239 ( .A(n15), .B(n3420), .C(n3433), .Y(n2228) );
  XOR2X1 U2240 ( .A(n2227), .B(n1780), .Y(fillcount[3]) );
  XNOR2X1 U2241 ( .A(n15), .B(wr_ptr[3]), .Y(n1780) );
  OAI21X1 U2242 ( .A(n14), .B(n3115), .C(n2230), .Y(n2227) );
  OAI21X1 U2243 ( .A(n3428), .B(n3421), .C(wr_ptr[2]), .Y(n2230) );
  XOR2X1 U2244 ( .A(n3421), .B(n1779), .Y(fillcount[2]) );
  XNOR2X1 U2245 ( .A(n14), .B(wr_ptr[2]), .Y(n1779) );
  AOI21X1 U2246 ( .A(n3427), .B(n3391), .C(n3116), .Y(n2229) );
  AOI21X1 U2247 ( .A(n13), .B(n2231), .C(n3431), .Y(n2232) );
  XNOR2X1 U2248 ( .A(n3391), .B(n1782), .Y(fillcount[1]) );
  XNOR2X1 U2249 ( .A(n13), .B(n3431), .Y(n1782) );
  OAI21X1 U2250 ( .A(n3399), .B(n3422), .C(n3391), .Y(fillcount[0]) );
  OR2X1 U3 ( .A(n2337), .B(n2401), .Y(n1587) );
  OR2X1 U4 ( .A(n2338), .B(n2402), .Y(n1588) );
  OR2X1 U5 ( .A(n2339), .B(n2403), .Y(n1589) );
  OR2X1 U6 ( .A(n2341), .B(n2405), .Y(n1553) );
  OR2X1 U7 ( .A(n2342), .B(n2406), .Y(n1554) );
  OR2X1 U8 ( .A(n2343), .B(n2407), .Y(n1555) );
  OR2X1 U9 ( .A(n2345), .B(n2409), .Y(n1519) );
  OR2X1 U10 ( .A(n2346), .B(n2410), .Y(n1520) );
  OR2X1 U11 ( .A(n2347), .B(n2411), .Y(n1521) );
  OR2X1 U12 ( .A(n2349), .B(n2413), .Y(n1485) );
  OR2X1 U13 ( .A(n2350), .B(n2414), .Y(n1486) );
  OR2X1 U14 ( .A(n2351), .B(n2415), .Y(n1487) );
  OR2X1 U15 ( .A(n2353), .B(n2417), .Y(n1451) );
  OR2X1 U16 ( .A(n2354), .B(n2418), .Y(n1452) );
  OR2X1 U17 ( .A(n2355), .B(n2419), .Y(n1453) );
  OR2X1 U18 ( .A(n2357), .B(n2421), .Y(n1417) );
  OR2X1 U19 ( .A(n2359), .B(n2423), .Y(n1419) );
  OR2X1 U20 ( .A(n2358), .B(n2422), .Y(n1418) );
  OR2X1 U21 ( .A(n2361), .B(n2425), .Y(n861) );
  OR2X1 U22 ( .A(n2363), .B(n2427), .Y(n863) );
  OR2X1 U23 ( .A(n2362), .B(n2426), .Y(n862) );
  OR2X1 U24 ( .A(n2365), .B(n2429), .Y(n827) );
  OR2X1 U25 ( .A(n2366), .B(n2430), .Y(n828) );
  OR2X1 U26 ( .A(n2367), .B(n2431), .Y(n829) );
  OR2X1 U27 ( .A(n2369), .B(n2433), .Y(n793) );
  OR2X1 U28 ( .A(n2370), .B(n2434), .Y(n794) );
  OR2X1 U29 ( .A(n2371), .B(n2435), .Y(n795) );
  OR2X1 U30 ( .A(n2373), .B(n2437), .Y(n759) );
  OR2X1 U31 ( .A(n2374), .B(n2438), .Y(n760) );
  OR2X1 U32 ( .A(n2375), .B(n2439), .Y(n761) );
  OR2X1 U33 ( .A(n2377), .B(n2441), .Y(n725) );
  OR2X1 U34 ( .A(n2378), .B(n2442), .Y(n726) );
  OR2X1 U35 ( .A(n2379), .B(n2443), .Y(n727) );
  OR2X1 U36 ( .A(n2381), .B(n2445), .Y(n691) );
  OR2X1 U37 ( .A(n2382), .B(n2446), .Y(n692) );
  OR2X1 U38 ( .A(n2383), .B(n2447), .Y(n693) );
  OR2X1 U39 ( .A(n2385), .B(n2449), .Y(n657) );
  OR2X1 U40 ( .A(n2386), .B(n2450), .Y(n658) );
  OR2X1 U41 ( .A(n2387), .B(n2451), .Y(n659) );
  OR2X1 U42 ( .A(n2389), .B(n2453), .Y(n623) );
  OR2X1 U43 ( .A(n2390), .B(n2454), .Y(n624) );
  OR2X1 U44 ( .A(n2391), .B(n2455), .Y(n625) );
  OR2X1 U45 ( .A(n2394), .B(n2458), .Y(n590) );
  OR2X1 U46 ( .A(n2395), .B(n2459), .Y(n591) );
  OR2X1 U47 ( .A(n2393), .B(n2457), .Y(n589) );
  OR2X1 U48 ( .A(n2397), .B(n2461), .Y(n545) );
  OR2X1 U49 ( .A(n2398), .B(n2462), .Y(n546) );
  OR2X1 U50 ( .A(n2399), .B(n2463), .Y(n547) );
  OR2X1 U51 ( .A(n2336), .B(n2400), .Y(n1585) );
  OR2X1 U52 ( .A(n2340), .B(n2404), .Y(n1551) );
  OR2X1 U53 ( .A(n2344), .B(n2408), .Y(n1517) );
  OR2X1 U54 ( .A(n2348), .B(n2412), .Y(n1483) );
  OR2X1 U55 ( .A(n2352), .B(n2416), .Y(n1449) );
  OR2X1 U56 ( .A(n2356), .B(n2420), .Y(n1415) );
  OR2X1 U57 ( .A(n2360), .B(n2424), .Y(n859) );
  OR2X1 U58 ( .A(n2364), .B(n2428), .Y(n825) );
  OR2X1 U59 ( .A(n2368), .B(n2432), .Y(n791) );
  OR2X1 U60 ( .A(n2372), .B(n2436), .Y(n757) );
  OR2X1 U61 ( .A(n2376), .B(n2440), .Y(n723) );
  OR2X1 U62 ( .A(n2380), .B(n2444), .Y(n689) );
  OR2X1 U63 ( .A(n2384), .B(n2448), .Y(n655) );
  OR2X1 U64 ( .A(n2388), .B(n2452), .Y(n621) );
  OR2X1 U65 ( .A(n2392), .B(n2456), .Y(n587) );
  OR2X1 U66 ( .A(n2396), .B(n2460), .Y(n543) );
  OR2X1 U67 ( .A(n3392), .B(n3300), .Y(n1791) );
  OR2X1 U68 ( .A(n3298), .B(n3422), .Y(n1766) );
  AND2X1 U69 ( .A(n3416), .B(n3247), .Y(n1610) );
  AND2X1 U70 ( .A(reset), .B(n3248), .Y(n1777) );
  AND2X1 U71 ( .A(n3415), .B(n3298), .Y(n1765) );
  BUFX2 U72 ( .A(n1412), .Y(n2316) );
  BUFX2 U73 ( .A(n2248), .Y(n2317) );
  BUFX2 U74 ( .A(n2247), .Y(n2318) );
  BUFX2 U75 ( .A(n2246), .Y(n2319) );
  BUFX2 U76 ( .A(n2245), .Y(n2320) );
  BUFX2 U77 ( .A(n2244), .Y(n2321) );
  BUFX2 U78 ( .A(n2243), .Y(n2322) );
  BUFX2 U79 ( .A(n2242), .Y(n2323) );
  BUFX2 U80 ( .A(n2241), .Y(n2324) );
  BUFX2 U81 ( .A(n2240), .Y(n2325) );
  BUFX2 U82 ( .A(n2239), .Y(n2326) );
  BUFX2 U83 ( .A(n2238), .Y(n2327) );
  BUFX2 U84 ( .A(n2237), .Y(n2328) );
  BUFX2 U85 ( .A(n2236), .Y(n2329) );
  BUFX2 U86 ( .A(n2235), .Y(n2330) );
  BUFX2 U87 ( .A(n2234), .Y(n2331) );
  BUFX2 U88 ( .A(n2233), .Y(n2332) );
  BUFX2 U89 ( .A(n1776), .Y(n2333) );
  BUFX2 U90 ( .A(n1773), .Y(n2334) );
  AND2X1 U91 ( .A(n1654), .B(n1950), .Y(n1951) );
  INVX1 U92 ( .A(n1951), .Y(n2335) );
  BUFX2 U93 ( .A(n1614), .Y(n2336) );
  BUFX2 U94 ( .A(n1606), .Y(n2337) );
  BUFX2 U95 ( .A(n1598), .Y(n2338) );
  BUFX2 U96 ( .A(n1590), .Y(n2339) );
  BUFX2 U97 ( .A(n1577), .Y(n2340) );
  BUFX2 U98 ( .A(n1570), .Y(n2341) );
  BUFX2 U99 ( .A(n1563), .Y(n2342) );
  BUFX2 U100 ( .A(n1556), .Y(n2343) );
  BUFX2 U101 ( .A(n1543), .Y(n2344) );
  BUFX2 U102 ( .A(n1536), .Y(n2345) );
  BUFX2 U103 ( .A(n1529), .Y(n2346) );
  BUFX2 U104 ( .A(n1522), .Y(n2347) );
  BUFX2 U105 ( .A(n1509), .Y(n2348) );
  BUFX2 U106 ( .A(n1502), .Y(n2349) );
  BUFX2 U107 ( .A(n1495), .Y(n2350) );
  BUFX2 U108 ( .A(n1488), .Y(n2351) );
  BUFX2 U109 ( .A(n1475), .Y(n2352) );
  BUFX2 U110 ( .A(n1468), .Y(n2353) );
  BUFX2 U111 ( .A(n1461), .Y(n2354) );
  BUFX2 U112 ( .A(n1454), .Y(n2355) );
  BUFX2 U113 ( .A(n1441), .Y(n2356) );
  BUFX2 U114 ( .A(n1434), .Y(n2357) );
  BUFX2 U115 ( .A(n1427), .Y(n2358) );
  BUFX2 U116 ( .A(n1420), .Y(n2359) );
  BUFX2 U117 ( .A(n885), .Y(n2360) );
  BUFX2 U118 ( .A(n878), .Y(n2361) );
  BUFX2 U119 ( .A(n871), .Y(n2362) );
  BUFX2 U120 ( .A(n864), .Y(n2363) );
  BUFX2 U121 ( .A(n851), .Y(n2364) );
  BUFX2 U122 ( .A(n844), .Y(n2365) );
  BUFX2 U123 ( .A(n837), .Y(n2366) );
  BUFX2 U124 ( .A(n830), .Y(n2367) );
  BUFX2 U125 ( .A(n817), .Y(n2368) );
  BUFX2 U126 ( .A(n810), .Y(n2369) );
  BUFX2 U127 ( .A(n803), .Y(n2370) );
  BUFX2 U128 ( .A(n796), .Y(n2371) );
  BUFX2 U129 ( .A(n783), .Y(n2372) );
  BUFX2 U130 ( .A(n776), .Y(n2373) );
  BUFX2 U131 ( .A(n769), .Y(n2374) );
  BUFX2 U132 ( .A(n762), .Y(n2375) );
  BUFX2 U133 ( .A(n749), .Y(n2376) );
  BUFX2 U134 ( .A(n742), .Y(n2377) );
  BUFX2 U135 ( .A(n735), .Y(n2378) );
  BUFX2 U136 ( .A(n728), .Y(n2379) );
  BUFX2 U137 ( .A(n715), .Y(n2380) );
  BUFX2 U138 ( .A(n708), .Y(n2381) );
  BUFX2 U139 ( .A(n701), .Y(n2382) );
  BUFX2 U140 ( .A(n694), .Y(n2383) );
  BUFX2 U141 ( .A(n681), .Y(n2384) );
  BUFX2 U142 ( .A(n674), .Y(n2385) );
  BUFX2 U143 ( .A(n667), .Y(n2386) );
  BUFX2 U144 ( .A(n660), .Y(n2387) );
  BUFX2 U145 ( .A(n647), .Y(n2388) );
  BUFX2 U146 ( .A(n640), .Y(n2389) );
  BUFX2 U147 ( .A(n633), .Y(n2390) );
  BUFX2 U148 ( .A(n626), .Y(n2391) );
  BUFX2 U149 ( .A(n613), .Y(n2392) );
  BUFX2 U150 ( .A(n606), .Y(n2393) );
  BUFX2 U151 ( .A(n599), .Y(n2394) );
  BUFX2 U152 ( .A(n592), .Y(n2395) );
  BUFX2 U153 ( .A(n578), .Y(n2396) );
  BUFX2 U154 ( .A(n570), .Y(n2397) );
  BUFX2 U155 ( .A(n562), .Y(n2398) );
  BUFX2 U156 ( .A(n548), .Y(n2399) );
  BUFX2 U157 ( .A(n1615), .Y(n2400) );
  BUFX2 U158 ( .A(n1607), .Y(n2401) );
  BUFX2 U159 ( .A(n1599), .Y(n2402) );
  BUFX2 U160 ( .A(n1591), .Y(n2403) );
  BUFX2 U161 ( .A(n1578), .Y(n2404) );
  BUFX2 U162 ( .A(n1571), .Y(n2405) );
  BUFX2 U163 ( .A(n1564), .Y(n2406) );
  BUFX2 U164 ( .A(n1557), .Y(n2407) );
  BUFX2 U165 ( .A(n1544), .Y(n2408) );
  BUFX2 U166 ( .A(n1537), .Y(n2409) );
  BUFX2 U167 ( .A(n1530), .Y(n2410) );
  BUFX2 U168 ( .A(n1523), .Y(n2411) );
  BUFX2 U169 ( .A(n1510), .Y(n2412) );
  BUFX2 U170 ( .A(n1503), .Y(n2413) );
  BUFX2 U171 ( .A(n1496), .Y(n2414) );
  BUFX2 U172 ( .A(n1489), .Y(n2415) );
  BUFX2 U173 ( .A(n1476), .Y(n2416) );
  BUFX2 U174 ( .A(n1469), .Y(n2417) );
  BUFX2 U175 ( .A(n1462), .Y(n2418) );
  BUFX2 U176 ( .A(n1455), .Y(n2419) );
  BUFX2 U177 ( .A(n1442), .Y(n2420) );
  BUFX2 U178 ( .A(n1435), .Y(n2421) );
  BUFX2 U179 ( .A(n1428), .Y(n2422) );
  BUFX2 U180 ( .A(n1421), .Y(n2423) );
  BUFX2 U181 ( .A(n886), .Y(n2424) );
  BUFX2 U182 ( .A(n879), .Y(n2425) );
  BUFX2 U183 ( .A(n872), .Y(n2426) );
  BUFX2 U184 ( .A(n865), .Y(n2427) );
  BUFX2 U185 ( .A(n852), .Y(n2428) );
  BUFX2 U186 ( .A(n845), .Y(n2429) );
  BUFX2 U187 ( .A(n838), .Y(n2430) );
  BUFX2 U188 ( .A(n831), .Y(n2431) );
  BUFX2 U189 ( .A(n818), .Y(n2432) );
  BUFX2 U190 ( .A(n811), .Y(n2433) );
  BUFX2 U191 ( .A(n804), .Y(n2434) );
  BUFX2 U192 ( .A(n797), .Y(n2435) );
  BUFX2 U193 ( .A(n784), .Y(n2436) );
  BUFX2 U194 ( .A(n777), .Y(n2437) );
  BUFX2 U195 ( .A(n770), .Y(n2438) );
  BUFX2 U196 ( .A(n763), .Y(n2439) );
  BUFX2 U197 ( .A(n750), .Y(n2440) );
  BUFX2 U198 ( .A(n743), .Y(n2441) );
  BUFX2 U199 ( .A(n736), .Y(n2442) );
  BUFX2 U200 ( .A(n729), .Y(n2443) );
  BUFX2 U201 ( .A(n716), .Y(n2444) );
  BUFX2 U202 ( .A(n709), .Y(n2445) );
  BUFX2 U203 ( .A(n702), .Y(n2446) );
  BUFX2 U204 ( .A(n695), .Y(n2447) );
  BUFX2 U205 ( .A(n682), .Y(n2448) );
  BUFX2 U206 ( .A(n675), .Y(n2449) );
  BUFX2 U207 ( .A(n668), .Y(n2450) );
  BUFX2 U208 ( .A(n661), .Y(n2451) );
  BUFX2 U209 ( .A(n648), .Y(n2452) );
  BUFX2 U210 ( .A(n641), .Y(n2453) );
  BUFX2 U211 ( .A(n634), .Y(n2454) );
  BUFX2 U212 ( .A(n627), .Y(n2455) );
  BUFX2 U213 ( .A(n614), .Y(n2456) );
  BUFX2 U214 ( .A(n607), .Y(n2457) );
  BUFX2 U215 ( .A(n600), .Y(n2458) );
  BUFX2 U216 ( .A(n593), .Y(n2459) );
  BUFX2 U217 ( .A(n579), .Y(n2460) );
  BUFX2 U218 ( .A(n571), .Y(n2461) );
  BUFX2 U219 ( .A(n563), .Y(n2462) );
  BUFX2 U220 ( .A(n549), .Y(n2463) );
  BUFX2 U221 ( .A(n1618), .Y(n2464) );
  BUFX2 U222 ( .A(n1611), .Y(n2465) );
  BUFX2 U223 ( .A(n1603), .Y(n2466) );
  BUFX2 U224 ( .A(n1595), .Y(n2467) );
  BUFX2 U225 ( .A(n1581), .Y(n2468) );
  BUFX2 U226 ( .A(n1574), .Y(n2469) );
  BUFX2 U227 ( .A(n1567), .Y(n2470) );
  BUFX2 U228 ( .A(n1560), .Y(n2471) );
  BUFX2 U229 ( .A(n1547), .Y(n2472) );
  BUFX2 U230 ( .A(n1540), .Y(n2473) );
  BUFX2 U231 ( .A(n1533), .Y(n2474) );
  BUFX2 U232 ( .A(n1526), .Y(n2475) );
  BUFX2 U233 ( .A(n1513), .Y(n2476) );
  BUFX2 U234 ( .A(n1506), .Y(n2477) );
  BUFX2 U235 ( .A(n1499), .Y(n2478) );
  BUFX2 U236 ( .A(n1492), .Y(n2479) );
  BUFX2 U237 ( .A(n1479), .Y(n2480) );
  BUFX2 U238 ( .A(n1472), .Y(n2481) );
  BUFX2 U239 ( .A(n1465), .Y(n2482) );
  BUFX2 U240 ( .A(n1458), .Y(n2483) );
  BUFX2 U241 ( .A(n1445), .Y(n2484) );
  BUFX2 U242 ( .A(n1438), .Y(n2485) );
  BUFX2 U243 ( .A(n1431), .Y(n2486) );
  BUFX2 U244 ( .A(n1424), .Y(n2487) );
  BUFX2 U245 ( .A(n889), .Y(n2488) );
  BUFX2 U246 ( .A(n882), .Y(n2489) );
  BUFX2 U247 ( .A(n875), .Y(n2490) );
  BUFX2 U248 ( .A(n868), .Y(n2491) );
  BUFX2 U249 ( .A(n855), .Y(n2492) );
  BUFX2 U250 ( .A(n848), .Y(n2493) );
  BUFX2 U251 ( .A(n841), .Y(n2494) );
  BUFX2 U252 ( .A(n834), .Y(n2495) );
  BUFX2 U253 ( .A(n821), .Y(n2496) );
  BUFX2 U254 ( .A(n814), .Y(n2497) );
  BUFX2 U255 ( .A(n807), .Y(n2498) );
  BUFX2 U256 ( .A(n800), .Y(n2499) );
  BUFX2 U257 ( .A(n787), .Y(n2500) );
  BUFX2 U258 ( .A(n780), .Y(n2501) );
  BUFX2 U259 ( .A(n773), .Y(n2502) );
  BUFX2 U260 ( .A(n766), .Y(n2503) );
  BUFX2 U261 ( .A(n753), .Y(n2504) );
  BUFX2 U262 ( .A(n746), .Y(n2505) );
  BUFX2 U263 ( .A(n739), .Y(n2506) );
  BUFX2 U264 ( .A(n732), .Y(n2507) );
  BUFX2 U265 ( .A(n719), .Y(n2508) );
  BUFX2 U266 ( .A(n712), .Y(n2509) );
  BUFX2 U267 ( .A(n705), .Y(n2510) );
  BUFX2 U268 ( .A(n698), .Y(n2511) );
  BUFX2 U269 ( .A(n685), .Y(n2512) );
  BUFX2 U270 ( .A(n678), .Y(n2513) );
  BUFX2 U271 ( .A(n671), .Y(n2514) );
  BUFX2 U272 ( .A(n664), .Y(n2515) );
  BUFX2 U273 ( .A(n651), .Y(n2516) );
  BUFX2 U274 ( .A(n644), .Y(n2517) );
  BUFX2 U275 ( .A(n637), .Y(n2518) );
  BUFX2 U276 ( .A(n630), .Y(n2519) );
  BUFX2 U277 ( .A(n617), .Y(n2520) );
  BUFX2 U278 ( .A(n610), .Y(n2521) );
  BUFX2 U279 ( .A(n603), .Y(n2522) );
  BUFX2 U280 ( .A(n596), .Y(n2523) );
  BUFX2 U281 ( .A(n583), .Y(n2524) );
  BUFX2 U282 ( .A(n575), .Y(n2525) );
  BUFX2 U283 ( .A(n567), .Y(n2526) );
  BUFX2 U284 ( .A(n554), .Y(n2527) );
  AND2X1 U285 ( .A(n3396), .B(n3400), .Y(n1768) );
  INVX1 U286 ( .A(n1768), .Y(n2528) );
  AND2X1 U287 ( .A(data_out[0]), .B(n1777), .Y(n1584) );
  INVX1 U288 ( .A(n1584), .Y(n2529) );
  AND2X1 U289 ( .A(data_out[1]), .B(n1777), .Y(n1550) );
  INVX1 U290 ( .A(n1550), .Y(n2530) );
  AND2X1 U291 ( .A(data_out[2]), .B(n1777), .Y(n1516) );
  INVX1 U292 ( .A(n1516), .Y(n2531) );
  AND2X1 U293 ( .A(data_out[3]), .B(n1777), .Y(n1482) );
  INVX1 U294 ( .A(n1482), .Y(n2532) );
  AND2X1 U295 ( .A(data_out[4]), .B(n1777), .Y(n1448) );
  INVX1 U296 ( .A(n1448), .Y(n2533) );
  AND2X1 U297 ( .A(data_out[5]), .B(n1777), .Y(n1414) );
  INVX1 U298 ( .A(n1414), .Y(n2534) );
  AND2X1 U299 ( .A(data_out[6]), .B(n1777), .Y(n858) );
  INVX1 U300 ( .A(n858), .Y(n2535) );
  AND2X1 U301 ( .A(data_out[7]), .B(n1777), .Y(n824) );
  INVX1 U302 ( .A(n824), .Y(n2536) );
  AND2X1 U303 ( .A(data_out[8]), .B(n1777), .Y(n790) );
  INVX1 U304 ( .A(n790), .Y(n2537) );
  AND2X1 U305 ( .A(data_out[9]), .B(n1777), .Y(n756) );
  INVX1 U306 ( .A(n756), .Y(n2538) );
  AND2X1 U307 ( .A(data_out[10]), .B(n1777), .Y(n722) );
  INVX1 U308 ( .A(n722), .Y(n2539) );
  AND2X1 U309 ( .A(data_out[11]), .B(n1777), .Y(n688) );
  INVX1 U310 ( .A(n688), .Y(n2540) );
  AND2X1 U311 ( .A(data_out[12]), .B(n1777), .Y(n654) );
  INVX1 U312 ( .A(n654), .Y(n2541) );
  AND2X1 U313 ( .A(data_out[13]), .B(n1777), .Y(n620) );
  INVX1 U314 ( .A(n620), .Y(n2542) );
  AND2X1 U315 ( .A(data_out[14]), .B(n1777), .Y(n586) );
  INVX1 U316 ( .A(n586), .Y(n2543) );
  AND2X1 U317 ( .A(data_out[15]), .B(n1777), .Y(n542) );
  INVX1 U318 ( .A(n542), .Y(n2544) );
  BUFX2 U319 ( .A(n1775), .Y(n2545) );
  AND2X1 U320 ( .A(n559), .B(n3753), .Y(n1619) );
  INVX1 U321 ( .A(n1619), .Y(n2546) );
  AND2X1 U322 ( .A(n3400), .B(n3705), .Y(n1616) );
  INVX1 U323 ( .A(n1616), .Y(n2547) );
  AND2X1 U324 ( .A(n559), .B(n3881), .Y(n1612) );
  INVX1 U325 ( .A(n1612), .Y(n2548) );
  AND2X1 U326 ( .A(n3400), .B(n3833), .Y(n1608) );
  INVX1 U327 ( .A(n1608), .Y(n2549) );
  AND2X1 U328 ( .A(n559), .B(n3497), .Y(n1604) );
  INVX1 U329 ( .A(n1604), .Y(n2550) );
  AND2X1 U330 ( .A(n3400), .B(n3449), .Y(n1600) );
  INVX1 U331 ( .A(n1600), .Y(n2551) );
  AND2X1 U332 ( .A(n559), .B(n3625), .Y(n1596) );
  INVX1 U333 ( .A(n1596), .Y(n2552) );
  AND2X1 U334 ( .A(n3400), .B(n3577), .Y(n1592) );
  INVX1 U335 ( .A(n1592), .Y(n2553) );
  AND2X1 U336 ( .A(n3405), .B(n3752), .Y(n1582) );
  INVX1 U337 ( .A(n1582), .Y(n2554) );
  AND2X1 U338 ( .A(n3400), .B(n3704), .Y(n1579) );
  INVX1 U339 ( .A(n1579), .Y(n2555) );
  AND2X1 U340 ( .A(n3405), .B(n3880), .Y(n1575) );
  INVX1 U341 ( .A(n1575), .Y(n2556) );
  AND2X1 U342 ( .A(n3400), .B(n3832), .Y(n1572) );
  INVX1 U343 ( .A(n1572), .Y(n2557) );
  AND2X1 U344 ( .A(n3405), .B(n3496), .Y(n1568) );
  INVX1 U345 ( .A(n1568), .Y(n2558) );
  AND2X1 U346 ( .A(n3400), .B(n3448), .Y(n1565) );
  INVX1 U347 ( .A(n1565), .Y(n2559) );
  AND2X1 U348 ( .A(n3405), .B(n3624), .Y(n1561) );
  INVX1 U349 ( .A(n1561), .Y(n2560) );
  AND2X1 U350 ( .A(n3400), .B(n3576), .Y(n1558) );
  INVX1 U351 ( .A(n1558), .Y(n2561) );
  AND2X1 U352 ( .A(n3405), .B(n3751), .Y(n1548) );
  INVX1 U353 ( .A(n1548), .Y(n2562) );
  AND2X1 U354 ( .A(n3400), .B(n3703), .Y(n1545) );
  INVX1 U355 ( .A(n1545), .Y(n2563) );
  AND2X1 U356 ( .A(n3405), .B(n3879), .Y(n1541) );
  INVX1 U357 ( .A(n1541), .Y(n2564) );
  AND2X1 U358 ( .A(n3400), .B(n3831), .Y(n1538) );
  INVX1 U359 ( .A(n1538), .Y(n2565) );
  AND2X1 U360 ( .A(n3405), .B(n3495), .Y(n1534) );
  INVX1 U361 ( .A(n1534), .Y(n2566) );
  AND2X1 U362 ( .A(n3400), .B(n3447), .Y(n1531) );
  INVX1 U363 ( .A(n1531), .Y(n2567) );
  AND2X1 U364 ( .A(n3405), .B(n3623), .Y(n1527) );
  INVX1 U365 ( .A(n1527), .Y(n2568) );
  AND2X1 U366 ( .A(n3400), .B(n3575), .Y(n1524) );
  INVX1 U367 ( .A(n1524), .Y(n2569) );
  AND2X1 U368 ( .A(n3405), .B(n3750), .Y(n1514) );
  INVX1 U369 ( .A(n1514), .Y(n2570) );
  AND2X1 U370 ( .A(n3400), .B(n3702), .Y(n1511) );
  INVX1 U371 ( .A(n1511), .Y(n2571) );
  AND2X1 U372 ( .A(n3405), .B(n3878), .Y(n1507) );
  INVX1 U373 ( .A(n1507), .Y(n2572) );
  AND2X1 U374 ( .A(n3400), .B(n3830), .Y(n1504) );
  INVX1 U375 ( .A(n1504), .Y(n2573) );
  AND2X1 U376 ( .A(n3405), .B(n3494), .Y(n1500) );
  INVX1 U377 ( .A(n1500), .Y(n2574) );
  AND2X1 U378 ( .A(n3400), .B(n3446), .Y(n1497) );
  INVX1 U379 ( .A(n1497), .Y(n2575) );
  AND2X1 U380 ( .A(n3405), .B(n3622), .Y(n1493) );
  INVX1 U381 ( .A(n1493), .Y(n2576) );
  AND2X1 U382 ( .A(n3400), .B(n3574), .Y(n1490) );
  INVX1 U383 ( .A(n1490), .Y(n2577) );
  AND2X1 U384 ( .A(n559), .B(n3749), .Y(n1480) );
  INVX1 U385 ( .A(n1480), .Y(n2578) );
  AND2X1 U386 ( .A(n3400), .B(n3701), .Y(n1477) );
  INVX1 U387 ( .A(n1477), .Y(n2579) );
  AND2X1 U388 ( .A(n559), .B(n3877), .Y(n1473) );
  INVX1 U389 ( .A(n1473), .Y(n2580) );
  AND2X1 U390 ( .A(n3400), .B(n3829), .Y(n1470) );
  INVX1 U391 ( .A(n1470), .Y(n2581) );
  AND2X1 U392 ( .A(n559), .B(n3493), .Y(n1466) );
  INVX1 U393 ( .A(n1466), .Y(n2582) );
  AND2X1 U394 ( .A(n3400), .B(n3445), .Y(n1463) );
  INVX1 U395 ( .A(n1463), .Y(n2583) );
  AND2X1 U396 ( .A(n559), .B(n3621), .Y(n1459) );
  INVX1 U397 ( .A(n1459), .Y(n2584) );
  AND2X1 U398 ( .A(n3400), .B(n3573), .Y(n1456) );
  INVX1 U399 ( .A(n1456), .Y(n2585) );
  AND2X1 U400 ( .A(n559), .B(n3748), .Y(n1446) );
  INVX1 U401 ( .A(n1446), .Y(n2586) );
  AND2X1 U402 ( .A(n3400), .B(n3700), .Y(n1443) );
  INVX1 U403 ( .A(n1443), .Y(n2587) );
  AND2X1 U404 ( .A(n559), .B(n3876), .Y(n1439) );
  INVX1 U405 ( .A(n1439), .Y(n2588) );
  AND2X1 U406 ( .A(n3400), .B(n3828), .Y(n1436) );
  INVX1 U407 ( .A(n1436), .Y(n2589) );
  AND2X1 U408 ( .A(n559), .B(n3492), .Y(n1432) );
  INVX1 U409 ( .A(n1432), .Y(n2590) );
  AND2X1 U410 ( .A(n3400), .B(n3444), .Y(n1429) );
  INVX1 U411 ( .A(n1429), .Y(n2591) );
  AND2X1 U412 ( .A(n559), .B(n3620), .Y(n1425) );
  INVX1 U413 ( .A(n1425), .Y(n2592) );
  AND2X1 U414 ( .A(n3400), .B(n3572), .Y(n1422) );
  INVX1 U415 ( .A(n1422), .Y(n2593) );
  AND2X1 U416 ( .A(n559), .B(n3747), .Y(n890) );
  INVX1 U417 ( .A(n890), .Y(n2594) );
  AND2X1 U418 ( .A(n3400), .B(n3699), .Y(n887) );
  INVX1 U419 ( .A(n887), .Y(n2595) );
  AND2X1 U420 ( .A(n559), .B(n3875), .Y(n883) );
  INVX1 U421 ( .A(n883), .Y(n2596) );
  AND2X1 U422 ( .A(n3400), .B(n3827), .Y(n880) );
  INVX1 U423 ( .A(n880), .Y(n2597) );
  AND2X1 U424 ( .A(n559), .B(n3491), .Y(n876) );
  INVX1 U425 ( .A(n876), .Y(n2598) );
  AND2X1 U426 ( .A(n3400), .B(n3443), .Y(n873) );
  INVX1 U427 ( .A(n873), .Y(n2599) );
  AND2X1 U428 ( .A(n559), .B(n3619), .Y(n869) );
  INVX1 U429 ( .A(n869), .Y(n2600) );
  AND2X1 U430 ( .A(n3400), .B(n3571), .Y(n866) );
  INVX1 U431 ( .A(n866), .Y(n2601) );
  AND2X1 U432 ( .A(n559), .B(n3746), .Y(n856) );
  INVX1 U433 ( .A(n856), .Y(n2602) );
  AND2X1 U434 ( .A(n3400), .B(n3698), .Y(n853) );
  INVX1 U435 ( .A(n853), .Y(n2603) );
  AND2X1 U436 ( .A(n559), .B(n3874), .Y(n849) );
  INVX1 U437 ( .A(n849), .Y(n2604) );
  AND2X1 U438 ( .A(n3400), .B(n3826), .Y(n846) );
  INVX1 U439 ( .A(n846), .Y(n2605) );
  AND2X1 U440 ( .A(n559), .B(n3490), .Y(n842) );
  INVX1 U441 ( .A(n842), .Y(n2606) );
  AND2X1 U442 ( .A(n3400), .B(n3442), .Y(n839) );
  INVX1 U443 ( .A(n839), .Y(n2607) );
  AND2X1 U444 ( .A(n559), .B(n3618), .Y(n835) );
  INVX1 U445 ( .A(n835), .Y(n2608) );
  AND2X1 U446 ( .A(n3400), .B(n3570), .Y(n832) );
  INVX1 U447 ( .A(n832), .Y(n2609) );
  AND2X1 U448 ( .A(n559), .B(n3745), .Y(n822) );
  INVX1 U449 ( .A(n822), .Y(n2610) );
  AND2X1 U450 ( .A(n3400), .B(n3697), .Y(n819) );
  INVX1 U451 ( .A(n819), .Y(n2611) );
  AND2X1 U452 ( .A(n559), .B(n3873), .Y(n815) );
  INVX1 U453 ( .A(n815), .Y(n2612) );
  AND2X1 U454 ( .A(n3400), .B(n3825), .Y(n812) );
  INVX1 U455 ( .A(n812), .Y(n2613) );
  AND2X1 U456 ( .A(n559), .B(n3489), .Y(n808) );
  INVX1 U457 ( .A(n808), .Y(n2614) );
  AND2X1 U458 ( .A(n3400), .B(n3441), .Y(n805) );
  INVX1 U459 ( .A(n805), .Y(n2615) );
  AND2X1 U460 ( .A(n559), .B(n3617), .Y(n801) );
  INVX1 U461 ( .A(n801), .Y(n2616) );
  AND2X1 U462 ( .A(n3400), .B(n3569), .Y(n798) );
  INVX1 U463 ( .A(n798), .Y(n2617) );
  AND2X1 U464 ( .A(n559), .B(n3744), .Y(n788) );
  INVX1 U465 ( .A(n788), .Y(n2618) );
  AND2X1 U466 ( .A(n3400), .B(n3696), .Y(n785) );
  INVX1 U467 ( .A(n785), .Y(n2619) );
  AND2X1 U468 ( .A(n559), .B(n3872), .Y(n781) );
  INVX1 U469 ( .A(n781), .Y(n2620) );
  AND2X1 U470 ( .A(n3400), .B(n3824), .Y(n778) );
  INVX1 U471 ( .A(n778), .Y(n2621) );
  AND2X1 U472 ( .A(n559), .B(n3488), .Y(n774) );
  INVX1 U473 ( .A(n774), .Y(n2622) );
  AND2X1 U474 ( .A(n3400), .B(n3440), .Y(n771) );
  INVX1 U475 ( .A(n771), .Y(n2623) );
  AND2X1 U476 ( .A(n559), .B(n3616), .Y(n767) );
  INVX1 U477 ( .A(n767), .Y(n2624) );
  AND2X1 U478 ( .A(n3400), .B(n3568), .Y(n764) );
  INVX1 U479 ( .A(n764), .Y(n2625) );
  AND2X1 U480 ( .A(n559), .B(n3743), .Y(n754) );
  INVX1 U481 ( .A(n754), .Y(n2626) );
  AND2X1 U482 ( .A(n3400), .B(n3695), .Y(n751) );
  INVX1 U483 ( .A(n751), .Y(n2627) );
  AND2X1 U484 ( .A(n559), .B(n3871), .Y(n747) );
  INVX1 U485 ( .A(n747), .Y(n2628) );
  AND2X1 U486 ( .A(n3400), .B(n3823), .Y(n744) );
  INVX1 U487 ( .A(n744), .Y(n2629) );
  AND2X1 U488 ( .A(n559), .B(n3487), .Y(n740) );
  INVX1 U489 ( .A(n740), .Y(n2630) );
  AND2X1 U490 ( .A(n3400), .B(n3439), .Y(n737) );
  INVX1 U491 ( .A(n737), .Y(n2631) );
  AND2X1 U492 ( .A(n559), .B(n3615), .Y(n733) );
  INVX1 U493 ( .A(n733), .Y(n2632) );
  AND2X1 U494 ( .A(n3400), .B(n3567), .Y(n730) );
  INVX1 U495 ( .A(n730), .Y(n2633) );
  AND2X1 U496 ( .A(n559), .B(n3742), .Y(n720) );
  INVX1 U497 ( .A(n720), .Y(n2634) );
  AND2X1 U498 ( .A(n3400), .B(n3694), .Y(n717) );
  INVX1 U499 ( .A(n717), .Y(n2635) );
  AND2X1 U500 ( .A(n559), .B(n3870), .Y(n713) );
  INVX1 U501 ( .A(n713), .Y(n2636) );
  AND2X1 U502 ( .A(n3400), .B(n3822), .Y(n710) );
  INVX1 U503 ( .A(n710), .Y(n2637) );
  AND2X1 U504 ( .A(n559), .B(n3486), .Y(n706) );
  INVX1 U505 ( .A(n706), .Y(n2638) );
  AND2X1 U506 ( .A(n3400), .B(n3438), .Y(n703) );
  INVX1 U507 ( .A(n703), .Y(n2639) );
  AND2X1 U508 ( .A(n559), .B(n3614), .Y(n699) );
  INVX1 U509 ( .A(n699), .Y(n2640) );
  AND2X1 U510 ( .A(n3400), .B(n3566), .Y(n696) );
  INVX1 U511 ( .A(n696), .Y(n2641) );
  AND2X1 U512 ( .A(n559), .B(n3741), .Y(n686) );
  INVX1 U513 ( .A(n686), .Y(n2642) );
  AND2X1 U514 ( .A(n3400), .B(n3693), .Y(n683) );
  INVX1 U515 ( .A(n683), .Y(n2643) );
  AND2X1 U516 ( .A(n559), .B(n3869), .Y(n679) );
  INVX1 U517 ( .A(n679), .Y(n2644) );
  AND2X1 U518 ( .A(n3400), .B(n3821), .Y(n676) );
  INVX1 U519 ( .A(n676), .Y(n2645) );
  AND2X1 U520 ( .A(n559), .B(n3485), .Y(n672) );
  INVX1 U521 ( .A(n672), .Y(n2646) );
  AND2X1 U522 ( .A(n3400), .B(n3437), .Y(n669) );
  INVX1 U523 ( .A(n669), .Y(n2647) );
  AND2X1 U524 ( .A(n559), .B(n3613), .Y(n665) );
  INVX1 U525 ( .A(n665), .Y(n2648) );
  AND2X1 U526 ( .A(n3400), .B(n3565), .Y(n662) );
  INVX1 U527 ( .A(n662), .Y(n2649) );
  AND2X1 U528 ( .A(n559), .B(n3740), .Y(n652) );
  INVX1 U529 ( .A(n652), .Y(n2650) );
  AND2X1 U530 ( .A(n3400), .B(n3692), .Y(n649) );
  INVX1 U531 ( .A(n649), .Y(n2651) );
  AND2X1 U532 ( .A(n559), .B(n3868), .Y(n645) );
  INVX1 U533 ( .A(n645), .Y(n2652) );
  AND2X1 U534 ( .A(n3400), .B(n3820), .Y(n642) );
  INVX1 U535 ( .A(n642), .Y(n2653) );
  AND2X1 U536 ( .A(n559), .B(n3484), .Y(n638) );
  INVX1 U537 ( .A(n638), .Y(n2654) );
  AND2X1 U538 ( .A(n3400), .B(n3436), .Y(n635) );
  INVX1 U539 ( .A(n635), .Y(n2655) );
  AND2X1 U540 ( .A(n559), .B(n3612), .Y(n631) );
  INVX1 U541 ( .A(n631), .Y(n2656) );
  AND2X1 U542 ( .A(n3400), .B(n3564), .Y(n628) );
  INVX1 U543 ( .A(n628), .Y(n2657) );
  AND2X1 U544 ( .A(n559), .B(n3739), .Y(n618) );
  INVX1 U545 ( .A(n618), .Y(n2658) );
  AND2X1 U546 ( .A(n3400), .B(n3691), .Y(n615) );
  INVX1 U547 ( .A(n615), .Y(n2659) );
  AND2X1 U548 ( .A(n559), .B(n3867), .Y(n611) );
  INVX1 U549 ( .A(n611), .Y(n2660) );
  AND2X1 U550 ( .A(n3400), .B(n3819), .Y(n608) );
  INVX1 U551 ( .A(n608), .Y(n2661) );
  AND2X1 U552 ( .A(n559), .B(n3483), .Y(n604) );
  INVX1 U553 ( .A(n604), .Y(n2662) );
  AND2X1 U554 ( .A(n3400), .B(n3435), .Y(n601) );
  INVX1 U555 ( .A(n601), .Y(n2663) );
  AND2X1 U556 ( .A(n559), .B(n3611), .Y(n597) );
  INVX1 U557 ( .A(n597), .Y(n2664) );
  AND2X1 U558 ( .A(n3400), .B(n3563), .Y(n594) );
  INVX1 U559 ( .A(n594), .Y(n2665) );
  AND2X1 U560 ( .A(n559), .B(n3738), .Y(n584) );
  INVX1 U561 ( .A(n584), .Y(n2666) );
  AND2X1 U562 ( .A(n3400), .B(n3690), .Y(n581) );
  INVX1 U563 ( .A(n581), .Y(n2667) );
  AND2X1 U564 ( .A(n559), .B(n3866), .Y(n576) );
  INVX1 U565 ( .A(n576), .Y(n2668) );
  AND2X1 U566 ( .A(n3400), .B(n3818), .Y(n573) );
  INVX1 U567 ( .A(n573), .Y(n2669) );
  AND2X1 U568 ( .A(n559), .B(n3482), .Y(n568) );
  INVX1 U569 ( .A(n568), .Y(n2670) );
  AND2X1 U570 ( .A(n3400), .B(n3434), .Y(n565) );
  INVX1 U571 ( .A(n565), .Y(n2671) );
  AND2X1 U572 ( .A(n559), .B(n3610), .Y(n555) );
  INVX1 U573 ( .A(n555), .Y(n2672) );
  AND2X1 U574 ( .A(n3400), .B(n3562), .Y(n550) );
  INVX1 U575 ( .A(n550), .Y(n2673) );
  BUFX2 U576 ( .A(n1769), .Y(n2674) );
  BUFX2 U577 ( .A(n1620), .Y(n2675) );
  BUFX2 U578 ( .A(n1617), .Y(n2676) );
  BUFX2 U579 ( .A(n1613), .Y(n2677) );
  BUFX2 U580 ( .A(n1609), .Y(n2678) );
  BUFX2 U581 ( .A(n1605), .Y(n2679) );
  BUFX2 U582 ( .A(n1601), .Y(n2680) );
  BUFX2 U585 ( .A(n1597), .Y(n2681) );
  BUFX2 U588 ( .A(n1593), .Y(n2682) );
  BUFX2 U591 ( .A(n1583), .Y(n2683) );
  BUFX2 U593 ( .A(n1580), .Y(n2684) );
  BUFX2 U596 ( .A(n1576), .Y(n2685) );
  BUFX2 U599 ( .A(n1573), .Y(n2686) );
  BUFX2 U601 ( .A(n1569), .Y(n2687) );
  BUFX2 U604 ( .A(n1566), .Y(n2688) );
  BUFX2 U607 ( .A(n1562), .Y(n2689) );
  BUFX2 U611 ( .A(n1559), .Y(n2690) );
  BUFX2 U614 ( .A(n1549), .Y(n2691) );
  BUFX2 U616 ( .A(n1546), .Y(n2692) );
  BUFX2 U619 ( .A(n1542), .Y(n2693) );
  BUFX2 U622 ( .A(n1539), .Y(n2694) );
  BUFX2 U625 ( .A(n1535), .Y(n2695) );
  BUFX2 U627 ( .A(n1532), .Y(n2696) );
  BUFX2 U630 ( .A(n1528), .Y(n2697) );
  BUFX2 U633 ( .A(n1525), .Y(n2698) );
  BUFX2 U635 ( .A(n1515), .Y(n2699) );
  BUFX2 U638 ( .A(n1512), .Y(n2700) );
  BUFX2 U641 ( .A(n1508), .Y(n2701) );
  BUFX2 U645 ( .A(n1505), .Y(n2702) );
  BUFX2 U648 ( .A(n1501), .Y(n2703) );
  BUFX2 U650 ( .A(n1498), .Y(n2704) );
  BUFX2 U653 ( .A(n1494), .Y(n2705) );
  BUFX2 U656 ( .A(n1491), .Y(n2706) );
  BUFX2 U659 ( .A(n1481), .Y(n2707) );
  BUFX2 U661 ( .A(n1478), .Y(n2708) );
  BUFX2 U664 ( .A(n1474), .Y(n2709) );
  BUFX2 U667 ( .A(n1471), .Y(n2710) );
  BUFX2 U669 ( .A(n1467), .Y(n2711) );
  BUFX2 U672 ( .A(n1464), .Y(n2712) );
  BUFX2 U675 ( .A(n1460), .Y(n2713) );
  BUFX2 U679 ( .A(n1457), .Y(n2714) );
  BUFX2 U682 ( .A(n1447), .Y(n2715) );
  BUFX2 U684 ( .A(n1444), .Y(n2716) );
  BUFX2 U687 ( .A(n1440), .Y(n2717) );
  BUFX2 U690 ( .A(n1437), .Y(n2718) );
  BUFX2 U693 ( .A(n1433), .Y(n2719) );
  BUFX2 U695 ( .A(n1430), .Y(n2720) );
  BUFX2 U698 ( .A(n1426), .Y(n2721) );
  BUFX2 U701 ( .A(n1423), .Y(n2722) );
  BUFX2 U703 ( .A(n891), .Y(n2723) );
  BUFX2 U706 ( .A(n888), .Y(n2724) );
  BUFX2 U709 ( .A(n884), .Y(n2725) );
  BUFX2 U713 ( .A(n881), .Y(n2726) );
  BUFX2 U716 ( .A(n877), .Y(n2727) );
  BUFX2 U718 ( .A(n874), .Y(n2728) );
  BUFX2 U721 ( .A(n870), .Y(n2729) );
  BUFX2 U724 ( .A(n867), .Y(n2730) );
  BUFX2 U727 ( .A(n857), .Y(n2731) );
  BUFX2 U729 ( .A(n854), .Y(n2732) );
  BUFX2 U732 ( .A(n850), .Y(n2733) );
  BUFX2 U735 ( .A(n847), .Y(n2734) );
  BUFX2 U737 ( .A(n843), .Y(n2735) );
  BUFX2 U740 ( .A(n840), .Y(n2736) );
  BUFX2 U743 ( .A(n836), .Y(n2737) );
  BUFX2 U747 ( .A(n833), .Y(n2738) );
  BUFX2 U750 ( .A(n823), .Y(n2739) );
  BUFX2 U752 ( .A(n820), .Y(n2740) );
  BUFX2 U755 ( .A(n816), .Y(n2741) );
  BUFX2 U758 ( .A(n813), .Y(n2742) );
  BUFX2 U761 ( .A(n809), .Y(n2743) );
  BUFX2 U763 ( .A(n806), .Y(n2744) );
  BUFX2 U766 ( .A(n802), .Y(n2745) );
  BUFX2 U769 ( .A(n799), .Y(n2746) );
  BUFX2 U771 ( .A(n789), .Y(n2747) );
  BUFX2 U774 ( .A(n786), .Y(n2748) );
  BUFX2 U777 ( .A(n782), .Y(n2749) );
  BUFX2 U781 ( .A(n779), .Y(n2750) );
  BUFX2 U784 ( .A(n775), .Y(n2751) );
  BUFX2 U786 ( .A(n772), .Y(n2752) );
  BUFX2 U789 ( .A(n768), .Y(n2753) );
  BUFX2 U792 ( .A(n765), .Y(n2754) );
  BUFX2 U795 ( .A(n755), .Y(n2755) );
  BUFX2 U797 ( .A(n752), .Y(n2756) );
  BUFX2 U800 ( .A(n748), .Y(n2757) );
  BUFX2 U803 ( .A(n745), .Y(n2758) );
  BUFX2 U805 ( .A(n741), .Y(n2759) );
  BUFX2 U808 ( .A(n738), .Y(n2760) );
  BUFX2 U811 ( .A(n734), .Y(n2761) );
  BUFX2 U815 ( .A(n731), .Y(n2762) );
  BUFX2 U818 ( .A(n721), .Y(n2763) );
  BUFX2 U820 ( .A(n718), .Y(n2764) );
  BUFX2 U823 ( .A(n714), .Y(n2765) );
  BUFX2 U826 ( .A(n711), .Y(n2766) );
  BUFX2 U829 ( .A(n707), .Y(n2767) );
  BUFX2 U831 ( .A(n704), .Y(n2768) );
  BUFX2 U834 ( .A(n700), .Y(n2769) );
  BUFX2 U837 ( .A(n697), .Y(n2770) );
  BUFX2 U839 ( .A(n687), .Y(n2771) );
  BUFX2 U842 ( .A(n684), .Y(n2772) );
  BUFX2 U845 ( .A(n680), .Y(n2773) );
  BUFX2 U849 ( .A(n677), .Y(n2774) );
  BUFX2 U852 ( .A(n673), .Y(n2775) );
  BUFX2 U854 ( .A(n670), .Y(n2776) );
  BUFX2 U857 ( .A(n666), .Y(n2777) );
  BUFX2 U860 ( .A(n663), .Y(n2778) );
  BUFX2 U863 ( .A(n653), .Y(n2779) );
  BUFX2 U865 ( .A(n650), .Y(n2780) );
  BUFX2 U868 ( .A(n646), .Y(n2781) );
  BUFX2 U871 ( .A(n643), .Y(n2782) );
  BUFX2 U873 ( .A(n639), .Y(n2783) );
  BUFX2 U876 ( .A(n636), .Y(n2784) );
  BUFX2 U879 ( .A(n632), .Y(n2785) );
  BUFX2 U883 ( .A(n629), .Y(n2786) );
  BUFX2 U886 ( .A(n619), .Y(n2787) );
  BUFX2 U888 ( .A(n616), .Y(n2788) );
  BUFX2 U891 ( .A(n612), .Y(n2789) );
  BUFX2 U894 ( .A(n609), .Y(n2790) );
  BUFX2 U897 ( .A(n605), .Y(n2791) );
  BUFX2 U899 ( .A(n602), .Y(n2792) );
  BUFX2 U902 ( .A(n598), .Y(n2793) );
  BUFX2 U905 ( .A(n595), .Y(n2794) );
  BUFX2 U907 ( .A(n585), .Y(n2795) );
  BUFX2 U910 ( .A(n582), .Y(n2796) );
  BUFX2 U913 ( .A(n577), .Y(n2797) );
  BUFX2 U917 ( .A(n574), .Y(n2798) );
  BUFX2 U920 ( .A(n569), .Y(n2799) );
  BUFX2 U922 ( .A(n566), .Y(n2800) );
  BUFX2 U925 ( .A(n556), .Y(n2801) );
  BUFX2 U928 ( .A(n551), .Y(n2802) );
  INVX1 U931 ( .A(n1587), .Y(n2803) );
  INVX1 U933 ( .A(n1553), .Y(n2804) );
  INVX1 U936 ( .A(n1519), .Y(n2805) );
  INVX1 U939 ( .A(n1485), .Y(n2806) );
  INVX1 U941 ( .A(n1451), .Y(n2807) );
  INVX1 U944 ( .A(n1417), .Y(n2808) );
  INVX1 U947 ( .A(n861), .Y(n2809) );
  INVX1 U951 ( .A(n827), .Y(n2810) );
  INVX1 U954 ( .A(n793), .Y(n2811) );
  INVX1 U956 ( .A(n759), .Y(n2812) );
  INVX1 U959 ( .A(n725), .Y(n2813) );
  INVX1 U962 ( .A(n691), .Y(n2814) );
  INVX1 U965 ( .A(n657), .Y(n2815) );
  INVX1 U967 ( .A(n623), .Y(n2816) );
  INVX1 U970 ( .A(n589), .Y(n2817) );
  INVX1 U973 ( .A(n545), .Y(n2818) );
  INVX1 U975 ( .A(n1588), .Y(n2819) );
  INVX1 U978 ( .A(n1554), .Y(n2820) );
  INVX1 U981 ( .A(n1520), .Y(n2821) );
  INVX1 U985 ( .A(n1486), .Y(n2822) );
  INVX1 U988 ( .A(n1452), .Y(n2823) );
  INVX1 U990 ( .A(n1418), .Y(n2824) );
  INVX1 U993 ( .A(n862), .Y(n2825) );
  INVX1 U996 ( .A(n828), .Y(n2826) );
  INVX1 U999 ( .A(n794), .Y(n2827) );
  INVX1 U1001 ( .A(n760), .Y(n2828) );
  INVX1 U1004 ( .A(n726), .Y(n2829) );
  INVX1 U1007 ( .A(n692), .Y(n2830) );
  INVX1 U1009 ( .A(n658), .Y(n2831) );
  INVX1 U1012 ( .A(n624), .Y(n2832) );
  INVX1 U1015 ( .A(n590), .Y(n2833) );
  INVX1 U1019 ( .A(n546), .Y(n2834) );
  INVX1 U1022 ( .A(n1589), .Y(n2835) );
  INVX1 U1024 ( .A(n1555), .Y(n2836) );
  INVX1 U1027 ( .A(n1521), .Y(n2837) );
  INVX1 U1030 ( .A(n1487), .Y(n2838) );
  INVX1 U1033 ( .A(n1453), .Y(n2839) );
  INVX1 U1035 ( .A(n1419), .Y(n2840) );
  INVX1 U1038 ( .A(n863), .Y(n2841) );
  INVX1 U1041 ( .A(n829), .Y(n2842) );
  INVX1 U1043 ( .A(n795), .Y(n2843) );
  INVX1 U1046 ( .A(n761), .Y(n2844) );
  INVX1 U1049 ( .A(n727), .Y(n2845) );
  INVX1 U1053 ( .A(n693), .Y(n2846) );
  INVX1 U1056 ( .A(n659), .Y(n2847) );
  INVX1 U1058 ( .A(n625), .Y(n2848) );
  INVX1 U1061 ( .A(n591), .Y(n2849) );
  INVX1 U1064 ( .A(n547), .Y(n2850) );
  AND2X1 U1067 ( .A(n1629), .B(n1794), .Y(n1799) );
  INVX1 U1069 ( .A(n1799), .Y(n2851) );
  AND2X1 U1072 ( .A(n1643), .B(n1794), .Y(n1806) );
  INVX1 U1075 ( .A(n1806), .Y(n2852) );
  AND2X1 U1077 ( .A(n1660), .B(n1812), .Y(n1816) );
  INVX1 U1080 ( .A(n1816), .Y(n2853) );
  AND2X1 U1083 ( .A(n1641), .B(n1812), .Y(n1823) );
  INVX1 U1087 ( .A(n1823), .Y(n2854) );
  AND2X1 U1090 ( .A(n1658), .B(n1830), .Y(n1833) );
  INVX1 U1092 ( .A(n1833), .Y(n2855) );
  AND2X1 U1095 ( .A(n1639), .B(n1830), .Y(n1840) );
  INVX1 U1098 ( .A(n1840), .Y(n2856) );
  AND2X1 U1101 ( .A(n1637), .B(n1847), .Y(n1856) );
  INVX1 U1103 ( .A(n1856), .Y(n2857) );
  AND2X1 U1106 ( .A(n1633), .B(n1864), .Y(n1871) );
  INVX1 U1109 ( .A(n1871), .Y(n2858) );
  AND2X1 U1111 ( .A(n1631), .B(n1881), .Y(n1887) );
  INVX1 U1114 ( .A(n1887), .Y(n2859) );
  AND2X1 U1118 ( .A(n1643), .B(n1881), .Y(n1893) );
  INVX1 U1123 ( .A(n1893), .Y(n2860) );
  AND2X1 U1126 ( .A(n1629), .B(n1898), .Y(n1903) );
  INVX1 U1128 ( .A(n1903), .Y(n2861) );
  AND2X1 U1132 ( .A(n1641), .B(n1898), .Y(n1909) );
  INVX1 U1134 ( .A(n1909), .Y(n2862) );
  AND2X1 U1136 ( .A(n1660), .B(n1915), .Y(n1919) );
  INVX1 U1138 ( .A(n1919), .Y(n2863) );
  AND2X1 U1140 ( .A(n1639), .B(n1915), .Y(n1925) );
  INVX1 U1142 ( .A(n1925), .Y(n2864) );
  AND2X1 U1144 ( .A(n1658), .B(n1932), .Y(n1935) );
  INVX1 U1146 ( .A(n1935), .Y(n2865) );
  AND2X1 U1148 ( .A(n1637), .B(n1932), .Y(n1941) );
  INVX1 U1150 ( .A(n1941), .Y(n2866) );
  AND2X1 U1152 ( .A(n1635), .B(n1950), .Y(n1958) );
  INVX1 U1154 ( .A(n1958), .Y(n2867) );
  AND2X1 U1156 ( .A(n1633), .B(n1967), .Y(n1974) );
  INVX1 U1158 ( .A(n1974), .Y(n2868) );
  AND2X1 U1160 ( .A(n1656), .B(n1984), .Y(n1986) );
  INVX1 U1162 ( .A(n1986), .Y(n2869) );
  AND2X1 U1164 ( .A(n1654), .B(n2001), .Y(n2002) );
  INVX1 U1166 ( .A(n2002), .Y(n2870) );
  AND2X1 U1168 ( .A(n1635), .B(n2087), .Y(n2095) );
  INVX1 U1170 ( .A(n2095), .Y(n2871) );
  AND2X1 U1172 ( .A(n1633), .B(n2104), .Y(n2111) );
  INVX1 U1174 ( .A(n2111), .Y(n2872) );
  AND2X1 U1176 ( .A(n1656), .B(n2121), .Y(n2123) );
  INVX1 U1178 ( .A(n2123), .Y(n2873) );
  AND2X1 U1180 ( .A(n1654), .B(n2138), .Y(n2139) );
  INVX1 U1182 ( .A(n2139), .Y(n2874) );
  AND2X1 U1184 ( .A(n1656), .B(n1652), .Y(n1655) );
  INVX1 U1186 ( .A(n1655), .Y(n2875) );
  AND2X1 U1189 ( .A(n1654), .B(n1675), .Y(n1676) );
  INVX1 U1191 ( .A(n1676), .Y(n2876) );
  AND2X1 U1193 ( .A(n1631), .B(n1794), .Y(n1800) );
  INVX1 U1195 ( .A(n1800), .Y(n2877) );
  AND2X1 U1197 ( .A(n1641), .B(n1794), .Y(n1805) );
  INVX1 U1199 ( .A(n1805), .Y(n2878) );
  AND2X1 U1201 ( .A(n1658), .B(n1812), .Y(n1815) );
  INVX1 U1203 ( .A(n1815), .Y(n2879) );
  AND2X1 U1205 ( .A(n1643), .B(n1812), .Y(n1824) );
  INVX1 U1207 ( .A(n1824), .Y(n2880) );
  AND2X1 U1209 ( .A(n1660), .B(n1830), .Y(n1834) );
  INVX1 U1211 ( .A(n1834), .Y(n2881) );
  AND2X1 U1213 ( .A(n1637), .B(n1830), .Y(n1839) );
  INVX1 U1215 ( .A(n1839), .Y(n2882) );
  AND2X1 U1217 ( .A(n1639), .B(n1847), .Y(n1857) );
  INVX1 U1219 ( .A(n1857), .Y(n2883) );
  AND2X1 U1222 ( .A(n1635), .B(n1864), .Y(n1872) );
  INVX1 U1224 ( .A(n1872), .Y(n2884) );
  AND2X1 U1226 ( .A(n1629), .B(n1881), .Y(n1886) );
  INVX1 U1228 ( .A(n1886), .Y(n2885) );
  AND2X1 U1230 ( .A(n1641), .B(n1881), .Y(n1892) );
  INVX1 U1232 ( .A(n1892), .Y(n2886) );
  AND2X1 U1234 ( .A(n1631), .B(n1898), .Y(n1904) );
  INVX1 U1236 ( .A(n1904), .Y(n2887) );
  AND2X1 U1238 ( .A(n1643), .B(n1898), .Y(n1910) );
  INVX1 U1240 ( .A(n1910), .Y(n2888) );
  AND2X1 U1242 ( .A(n1658), .B(n1915), .Y(n1918) );
  INVX1 U1244 ( .A(n1918), .Y(n2889) );
  AND2X1 U1246 ( .A(n1637), .B(n1915), .Y(n1924) );
  INVX1 U1248 ( .A(n1924), .Y(n2890) );
  AND2X1 U1250 ( .A(n1660), .B(n1932), .Y(n1936) );
  INVX1 U1252 ( .A(n1936), .Y(n2891) );
  AND2X1 U1255 ( .A(n1639), .B(n1932), .Y(n1942) );
  INVX1 U1257 ( .A(n1942), .Y(n2892) );
  AND2X1 U1259 ( .A(n1633), .B(n1950), .Y(n1957) );
  INVX1 U1261 ( .A(n1957), .Y(n2893) );
  AND2X1 U1263 ( .A(n1635), .B(n1967), .Y(n1975) );
  INVX1 U1265 ( .A(n1975), .Y(n2894) );
  AND2X1 U1267 ( .A(n1654), .B(n1984), .Y(n1985) );
  INVX1 U1269 ( .A(n1985), .Y(n2895) );
  AND2X1 U1271 ( .A(n1656), .B(n2001), .Y(n2003) );
  INVX1 U1273 ( .A(n2003), .Y(n2896) );
  AND2X1 U1275 ( .A(n1633), .B(n2087), .Y(n2094) );
  INVX1 U1277 ( .A(n2094), .Y(n2897) );
  AND2X1 U1279 ( .A(n1635), .B(n2104), .Y(n2112) );
  INVX1 U1281 ( .A(n2112), .Y(n2898) );
  AND2X1 U1283 ( .A(n1654), .B(n2121), .Y(n2122) );
  INVX1 U1285 ( .A(n2122), .Y(n2899) );
  AND2X1 U1288 ( .A(n1656), .B(n2138), .Y(n2140) );
  INVX1 U1290 ( .A(n2140), .Y(n2900) );
  AND2X1 U1292 ( .A(n1654), .B(n1652), .Y(n1653) );
  INVX1 U1294 ( .A(n1653), .Y(n2901) );
  AND2X1 U1296 ( .A(n1656), .B(n1675), .Y(n1677) );
  INVX1 U1298 ( .A(n1677), .Y(n2902) );
  AND2X1 U1300 ( .A(n1660), .B(n1794), .Y(n1798) );
  INVX1 U1302 ( .A(n1798), .Y(n2903) );
  AND2X1 U1304 ( .A(n1639), .B(n1794), .Y(n1804) );
  INVX1 U1306 ( .A(n1804), .Y(n2904) );
  AND2X1 U1308 ( .A(n1631), .B(n1812), .Y(n1818) );
  INVX1 U1310 ( .A(n1818), .Y(n2905) );
  AND2X1 U1312 ( .A(n1637), .B(n1812), .Y(n1821) );
  INVX1 U1314 ( .A(n1821), .Y(n2906) );
  AND2X1 U1316 ( .A(n1629), .B(n1830), .Y(n1835) );
  INVX1 U1318 ( .A(n1835), .Y(n2907) );
  AND2X1 U1321 ( .A(n1643), .B(n1830), .Y(n1842) );
  INVX1 U1323 ( .A(n1842), .Y(n2908) );
  AND2X1 U1325 ( .A(n1658), .B(n1847), .Y(n1850) );
  INVX1 U1327 ( .A(n1850), .Y(n2909) );
  AND2X1 U1329 ( .A(n1641), .B(n1847), .Y(n1858) );
  INVX1 U1331 ( .A(n1858), .Y(n2910) );
  AND2X1 U1333 ( .A(n1654), .B(n1864), .Y(n1865) );
  INVX1 U1335 ( .A(n1865), .Y(n2911) );
  AND2X1 U1337 ( .A(n1639), .B(n1881), .Y(n1891) );
  INVX1 U1339 ( .A(n1891), .Y(n2912) );
  AND2X1 U1341 ( .A(n1658), .B(n1898), .Y(n1901) );
  INVX1 U1343 ( .A(n1901), .Y(n2913) );
  AND2X1 U1345 ( .A(n1637), .B(n1898), .Y(n1907) );
  INVX1 U1347 ( .A(n1907), .Y(n2914) );
  AND2X1 U1349 ( .A(n1631), .B(n1915), .Y(n1921) );
  INVX1 U1351 ( .A(n1921), .Y(n2915) );
  AND2X1 U1357 ( .A(n1643), .B(n1915), .Y(n1927) );
  INVX1 U1358 ( .A(n1927), .Y(n2916) );
  AND2X1 U1361 ( .A(n1629), .B(n1932), .Y(n1937) );
  INVX1 U1371 ( .A(n1937), .Y(n2917) );
  AND2X1 U1372 ( .A(n1641), .B(n1932), .Y(n1943) );
  INVX1 U1373 ( .A(n1943), .Y(n2918) );
  AND2X1 U1378 ( .A(n1656), .B(n1967), .Y(n1969) );
  INVX1 U1388 ( .A(n1969), .Y(n2919) );
  AND2X1 U1389 ( .A(n1635), .B(n1984), .Y(n1992) );
  INVX1 U1391 ( .A(n1992), .Y(n2920) );
  AND2X1 U1393 ( .A(n1633), .B(n2001), .Y(n2008) );
  INVX1 U1395 ( .A(n2008), .Y(n2921) );
  AND2X1 U1397 ( .A(n1654), .B(n2018), .Y(n2019) );
  INVX1 U1399 ( .A(n2019), .Y(n2922) );
  AND2X1 U1401 ( .A(n1656), .B(n2104), .Y(n2106) );
  INVX1 U1403 ( .A(n2106), .Y(n2923) );
  AND2X1 U1405 ( .A(n1635), .B(n2121), .Y(n2129) );
  INVX1 U1407 ( .A(n2129), .Y(n2924) );
  AND2X1 U1409 ( .A(n1633), .B(n2138), .Y(n2145) );
  INVX1 U1411 ( .A(n2145), .Y(n2925) );
  AND2X1 U1413 ( .A(n1654), .B(n1627), .Y(n2223) );
  INVX1 U1415 ( .A(n2223), .Y(n2926) );
  AND2X1 U1417 ( .A(n1635), .B(n1652), .Y(n1664) );
  INVX1 U1419 ( .A(n1664), .Y(n2927) );
  AND2X1 U1421 ( .A(n1633), .B(n1675), .Y(n1682) );
  INVX1 U1424 ( .A(n1682), .Y(n2928) );
  AND2X1 U1426 ( .A(n1658), .B(n1794), .Y(n1797) );
  INVX1 U1428 ( .A(n1797), .Y(n2929) );
  AND2X1 U1430 ( .A(n1637), .B(n1794), .Y(n1803) );
  INVX1 U1432 ( .A(n1803), .Y(n2930) );
  AND2X1 U1434 ( .A(n1629), .B(n1812), .Y(n1817) );
  INVX1 U1436 ( .A(n1817), .Y(n2931) );
  AND2X1 U1438 ( .A(n1639), .B(n1812), .Y(n1822) );
  INVX1 U1440 ( .A(n1822), .Y(n2932) );
  AND2X1 U1442 ( .A(n1631), .B(n1830), .Y(n1836) );
  INVX1 U1444 ( .A(n1836), .Y(n2933) );
  AND2X1 U1446 ( .A(n1641), .B(n1830), .Y(n1841) );
  INVX1 U1448 ( .A(n1841), .Y(n2934) );
  AND2X1 U1450 ( .A(n1660), .B(n1847), .Y(n1851) );
  INVX1 U1452 ( .A(n1851), .Y(n2935) );
  AND2X1 U1454 ( .A(n1643), .B(n1847), .Y(n1859) );
  INVX1 U1457 ( .A(n1859), .Y(n2936) );
  AND2X1 U1459 ( .A(n1656), .B(n1864), .Y(n1866) );
  INVX1 U1461 ( .A(n1866), .Y(n2937) );
  AND2X1 U1463 ( .A(n1637), .B(n1881), .Y(n1890) );
  INVX1 U1465 ( .A(n1890), .Y(n2938) );
  AND2X1 U1467 ( .A(n1660), .B(n1898), .Y(n1902) );
  INVX1 U1469 ( .A(n1902), .Y(n2939) );
  AND2X1 U1471 ( .A(n1639), .B(n1898), .Y(n1908) );
  INVX1 U1473 ( .A(n1908), .Y(n2940) );
  AND2X1 U1475 ( .A(n1629), .B(n1915), .Y(n1920) );
  INVX1 U1477 ( .A(n1920), .Y(n2941) );
  AND2X1 U1479 ( .A(n1641), .B(n1915), .Y(n1926) );
  INVX1 U1481 ( .A(n1926), .Y(n2942) );
  AND2X1 U1483 ( .A(n1631), .B(n1932), .Y(n1938) );
  INVX1 U1485 ( .A(n1938), .Y(n2943) );
  AND2X1 U1487 ( .A(n1643), .B(n1932), .Y(n1944) );
  INVX1 U1490 ( .A(n1944), .Y(n2944) );
  AND2X1 U1492 ( .A(n1654), .B(n1967), .Y(n1968) );
  INVX1 U1494 ( .A(n1968), .Y(n2945) );
  AND2X1 U1496 ( .A(n1633), .B(n1984), .Y(n1991) );
  INVX1 U1498 ( .A(n1991), .Y(n2946) );
  AND2X1 U1500 ( .A(n1635), .B(n2001), .Y(n2009) );
  INVX1 U1502 ( .A(n2009), .Y(n2947) );
  AND2X1 U1504 ( .A(n1656), .B(n2018), .Y(n2020) );
  INVX1 U1506 ( .A(n2020), .Y(n2948) );
  AND2X1 U1508 ( .A(n1654), .B(n2104), .Y(n2105) );
  INVX1 U1510 ( .A(n2105), .Y(n2949) );
  AND2X1 U1512 ( .A(n1633), .B(n2121), .Y(n2128) );
  INVX1 U1514 ( .A(n2128), .Y(n2950) );
  AND2X1 U1516 ( .A(n1635), .B(n2138), .Y(n2146) );
  INVX1 U1518 ( .A(n2146), .Y(n2951) );
  AND2X1 U1520 ( .A(n1656), .B(n1627), .Y(n2224) );
  INVX1 U1523 ( .A(n2224), .Y(n2952) );
  AND2X1 U1525 ( .A(n1633), .B(n1652), .Y(n1663) );
  INVX1 U1527 ( .A(n1663), .Y(n2953) );
  AND2X1 U1529 ( .A(n1635), .B(n1675), .Y(n1683) );
  INVX1 U1531 ( .A(n1683), .Y(n2954) );
  AND2X1 U1533 ( .A(n1651), .B(n1794), .Y(n1810) );
  INVX1 U1535 ( .A(n1810), .Y(n2955) );
  AND2X1 U1537 ( .A(n1649), .B(n1812), .Y(n1827) );
  INVX1 U1539 ( .A(n1827), .Y(n2956) );
  AND2X1 U1541 ( .A(n1647), .B(n1830), .Y(n1844) );
  INVX1 U1543 ( .A(n1844), .Y(n2957) );
  AND2X1 U1545 ( .A(n1645), .B(n1847), .Y(n1860) );
  INVX1 U1547 ( .A(n1860), .Y(n2958) );
  AND2X1 U1549 ( .A(n1651), .B(n1881), .Y(n1897) );
  INVX1 U1551 ( .A(n1897), .Y(n2959) );
  AND2X1 U1553 ( .A(n1649), .B(n1898), .Y(n1913) );
  INVX1 U1556 ( .A(n1913), .Y(n2960) );
  AND2X1 U1558 ( .A(n1647), .B(n1915), .Y(n1929) );
  INVX1 U1560 ( .A(n1929), .Y(n2961) );
  AND2X1 U1562 ( .A(n1645), .B(n1932), .Y(n1945) );
  INVX1 U1564 ( .A(n1945), .Y(n2962) );
  AND2X1 U1566 ( .A(n1635), .B(n2018), .Y(n2026) );
  INVX1 U1568 ( .A(n2026), .Y(n2963) );
  AND2X1 U1570 ( .A(n1633), .B(n2035), .Y(n2042) );
  INVX1 U1572 ( .A(n2042), .Y(n2964) );
  AND2X1 U1574 ( .A(n1656), .B(n2052), .Y(n2054) );
  INVX1 U1576 ( .A(n2054), .Y(n2965) );
  AND2X1 U1578 ( .A(n1654), .B(n2069), .Y(n2070) );
  INVX1 U1580 ( .A(n2070), .Y(n2966) );
  AND2X1 U1582 ( .A(n1635), .B(n2155), .Y(n2163) );
  INVX1 U1584 ( .A(n2163), .Y(n2967) );
  AND2X1 U1586 ( .A(n1633), .B(n2172), .Y(n2179) );
  INVX1 U1589 ( .A(n2179), .Y(n2968) );
  AND2X1 U1591 ( .A(n1656), .B(n2189), .Y(n2191) );
  INVX1 U1593 ( .A(n2191), .Y(n2969) );
  AND2X1 U1595 ( .A(n1654), .B(n2206), .Y(n2207) );
  INVX1 U1597 ( .A(n2207), .Y(n2970) );
  AND2X1 U1599 ( .A(n1658), .B(n1627), .Y(n2225) );
  INVX1 U1601 ( .A(n2225), .Y(n2971) );
  AND2X1 U1603 ( .A(n1635), .B(n1693), .Y(n1701) );
  INVX1 U1605 ( .A(n1701), .Y(n2972) );
  AND2X1 U1607 ( .A(n1633), .B(n1711), .Y(n1718) );
  INVX1 U1609 ( .A(n1718), .Y(n2973) );
  AND2X1 U1611 ( .A(n1656), .B(n1729), .Y(n1731) );
  INVX1 U1613 ( .A(n1731), .Y(n2974) );
  AND2X1 U1615 ( .A(n1654), .B(n1747), .Y(n1748) );
  INVX1 U1617 ( .A(n1748), .Y(n2975) );
  AND2X1 U1619 ( .A(n1649), .B(n1794), .Y(n1809) );
  INVX1 U1622 ( .A(n1809), .Y(n2976) );
  AND2X1 U1624 ( .A(n1651), .B(n1812), .Y(n1828) );
  INVX1 U1626 ( .A(n1828), .Y(n2977) );
  AND2X1 U1628 ( .A(n1645), .B(n1830), .Y(n1843) );
  INVX1 U1630 ( .A(n1843), .Y(n2978) );
  AND2X1 U1632 ( .A(n1647), .B(n1847), .Y(n1861) );
  INVX1 U1634 ( .A(n1861), .Y(n2979) );
  AND2X1 U1636 ( .A(n1649), .B(n1881), .Y(n1896) );
  INVX1 U1638 ( .A(n1896), .Y(n2980) );
  AND2X1 U1640 ( .A(n1651), .B(n1898), .Y(n1914) );
  INVX1 U1642 ( .A(n1914), .Y(n2981) );
  AND2X1 U1644 ( .A(n1645), .B(n1915), .Y(n1928) );
  INVX1 U1646 ( .A(n1928), .Y(n2982) );
  AND2X1 U1648 ( .A(n1647), .B(n1932), .Y(n1946) );
  INVX1 U1650 ( .A(n1946), .Y(n2983) );
  AND2X1 U1652 ( .A(n1633), .B(n2018), .Y(n2025) );
  INVX1 U1656 ( .A(n2025), .Y(n2984) );
  AND2X1 U1658 ( .A(n1635), .B(n2035), .Y(n2043) );
  INVX1 U1660 ( .A(n2043), .Y(n2985) );
  AND2X1 U1662 ( .A(n1654), .B(n2052), .Y(n2053) );
  INVX1 U1664 ( .A(n2053), .Y(n2986) );
  AND2X1 U1666 ( .A(n1656), .B(n2069), .Y(n2071) );
  INVX1 U1668 ( .A(n2071), .Y(n2987) );
  AND2X1 U1670 ( .A(n1633), .B(n2155), .Y(n2162) );
  INVX1 U1672 ( .A(n2162), .Y(n2988) );
  AND2X1 U1674 ( .A(n1635), .B(n2172), .Y(n2180) );
  INVX1 U1676 ( .A(n2180), .Y(n2989) );
  AND2X1 U1678 ( .A(n1654), .B(n2189), .Y(n2190) );
  INVX1 U1680 ( .A(n2190), .Y(n2990) );
  AND2X1 U1682 ( .A(n1656), .B(n2206), .Y(n2208) );
  INVX1 U1684 ( .A(n2208), .Y(n2991) );
  AND2X1 U1686 ( .A(n1660), .B(n1627), .Y(n2226) );
  INVX1 U1689 ( .A(n2226), .Y(n2992) );
  AND2X1 U1691 ( .A(n1633), .B(n1693), .Y(n1700) );
  INVX1 U1693 ( .A(n1700), .Y(n2993) );
  AND2X1 U1695 ( .A(n1635), .B(n1711), .Y(n1719) );
  INVX1 U1697 ( .A(n1719), .Y(n2994) );
  AND2X1 U1699 ( .A(n1654), .B(n1729), .Y(n1730) );
  INVX1 U1701 ( .A(n1730), .Y(n2995) );
  AND2X1 U1703 ( .A(n1656), .B(n1747), .Y(n1749) );
  INVX1 U1705 ( .A(n1749), .Y(n2996) );
  AND2X1 U1707 ( .A(n1647), .B(n1794), .Y(n1808) );
  INVX1 U1709 ( .A(n1808), .Y(n2997) );
  AND2X1 U1711 ( .A(n1645), .B(n1812), .Y(n1825) );
  INVX1 U1713 ( .A(n1825), .Y(n2998) );
  AND2X1 U1715 ( .A(n1651), .B(n1830), .Y(n1846) );
  INVX1 U1717 ( .A(n1846), .Y(n2999) );
  AND2X1 U1719 ( .A(n1649), .B(n1847), .Y(n1862) );
  INVX1 U1722 ( .A(n1862), .Y(n3000) );
  AND2X1 U1724 ( .A(n1647), .B(n1881), .Y(n1895) );
  INVX1 U1726 ( .A(n1895), .Y(n3001) );
  AND2X1 U1728 ( .A(n1645), .B(n1898), .Y(n1911) );
  INVX1 U1730 ( .A(n1911), .Y(n3002) );
  AND2X1 U1732 ( .A(n1651), .B(n1915), .Y(n1931) );
  INVX1 U1734 ( .A(n1931), .Y(n3003) );
  AND2X1 U1736 ( .A(n1649), .B(n1932), .Y(n1947) );
  INVX1 U1738 ( .A(n1947), .Y(n3004) );
  AND2X1 U1740 ( .A(n1658), .B(n1950), .Y(n1953) );
  INVX1 U1742 ( .A(n1953), .Y(n3005) );
  AND2X1 U1744 ( .A(n1656), .B(n2035), .Y(n2037) );
  INVX1 U1746 ( .A(n2037), .Y(n3006) );
  AND2X1 U1748 ( .A(n1635), .B(n2052), .Y(n2060) );
  INVX1 U1750 ( .A(n2060), .Y(n3007) );
  AND2X1 U1752 ( .A(n1633), .B(n2069), .Y(n2076) );
  INVX1 U1755 ( .A(n2076), .Y(n3008) );
  AND2X1 U1757 ( .A(n1654), .B(n2087), .Y(n2088) );
  INVX1 U1759 ( .A(n2088), .Y(n3009) );
  AND2X1 U1761 ( .A(n1656), .B(n2155), .Y(n2157) );
  INVX1 U1763 ( .A(n2157), .Y(n3010) );
  AND2X1 U1765 ( .A(n1654), .B(n2172), .Y(n2173) );
  INVX1 U1767 ( .A(n2173), .Y(n3011) );
  AND2X1 U1769 ( .A(n1635), .B(n2189), .Y(n2197) );
  INVX1 U1771 ( .A(n2197), .Y(n3012) );
  AND2X1 U1773 ( .A(n1633), .B(n2206), .Y(n2213) );
  INVX1 U1775 ( .A(n2213), .Y(n3013) );
  AND2X1 U1777 ( .A(n1629), .B(n1627), .Y(n1628) );
  INVX1 U1779 ( .A(n1628), .Y(n3014) );
  AND2X1 U1781 ( .A(n1656), .B(n1693), .Y(n1695) );
  INVX1 U1783 ( .A(n1695), .Y(n3015) );
  AND2X1 U1785 ( .A(n1654), .B(n1711), .Y(n1712) );
  INVX1 U1788 ( .A(n1712), .Y(n3016) );
  AND2X1 U1790 ( .A(n1635), .B(n1729), .Y(n1737) );
  INVX1 U1792 ( .A(n1737), .Y(n3017) );
  AND2X1 U1794 ( .A(n1633), .B(n1747), .Y(n1754) );
  INVX1 U1796 ( .A(n1754), .Y(n3018) );
  AND2X1 U1798 ( .A(n1645), .B(n1794), .Y(n1807) );
  INVX1 U1800 ( .A(n1807), .Y(n3019) );
  AND2X1 U1802 ( .A(n1647), .B(n1812), .Y(n1826) );
  INVX1 U1804 ( .A(n1826), .Y(n3020) );
  AND2X1 U1806 ( .A(n1649), .B(n1830), .Y(n1845) );
  INVX1 U1808 ( .A(n1845), .Y(n3021) );
  AND2X1 U1810 ( .A(n1651), .B(n1847), .Y(n1863) );
  INVX1 U1812 ( .A(n1863), .Y(n3022) );
  AND2X1 U1814 ( .A(n1645), .B(n1881), .Y(n1894) );
  INVX1 U1816 ( .A(n1894), .Y(n3023) );
  AND2X1 U1818 ( .A(n1647), .B(n1898), .Y(n1912) );
  INVX1 U1821 ( .A(n1912), .Y(n3024) );
  AND2X1 U1823 ( .A(n1649), .B(n1915), .Y(n1930) );
  INVX1 U1825 ( .A(n1930), .Y(n3025) );
  AND2X1 U1827 ( .A(n1651), .B(n1932), .Y(n1948) );
  INVX1 U1829 ( .A(n1948), .Y(n3026) );
  AND2X1 U1831 ( .A(n1660), .B(n1950), .Y(n1954) );
  INVX1 U1833 ( .A(n1954), .Y(n3027) );
  AND2X1 U1835 ( .A(n1654), .B(n2035), .Y(n2036) );
  INVX1 U1837 ( .A(n2036), .Y(n3028) );
  AND2X1 U1839 ( .A(n1633), .B(n2052), .Y(n2059) );
  INVX1 U1841 ( .A(n2059), .Y(n3029) );
  AND2X1 U1843 ( .A(n1635), .B(n2069), .Y(n2077) );
  INVX1 U1845 ( .A(n2077), .Y(n3030) );
  AND2X1 U1847 ( .A(n1656), .B(n2087), .Y(n2089) );
  INVX1 U1849 ( .A(n2089), .Y(n3031) );
  AND2X1 U1851 ( .A(n1654), .B(n2155), .Y(n2156) );
  INVX1 U1854 ( .A(n2156), .Y(n3032) );
  AND2X1 U1856 ( .A(n1656), .B(n2172), .Y(n2174) );
  INVX1 U1858 ( .A(n2174), .Y(n3033) );
  AND2X1 U1860 ( .A(n1633), .B(n2189), .Y(n2196) );
  INVX1 U1862 ( .A(n2196), .Y(n3034) );
  AND2X1 U1864 ( .A(n1635), .B(n2206), .Y(n2214) );
  INVX1 U1866 ( .A(n2214), .Y(n3035) );
  AND2X1 U1868 ( .A(n1631), .B(n1627), .Y(n1630) );
  INVX1 U1870 ( .A(n1630), .Y(n3036) );
  AND2X1 U1872 ( .A(n1654), .B(n1693), .Y(n1694) );
  INVX1 U1874 ( .A(n1694), .Y(n3037) );
  AND2X1 U1876 ( .A(n1656), .B(n1711), .Y(n1713) );
  INVX1 U1878 ( .A(n1713), .Y(n3038) );
  AND2X1 U1880 ( .A(n1633), .B(n1729), .Y(n1736) );
  INVX1 U1882 ( .A(n1736), .Y(n3039) );
  AND2X1 U1884 ( .A(n1635), .B(n1747), .Y(n1755) );
  INVX1 U1887 ( .A(n1755), .Y(n3040) );
  BUFX2 U1889 ( .A(n1788), .Y(n3041) );
  AND2X1 U1891 ( .A(n1651), .B(n1864), .Y(n1880) );
  INVX1 U1893 ( .A(n1880), .Y(n3042) );
  AND2X1 U1895 ( .A(n1651), .B(n1950), .Y(n1966) );
  INVX1 U1897 ( .A(n1966), .Y(n3043) );
  AND2X1 U1899 ( .A(n1649), .B(n1967), .Y(n1982) );
  INVX1 U1901 ( .A(n1982), .Y(n3044) );
  AND2X1 U1903 ( .A(n1647), .B(n1984), .Y(n1998) );
  INVX1 U1905 ( .A(n1998), .Y(n3045) );
  AND2X1 U1907 ( .A(n1645), .B(n2001), .Y(n2014) );
  INVX1 U1909 ( .A(n2014), .Y(n3046) );
  AND2X1 U1911 ( .A(n1631), .B(n2018), .Y(n2024) );
  INVX1 U1913 ( .A(n2024), .Y(n3047) );
  AND2X1 U1915 ( .A(n1643), .B(n2018), .Y(n2030) );
  INVX1 U1917 ( .A(n2030), .Y(n3048) );
  AND2X1 U1921 ( .A(n1629), .B(n2035), .Y(n2040) );
  INVX1 U1923 ( .A(n2040), .Y(n3049) );
  AND2X1 U1925 ( .A(n1641), .B(n2035), .Y(n2046) );
  INVX1 U1927 ( .A(n2046), .Y(n3050) );
  AND2X1 U1929 ( .A(n1660), .B(n2052), .Y(n2056) );
  INVX1 U1931 ( .A(n2056), .Y(n3051) );
  AND2X1 U1933 ( .A(n1639), .B(n2052), .Y(n2062) );
  INVX1 U1935 ( .A(n2062), .Y(n3052) );
  AND2X1 U1937 ( .A(n1658), .B(n2069), .Y(n2072) );
  INVX1 U1939 ( .A(n2072), .Y(n3053) );
  AND2X1 U1941 ( .A(n1637), .B(n2069), .Y(n2078) );
  INVX1 U1943 ( .A(n2078), .Y(n3054) );
  AND2X1 U1945 ( .A(n1651), .B(n2087), .Y(n2103) );
  INVX1 U1947 ( .A(n2103), .Y(n3055) );
  AND2X1 U1949 ( .A(n1649), .B(n2104), .Y(n2119) );
  INVX1 U1951 ( .A(n2119), .Y(n3056) );
  AND2X1 U1954 ( .A(n1647), .B(n2121), .Y(n2135) );
  INVX1 U1956 ( .A(n2135), .Y(n3057) );
  AND2X1 U1958 ( .A(n1645), .B(n2138), .Y(n2151) );
  INVX1 U1960 ( .A(n2151), .Y(n3058) );
  AND2X1 U1962 ( .A(n1631), .B(n2155), .Y(n2161) );
  INVX1 U1964 ( .A(n2161), .Y(n3059) );
  AND2X1 U1966 ( .A(n1643), .B(n2155), .Y(n2167) );
  INVX1 U1968 ( .A(n2167), .Y(n3060) );
  AND2X1 U1970 ( .A(n1629), .B(n2172), .Y(n2177) );
  INVX1 U1972 ( .A(n2177), .Y(n3061) );
  AND2X1 U1974 ( .A(n1641), .B(n2172), .Y(n2183) );
  INVX1 U1976 ( .A(n2183), .Y(n3062) );
  AND2X1 U1978 ( .A(n1660), .B(n2189), .Y(n2193) );
  INVX1 U1980 ( .A(n2193), .Y(n3063) );
  AND2X1 U1982 ( .A(n1639), .B(n2189), .Y(n2199) );
  INVX1 U1984 ( .A(n2199), .Y(n3064) );
  AND2X1 U1987 ( .A(n1658), .B(n2206), .Y(n2209) );
  INVX1 U1989 ( .A(n2209), .Y(n3065) );
  AND2X1 U1991 ( .A(n1637), .B(n2206), .Y(n2215) );
  INVX1 U1993 ( .A(n2215), .Y(n3066) );
  AND2X1 U1995 ( .A(n1649), .B(n1627), .Y(n1648) );
  INVX1 U1997 ( .A(n1648), .Y(n3067) );
  AND2X1 U1999 ( .A(n1647), .B(n1652), .Y(n1670) );
  INVX1 U2001 ( .A(n1670), .Y(n3068) );
  AND2X1 U2003 ( .A(n1645), .B(n1675), .Y(n1688) );
  INVX1 U2005 ( .A(n1688), .Y(n3069) );
  AND2X1 U2007 ( .A(n1631), .B(n1693), .Y(n1699) );
  INVX1 U2009 ( .A(n1699), .Y(n3070) );
  AND2X1 U2011 ( .A(n1643), .B(n1693), .Y(n1705) );
  INVX1 U2013 ( .A(n1705), .Y(n3071) );
  AND2X1 U2015 ( .A(n1629), .B(n1711), .Y(n1716) );
  INVX1 U2017 ( .A(n1716), .Y(n3072) );
  AND2X1 U2021 ( .A(n1641), .B(n1711), .Y(n1722) );
  INVX1 U2023 ( .A(n1722), .Y(n3073) );
  AND2X1 U2025 ( .A(n1660), .B(n1729), .Y(n1733) );
  INVX1 U2027 ( .A(n1733), .Y(n3074) );
  AND2X1 U2029 ( .A(n1639), .B(n1729), .Y(n1739) );
  INVX1 U2031 ( .A(n1739), .Y(n3075) );
  AND2X1 U2033 ( .A(n1658), .B(n1747), .Y(n1750) );
  INVX1 U2035 ( .A(n1750), .Y(n3076) );
  AND2X1 U2037 ( .A(n1637), .B(n1747), .Y(n1756) );
  INVX1 U2039 ( .A(n1756), .Y(n3077) );
  BUFX2 U2041 ( .A(n1790), .Y(n3078) );
  AND2X1 U2043 ( .A(n1649), .B(n1864), .Y(n1879) );
  INVX1 U2045 ( .A(n1879), .Y(n3079) );
  AND2X1 U2047 ( .A(n1649), .B(n1950), .Y(n1965) );
  INVX1 U2049 ( .A(n1965), .Y(n3080) );
  AND2X1 U2051 ( .A(n1651), .B(n1967), .Y(n1983) );
  INVX1 U2055 ( .A(n1983), .Y(n3081) );
  AND2X1 U2057 ( .A(n1645), .B(n1984), .Y(n1997) );
  INVX1 U2059 ( .A(n1997), .Y(n3082) );
  AND2X1 U2061 ( .A(n1647), .B(n2001), .Y(n2015) );
  INVX1 U2063 ( .A(n2015), .Y(n3083) );
  AND2X1 U2065 ( .A(n1629), .B(n2018), .Y(n2023) );
  INVX1 U2067 ( .A(n2023), .Y(n3084) );
  AND2X1 U2069 ( .A(n1641), .B(n2018), .Y(n2029) );
  INVX1 U2071 ( .A(n2029), .Y(n3085) );
  AND2X1 U2073 ( .A(n1631), .B(n2035), .Y(n2041) );
  INVX1 U2075 ( .A(n2041), .Y(n3086) );
  AND2X1 U2077 ( .A(n1643), .B(n2035), .Y(n2047) );
  INVX1 U2079 ( .A(n2047), .Y(n3087) );
  AND2X1 U2081 ( .A(n1658), .B(n2052), .Y(n2055) );
  INVX1 U2083 ( .A(n2055), .Y(n3088) );
  AND2X1 U2085 ( .A(n1637), .B(n2052), .Y(n2061) );
  INVX1 U2089 ( .A(n2061), .Y(n3089) );
  AND2X1 U2091 ( .A(n1660), .B(n2069), .Y(n2073) );
  INVX1 U2093 ( .A(n2073), .Y(n3090) );
  AND2X1 U2095 ( .A(n1639), .B(n2069), .Y(n2079) );
  INVX1 U2097 ( .A(n2079), .Y(n3091) );
  AND2X1 U2099 ( .A(n1649), .B(n2087), .Y(n2102) );
  INVX1 U2101 ( .A(n2102), .Y(n3092) );
  AND2X1 U2103 ( .A(n1651), .B(n2104), .Y(n2120) );
  INVX1 U2105 ( .A(n2120), .Y(n3093) );
  AND2X1 U2107 ( .A(n1645), .B(n2121), .Y(n2134) );
  INVX1 U2109 ( .A(n2134), .Y(n3094) );
  AND2X1 U2111 ( .A(n1647), .B(n2138), .Y(n2152) );
  INVX1 U2113 ( .A(n2152), .Y(n3095) );
  AND2X1 U2115 ( .A(n1629), .B(n2155), .Y(n2160) );
  INVX1 U2117 ( .A(n2160), .Y(n3096) );
  AND2X1 U2119 ( .A(n1641), .B(n2155), .Y(n2166) );
  INVX1 U2123 ( .A(n2166), .Y(n3097) );
  AND2X1 U2125 ( .A(n1631), .B(n2172), .Y(n2178) );
  INVX1 U2127 ( .A(n2178), .Y(n3098) );
  AND2X1 U2129 ( .A(n1643), .B(n2172), .Y(n2184) );
  INVX1 U2131 ( .A(n2184), .Y(n3099) );
  AND2X1 U2133 ( .A(n1658), .B(n2189), .Y(n2192) );
  INVX1 U2135 ( .A(n2192), .Y(n3100) );
  AND2X1 U2137 ( .A(n1637), .B(n2189), .Y(n2198) );
  INVX1 U2139 ( .A(n2198), .Y(n3101) );
  AND2X1 U2141 ( .A(n1660), .B(n2206), .Y(n2210) );
  INVX1 U2143 ( .A(n2210), .Y(n3102) );
  AND2X1 U2145 ( .A(n1639), .B(n2206), .Y(n2216) );
  INVX1 U2147 ( .A(n2216), .Y(n3103) );
  AND2X1 U2149 ( .A(n1651), .B(n1627), .Y(n1650) );
  INVX1 U2151 ( .A(n1650), .Y(n3104) );
  AND2X1 U2153 ( .A(n1645), .B(n1652), .Y(n1669) );
  INVX1 U2157 ( .A(n1669), .Y(n3105) );
  AND2X1 U2159 ( .A(n1647), .B(n1675), .Y(n1689) );
  INVX1 U2161 ( .A(n1689), .Y(n3106) );
  AND2X1 U2163 ( .A(n1629), .B(n1693), .Y(n1698) );
  INVX1 U2165 ( .A(n1698), .Y(n3107) );
  AND2X1 U2167 ( .A(n1641), .B(n1693), .Y(n1704) );
  INVX1 U2169 ( .A(n1704), .Y(n3108) );
  AND2X1 U2171 ( .A(n1631), .B(n1711), .Y(n1717) );
  INVX1 U2173 ( .A(n1717), .Y(n3109) );
  AND2X1 U2175 ( .A(n1643), .B(n1711), .Y(n1723) );
  INVX1 U2177 ( .A(n1723), .Y(n3110) );
  AND2X1 U2179 ( .A(n1658), .B(n1729), .Y(n1732) );
  INVX1 U2181 ( .A(n1732), .Y(n3111) );
  AND2X1 U2183 ( .A(n1637), .B(n1729), .Y(n1738) );
  INVX1 U2185 ( .A(n1738), .Y(n3112) );
  AND2X1 U2187 ( .A(n1660), .B(n1747), .Y(n1751) );
  INVX1 U2192 ( .A(n1751), .Y(n3113) );
  AND2X1 U2194 ( .A(n1639), .B(n1747), .Y(n1757) );
  INVX1 U2196 ( .A(n1757), .Y(n3114) );
  BUFX2 U2198 ( .A(n2229), .Y(n3115) );
  BUFX2 U2200 ( .A(n2232), .Y(n3116) );
  AND2X1 U2202 ( .A(n1656), .B(n1847), .Y(n1849) );
  INVX1 U2204 ( .A(n1849), .Y(n3117) );
  AND2X1 U2206 ( .A(n1647), .B(n1864), .Y(n1878) );
  INVX1 U2208 ( .A(n1878), .Y(n3118) );
  AND2X1 U2210 ( .A(n1654), .B(n1881), .Y(n1882) );
  INVX1 U2212 ( .A(n1882), .Y(n3119) );
  AND2X1 U2214 ( .A(n1647), .B(n1950), .Y(n1964) );
  INVX1 U2216 ( .A(n1964), .Y(n3120) );
  AND2X1 U2218 ( .A(n1645), .B(n1967), .Y(n1980) );
  INVX1 U2220 ( .A(n1980), .Y(n3121) );
  AND2X1 U2222 ( .A(n1651), .B(n1984), .Y(n2000) );
  INVX1 U2226 ( .A(n2000), .Y(n3122) );
  AND2X1 U2228 ( .A(n1649), .B(n2001), .Y(n2016) );
  INVX1 U2230 ( .A(n2016), .Y(n3123) );
  AND2X1 U2232 ( .A(n1660), .B(n2018), .Y(n2022) );
  INVX1 U2251 ( .A(n2022), .Y(n3124) );
  AND2X1 U2252 ( .A(n1639), .B(n2018), .Y(n2028) );
  INVX1 U2253 ( .A(n2028), .Y(n3125) );
  AND2X1 U2254 ( .A(n1658), .B(n2035), .Y(n2038) );
  INVX1 U2255 ( .A(n2038), .Y(n3126) );
  AND2X1 U2256 ( .A(n1637), .B(n2035), .Y(n2044) );
  INVX1 U2257 ( .A(n2044), .Y(n3127) );
  AND2X1 U2258 ( .A(n1631), .B(n2052), .Y(n2058) );
  INVX1 U2259 ( .A(n2058), .Y(n3128) );
  AND2X1 U2260 ( .A(n1643), .B(n2052), .Y(n2064) );
  INVX1 U2261 ( .A(n2064), .Y(n3129) );
  AND2X1 U2262 ( .A(n1629), .B(n2069), .Y(n2074) );
  INVX1 U2263 ( .A(n2074), .Y(n3130) );
  AND2X1 U2264 ( .A(n1641), .B(n2069), .Y(n2080) );
  INVX1 U2265 ( .A(n2080), .Y(n3131) );
  AND2X1 U2266 ( .A(n1647), .B(n2087), .Y(n2101) );
  INVX1 U2267 ( .A(n2101), .Y(n3132) );
  AND2X1 U2268 ( .A(n1645), .B(n2104), .Y(n2117) );
  INVX1 U2269 ( .A(n2117), .Y(n3133) );
  AND2X1 U2270 ( .A(n1651), .B(n2121), .Y(n2137) );
  INVX1 U2271 ( .A(n2137), .Y(n3134) );
  AND2X1 U2272 ( .A(n1649), .B(n2138), .Y(n2153) );
  INVX1 U2273 ( .A(n2153), .Y(n3135) );
  AND2X1 U2274 ( .A(n1660), .B(n2155), .Y(n2159) );
  INVX1 U2275 ( .A(n2159), .Y(n3136) );
  AND2X1 U2276 ( .A(n1639), .B(n2155), .Y(n2165) );
  INVX1 U2277 ( .A(n2165), .Y(n3137) );
  AND2X1 U2278 ( .A(n1658), .B(n2172), .Y(n2175) );
  INVX1 U2279 ( .A(n2175), .Y(n3138) );
  AND2X1 U2280 ( .A(n1637), .B(n2172), .Y(n2181) );
  INVX1 U2281 ( .A(n2181), .Y(n3139) );
  AND2X1 U2282 ( .A(n1631), .B(n2189), .Y(n2195) );
  INVX1 U2283 ( .A(n2195), .Y(n3140) );
  AND2X1 U2284 ( .A(n1643), .B(n2189), .Y(n2201) );
  INVX1 U2285 ( .A(n2201), .Y(n3141) );
  AND2X1 U2286 ( .A(n1629), .B(n2206), .Y(n2211) );
  INVX1 U2287 ( .A(n2211), .Y(n3142) );
  AND2X1 U2288 ( .A(n1641), .B(n2206), .Y(n2217) );
  INVX1 U2289 ( .A(n2217), .Y(n3143) );
  AND2X1 U2290 ( .A(n1633), .B(n1627), .Y(n1632) );
  INVX1 U2291 ( .A(n1632), .Y(n3144) );
  AND2X1 U2292 ( .A(n1645), .B(n1627), .Y(n1644) );
  INVX1 U2293 ( .A(n1644), .Y(n3145) );
  AND2X1 U2294 ( .A(n1651), .B(n1652), .Y(n1672) );
  INVX1 U2295 ( .A(n1672), .Y(n3146) );
  AND2X1 U2296 ( .A(n1649), .B(n1675), .Y(n1690) );
  INVX1 U2297 ( .A(n1690), .Y(n3147) );
  AND2X1 U2298 ( .A(n1660), .B(n1693), .Y(n1697) );
  INVX1 U2299 ( .A(n1697), .Y(n3148) );
  AND2X1 U2300 ( .A(n1639), .B(n1693), .Y(n1703) );
  INVX1 U2301 ( .A(n1703), .Y(n3149) );
  AND2X1 U2302 ( .A(n1658), .B(n1711), .Y(n1714) );
  INVX1 U2303 ( .A(n1714), .Y(n3150) );
  AND2X1 U2304 ( .A(n1637), .B(n1711), .Y(n1720) );
  INVX1 U2305 ( .A(n1720), .Y(n3151) );
  AND2X1 U2306 ( .A(n1631), .B(n1729), .Y(n1735) );
  INVX1 U2307 ( .A(n1735), .Y(n3152) );
  AND2X1 U2308 ( .A(n1643), .B(n1729), .Y(n1741) );
  INVX1 U2309 ( .A(n1741), .Y(n3153) );
  AND2X1 U2310 ( .A(n1629), .B(n1747), .Y(n1752) );
  INVX1 U2311 ( .A(n1752), .Y(n3154) );
  AND2X1 U2312 ( .A(n1641), .B(n1747), .Y(n1758) );
  INVX1 U2313 ( .A(n1758), .Y(n3155) );
  BUFX2 U2314 ( .A(n1792), .Y(n3156) );
  BUFX2 U2315 ( .A(n1674), .Y(n3157) );
  BUFX2 U2316 ( .A(n1728), .Y(n3158) );
  AND2X1 U2317 ( .A(n1654), .B(n1847), .Y(n1848) );
  INVX1 U2318 ( .A(n1848), .Y(n3159) );
  AND2X1 U2319 ( .A(n1645), .B(n1864), .Y(n1877) );
  INVX1 U2320 ( .A(n1877), .Y(n3160) );
  AND2X1 U2321 ( .A(n1656), .B(n1881), .Y(n1883) );
  INVX1 U2322 ( .A(n1883), .Y(n3161) );
  AND2X1 U2323 ( .A(n1645), .B(n1950), .Y(n1963) );
  INVX1 U2324 ( .A(n1963), .Y(n3162) );
  AND2X1 U2325 ( .A(n1647), .B(n1967), .Y(n1981) );
  INVX1 U2326 ( .A(n1981), .Y(n3163) );
  AND2X1 U2327 ( .A(n1649), .B(n1984), .Y(n1999) );
  INVX1 U2328 ( .A(n1999), .Y(n3164) );
  AND2X1 U2329 ( .A(n1651), .B(n2001), .Y(n2017) );
  INVX1 U2330 ( .A(n2017), .Y(n3165) );
  AND2X1 U2331 ( .A(n1658), .B(n2018), .Y(n2021) );
  INVX1 U2332 ( .A(n2021), .Y(n3166) );
  AND2X1 U2333 ( .A(n1637), .B(n2018), .Y(n2027) );
  INVX1 U2334 ( .A(n2027), .Y(n3167) );
  AND2X1 U2335 ( .A(n1660), .B(n2035), .Y(n2039) );
  INVX1 U2336 ( .A(n2039), .Y(n3168) );
  AND2X1 U2337 ( .A(n1639), .B(n2035), .Y(n2045) );
  INVX1 U2338 ( .A(n2045), .Y(n3169) );
  AND2X1 U2339 ( .A(n1629), .B(n2052), .Y(n2057) );
  INVX1 U2340 ( .A(n2057), .Y(n3170) );
  AND2X1 U2341 ( .A(n1641), .B(n2052), .Y(n2063) );
  INVX1 U2342 ( .A(n2063), .Y(n3171) );
  AND2X1 U2343 ( .A(n1631), .B(n2069), .Y(n2075) );
  INVX1 U2344 ( .A(n2075), .Y(n3172) );
  AND2X1 U2345 ( .A(n1643), .B(n2069), .Y(n2081) );
  INVX1 U2346 ( .A(n2081), .Y(n3173) );
  AND2X1 U2347 ( .A(n1645), .B(n2087), .Y(n2100) );
  INVX1 U2348 ( .A(n2100), .Y(n3174) );
  AND2X1 U2349 ( .A(n1647), .B(n2104), .Y(n2118) );
  INVX1 U2350 ( .A(n2118), .Y(n3175) );
  AND2X1 U2351 ( .A(n1649), .B(n2121), .Y(n2136) );
  INVX1 U2352 ( .A(n2136), .Y(n3176) );
  AND2X1 U2353 ( .A(n1651), .B(n2138), .Y(n2154) );
  INVX1 U2354 ( .A(n2154), .Y(n3177) );
  AND2X1 U2355 ( .A(n1658), .B(n2155), .Y(n2158) );
  INVX1 U2356 ( .A(n2158), .Y(n3178) );
  AND2X1 U2357 ( .A(n1637), .B(n2155), .Y(n2164) );
  INVX1 U2358 ( .A(n2164), .Y(n3179) );
  AND2X1 U2359 ( .A(n1660), .B(n2172), .Y(n2176) );
  INVX1 U2360 ( .A(n2176), .Y(n3180) );
  AND2X1 U2361 ( .A(n1639), .B(n2172), .Y(n2182) );
  INVX1 U2362 ( .A(n2182), .Y(n3181) );
  AND2X1 U2363 ( .A(n1629), .B(n2189), .Y(n2194) );
  INVX1 U2364 ( .A(n2194), .Y(n3182) );
  AND2X1 U2365 ( .A(n1641), .B(n2189), .Y(n2200) );
  INVX1 U2366 ( .A(n2200), .Y(n3183) );
  AND2X1 U2367 ( .A(n1631), .B(n2206), .Y(n2212) );
  INVX1 U2368 ( .A(n2212), .Y(n3184) );
  AND2X1 U2369 ( .A(n1643), .B(n2206), .Y(n2218) );
  INVX1 U2370 ( .A(n2218), .Y(n3185) );
  AND2X1 U2371 ( .A(n1635), .B(n1627), .Y(n1634) );
  INVX1 U2372 ( .A(n1634), .Y(n3186) );
  AND2X1 U2373 ( .A(n1647), .B(n1627), .Y(n1646) );
  INVX1 U2374 ( .A(n1646), .Y(n3187) );
  AND2X1 U2375 ( .A(n1649), .B(n1652), .Y(n1671) );
  INVX1 U2376 ( .A(n1671), .Y(n3188) );
  AND2X1 U2377 ( .A(n1651), .B(n1675), .Y(n1691) );
  INVX1 U2378 ( .A(n1691), .Y(n3189) );
  AND2X1 U2379 ( .A(n1658), .B(n1693), .Y(n1696) );
  INVX1 U2380 ( .A(n1696), .Y(n3190) );
  AND2X1 U2381 ( .A(n1637), .B(n1693), .Y(n1702) );
  INVX1 U2382 ( .A(n1702), .Y(n3191) );
  AND2X1 U2383 ( .A(n1660), .B(n1711), .Y(n1715) );
  INVX1 U2384 ( .A(n1715), .Y(n3192) );
  AND2X1 U2385 ( .A(n1639), .B(n1711), .Y(n1721) );
  INVX1 U2386 ( .A(n1721), .Y(n3193) );
  AND2X1 U2387 ( .A(n1629), .B(n1729), .Y(n1734) );
  INVX1 U2388 ( .A(n1734), .Y(n3194) );
  AND2X1 U2389 ( .A(n1641), .B(n1729), .Y(n1740) );
  INVX1 U2390 ( .A(n1740), .Y(n3195) );
  AND2X1 U2391 ( .A(n1631), .B(n1747), .Y(n1753) );
  INVX1 U2392 ( .A(n1753), .Y(n3196) );
  AND2X1 U2393 ( .A(n1643), .B(n1747), .Y(n1759) );
  INVX1 U2394 ( .A(n1759), .Y(n3197) );
  AND2X1 U2395 ( .A(n1777), .B(n3399), .Y(n1771) );
  INVX1 U2396 ( .A(n1771), .Y(n3198) );
  BUFX2 U2397 ( .A(n1785), .Y(n3199) );
  BUFX2 U2398 ( .A(n1784), .Y(n3200) );
  OR2X1 U2399 ( .A(n3433), .B(wr_ptr[4]), .Y(n1786) );
  INVX1 U2400 ( .A(n1786), .Y(n3201) );
  BUFX2 U2401 ( .A(n1829), .Y(n3202) );
  BUFX2 U2402 ( .A(n1746), .Y(n3203) );
  AND2X1 U2403 ( .A(n1635), .B(n1794), .Y(n1802) );
  INVX1 U2404 ( .A(n1802), .Y(n3204) );
  AND2X1 U2405 ( .A(n1633), .B(n1812), .Y(n1819) );
  INVX1 U2406 ( .A(n1819), .Y(n3205) );
  AND2X1 U2407 ( .A(n1654), .B(n1830), .Y(n1831) );
  INVX1 U2408 ( .A(n1831), .Y(n3206) );
  AND2X1 U2409 ( .A(n1631), .B(n1847), .Y(n1853) );
  INVX1 U2410 ( .A(n1853), .Y(n3207) );
  AND2X1 U2411 ( .A(n1629), .B(n1864), .Y(n1869) );
  INVX1 U2412 ( .A(n1869), .Y(n3208) );
  AND2X1 U2413 ( .A(n1643), .B(n1864), .Y(n1876) );
  INVX1 U2414 ( .A(n1876), .Y(n3209) );
  AND2X1 U2415 ( .A(n1635), .B(n1881), .Y(n1889) );
  INVX1 U2416 ( .A(n1889), .Y(n3210) );
  AND2X1 U2417 ( .A(n1633), .B(n1898), .Y(n1905) );
  INVX1 U2418 ( .A(n1905), .Y(n3211) );
  AND2X1 U2419 ( .A(n1656), .B(n1915), .Y(n1917) );
  INVX1 U2420 ( .A(n1917), .Y(n3212) );
  AND2X1 U2421 ( .A(n1654), .B(n1932), .Y(n1933) );
  INVX1 U2422 ( .A(n1933), .Y(n3213) );
  AND2X1 U2423 ( .A(n1631), .B(n1950), .Y(n1956) );
  INVX1 U2424 ( .A(n1956), .Y(n3214) );
  AND2X1 U2425 ( .A(n1643), .B(n1950), .Y(n1962) );
  INVX1 U2426 ( .A(n1962), .Y(n3215) );
  AND2X1 U2427 ( .A(n1629), .B(n1967), .Y(n1972) );
  INVX1 U2428 ( .A(n1972), .Y(n3216) );
  AND2X1 U2429 ( .A(n1641), .B(n1967), .Y(n1978) );
  INVX1 U2430 ( .A(n1978), .Y(n3217) );
  AND2X1 U2431 ( .A(n1660), .B(n1984), .Y(n1988) );
  INVX1 U2432 ( .A(n1988), .Y(n3218) );
  AND2X1 U2433 ( .A(n1639), .B(n1984), .Y(n1994) );
  INVX1 U2434 ( .A(n1994), .Y(n3219) );
  AND2X1 U2435 ( .A(n1658), .B(n2001), .Y(n2004) );
  INVX1 U2436 ( .A(n2004), .Y(n3220) );
  AND2X1 U2437 ( .A(n1637), .B(n2001), .Y(n2010) );
  INVX1 U2438 ( .A(n2010), .Y(n3221) );
  AND2X1 U2439 ( .A(n1651), .B(n2018), .Y(n2034) );
  INVX1 U2440 ( .A(n2034), .Y(n3222) );
  AND2X1 U2441 ( .A(n1649), .B(n2035), .Y(n2050) );
  INVX1 U2442 ( .A(n2050), .Y(n3223) );
  AND2X1 U2443 ( .A(n1647), .B(n2052), .Y(n2066) );
  INVX1 U2444 ( .A(n2066), .Y(n3224) );
  AND2X1 U2445 ( .A(n1645), .B(n2069), .Y(n2082) );
  INVX1 U2446 ( .A(n2082), .Y(n3225) );
  AND2X1 U2447 ( .A(n1631), .B(n2087), .Y(n2093) );
  INVX1 U2448 ( .A(n2093), .Y(n3226) );
  AND2X1 U2449 ( .A(n1643), .B(n2087), .Y(n2099) );
  INVX1 U2450 ( .A(n2099), .Y(n3227) );
  AND2X1 U2451 ( .A(n1629), .B(n2104), .Y(n2109) );
  INVX1 U2452 ( .A(n2109), .Y(n3228) );
  AND2X1 U2453 ( .A(n1641), .B(n2104), .Y(n2115) );
  INVX1 U2454 ( .A(n2115), .Y(n3229) );
  AND2X1 U2455 ( .A(n1660), .B(n2121), .Y(n2125) );
  INVX1 U2456 ( .A(n2125), .Y(n3230) );
  AND2X1 U2457 ( .A(n1639), .B(n2121), .Y(n2131) );
  INVX1 U2458 ( .A(n2131), .Y(n3231) );
  AND2X1 U2459 ( .A(n1658), .B(n2138), .Y(n2141) );
  INVX1 U2460 ( .A(n2141), .Y(n3232) );
  AND2X1 U2461 ( .A(n1637), .B(n2138), .Y(n2147) );
  INVX1 U2462 ( .A(n2147), .Y(n3233) );
  AND2X1 U2463 ( .A(n1651), .B(n2155), .Y(n2171) );
  INVX1 U2464 ( .A(n2171), .Y(n3234) );
  AND2X1 U2465 ( .A(n1649), .B(n2172), .Y(n2187) );
  INVX1 U2466 ( .A(n2187), .Y(n3235) );
  AND2X1 U2467 ( .A(n1647), .B(n2189), .Y(n2203) );
  INVX1 U2468 ( .A(n2203), .Y(n3236) );
  AND2X1 U2469 ( .A(n1645), .B(n2206), .Y(n2219) );
  INVX1 U2470 ( .A(n2219), .Y(n3237) );
  AND2X1 U2471 ( .A(n1641), .B(n1627), .Y(n1640) );
  INVX1 U2472 ( .A(n1640), .Y(n3238) );
  AND2X1 U2473 ( .A(n1660), .B(n1652), .Y(n1659) );
  INVX1 U2474 ( .A(n1659), .Y(n3239) );
  AND2X1 U2475 ( .A(n1639), .B(n1652), .Y(n1666) );
  INVX1 U2476 ( .A(n1666), .Y(n3240) );
  AND2X1 U2477 ( .A(n1658), .B(n1675), .Y(n1678) );
  INVX1 U2478 ( .A(n1678), .Y(n3241) );
  AND2X1 U2479 ( .A(n1637), .B(n1675), .Y(n1684) );
  INVX1 U2480 ( .A(n1684), .Y(n3242) );
  AND2X1 U2481 ( .A(n1651), .B(n1693), .Y(n1709) );
  INVX1 U2482 ( .A(n1709), .Y(n3243) );
  AND2X1 U2483 ( .A(n1649), .B(n1711), .Y(n1726) );
  INVX1 U2484 ( .A(n1726), .Y(n3244) );
  AND2X1 U2485 ( .A(n1647), .B(n1729), .Y(n1743) );
  INVX1 U2486 ( .A(n1743), .Y(n3245) );
  AND2X1 U2487 ( .A(n1645), .B(n1747), .Y(n1760) );
  INVX1 U2488 ( .A(n1760), .Y(n3246) );
  INVX1 U2489 ( .A(n1777), .Y(n3247) );
  AND2X1 U2490 ( .A(get), .B(empty_bar), .Y(n1778) );
  INVX1 U2491 ( .A(n1778), .Y(n3248) );
  BUFX2 U2492 ( .A(n1764), .Y(n3249) );
  BUFX2 U2493 ( .A(n1793), .Y(n3250) );
  AND2X1 U2494 ( .A(n1633), .B(n1794), .Y(n1801) );
  INVX1 U2495 ( .A(n1801), .Y(n3251) );
  AND2X1 U2496 ( .A(n1635), .B(n1812), .Y(n1820) );
  INVX1 U2497 ( .A(n1820), .Y(n3252) );
  AND2X1 U2498 ( .A(n1656), .B(n1830), .Y(n1832) );
  INVX1 U2499 ( .A(n1832), .Y(n3253) );
  AND2X1 U2500 ( .A(n1629), .B(n1847), .Y(n1852) );
  INVX1 U2501 ( .A(n1852), .Y(n3254) );
  AND2X1 U2502 ( .A(n1631), .B(n1864), .Y(n1870) );
  INVX1 U2503 ( .A(n1870), .Y(n3255) );
  AND2X1 U2504 ( .A(n1641), .B(n1864), .Y(n1875) );
  INVX1 U2505 ( .A(n1875), .Y(n3256) );
  AND2X1 U2506 ( .A(n1633), .B(n1881), .Y(n1888) );
  INVX1 U2507 ( .A(n1888), .Y(n3257) );
  AND2X1 U2508 ( .A(n1635), .B(n1898), .Y(n1906) );
  INVX1 U2509 ( .A(n1906), .Y(n3258) );
  AND2X1 U2510 ( .A(n1654), .B(n1915), .Y(n1916) );
  INVX1 U2511 ( .A(n1916), .Y(n3259) );
  AND2X1 U2512 ( .A(n1656), .B(n1932), .Y(n1934) );
  INVX1 U2513 ( .A(n1934), .Y(n3260) );
  AND2X1 U2514 ( .A(n1629), .B(n1950), .Y(n1955) );
  INVX1 U2515 ( .A(n1955), .Y(n3261) );
  AND2X1 U2516 ( .A(n1641), .B(n1950), .Y(n1961) );
  INVX1 U2517 ( .A(n1961), .Y(n3262) );
  AND2X1 U2518 ( .A(n1631), .B(n1967), .Y(n1973) );
  INVX1 U2519 ( .A(n1973), .Y(n3263) );
  AND2X1 U2520 ( .A(n1643), .B(n1967), .Y(n1979) );
  INVX1 U2521 ( .A(n1979), .Y(n3264) );
  AND2X1 U2522 ( .A(n1658), .B(n1984), .Y(n1987) );
  INVX1 U2523 ( .A(n1987), .Y(n3265) );
  AND2X1 U2524 ( .A(n1637), .B(n1984), .Y(n1993) );
  INVX1 U2525 ( .A(n1993), .Y(n3266) );
  AND2X1 U2526 ( .A(n1660), .B(n2001), .Y(n2005) );
  INVX1 U2527 ( .A(n2005), .Y(n3267) );
  AND2X1 U2528 ( .A(n1639), .B(n2001), .Y(n2011) );
  INVX1 U2529 ( .A(n2011), .Y(n3268) );
  AND2X1 U2530 ( .A(n1649), .B(n2018), .Y(n2033) );
  INVX1 U2531 ( .A(n2033), .Y(n3269) );
  AND2X1 U2532 ( .A(n1651), .B(n2035), .Y(n2051) );
  INVX1 U2533 ( .A(n2051), .Y(n3270) );
  AND2X1 U2534 ( .A(n1645), .B(n2052), .Y(n2065) );
  INVX1 U2535 ( .A(n2065), .Y(n3271) );
  AND2X1 U2536 ( .A(n1647), .B(n2069), .Y(n2083) );
  INVX1 U2537 ( .A(n2083), .Y(n3272) );
  AND2X1 U2538 ( .A(n1629), .B(n2087), .Y(n2092) );
  INVX1 U2539 ( .A(n2092), .Y(n3273) );
  AND2X1 U2540 ( .A(n1641), .B(n2087), .Y(n2098) );
  INVX1 U2541 ( .A(n2098), .Y(n3274) );
  AND2X1 U2542 ( .A(n1631), .B(n2104), .Y(n2110) );
  INVX1 U2543 ( .A(n2110), .Y(n3275) );
  AND2X1 U2544 ( .A(n1643), .B(n2104), .Y(n2116) );
  INVX1 U2545 ( .A(n2116), .Y(n3276) );
  AND2X1 U2546 ( .A(n1658), .B(n2121), .Y(n2124) );
  INVX1 U2547 ( .A(n2124), .Y(n3277) );
  AND2X1 U2548 ( .A(n1637), .B(n2121), .Y(n2130) );
  INVX1 U2549 ( .A(n2130), .Y(n3278) );
  AND2X1 U2550 ( .A(n1660), .B(n2138), .Y(n2142) );
  INVX1 U2551 ( .A(n2142), .Y(n3279) );
  AND2X1 U2552 ( .A(n1639), .B(n2138), .Y(n2148) );
  INVX1 U2553 ( .A(n2148), .Y(n3280) );
  AND2X1 U2554 ( .A(n1649), .B(n2155), .Y(n2170) );
  INVX1 U2555 ( .A(n2170), .Y(n3281) );
  AND2X1 U2556 ( .A(n1651), .B(n2172), .Y(n2188) );
  INVX1 U2557 ( .A(n2188), .Y(n3282) );
  AND2X1 U2558 ( .A(n1645), .B(n2189), .Y(n2202) );
  INVX1 U2559 ( .A(n2202), .Y(n3283) );
  AND2X1 U2560 ( .A(n1647), .B(n2206), .Y(n2220) );
  INVX1 U2561 ( .A(n2220), .Y(n3284) );
  AND2X1 U2562 ( .A(n1643), .B(n1627), .Y(n1642) );
  INVX1 U2563 ( .A(n1642), .Y(n3285) );
  AND2X1 U2564 ( .A(n1658), .B(n1652), .Y(n1657) );
  INVX1 U2565 ( .A(n1657), .Y(n3286) );
  AND2X1 U2566 ( .A(n1637), .B(n1652), .Y(n1665) );
  INVX1 U2567 ( .A(n1665), .Y(n3287) );
  AND2X1 U2568 ( .A(n1660), .B(n1675), .Y(n1679) );
  INVX1 U2569 ( .A(n1679), .Y(n3288) );
  AND2X1 U2570 ( .A(n1639), .B(n1675), .Y(n1685) );
  INVX1 U2571 ( .A(n1685), .Y(n3289) );
  AND2X1 U2572 ( .A(n1649), .B(n1693), .Y(n1708) );
  INVX1 U2573 ( .A(n1708), .Y(n3290) );
  AND2X1 U2574 ( .A(n1651), .B(n1711), .Y(n1727) );
  INVX1 U2575 ( .A(n1727), .Y(n3291) );
  AND2X1 U2576 ( .A(n1645), .B(n1729), .Y(n1742) );
  INVX1 U2577 ( .A(n1742), .Y(n3292) );
  AND2X1 U2578 ( .A(n1647), .B(n1747), .Y(n1761) );
  INVX1 U2579 ( .A(n1761), .Y(n3293) );
  BUFX2 U2580 ( .A(n2314), .Y(empty_bar) );
  BUFX2 U2581 ( .A(n1772), .Y(n3295) );
  BUFX2 U2582 ( .A(n1625), .Y(n3296) );
  BUFX2 U2583 ( .A(n2228), .Y(n3297) );
  AND2X1 U2584 ( .A(n3415), .B(n3946), .Y(n1767) );
  INVX1 U2585 ( .A(n1767), .Y(n3298) );
  BUFX2 U2586 ( .A(n1692), .Y(n3299) );
  BUFX2 U2587 ( .A(n1710), .Y(n3300) );
  AND2X1 U2588 ( .A(n1656), .B(n1794), .Y(n1796) );
  INVX1 U2589 ( .A(n1796), .Y(n3301) );
  AND2X1 U2590 ( .A(n1654), .B(n1812), .Y(n1813) );
  INVX1 U2591 ( .A(n1813), .Y(n3302) );
  AND2X1 U2592 ( .A(n1635), .B(n1830), .Y(n1838) );
  INVX1 U2593 ( .A(n1838), .Y(n3303) );
  AND2X1 U2594 ( .A(n1633), .B(n1847), .Y(n1854) );
  INVX1 U2595 ( .A(n1854), .Y(n3304) );
  AND2X1 U2596 ( .A(n1660), .B(n1864), .Y(n1868) );
  INVX1 U2597 ( .A(n1868), .Y(n3305) );
  AND2X1 U2598 ( .A(n1639), .B(n1864), .Y(n1874) );
  INVX1 U2599 ( .A(n1874), .Y(n3306) );
  AND2X1 U2600 ( .A(n1658), .B(n1881), .Y(n1884) );
  INVX1 U2601 ( .A(n1884), .Y(n3307) );
  AND2X1 U2602 ( .A(n1656), .B(n1898), .Y(n1900) );
  INVX1 U2603 ( .A(n1900), .Y(n3308) );
  AND2X1 U2604 ( .A(n1635), .B(n1915), .Y(n1923) );
  INVX1 U2605 ( .A(n1923), .Y(n3309) );
  AND2X1 U2606 ( .A(n1633), .B(n1932), .Y(n1939) );
  INVX1 U2607 ( .A(n1939), .Y(n3310) );
  AND2X1 U2608 ( .A(n1639), .B(n1950), .Y(n1960) );
  INVX1 U2609 ( .A(n1960), .Y(n3311) );
  AND2X1 U2610 ( .A(n1660), .B(n1967), .Y(n1971) );
  INVX1 U2611 ( .A(n1971), .Y(n3312) );
  AND2X1 U2612 ( .A(n1637), .B(n1967), .Y(n1976) );
  INVX1 U2613 ( .A(n1976), .Y(n3313) );
  AND2X1 U2614 ( .A(n1631), .B(n1984), .Y(n1990) );
  INVX1 U2615 ( .A(n1990), .Y(n3314) );
  AND2X1 U2616 ( .A(n1643), .B(n1984), .Y(n1996) );
  INVX1 U2617 ( .A(n1996), .Y(n3315) );
  AND2X1 U2618 ( .A(n1629), .B(n2001), .Y(n2006) );
  INVX1 U2619 ( .A(n2006), .Y(n3316) );
  AND2X1 U2620 ( .A(n1641), .B(n2001), .Y(n2012) );
  INVX1 U2621 ( .A(n2012), .Y(n3317) );
  AND2X1 U2622 ( .A(n1647), .B(n2018), .Y(n2032) );
  INVX1 U2623 ( .A(n2032), .Y(n3318) );
  AND2X1 U2624 ( .A(n1645), .B(n2035), .Y(n2048) );
  INVX1 U2625 ( .A(n2048), .Y(n3319) );
  AND2X1 U2626 ( .A(n1651), .B(n2052), .Y(n2068) );
  INVX1 U2627 ( .A(n2068), .Y(n3320) );
  AND2X1 U2628 ( .A(n1649), .B(n2069), .Y(n2084) );
  INVX1 U2629 ( .A(n2084), .Y(n3321) );
  AND2X1 U2630 ( .A(n1658), .B(n2087), .Y(n2090) );
  INVX1 U2631 ( .A(n2090), .Y(n3322) );
  AND2X1 U2632 ( .A(n1639), .B(n2087), .Y(n2097) );
  INVX1 U2633 ( .A(n2097), .Y(n3323) );
  AND2X1 U2634 ( .A(n1658), .B(n2104), .Y(n2107) );
  INVX1 U2635 ( .A(n2107), .Y(n3324) );
  AND2X1 U2636 ( .A(n1637), .B(n2104), .Y(n2113) );
  INVX1 U2637 ( .A(n2113), .Y(n3325) );
  AND2X1 U2638 ( .A(n1631), .B(n2121), .Y(n2127) );
  INVX1 U2639 ( .A(n2127), .Y(n3326) );
  AND2X1 U2640 ( .A(n1643), .B(n2121), .Y(n2133) );
  INVX1 U2641 ( .A(n2133), .Y(n3327) );
  AND2X1 U2642 ( .A(n1629), .B(n2138), .Y(n2143) );
  INVX1 U2643 ( .A(n2143), .Y(n3328) );
  AND2X1 U2644 ( .A(n1641), .B(n2138), .Y(n2149) );
  INVX1 U2645 ( .A(n2149), .Y(n3329) );
  AND2X1 U2646 ( .A(n1647), .B(n2155), .Y(n2169) );
  INVX1 U2647 ( .A(n2169), .Y(n3330) );
  AND2X1 U2648 ( .A(n1645), .B(n2172), .Y(n2185) );
  INVX1 U2649 ( .A(n2185), .Y(n3331) );
  AND2X1 U2650 ( .A(n1651), .B(n2189), .Y(n2205) );
  INVX1 U2651 ( .A(n2205), .Y(n3332) );
  AND2X1 U2652 ( .A(n1649), .B(n2206), .Y(n2221) );
  INVX1 U2653 ( .A(n2221), .Y(n3333) );
  AND2X1 U2654 ( .A(n1637), .B(n1627), .Y(n1636) );
  INVX1 U2655 ( .A(n1636), .Y(n3334) );
  AND2X1 U2656 ( .A(n1631), .B(n1652), .Y(n1662) );
  INVX1 U2657 ( .A(n1662), .Y(n3335) );
  AND2X1 U2658 ( .A(n1643), .B(n1652), .Y(n1668) );
  INVX1 U2659 ( .A(n1668), .Y(n3336) );
  AND2X1 U2660 ( .A(n1629), .B(n1675), .Y(n1680) );
  INVX1 U2661 ( .A(n1680), .Y(n3337) );
  AND2X1 U2662 ( .A(n1641), .B(n1675), .Y(n1686) );
  INVX1 U2663 ( .A(n1686), .Y(n3338) );
  AND2X1 U2664 ( .A(n1647), .B(n1693), .Y(n1707) );
  INVX1 U2665 ( .A(n1707), .Y(n3339) );
  AND2X1 U2666 ( .A(n1645), .B(n1711), .Y(n1724) );
  INVX1 U2667 ( .A(n1724), .Y(n3340) );
  AND2X1 U2668 ( .A(n1651), .B(n1729), .Y(n1745) );
  INVX1 U2669 ( .A(n1745), .Y(n3341) );
  AND2X1 U2670 ( .A(n1649), .B(n1747), .Y(n1762) );
  INVX1 U2671 ( .A(n1762), .Y(n3342) );
  BUFX2 U2672 ( .A(n1770), .Y(n3343) );
  INVX1 U2673 ( .A(n1610), .Y(n3344) );
  BUFX2 U2674 ( .A(n1673), .Y(n3345) );
  BUFX2 U2675 ( .A(n1811), .Y(n3346) );
  AND2X1 U2676 ( .A(n1654), .B(n1794), .Y(n1795) );
  INVX1 U2677 ( .A(n1795), .Y(n3347) );
  AND2X1 U2678 ( .A(n1656), .B(n1812), .Y(n1814) );
  INVX1 U2679 ( .A(n1814), .Y(n3348) );
  AND2X1 U2680 ( .A(n1633), .B(n1830), .Y(n1837) );
  INVX1 U2681 ( .A(n1837), .Y(n3349) );
  AND2X1 U2682 ( .A(n1635), .B(n1847), .Y(n1855) );
  INVX1 U2683 ( .A(n1855), .Y(n3350) );
  AND2X1 U2684 ( .A(n1658), .B(n1864), .Y(n1867) );
  INVX1 U2685 ( .A(n1867), .Y(n3351) );
  AND2X1 U2686 ( .A(n1637), .B(n1864), .Y(n1873) );
  INVX1 U2687 ( .A(n1873), .Y(n3352) );
  AND2X1 U2688 ( .A(n1660), .B(n1881), .Y(n1885) );
  INVX1 U2689 ( .A(n1885), .Y(n3353) );
  AND2X1 U2690 ( .A(n1654), .B(n1898), .Y(n1899) );
  INVX1 U2691 ( .A(n1899), .Y(n3354) );
  AND2X1 U2692 ( .A(n1633), .B(n1915), .Y(n1922) );
  INVX1 U2693 ( .A(n1922), .Y(n3355) );
  AND2X1 U2694 ( .A(n1635), .B(n1932), .Y(n1940) );
  INVX1 U2695 ( .A(n1940), .Y(n3356) );
  AND2X1 U2696 ( .A(n1656), .B(n1950), .Y(n1952) );
  INVX1 U2697 ( .A(n1952), .Y(n3357) );
  AND2X1 U2698 ( .A(n1637), .B(n1950), .Y(n1959) );
  INVX1 U2699 ( .A(n1959), .Y(n3358) );
  AND2X1 U2700 ( .A(n1658), .B(n1967), .Y(n1970) );
  INVX1 U2701 ( .A(n1970), .Y(n3359) );
  AND2X1 U2702 ( .A(n1639), .B(n1967), .Y(n1977) );
  INVX1 U2703 ( .A(n1977), .Y(n3360) );
  AND2X1 U2704 ( .A(n1629), .B(n1984), .Y(n1989) );
  INVX1 U2705 ( .A(n1989), .Y(n3361) );
  AND2X1 U2706 ( .A(n1641), .B(n1984), .Y(n1995) );
  INVX1 U2707 ( .A(n1995), .Y(n3362) );
  AND2X1 U2708 ( .A(n1631), .B(n2001), .Y(n2007) );
  INVX1 U2709 ( .A(n2007), .Y(n3363) );
  AND2X1 U2710 ( .A(n1643), .B(n2001), .Y(n2013) );
  INVX1 U2711 ( .A(n2013), .Y(n3364) );
  AND2X1 U2712 ( .A(n1645), .B(n2018), .Y(n2031) );
  INVX1 U2713 ( .A(n2031), .Y(n3365) );
  AND2X1 U2714 ( .A(n1647), .B(n2035), .Y(n2049) );
  INVX1 U2715 ( .A(n2049), .Y(n3366) );
  AND2X1 U2716 ( .A(n1649), .B(n2052), .Y(n2067) );
  INVX1 U2717 ( .A(n2067), .Y(n3367) );
  AND2X1 U2718 ( .A(n1651), .B(n2069), .Y(n2085) );
  INVX1 U2719 ( .A(n2085), .Y(n3368) );
  AND2X1 U2720 ( .A(n1660), .B(n2087), .Y(n2091) );
  INVX1 U2721 ( .A(n2091), .Y(n3369) );
  AND2X1 U2722 ( .A(n1637), .B(n2087), .Y(n2096) );
  INVX1 U2723 ( .A(n2096), .Y(n3370) );
  AND2X1 U2724 ( .A(n1660), .B(n2104), .Y(n2108) );
  INVX1 U2725 ( .A(n2108), .Y(n3371) );
  AND2X1 U2726 ( .A(n1639), .B(n2104), .Y(n2114) );
  INVX1 U2727 ( .A(n2114), .Y(n3372) );
  AND2X1 U2728 ( .A(n1629), .B(n2121), .Y(n2126) );
  INVX1 U2729 ( .A(n2126), .Y(n3373) );
  AND2X1 U2730 ( .A(n1641), .B(n2121), .Y(n2132) );
  INVX1 U2731 ( .A(n2132), .Y(n3374) );
  AND2X1 U2732 ( .A(n1631), .B(n2138), .Y(n2144) );
  INVX1 U2733 ( .A(n2144), .Y(n3375) );
  AND2X1 U2734 ( .A(n1643), .B(n2138), .Y(n2150) );
  INVX1 U2735 ( .A(n2150), .Y(n3376) );
  AND2X1 U2736 ( .A(n1645), .B(n2155), .Y(n2168) );
  INVX1 U2737 ( .A(n2168), .Y(n3377) );
  AND2X1 U2738 ( .A(n1647), .B(n2172), .Y(n2186) );
  INVX1 U2739 ( .A(n2186), .Y(n3378) );
  AND2X1 U2740 ( .A(n1649), .B(n2189), .Y(n2204) );
  INVX1 U2741 ( .A(n2204), .Y(n3379) );
  AND2X1 U2742 ( .A(n1651), .B(n2206), .Y(n2222) );
  INVX1 U2743 ( .A(n2222), .Y(n3380) );
  AND2X1 U2744 ( .A(n1639), .B(n1627), .Y(n1638) );
  INVX1 U2745 ( .A(n1638), .Y(n3381) );
  AND2X1 U2746 ( .A(n1629), .B(n1652), .Y(n1661) );
  INVX1 U2747 ( .A(n1661), .Y(n3382) );
  AND2X1 U2748 ( .A(n1641), .B(n1652), .Y(n1667) );
  INVX1 U2749 ( .A(n1667), .Y(n3383) );
  AND2X1 U2750 ( .A(n1631), .B(n1675), .Y(n1681) );
  INVX1 U2751 ( .A(n1681), .Y(n3384) );
  AND2X1 U2752 ( .A(n1643), .B(n1675), .Y(n1687) );
  INVX1 U2753 ( .A(n1687), .Y(n3385) );
  AND2X1 U2754 ( .A(n1645), .B(n1693), .Y(n1706) );
  INVX1 U2755 ( .A(n1706), .Y(n3386) );
  AND2X1 U2756 ( .A(n1647), .B(n1711), .Y(n1725) );
  INVX1 U2757 ( .A(n1725), .Y(n3387) );
  AND2X1 U2758 ( .A(n1649), .B(n1729), .Y(n1744) );
  INVX1 U2759 ( .A(n1744), .Y(n3388) );
  AND2X1 U2760 ( .A(n1651), .B(n1747), .Y(n1763) );
  INVX1 U2761 ( .A(n1763), .Y(n3389) );
  AND2X1 U2762 ( .A(n1602), .B(n3429), .Y(n1594) );
  INVX1 U2763 ( .A(n1594), .Y(n3390) );
  AND2X1 U2764 ( .A(n3399), .B(n3422), .Y(n2231) );
  INVX1 U2765 ( .A(n2231), .Y(n3391) );
  INVX1 U2766 ( .A(n1765), .Y(n3392) );
  BUFX2 U2767 ( .A(n1949), .Y(n3393) );
  BUFX2 U2768 ( .A(n2086), .Y(n3394) );
  INVX1 U2769 ( .A(n3404), .Y(n3403) );
  INVX1 U2770 ( .A(n560), .Y(n3404) );
  INVX1 U2771 ( .A(n3414), .Y(n3413) );
  INVX1 U2772 ( .A(n3410), .Y(n3409) );
  INVX1 U2773 ( .A(n3408), .Y(n3407) );
  INVX1 U2774 ( .A(n3402), .Y(n3401) );
  INVX1 U2775 ( .A(n3343), .Y(n3400) );
  INVX1 U2776 ( .A(n3406), .Y(n3405) );
  INVX1 U2777 ( .A(n3412), .Y(n3411) );
  INVX1 U2778 ( .A(n3417), .Y(n3415) );
  INVX1 U2779 ( .A(n3417), .Y(n3416) );
  INVX1 U2780 ( .A(reset), .Y(n3417) );
  AND2X1 U2781 ( .A(n1622), .B(n3426), .Y(n560) );
  INVX1 U2782 ( .A(n552), .Y(n3414) );
  INVX1 U2783 ( .A(n558), .Y(n3408) );
  INVX1 U2784 ( .A(n557), .Y(n3410) );
  INVX1 U2785 ( .A(n561), .Y(n3402) );
  INVX1 U2786 ( .A(n559), .Y(n3406) );
  INVX1 U2787 ( .A(n553), .Y(n3412) );
  INVX1 U2788 ( .A(n3115), .Y(n3421) );
  AND2X1 U2789 ( .A(n1623), .B(n3399), .Y(n552) );
  AND2X1 U2790 ( .A(n1622), .B(n3399), .Y(n557) );
  AND2X1 U2791 ( .A(n1621), .B(n3399), .Y(n558) );
  AND2X1 U2792 ( .A(n1623), .B(n3426), .Y(n561) );
  AND2X1 U2793 ( .A(n1621), .B(n3426), .Y(n559) );
  INVX1 U2794 ( .A(n1787), .Y(n3424) );
  INVX1 U2795 ( .A(n3250), .Y(n3425) );
  BUFX2 U2796 ( .A(n580), .Y(n3396) );
  BUFX2 U2797 ( .A(n580), .Y(n3395) );
  BUFX2 U2798 ( .A(n572), .Y(n3397) );
  BUFX2 U2799 ( .A(n572), .Y(n3398) );
  INVX1 U2800 ( .A(n3399), .Y(n3426) );
  AND2X1 U2801 ( .A(n3427), .B(n3428), .Y(n1622) );
  AND2X1 U2802 ( .A(n1602), .B(n15), .Y(n564) );
  INVX1 U2803 ( .A(wr_ptr[0]), .Y(n3422) );
  BUFX2 U2804 ( .A(n12), .Y(n3399) );
  INVX1 U2805 ( .A(n2227), .Y(n3420) );
  AND2X1 U2806 ( .A(n1610), .B(n16), .Y(n1602) );
  INVX1 U2807 ( .A(n1624), .Y(fillcount[5]) );
  INVX1 U2808 ( .A(n1626), .Y(n3419) );
  INVX1 U2809 ( .A(put), .Y(n3946) );
  INVX1 U2810 ( .A(wr_ptr[3]), .Y(n3433) );
  INVX1 U2811 ( .A(n1789), .Y(n3423) );
  INVX1 U2812 ( .A(wr_ptr[2]), .Y(n3432) );
  INVX1 U2813 ( .A(n13), .Y(n3427) );
  INVX1 U2814 ( .A(wr_ptr[4]), .Y(n3430) );
  INVX1 U2815 ( .A(n15), .Y(n3429) );
  INVX1 U2816 ( .A(n14), .Y(n3428) );
  INVX1 U2817 ( .A(wr_ptr[1]), .Y(n3431) );
  AND2X1 U2818 ( .A(data_in[9]), .B(n3416), .Y(n1633) );
  AND2X1 U2819 ( .A(data_in[10]), .B(n3416), .Y(n1631) );
  AND2X1 U2820 ( .A(data_in[11]), .B(n3416), .Y(n1629) );
  AND2X1 U2821 ( .A(n14), .B(n3427), .Y(n1621) );
  AND2X1 U2822 ( .A(data_in[0]), .B(n3415), .Y(n1651) );
  AND2X1 U2823 ( .A(data_in[1]), .B(n3416), .Y(n1649) );
  AND2X1 U2824 ( .A(data_in[2]), .B(n3415), .Y(n1647) );
  AND2X1 U2825 ( .A(data_in[3]), .B(n3416), .Y(n1645) );
  AND2X1 U2826 ( .A(data_in[4]), .B(n3415), .Y(n1643) );
  AND2X1 U2827 ( .A(data_in[5]), .B(n3416), .Y(n1641) );
  AND2X1 U2828 ( .A(data_in[6]), .B(n3415), .Y(n1639) );
  AND2X1 U2829 ( .A(data_in[7]), .B(n3416), .Y(n1637) );
  AND2X1 U2830 ( .A(data_in[8]), .B(n3415), .Y(n1635) );
  AND2X1 U2831 ( .A(data_in[12]), .B(n3416), .Y(n1660) );
  AND2X1 U2832 ( .A(data_in[13]), .B(n3415), .Y(n1658) );
  AND2X1 U2833 ( .A(data_in[14]), .B(n3416), .Y(n1656) );
  AND2X1 U2834 ( .A(data_in[15]), .B(n3415), .Y(n1654) );
  AND2X1 U2835 ( .A(n13), .B(n3428), .Y(n1623) );
  INVX1 U2836 ( .A(mem[480]), .Y(n3465) );
  INVX1 U2837 ( .A(mem[416]), .Y(n3529) );
  INVX1 U2838 ( .A(mem[464]), .Y(n3481) );
  INVX1 U2839 ( .A(mem[352]), .Y(n3593) );
  INVX1 U2840 ( .A(mem[288]), .Y(n3657) );
  INVX1 U2841 ( .A(mem[336]), .Y(n3609) );
  INVX1 U2842 ( .A(mem[96]), .Y(n3849) );
  INVX1 U2843 ( .A(mem[32]), .Y(n3913) );
  INVX1 U2844 ( .A(mem[80]), .Y(n3865) );
  INVX1 U2845 ( .A(mem[481]), .Y(n3464) );
  INVX1 U2846 ( .A(mem[417]), .Y(n3528) );
  INVX1 U2847 ( .A(mem[465]), .Y(n3480) );
  INVX1 U2848 ( .A(mem[353]), .Y(n3592) );
  INVX1 U2849 ( .A(mem[289]), .Y(n3656) );
  INVX1 U2850 ( .A(mem[337]), .Y(n3608) );
  INVX1 U2851 ( .A(mem[97]), .Y(n3848) );
  INVX1 U2852 ( .A(mem[33]), .Y(n3912) );
  INVX1 U2853 ( .A(mem[81]), .Y(n3864) );
  INVX1 U2854 ( .A(mem[482]), .Y(n3463) );
  INVX1 U2855 ( .A(mem[418]), .Y(n3527) );
  INVX1 U2856 ( .A(mem[466]), .Y(n3479) );
  INVX1 U2857 ( .A(mem[354]), .Y(n3591) );
  INVX1 U2858 ( .A(mem[290]), .Y(n3655) );
  INVX1 U2859 ( .A(mem[338]), .Y(n3607) );
  INVX1 U2860 ( .A(mem[98]), .Y(n3847) );
  INVX1 U2861 ( .A(mem[34]), .Y(n3911) );
  INVX1 U2862 ( .A(mem[82]), .Y(n3863) );
  INVX1 U2863 ( .A(mem[483]), .Y(n3462) );
  INVX1 U2864 ( .A(mem[419]), .Y(n3526) );
  INVX1 U2865 ( .A(mem[467]), .Y(n3478) );
  INVX1 U2866 ( .A(mem[355]), .Y(n3590) );
  INVX1 U2867 ( .A(mem[291]), .Y(n3654) );
  INVX1 U2868 ( .A(mem[339]), .Y(n3606) );
  INVX1 U2869 ( .A(mem[99]), .Y(n3846) );
  INVX1 U2870 ( .A(mem[35]), .Y(n3910) );
  INVX1 U2871 ( .A(mem[83]), .Y(n3862) );
  INVX1 U2872 ( .A(mem[484]), .Y(n3461) );
  INVX1 U2873 ( .A(mem[420]), .Y(n3525) );
  INVX1 U2874 ( .A(mem[468]), .Y(n3477) );
  INVX1 U2875 ( .A(mem[356]), .Y(n3589) );
  INVX1 U2876 ( .A(mem[292]), .Y(n3653) );
  INVX1 U2877 ( .A(mem[340]), .Y(n3605) );
  INVX1 U2878 ( .A(mem[100]), .Y(n3845) );
  INVX1 U2879 ( .A(mem[36]), .Y(n3909) );
  INVX1 U2880 ( .A(mem[84]), .Y(n3861) );
  INVX1 U2881 ( .A(mem[485]), .Y(n3460) );
  INVX1 U2882 ( .A(mem[421]), .Y(n3524) );
  INVX1 U2883 ( .A(mem[469]), .Y(n3476) );
  INVX1 U2884 ( .A(mem[357]), .Y(n3588) );
  INVX1 U2885 ( .A(mem[293]), .Y(n3652) );
  INVX1 U2886 ( .A(mem[341]), .Y(n3604) );
  INVX1 U2887 ( .A(mem[101]), .Y(n3844) );
  INVX1 U2888 ( .A(mem[37]), .Y(n3908) );
  INVX1 U2889 ( .A(mem[85]), .Y(n3860) );
  INVX1 U2890 ( .A(mem[486]), .Y(n3459) );
  INVX1 U2891 ( .A(mem[422]), .Y(n3523) );
  INVX1 U2892 ( .A(mem[470]), .Y(n3475) );
  INVX1 U2893 ( .A(mem[358]), .Y(n3587) );
  INVX1 U2894 ( .A(mem[294]), .Y(n3651) );
  INVX1 U2895 ( .A(mem[342]), .Y(n3603) );
  INVX1 U2896 ( .A(mem[102]), .Y(n3843) );
  INVX1 U2897 ( .A(mem[38]), .Y(n3907) );
  INVX1 U2898 ( .A(mem[86]), .Y(n3859) );
  INVX1 U2899 ( .A(mem[487]), .Y(n3458) );
  INVX1 U2900 ( .A(mem[423]), .Y(n3522) );
  INVX1 U2901 ( .A(mem[471]), .Y(n3474) );
  INVX1 U2902 ( .A(mem[359]), .Y(n3586) );
  INVX1 U2903 ( .A(mem[295]), .Y(n3650) );
  INVX1 U2904 ( .A(mem[343]), .Y(n3602) );
  INVX1 U2905 ( .A(mem[103]), .Y(n3842) );
  INVX1 U2906 ( .A(mem[39]), .Y(n3906) );
  INVX1 U2907 ( .A(mem[87]), .Y(n3858) );
  INVX1 U2908 ( .A(mem[488]), .Y(n3457) );
  INVX1 U2909 ( .A(mem[424]), .Y(n3521) );
  INVX1 U2910 ( .A(mem[472]), .Y(n3473) );
  INVX1 U2911 ( .A(mem[360]), .Y(n3585) );
  INVX1 U2912 ( .A(mem[296]), .Y(n3649) );
  INVX1 U2913 ( .A(mem[344]), .Y(n3601) );
  INVX1 U2914 ( .A(mem[104]), .Y(n3841) );
  INVX1 U2915 ( .A(mem[40]), .Y(n3905) );
  INVX1 U2916 ( .A(mem[88]), .Y(n3857) );
  INVX1 U2917 ( .A(mem[489]), .Y(n3456) );
  INVX1 U2918 ( .A(mem[425]), .Y(n3520) );
  INVX1 U2919 ( .A(mem[473]), .Y(n3472) );
  INVX1 U2920 ( .A(mem[361]), .Y(n3584) );
  INVX1 U2921 ( .A(mem[297]), .Y(n3648) );
  INVX1 U2922 ( .A(mem[345]), .Y(n3600) );
  INVX1 U2923 ( .A(mem[105]), .Y(n3840) );
  INVX1 U2924 ( .A(mem[41]), .Y(n3904) );
  INVX1 U2925 ( .A(mem[89]), .Y(n3856) );
  INVX1 U2926 ( .A(mem[490]), .Y(n3455) );
  INVX1 U2927 ( .A(mem[426]), .Y(n3519) );
  INVX1 U2928 ( .A(mem[474]), .Y(n3471) );
  INVX1 U2929 ( .A(mem[362]), .Y(n3583) );
  INVX1 U2930 ( .A(mem[298]), .Y(n3647) );
  INVX1 U2931 ( .A(mem[346]), .Y(n3599) );
  INVX1 U2932 ( .A(mem[106]), .Y(n3839) );
  INVX1 U2933 ( .A(mem[42]), .Y(n3903) );
  INVX1 U2934 ( .A(mem[90]), .Y(n3855) );
  INVX1 U2935 ( .A(mem[491]), .Y(n3454) );
  INVX1 U2936 ( .A(mem[427]), .Y(n3518) );
  INVX1 U2937 ( .A(mem[475]), .Y(n3470) );
  INVX1 U2938 ( .A(mem[363]), .Y(n3582) );
  INVX1 U2939 ( .A(mem[299]), .Y(n3646) );
  INVX1 U2940 ( .A(mem[347]), .Y(n3598) );
  INVX1 U2941 ( .A(mem[107]), .Y(n3838) );
  INVX1 U2942 ( .A(mem[43]), .Y(n3902) );
  INVX1 U2943 ( .A(mem[91]), .Y(n3854) );
  INVX1 U2944 ( .A(mem[492]), .Y(n3453) );
  INVX1 U2945 ( .A(mem[428]), .Y(n3517) );
  INVX1 U2946 ( .A(mem[476]), .Y(n3469) );
  INVX1 U2947 ( .A(mem[364]), .Y(n3581) );
  INVX1 U2948 ( .A(mem[300]), .Y(n3645) );
  INVX1 U2949 ( .A(mem[348]), .Y(n3597) );
  INVX1 U2950 ( .A(mem[108]), .Y(n3837) );
  INVX1 U2951 ( .A(mem[44]), .Y(n3901) );
  INVX1 U2952 ( .A(mem[92]), .Y(n3853) );
  INVX1 U2953 ( .A(mem[493]), .Y(n3452) );
  INVX1 U2954 ( .A(mem[429]), .Y(n3516) );
  INVX1 U2955 ( .A(mem[477]), .Y(n3468) );
  INVX1 U2956 ( .A(mem[365]), .Y(n3580) );
  INVX1 U2957 ( .A(mem[301]), .Y(n3644) );
  INVX1 U2958 ( .A(mem[349]), .Y(n3596) );
  INVX1 U2959 ( .A(mem[109]), .Y(n3836) );
  INVX1 U2960 ( .A(mem[45]), .Y(n3900) );
  INVX1 U2961 ( .A(mem[93]), .Y(n3852) );
  INVX1 U2962 ( .A(mem[494]), .Y(n3451) );
  INVX1 U2963 ( .A(mem[430]), .Y(n3515) );
  INVX1 U2964 ( .A(mem[478]), .Y(n3467) );
  INVX1 U2965 ( .A(mem[366]), .Y(n3579) );
  INVX1 U2966 ( .A(mem[302]), .Y(n3643) );
  INVX1 U2967 ( .A(mem[350]), .Y(n3595) );
  INVX1 U2968 ( .A(mem[110]), .Y(n3835) );
  INVX1 U2969 ( .A(mem[46]), .Y(n3899) );
  INVX1 U2970 ( .A(mem[94]), .Y(n3851) );
  INVX1 U2971 ( .A(mem[495]), .Y(n3450) );
  INVX1 U2972 ( .A(mem[431]), .Y(n3514) );
  INVX1 U2973 ( .A(mem[479]), .Y(n3466) );
  INVX1 U2974 ( .A(mem[367]), .Y(n3578) );
  INVX1 U2975 ( .A(mem[303]), .Y(n3642) );
  INVX1 U2976 ( .A(mem[351]), .Y(n3594) );
  INVX1 U2977 ( .A(mem[111]), .Y(n3834) );
  INVX1 U2978 ( .A(mem[47]), .Y(n3898) );
  INVX1 U2979 ( .A(mem[95]), .Y(n3850) );
  INVX1 U2980 ( .A(mem[224]), .Y(n3721) );
  INVX1 U2981 ( .A(mem[160]), .Y(n3785) );
  INVX1 U2982 ( .A(mem[208]), .Y(n3737) );
  INVX1 U2983 ( .A(mem[225]), .Y(n3720) );
  INVX1 U2984 ( .A(mem[161]), .Y(n3784) );
  INVX1 U2985 ( .A(mem[209]), .Y(n3736) );
  INVX1 U2986 ( .A(mem[226]), .Y(n3719) );
  INVX1 U2987 ( .A(mem[162]), .Y(n3783) );
  INVX1 U2988 ( .A(mem[210]), .Y(n3735) );
  INVX1 U2989 ( .A(mem[227]), .Y(n3718) );
  INVX1 U2990 ( .A(mem[163]), .Y(n3782) );
  INVX1 U2991 ( .A(mem[211]), .Y(n3734) );
  INVX1 U2992 ( .A(mem[228]), .Y(n3717) );
  INVX1 U2993 ( .A(mem[164]), .Y(n3781) );
  INVX1 U2994 ( .A(mem[212]), .Y(n3733) );
  INVX1 U2995 ( .A(mem[229]), .Y(n3716) );
  INVX1 U2996 ( .A(mem[165]), .Y(n3780) );
  INVX1 U2997 ( .A(mem[213]), .Y(n3732) );
  INVX1 U2998 ( .A(mem[230]), .Y(n3715) );
  INVX1 U2999 ( .A(mem[166]), .Y(n3779) );
  INVX1 U3000 ( .A(mem[214]), .Y(n3731) );
  INVX1 U3001 ( .A(mem[231]), .Y(n3714) );
  INVX1 U3002 ( .A(mem[167]), .Y(n3778) );
  INVX1 U3003 ( .A(mem[215]), .Y(n3730) );
  INVX1 U3004 ( .A(mem[232]), .Y(n3713) );
  INVX1 U3005 ( .A(mem[168]), .Y(n3777) );
  INVX1 U3006 ( .A(mem[216]), .Y(n3729) );
  INVX1 U3007 ( .A(mem[233]), .Y(n3712) );
  INVX1 U3008 ( .A(mem[169]), .Y(n3776) );
  INVX1 U3009 ( .A(mem[217]), .Y(n3728) );
  INVX1 U3010 ( .A(mem[234]), .Y(n3711) );
  INVX1 U3011 ( .A(mem[170]), .Y(n3775) );
  INVX1 U3012 ( .A(mem[218]), .Y(n3727) );
  INVX1 U3013 ( .A(mem[235]), .Y(n3710) );
  INVX1 U3014 ( .A(mem[171]), .Y(n3774) );
  INVX1 U3015 ( .A(mem[219]), .Y(n3726) );
  INVX1 U3016 ( .A(mem[236]), .Y(n3709) );
  INVX1 U3017 ( .A(mem[172]), .Y(n3773) );
  INVX1 U3018 ( .A(mem[220]), .Y(n3725) );
  INVX1 U3019 ( .A(mem[237]), .Y(n3708) );
  INVX1 U3020 ( .A(mem[173]), .Y(n3772) );
  INVX1 U3021 ( .A(mem[221]), .Y(n3724) );
  INVX1 U3022 ( .A(mem[238]), .Y(n3707) );
  INVX1 U3023 ( .A(mem[174]), .Y(n3771) );
  INVX1 U3024 ( .A(mem[222]), .Y(n3723) );
  INVX1 U3025 ( .A(mem[239]), .Y(n3706) );
  INVX1 U3026 ( .A(mem[175]), .Y(n3770) );
  INVX1 U3027 ( .A(mem[223]), .Y(n3722) );
  INVX1 U3028 ( .A(mem[432]), .Y(n3513) );
  INVX1 U3029 ( .A(mem[384]), .Y(n3561) );
  INVX1 U3030 ( .A(mem[400]), .Y(n3545) );
  INVX1 U3031 ( .A(mem[304]), .Y(n3641) );
  INVX1 U3032 ( .A(mem[256]), .Y(n3689) );
  INVX1 U3033 ( .A(mem[272]), .Y(n3673) );
  INVX1 U3034 ( .A(mem[48]), .Y(n3897) );
  INVX1 U3035 ( .A(mem[0]), .Y(n3945) );
  INVX1 U3036 ( .A(mem[16]), .Y(n3929) );
  INVX1 U3037 ( .A(mem[433]), .Y(n3512) );
  INVX1 U3038 ( .A(mem[385]), .Y(n3560) );
  INVX1 U3039 ( .A(mem[401]), .Y(n3544) );
  INVX1 U3040 ( .A(mem[305]), .Y(n3640) );
  INVX1 U3041 ( .A(mem[257]), .Y(n3688) );
  INVX1 U3042 ( .A(mem[273]), .Y(n3672) );
  INVX1 U3043 ( .A(mem[49]), .Y(n3896) );
  INVX1 U3044 ( .A(mem[1]), .Y(n3944) );
  INVX1 U3045 ( .A(mem[17]), .Y(n3928) );
  INVX1 U3046 ( .A(mem[434]), .Y(n3511) );
  INVX1 U3047 ( .A(mem[386]), .Y(n3559) );
  INVX1 U3048 ( .A(mem[402]), .Y(n3543) );
  INVX1 U3049 ( .A(mem[306]), .Y(n3639) );
  INVX1 U3050 ( .A(mem[258]), .Y(n3687) );
  INVX1 U3051 ( .A(mem[274]), .Y(n3671) );
  INVX1 U3052 ( .A(mem[50]), .Y(n3895) );
  INVX1 U3053 ( .A(mem[2]), .Y(n3943) );
  INVX1 U3054 ( .A(mem[18]), .Y(n3927) );
  INVX1 U3055 ( .A(mem[435]), .Y(n3510) );
  INVX1 U3056 ( .A(mem[387]), .Y(n3558) );
  INVX1 U3057 ( .A(mem[403]), .Y(n3542) );
  INVX1 U3058 ( .A(mem[307]), .Y(n3638) );
  INVX1 U3059 ( .A(mem[259]), .Y(n3686) );
  INVX1 U3060 ( .A(mem[275]), .Y(n3670) );
  INVX1 U3061 ( .A(mem[51]), .Y(n3894) );
  INVX1 U3062 ( .A(mem[3]), .Y(n3942) );
  INVX1 U3063 ( .A(mem[19]), .Y(n3926) );
  INVX1 U3064 ( .A(mem[436]), .Y(n3509) );
  INVX1 U3065 ( .A(mem[388]), .Y(n3557) );
  INVX1 U3066 ( .A(mem[404]), .Y(n3541) );
  INVX1 U3067 ( .A(mem[308]), .Y(n3637) );
  INVX1 U3068 ( .A(mem[260]), .Y(n3685) );
  INVX1 U3069 ( .A(mem[276]), .Y(n3669) );
  INVX1 U3070 ( .A(mem[52]), .Y(n3893) );
  INVX1 U3071 ( .A(mem[4]), .Y(n3941) );
  INVX1 U3072 ( .A(mem[20]), .Y(n3925) );
  INVX1 U3073 ( .A(mem[437]), .Y(n3508) );
  INVX1 U3074 ( .A(mem[389]), .Y(n3556) );
  INVX1 U3075 ( .A(mem[405]), .Y(n3540) );
  INVX1 U3076 ( .A(mem[309]), .Y(n3636) );
  INVX1 U3077 ( .A(mem[261]), .Y(n3684) );
  INVX1 U3078 ( .A(mem[277]), .Y(n3668) );
  INVX1 U3079 ( .A(mem[53]), .Y(n3892) );
  INVX1 U3080 ( .A(mem[5]), .Y(n3940) );
  INVX1 U3081 ( .A(mem[21]), .Y(n3924) );
  INVX1 U3082 ( .A(mem[438]), .Y(n3507) );
  INVX1 U3083 ( .A(mem[390]), .Y(n3555) );
  INVX1 U3084 ( .A(mem[406]), .Y(n3539) );
  INVX1 U3085 ( .A(mem[310]), .Y(n3635) );
  INVX1 U3086 ( .A(mem[262]), .Y(n3683) );
  INVX1 U3087 ( .A(mem[278]), .Y(n3667) );
  INVX1 U3088 ( .A(mem[54]), .Y(n3891) );
  INVX1 U3089 ( .A(mem[6]), .Y(n3939) );
  INVX1 U3090 ( .A(mem[22]), .Y(n3923) );
  INVX1 U3091 ( .A(mem[439]), .Y(n3506) );
  INVX1 U3092 ( .A(mem[391]), .Y(n3554) );
  INVX1 U3093 ( .A(mem[407]), .Y(n3538) );
  INVX1 U3094 ( .A(mem[311]), .Y(n3634) );
  INVX1 U3095 ( .A(mem[263]), .Y(n3682) );
  INVX1 U3096 ( .A(mem[279]), .Y(n3666) );
  INVX1 U3097 ( .A(mem[55]), .Y(n3890) );
  INVX1 U3098 ( .A(mem[7]), .Y(n3938) );
  INVX1 U3099 ( .A(mem[23]), .Y(n3922) );
  INVX1 U3100 ( .A(mem[440]), .Y(n3505) );
  INVX1 U3101 ( .A(mem[392]), .Y(n3553) );
  INVX1 U3102 ( .A(mem[408]), .Y(n3537) );
  INVX1 U3103 ( .A(mem[312]), .Y(n3633) );
  INVX1 U3104 ( .A(mem[264]), .Y(n3681) );
  INVX1 U3105 ( .A(mem[280]), .Y(n3665) );
  INVX1 U3106 ( .A(mem[56]), .Y(n3889) );
  INVX1 U3107 ( .A(mem[8]), .Y(n3937) );
  INVX1 U3108 ( .A(mem[24]), .Y(n3921) );
  INVX1 U3109 ( .A(mem[441]), .Y(n3504) );
  INVX1 U3110 ( .A(mem[393]), .Y(n3552) );
  INVX1 U3111 ( .A(mem[409]), .Y(n3536) );
  INVX1 U3112 ( .A(mem[313]), .Y(n3632) );
  INVX1 U3113 ( .A(mem[265]), .Y(n3680) );
  INVX1 U3114 ( .A(mem[281]), .Y(n3664) );
  INVX1 U3115 ( .A(mem[57]), .Y(n3888) );
  INVX1 U3116 ( .A(mem[9]), .Y(n3936) );
  INVX1 U3117 ( .A(mem[25]), .Y(n3920) );
  INVX1 U3118 ( .A(mem[442]), .Y(n3503) );
  INVX1 U3119 ( .A(mem[394]), .Y(n3551) );
  INVX1 U3120 ( .A(mem[410]), .Y(n3535) );
  INVX1 U3121 ( .A(mem[314]), .Y(n3631) );
  INVX1 U3122 ( .A(mem[266]), .Y(n3679) );
  INVX1 U3123 ( .A(mem[282]), .Y(n3663) );
  INVX1 U3124 ( .A(mem[58]), .Y(n3887) );
  INVX1 U3125 ( .A(mem[10]), .Y(n3935) );
  INVX1 U3126 ( .A(mem[26]), .Y(n3919) );
  INVX1 U3127 ( .A(mem[443]), .Y(n3502) );
  INVX1 U3128 ( .A(mem[395]), .Y(n3550) );
  INVX1 U3129 ( .A(mem[411]), .Y(n3534) );
  INVX1 U3130 ( .A(mem[315]), .Y(n3630) );
  INVX1 U3131 ( .A(mem[267]), .Y(n3678) );
  INVX1 U3132 ( .A(mem[283]), .Y(n3662) );
  INVX1 U3133 ( .A(mem[59]), .Y(n3886) );
  INVX1 U3134 ( .A(mem[11]), .Y(n3934) );
  INVX1 U3135 ( .A(mem[27]), .Y(n3918) );
  INVX1 U3136 ( .A(mem[444]), .Y(n3501) );
  INVX1 U3137 ( .A(mem[396]), .Y(n3549) );
  INVX1 U3138 ( .A(mem[412]), .Y(n3533) );
  INVX1 U3139 ( .A(mem[316]), .Y(n3629) );
  INVX1 U3140 ( .A(mem[268]), .Y(n3677) );
  INVX1 U3141 ( .A(mem[284]), .Y(n3661) );
  INVX1 U3142 ( .A(mem[60]), .Y(n3885) );
  INVX1 U3143 ( .A(mem[12]), .Y(n3933) );
  INVX1 U3144 ( .A(mem[28]), .Y(n3917) );
  INVX1 U3145 ( .A(mem[445]), .Y(n3500) );
  INVX1 U3146 ( .A(mem[397]), .Y(n3548) );
  INVX1 U3147 ( .A(mem[413]), .Y(n3532) );
  INVX1 U3148 ( .A(mem[317]), .Y(n3628) );
  INVX1 U3149 ( .A(mem[269]), .Y(n3676) );
  INVX1 U3150 ( .A(mem[285]), .Y(n3660) );
  INVX1 U3151 ( .A(mem[61]), .Y(n3884) );
  INVX1 U3152 ( .A(mem[13]), .Y(n3932) );
  INVX1 U3153 ( .A(mem[29]), .Y(n3916) );
  INVX1 U3154 ( .A(mem[446]), .Y(n3499) );
  INVX1 U3155 ( .A(mem[398]), .Y(n3547) );
  INVX1 U3156 ( .A(mem[414]), .Y(n3531) );
  INVX1 U3157 ( .A(mem[318]), .Y(n3627) );
  INVX1 U3158 ( .A(mem[270]), .Y(n3675) );
  INVX1 U3159 ( .A(mem[286]), .Y(n3659) );
  INVX1 U3160 ( .A(mem[62]), .Y(n3883) );
  INVX1 U3161 ( .A(mem[14]), .Y(n3931) );
  INVX1 U3162 ( .A(mem[30]), .Y(n3915) );
  INVX1 U3163 ( .A(mem[447]), .Y(n3498) );
  INVX1 U3164 ( .A(mem[399]), .Y(n3546) );
  INVX1 U3165 ( .A(mem[415]), .Y(n3530) );
  INVX1 U3166 ( .A(mem[319]), .Y(n3626) );
  INVX1 U3167 ( .A(mem[271]), .Y(n3674) );
  INVX1 U3168 ( .A(mem[287]), .Y(n3658) );
  INVX1 U3169 ( .A(mem[63]), .Y(n3882) );
  INVX1 U3170 ( .A(mem[15]), .Y(n3930) );
  INVX1 U3171 ( .A(mem[31]), .Y(n3914) );
  INVX1 U3172 ( .A(mem[176]), .Y(n3769) );
  INVX1 U3173 ( .A(mem[128]), .Y(n3817) );
  INVX1 U3174 ( .A(mem[144]), .Y(n3801) );
  INVX1 U3175 ( .A(mem[177]), .Y(n3768) );
  INVX1 U3176 ( .A(mem[129]), .Y(n3816) );
  INVX1 U3177 ( .A(mem[145]), .Y(n3800) );
  INVX1 U3178 ( .A(mem[178]), .Y(n3767) );
  INVX1 U3179 ( .A(mem[130]), .Y(n3815) );
  INVX1 U3180 ( .A(mem[146]), .Y(n3799) );
  INVX1 U3181 ( .A(mem[179]), .Y(n3766) );
  INVX1 U3182 ( .A(mem[131]), .Y(n3814) );
  INVX1 U3183 ( .A(mem[147]), .Y(n3798) );
  INVX1 U3184 ( .A(mem[180]), .Y(n3765) );
  INVX1 U3185 ( .A(mem[132]), .Y(n3813) );
  INVX1 U3186 ( .A(mem[148]), .Y(n3797) );
  INVX1 U3187 ( .A(mem[181]), .Y(n3764) );
  INVX1 U3188 ( .A(mem[133]), .Y(n3812) );
  INVX1 U3189 ( .A(mem[149]), .Y(n3796) );
  INVX1 U3190 ( .A(mem[182]), .Y(n3763) );
  INVX1 U3191 ( .A(mem[134]), .Y(n3811) );
  INVX1 U3192 ( .A(mem[150]), .Y(n3795) );
  INVX1 U3193 ( .A(mem[183]), .Y(n3762) );
  INVX1 U3194 ( .A(mem[135]), .Y(n3810) );
  INVX1 U3195 ( .A(mem[151]), .Y(n3794) );
  INVX1 U3196 ( .A(mem[184]), .Y(n3761) );
  INVX1 U3197 ( .A(mem[136]), .Y(n3809) );
  INVX1 U3198 ( .A(mem[152]), .Y(n3793) );
  INVX1 U3199 ( .A(mem[185]), .Y(n3760) );
  INVX1 U3200 ( .A(mem[137]), .Y(n3808) );
  INVX1 U3201 ( .A(mem[153]), .Y(n3792) );
  INVX1 U3202 ( .A(mem[186]), .Y(n3759) );
  INVX1 U3203 ( .A(mem[138]), .Y(n3807) );
  INVX1 U3204 ( .A(mem[154]), .Y(n3791) );
  INVX1 U3205 ( .A(mem[187]), .Y(n3758) );
  INVX1 U3206 ( .A(mem[139]), .Y(n3806) );
  INVX1 U3207 ( .A(mem[155]), .Y(n3790) );
  INVX1 U3208 ( .A(mem[188]), .Y(n3757) );
  INVX1 U3209 ( .A(mem[140]), .Y(n3805) );
  INVX1 U3210 ( .A(mem[156]), .Y(n3789) );
  INVX1 U3211 ( .A(mem[189]), .Y(n3756) );
  INVX1 U3212 ( .A(mem[141]), .Y(n3804) );
  INVX1 U3213 ( .A(mem[157]), .Y(n3788) );
  INVX1 U3214 ( .A(mem[190]), .Y(n3755) );
  INVX1 U3215 ( .A(mem[142]), .Y(n3803) );
  INVX1 U3216 ( .A(mem[158]), .Y(n3787) );
  INVX1 U3217 ( .A(mem[191]), .Y(n3754) );
  INVX1 U3218 ( .A(mem[143]), .Y(n3802) );
  INVX1 U3219 ( .A(mem[159]), .Y(n3786) );
  INVX1 U3220 ( .A(mem[496]), .Y(n3449) );
  INVX1 U3221 ( .A(mem[448]), .Y(n3497) );
  INVX1 U3222 ( .A(mem[368]), .Y(n3577) );
  INVX1 U3223 ( .A(mem[320]), .Y(n3625) );
  INVX1 U3224 ( .A(mem[112]), .Y(n3833) );
  INVX1 U3225 ( .A(mem[64]), .Y(n3881) );
  INVX1 U3226 ( .A(mem[497]), .Y(n3448) );
  INVX1 U3227 ( .A(mem[449]), .Y(n3496) );
  INVX1 U3228 ( .A(mem[369]), .Y(n3576) );
  INVX1 U3229 ( .A(mem[321]), .Y(n3624) );
  INVX1 U3230 ( .A(mem[113]), .Y(n3832) );
  INVX1 U3231 ( .A(mem[65]), .Y(n3880) );
  INVX1 U3232 ( .A(mem[498]), .Y(n3447) );
  INVX1 U3233 ( .A(mem[450]), .Y(n3495) );
  INVX1 U3234 ( .A(mem[370]), .Y(n3575) );
  INVX1 U3235 ( .A(mem[322]), .Y(n3623) );
  INVX1 U3236 ( .A(mem[114]), .Y(n3831) );
  INVX1 U3237 ( .A(mem[66]), .Y(n3879) );
  INVX1 U3238 ( .A(mem[499]), .Y(n3446) );
  INVX1 U3239 ( .A(mem[451]), .Y(n3494) );
  INVX1 U3240 ( .A(mem[371]), .Y(n3574) );
  INVX1 U3241 ( .A(mem[323]), .Y(n3622) );
  INVX1 U3242 ( .A(mem[115]), .Y(n3830) );
  INVX1 U3243 ( .A(mem[67]), .Y(n3878) );
  INVX1 U3244 ( .A(mem[500]), .Y(n3445) );
  INVX1 U3245 ( .A(mem[452]), .Y(n3493) );
  INVX1 U3246 ( .A(mem[372]), .Y(n3573) );
  INVX1 U3247 ( .A(mem[324]), .Y(n3621) );
  INVX1 U3248 ( .A(mem[116]), .Y(n3829) );
  INVX1 U3249 ( .A(mem[68]), .Y(n3877) );
  INVX1 U3250 ( .A(mem[501]), .Y(n3444) );
  INVX1 U3251 ( .A(mem[453]), .Y(n3492) );
  INVX1 U3252 ( .A(mem[373]), .Y(n3572) );
  INVX1 U3253 ( .A(mem[325]), .Y(n3620) );
  INVX1 U3254 ( .A(mem[117]), .Y(n3828) );
  INVX1 U3255 ( .A(mem[69]), .Y(n3876) );
  INVX1 U3256 ( .A(mem[502]), .Y(n3443) );
  INVX1 U3257 ( .A(mem[454]), .Y(n3491) );
  INVX1 U3258 ( .A(mem[374]), .Y(n3571) );
  INVX1 U3259 ( .A(mem[326]), .Y(n3619) );
  INVX1 U3260 ( .A(mem[118]), .Y(n3827) );
  INVX1 U3261 ( .A(mem[70]), .Y(n3875) );
  INVX1 U3262 ( .A(mem[503]), .Y(n3442) );
  INVX1 U3263 ( .A(mem[455]), .Y(n3490) );
  INVX1 U3264 ( .A(mem[375]), .Y(n3570) );
  INVX1 U3265 ( .A(mem[327]), .Y(n3618) );
  INVX1 U3266 ( .A(mem[119]), .Y(n3826) );
  INVX1 U3267 ( .A(mem[71]), .Y(n3874) );
  INVX1 U3268 ( .A(mem[504]), .Y(n3441) );
  INVX1 U3269 ( .A(mem[456]), .Y(n3489) );
  INVX1 U3270 ( .A(mem[376]), .Y(n3569) );
  INVX1 U3271 ( .A(mem[328]), .Y(n3617) );
  INVX1 U3272 ( .A(mem[120]), .Y(n3825) );
  INVX1 U3273 ( .A(mem[72]), .Y(n3873) );
  INVX1 U3274 ( .A(mem[505]), .Y(n3440) );
  INVX1 U3275 ( .A(mem[457]), .Y(n3488) );
  INVX1 U3276 ( .A(mem[377]), .Y(n3568) );
  INVX1 U3277 ( .A(mem[329]), .Y(n3616) );
  INVX1 U3278 ( .A(mem[121]), .Y(n3824) );
  INVX1 U3279 ( .A(mem[73]), .Y(n3872) );
  INVX1 U3280 ( .A(mem[506]), .Y(n3439) );
  INVX1 U3281 ( .A(mem[458]), .Y(n3487) );
  INVX1 U3282 ( .A(mem[378]), .Y(n3567) );
  INVX1 U3283 ( .A(mem[330]), .Y(n3615) );
  INVX1 U3284 ( .A(mem[122]), .Y(n3823) );
  INVX1 U3285 ( .A(mem[74]), .Y(n3871) );
  INVX1 U3286 ( .A(mem[507]), .Y(n3438) );
  INVX1 U3287 ( .A(mem[459]), .Y(n3486) );
  INVX1 U3288 ( .A(mem[379]), .Y(n3566) );
  INVX1 U3289 ( .A(mem[331]), .Y(n3614) );
  INVX1 U3290 ( .A(mem[123]), .Y(n3822) );
  INVX1 U3291 ( .A(mem[75]), .Y(n3870) );
  INVX1 U3292 ( .A(mem[508]), .Y(n3437) );
  INVX1 U3293 ( .A(mem[460]), .Y(n3485) );
  INVX1 U3294 ( .A(mem[380]), .Y(n3565) );
  INVX1 U3295 ( .A(mem[332]), .Y(n3613) );
  INVX1 U3296 ( .A(mem[124]), .Y(n3821) );
  INVX1 U3297 ( .A(mem[76]), .Y(n3869) );
  INVX1 U3298 ( .A(mem[509]), .Y(n3436) );
  INVX1 U3299 ( .A(mem[461]), .Y(n3484) );
  INVX1 U3300 ( .A(mem[381]), .Y(n3564) );
  INVX1 U3301 ( .A(mem[333]), .Y(n3612) );
  INVX1 U3302 ( .A(mem[125]), .Y(n3820) );
  INVX1 U3303 ( .A(mem[77]), .Y(n3868) );
  INVX1 U3304 ( .A(mem[510]), .Y(n3435) );
  INVX1 U3305 ( .A(mem[462]), .Y(n3483) );
  INVX1 U3306 ( .A(mem[382]), .Y(n3563) );
  INVX1 U3307 ( .A(mem[334]), .Y(n3611) );
  INVX1 U3308 ( .A(mem[126]), .Y(n3819) );
  INVX1 U3309 ( .A(mem[78]), .Y(n3867) );
  INVX1 U3310 ( .A(mem[511]), .Y(n3434) );
  INVX1 U3311 ( .A(mem[463]), .Y(n3482) );
  INVX1 U3312 ( .A(mem[383]), .Y(n3562) );
  INVX1 U3313 ( .A(mem[335]), .Y(n3610) );
  INVX1 U3314 ( .A(mem[127]), .Y(n3818) );
  INVX1 U3315 ( .A(mem[79]), .Y(n3866) );
  INVX1 U3316 ( .A(mem[240]), .Y(n3705) );
  INVX1 U3317 ( .A(mem[192]), .Y(n3753) );
  INVX1 U3318 ( .A(mem[241]), .Y(n3704) );
  INVX1 U3319 ( .A(mem[193]), .Y(n3752) );
  INVX1 U3320 ( .A(mem[242]), .Y(n3703) );
  INVX1 U3321 ( .A(mem[194]), .Y(n3751) );
  INVX1 U3322 ( .A(mem[243]), .Y(n3702) );
  INVX1 U3323 ( .A(mem[195]), .Y(n3750) );
  INVX1 U3324 ( .A(mem[244]), .Y(n3701) );
  INVX1 U3325 ( .A(mem[196]), .Y(n3749) );
  INVX1 U3326 ( .A(mem[245]), .Y(n3700) );
  INVX1 U3327 ( .A(mem[197]), .Y(n3748) );
  INVX1 U3328 ( .A(mem[246]), .Y(n3699) );
  INVX1 U3329 ( .A(mem[198]), .Y(n3747) );
  INVX1 U3330 ( .A(mem[247]), .Y(n3698) );
  INVX1 U3331 ( .A(mem[199]), .Y(n3746) );
  INVX1 U3332 ( .A(mem[248]), .Y(n3697) );
  INVX1 U3333 ( .A(mem[200]), .Y(n3745) );
  INVX1 U3334 ( .A(mem[249]), .Y(n3696) );
  INVX1 U3335 ( .A(mem[201]), .Y(n3744) );
  INVX1 U3336 ( .A(mem[250]), .Y(n3695) );
  INVX1 U3337 ( .A(mem[202]), .Y(n3743) );
  INVX1 U3338 ( .A(mem[251]), .Y(n3694) );
  INVX1 U3339 ( .A(mem[203]), .Y(n3742) );
  INVX1 U3340 ( .A(mem[252]), .Y(n3693) );
  INVX1 U3341 ( .A(mem[204]), .Y(n3741) );
  INVX1 U3342 ( .A(mem[253]), .Y(n3692) );
  INVX1 U3343 ( .A(mem[205]), .Y(n3740) );
  INVX1 U3344 ( .A(mem[254]), .Y(n3691) );
  INVX1 U3345 ( .A(mem[206]), .Y(n3739) );
  INVX1 U3346 ( .A(mem[255]), .Y(n3690) );
  INVX1 U3347 ( .A(mem[207]), .Y(n3738) );
endmodule


module FIFO_DEPTH_P25_WIDTH33 ( clk, reset, data_in, put, get, data_out, 
        empty_bar, full_bar, fillcount );
  input [32:0] data_in;
  output [32:0] data_out;
  output [5:0] fillcount;
  input clk, reset, put, get;
  output empty_bar, full_bar;
  wire   n12, n13, n14, n15, n16, n4624, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
         n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
         n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
         n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
         n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
         n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
         n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
         n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
         n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
         n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
         n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
         n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
         n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
         n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
         n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
         n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
         n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
         n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
         n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
         n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
         n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
         n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
         n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
         n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
         n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
         n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
         n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
         n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
         n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
         n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
         n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
         n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
         n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
         n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
         n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
         n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
         n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917;
  wire   [4:0] wr_ptr;
  wire   [1055:0] mem;
  assign full_bar = 1'b1;

  DFFPOSX1 wr_ptr_reg_0_ ( .D(n2603), .CLK(clk), .Q(wr_ptr[0]) );
  DFFPOSX1 rd_ptr_reg_4_ ( .D(n4626), .CLK(clk), .Q(n16) );
  DFFPOSX1 rd_ptr_reg_0_ ( .D(n2601), .CLK(clk), .Q(n12) );
  DFFPOSX1 rd_ptr_reg_1_ ( .D(n2600), .CLK(clk), .Q(n13) );
  DFFPOSX1 rd_ptr_reg_2_ ( .D(n2599), .CLK(clk), .Q(n14) );
  DFFPOSX1 rd_ptr_reg_3_ ( .D(n2598), .CLK(clk), .Q(n15) );
  DFFPOSX1 wr_ptr_reg_4_ ( .D(n2597), .CLK(clk), .Q(wr_ptr[4]) );
  DFFPOSX1 wr_ptr_reg_1_ ( .D(n2596), .CLK(clk), .Q(wr_ptr[1]) );
  DFFPOSX1 wr_ptr_reg_2_ ( .D(n2595), .CLK(clk), .Q(wr_ptr[2]) );
  DFFPOSX1 wr_ptr_reg_3_ ( .D(n2594), .CLK(clk), .Q(wr_ptr[3]) );
  DFFPOSX1 data_out_reg_32_ ( .D(n4643), .CLK(clk), .Q(data_out[32]) );
  DFFPOSX1 data_out_reg_31_ ( .D(n4659), .CLK(clk), .Q(data_out[31]) );
  DFFPOSX1 data_out_reg_30_ ( .D(n4642), .CLK(clk), .Q(data_out[30]) );
  DFFPOSX1 data_out_reg_29_ ( .D(n4658), .CLK(clk), .Q(data_out[29]) );
  DFFPOSX1 data_out_reg_28_ ( .D(n4641), .CLK(clk), .Q(data_out[28]) );
  DFFPOSX1 data_out_reg_27_ ( .D(n4657), .CLK(clk), .Q(data_out[27]) );
  DFFPOSX1 data_out_reg_26_ ( .D(n4640), .CLK(clk), .Q(data_out[26]) );
  DFFPOSX1 data_out_reg_25_ ( .D(n4656), .CLK(clk), .Q(data_out[25]) );
  DFFPOSX1 data_out_reg_24_ ( .D(n4639), .CLK(clk), .Q(data_out[24]) );
  DFFPOSX1 data_out_reg_23_ ( .D(n4655), .CLK(clk), .Q(data_out[23]) );
  DFFPOSX1 data_out_reg_22_ ( .D(n4654), .CLK(clk), .Q(data_out[22]) );
  DFFPOSX1 data_out_reg_21_ ( .D(n4653), .CLK(clk), .Q(data_out[21]) );
  DFFPOSX1 data_out_reg_20_ ( .D(n4652), .CLK(clk), .Q(data_out[20]) );
  DFFPOSX1 data_out_reg_19_ ( .D(n4651), .CLK(clk), .Q(data_out[19]) );
  DFFPOSX1 data_out_reg_18_ ( .D(n4650), .CLK(clk), .Q(data_out[18]) );
  DFFPOSX1 data_out_reg_17_ ( .D(n4649), .CLK(clk), .Q(data_out[17]) );
  DFFPOSX1 data_out_reg_16_ ( .D(n4648), .CLK(clk), .Q(data_out[16]) );
  DFFPOSX1 data_out_reg_15_ ( .D(n4647), .CLK(clk), .Q(data_out[15]) );
  DFFPOSX1 data_out_reg_14_ ( .D(n4646), .CLK(clk), .Q(data_out[14]) );
  DFFPOSX1 data_out_reg_13_ ( .D(n4645), .CLK(clk), .Q(data_out[13]) );
  DFFPOSX1 data_out_reg_12_ ( .D(n4644), .CLK(clk), .Q(data_out[12]) );
  DFFPOSX1 data_out_reg_11_ ( .D(n4638), .CLK(clk), .Q(data_out[11]) );
  DFFPOSX1 data_out_reg_10_ ( .D(n4637), .CLK(clk), .Q(data_out[10]) );
  DFFPOSX1 data_out_reg_9_ ( .D(n4636), .CLK(clk), .Q(data_out[9]) );
  DFFPOSX1 data_out_reg_8_ ( .D(n4635), .CLK(clk), .Q(data_out[8]) );
  DFFPOSX1 data_out_reg_7_ ( .D(n4634), .CLK(clk), .Q(data_out[7]) );
  DFFPOSX1 data_out_reg_6_ ( .D(n4633), .CLK(clk), .Q(data_out[6]) );
  DFFPOSX1 data_out_reg_5_ ( .D(n4632), .CLK(clk), .Q(data_out[5]) );
  DFFPOSX1 data_out_reg_4_ ( .D(n4631), .CLK(clk), .Q(data_out[4]) );
  DFFPOSX1 data_out_reg_3_ ( .D(n4630), .CLK(clk), .Q(data_out[3]) );
  DFFPOSX1 data_out_reg_2_ ( .D(n4629), .CLK(clk), .Q(data_out[2]) );
  DFFPOSX1 data_out_reg_1_ ( .D(n4628), .CLK(clk), .Q(data_out[1]) );
  DFFPOSX1 data_out_reg_0_ ( .D(n4627), .CLK(clk), .Q(data_out[0]) );
  DFFPOSX1 mem_reg_31__32_ ( .D(n2593), .CLK(clk), .Q(mem[1055]) );
  DFFPOSX1 mem_reg_31__31_ ( .D(n2592), .CLK(clk), .Q(mem[1054]) );
  DFFPOSX1 mem_reg_31__30_ ( .D(n2591), .CLK(clk), .Q(mem[1053]) );
  DFFPOSX1 mem_reg_31__29_ ( .D(n2590), .CLK(clk), .Q(mem[1052]) );
  DFFPOSX1 mem_reg_31__28_ ( .D(n2589), .CLK(clk), .Q(mem[1051]) );
  DFFPOSX1 mem_reg_31__27_ ( .D(n2588), .CLK(clk), .Q(mem[1050]) );
  DFFPOSX1 mem_reg_31__26_ ( .D(n2587), .CLK(clk), .Q(mem[1049]) );
  DFFPOSX1 mem_reg_31__25_ ( .D(n2586), .CLK(clk), .Q(mem[1048]) );
  DFFPOSX1 mem_reg_31__24_ ( .D(n2585), .CLK(clk), .Q(mem[1047]) );
  DFFPOSX1 mem_reg_31__23_ ( .D(n2584), .CLK(clk), .Q(mem[1046]) );
  DFFPOSX1 mem_reg_31__22_ ( .D(n2583), .CLK(clk), .Q(mem[1045]) );
  DFFPOSX1 mem_reg_31__21_ ( .D(n2582), .CLK(clk), .Q(mem[1044]) );
  DFFPOSX1 mem_reg_31__20_ ( .D(n2581), .CLK(clk), .Q(mem[1043]) );
  DFFPOSX1 mem_reg_31__19_ ( .D(n2580), .CLK(clk), .Q(mem[1042]) );
  DFFPOSX1 mem_reg_31__18_ ( .D(n2579), .CLK(clk), .Q(mem[1041]) );
  DFFPOSX1 mem_reg_31__17_ ( .D(n2578), .CLK(clk), .Q(mem[1040]) );
  DFFPOSX1 mem_reg_31__16_ ( .D(n2577), .CLK(clk), .Q(mem[1039]) );
  DFFPOSX1 mem_reg_31__15_ ( .D(n2576), .CLK(clk), .Q(mem[1038]) );
  DFFPOSX1 mem_reg_31__14_ ( .D(n2575), .CLK(clk), .Q(mem[1037]) );
  DFFPOSX1 mem_reg_31__13_ ( .D(n2574), .CLK(clk), .Q(mem[1036]) );
  DFFPOSX1 mem_reg_31__12_ ( .D(n2573), .CLK(clk), .Q(mem[1035]) );
  DFFPOSX1 mem_reg_31__11_ ( .D(n2572), .CLK(clk), .Q(mem[1034]) );
  DFFPOSX1 mem_reg_31__10_ ( .D(n2571), .CLK(clk), .Q(mem[1033]) );
  DFFPOSX1 mem_reg_31__9_ ( .D(n2570), .CLK(clk), .Q(mem[1032]) );
  DFFPOSX1 mem_reg_31__8_ ( .D(n2569), .CLK(clk), .Q(mem[1031]) );
  DFFPOSX1 mem_reg_31__7_ ( .D(n2568), .CLK(clk), .Q(mem[1030]) );
  DFFPOSX1 mem_reg_31__6_ ( .D(n2567), .CLK(clk), .Q(mem[1029]) );
  DFFPOSX1 mem_reg_31__5_ ( .D(n2566), .CLK(clk), .Q(mem[1028]) );
  DFFPOSX1 mem_reg_31__4_ ( .D(n2565), .CLK(clk), .Q(mem[1027]) );
  DFFPOSX1 mem_reg_31__3_ ( .D(n2564), .CLK(clk), .Q(mem[1026]) );
  DFFPOSX1 mem_reg_31__2_ ( .D(n2563), .CLK(clk), .Q(mem[1025]) );
  DFFPOSX1 mem_reg_31__1_ ( .D(n2562), .CLK(clk), .Q(mem[1024]) );
  DFFPOSX1 mem_reg_31__0_ ( .D(n2561), .CLK(clk), .Q(mem[1023]) );
  DFFPOSX1 mem_reg_30__32_ ( .D(n2560), .CLK(clk), .Q(mem[1022]) );
  DFFPOSX1 mem_reg_30__31_ ( .D(n2559), .CLK(clk), .Q(mem[1021]) );
  DFFPOSX1 mem_reg_30__30_ ( .D(n2558), .CLK(clk), .Q(mem[1020]) );
  DFFPOSX1 mem_reg_30__29_ ( .D(n2557), .CLK(clk), .Q(mem[1019]) );
  DFFPOSX1 mem_reg_30__28_ ( .D(n2556), .CLK(clk), .Q(mem[1018]) );
  DFFPOSX1 mem_reg_30__27_ ( .D(n2555), .CLK(clk), .Q(mem[1017]) );
  DFFPOSX1 mem_reg_30__26_ ( .D(n2554), .CLK(clk), .Q(mem[1016]) );
  DFFPOSX1 mem_reg_30__25_ ( .D(n2553), .CLK(clk), .Q(mem[1015]) );
  DFFPOSX1 mem_reg_30__24_ ( .D(n2552), .CLK(clk), .Q(mem[1014]) );
  DFFPOSX1 mem_reg_30__23_ ( .D(n2551), .CLK(clk), .Q(mem[1013]) );
  DFFPOSX1 mem_reg_30__22_ ( .D(n2550), .CLK(clk), .Q(mem[1012]) );
  DFFPOSX1 mem_reg_30__21_ ( .D(n2549), .CLK(clk), .Q(mem[1011]) );
  DFFPOSX1 mem_reg_30__20_ ( .D(n2548), .CLK(clk), .Q(mem[1010]) );
  DFFPOSX1 mem_reg_30__19_ ( .D(n2547), .CLK(clk), .Q(mem[1009]) );
  DFFPOSX1 mem_reg_30__18_ ( .D(n2546), .CLK(clk), .Q(mem[1008]) );
  DFFPOSX1 mem_reg_30__17_ ( .D(n2545), .CLK(clk), .Q(mem[1007]) );
  DFFPOSX1 mem_reg_30__16_ ( .D(n2544), .CLK(clk), .Q(mem[1006]) );
  DFFPOSX1 mem_reg_30__15_ ( .D(n2543), .CLK(clk), .Q(mem[1005]) );
  DFFPOSX1 mem_reg_30__14_ ( .D(n2542), .CLK(clk), .Q(mem[1004]) );
  DFFPOSX1 mem_reg_30__13_ ( .D(n2541), .CLK(clk), .Q(mem[1003]) );
  DFFPOSX1 mem_reg_30__12_ ( .D(n2540), .CLK(clk), .Q(mem[1002]) );
  DFFPOSX1 mem_reg_30__11_ ( .D(n2539), .CLK(clk), .Q(mem[1001]) );
  DFFPOSX1 mem_reg_30__10_ ( .D(n2538), .CLK(clk), .Q(mem[1000]) );
  DFFPOSX1 mem_reg_30__9_ ( .D(n2537), .CLK(clk), .Q(mem[999]) );
  DFFPOSX1 mem_reg_30__8_ ( .D(n2536), .CLK(clk), .Q(mem[998]) );
  DFFPOSX1 mem_reg_30__7_ ( .D(n2535), .CLK(clk), .Q(mem[997]) );
  DFFPOSX1 mem_reg_30__6_ ( .D(n2534), .CLK(clk), .Q(mem[996]) );
  DFFPOSX1 mem_reg_30__5_ ( .D(n2533), .CLK(clk), .Q(mem[995]) );
  DFFPOSX1 mem_reg_30__4_ ( .D(n2532), .CLK(clk), .Q(mem[994]) );
  DFFPOSX1 mem_reg_30__3_ ( .D(n2531), .CLK(clk), .Q(mem[993]) );
  DFFPOSX1 mem_reg_30__2_ ( .D(n2530), .CLK(clk), .Q(mem[992]) );
  DFFPOSX1 mem_reg_30__1_ ( .D(n2529), .CLK(clk), .Q(mem[991]) );
  DFFPOSX1 mem_reg_30__0_ ( .D(n2528), .CLK(clk), .Q(mem[990]) );
  DFFPOSX1 mem_reg_29__32_ ( .D(n2527), .CLK(clk), .Q(mem[989]) );
  DFFPOSX1 mem_reg_29__31_ ( .D(n2526), .CLK(clk), .Q(mem[988]) );
  DFFPOSX1 mem_reg_29__30_ ( .D(n2525), .CLK(clk), .Q(mem[987]) );
  DFFPOSX1 mem_reg_29__29_ ( .D(n2524), .CLK(clk), .Q(mem[986]) );
  DFFPOSX1 mem_reg_29__28_ ( .D(n2523), .CLK(clk), .Q(mem[985]) );
  DFFPOSX1 mem_reg_29__27_ ( .D(n2522), .CLK(clk), .Q(mem[984]) );
  DFFPOSX1 mem_reg_29__26_ ( .D(n2521), .CLK(clk), .Q(mem[983]) );
  DFFPOSX1 mem_reg_29__25_ ( .D(n2520), .CLK(clk), .Q(mem[982]) );
  DFFPOSX1 mem_reg_29__24_ ( .D(n2519), .CLK(clk), .Q(mem[981]) );
  DFFPOSX1 mem_reg_29__23_ ( .D(n2518), .CLK(clk), .Q(mem[980]) );
  DFFPOSX1 mem_reg_29__22_ ( .D(n2517), .CLK(clk), .Q(mem[979]) );
  DFFPOSX1 mem_reg_29__21_ ( .D(n2516), .CLK(clk), .Q(mem[978]) );
  DFFPOSX1 mem_reg_29__20_ ( .D(n2515), .CLK(clk), .Q(mem[977]) );
  DFFPOSX1 mem_reg_29__19_ ( .D(n2514), .CLK(clk), .Q(mem[976]) );
  DFFPOSX1 mem_reg_29__18_ ( .D(n2513), .CLK(clk), .Q(mem[975]) );
  DFFPOSX1 mem_reg_29__17_ ( .D(n2512), .CLK(clk), .Q(mem[974]) );
  DFFPOSX1 mem_reg_29__16_ ( .D(n2511), .CLK(clk), .Q(mem[973]) );
  DFFPOSX1 mem_reg_29__15_ ( .D(n2510), .CLK(clk), .Q(mem[972]) );
  DFFPOSX1 mem_reg_29__14_ ( .D(n2509), .CLK(clk), .Q(mem[971]) );
  DFFPOSX1 mem_reg_29__13_ ( .D(n2508), .CLK(clk), .Q(mem[970]) );
  DFFPOSX1 mem_reg_29__12_ ( .D(n2507), .CLK(clk), .Q(mem[969]) );
  DFFPOSX1 mem_reg_29__11_ ( .D(n2506), .CLK(clk), .Q(mem[968]) );
  DFFPOSX1 mem_reg_29__10_ ( .D(n2505), .CLK(clk), .Q(mem[967]) );
  DFFPOSX1 mem_reg_29__9_ ( .D(n2504), .CLK(clk), .Q(mem[966]) );
  DFFPOSX1 mem_reg_29__8_ ( .D(n2503), .CLK(clk), .Q(mem[965]) );
  DFFPOSX1 mem_reg_29__7_ ( .D(n2502), .CLK(clk), .Q(mem[964]) );
  DFFPOSX1 mem_reg_29__6_ ( .D(n2501), .CLK(clk), .Q(mem[963]) );
  DFFPOSX1 mem_reg_29__5_ ( .D(n2500), .CLK(clk), .Q(mem[962]) );
  DFFPOSX1 mem_reg_29__4_ ( .D(n2499), .CLK(clk), .Q(mem[961]) );
  DFFPOSX1 mem_reg_29__3_ ( .D(n2498), .CLK(clk), .Q(mem[960]) );
  DFFPOSX1 mem_reg_29__2_ ( .D(n2497), .CLK(clk), .Q(mem[959]) );
  DFFPOSX1 mem_reg_29__1_ ( .D(n2496), .CLK(clk), .Q(mem[958]) );
  DFFPOSX1 mem_reg_29__0_ ( .D(n2495), .CLK(clk), .Q(mem[957]) );
  DFFPOSX1 mem_reg_28__32_ ( .D(n2494), .CLK(clk), .Q(mem[956]) );
  DFFPOSX1 mem_reg_28__31_ ( .D(n2493), .CLK(clk), .Q(mem[955]) );
  DFFPOSX1 mem_reg_28__30_ ( .D(n2492), .CLK(clk), .Q(mem[954]) );
  DFFPOSX1 mem_reg_28__29_ ( .D(n2491), .CLK(clk), .Q(mem[953]) );
  DFFPOSX1 mem_reg_28__28_ ( .D(n2490), .CLK(clk), .Q(mem[952]) );
  DFFPOSX1 mem_reg_28__27_ ( .D(n2489), .CLK(clk), .Q(mem[951]) );
  DFFPOSX1 mem_reg_28__26_ ( .D(n2488), .CLK(clk), .Q(mem[950]) );
  DFFPOSX1 mem_reg_28__25_ ( .D(n2487), .CLK(clk), .Q(mem[949]) );
  DFFPOSX1 mem_reg_28__24_ ( .D(n2486), .CLK(clk), .Q(mem[948]) );
  DFFPOSX1 mem_reg_28__23_ ( .D(n2485), .CLK(clk), .Q(mem[947]) );
  DFFPOSX1 mem_reg_28__22_ ( .D(n2484), .CLK(clk), .Q(mem[946]) );
  DFFPOSX1 mem_reg_28__21_ ( .D(n2483), .CLK(clk), .Q(mem[945]) );
  DFFPOSX1 mem_reg_28__20_ ( .D(n2482), .CLK(clk), .Q(mem[944]) );
  DFFPOSX1 mem_reg_28__19_ ( .D(n2481), .CLK(clk), .Q(mem[943]) );
  DFFPOSX1 mem_reg_28__18_ ( .D(n2480), .CLK(clk), .Q(mem[942]) );
  DFFPOSX1 mem_reg_28__17_ ( .D(n2479), .CLK(clk), .Q(mem[941]) );
  DFFPOSX1 mem_reg_28__16_ ( .D(n2478), .CLK(clk), .Q(mem[940]) );
  DFFPOSX1 mem_reg_28__15_ ( .D(n2477), .CLK(clk), .Q(mem[939]) );
  DFFPOSX1 mem_reg_28__14_ ( .D(n2476), .CLK(clk), .Q(mem[938]) );
  DFFPOSX1 mem_reg_28__13_ ( .D(n2475), .CLK(clk), .Q(mem[937]) );
  DFFPOSX1 mem_reg_28__12_ ( .D(n2474), .CLK(clk), .Q(mem[936]) );
  DFFPOSX1 mem_reg_28__11_ ( .D(n2473), .CLK(clk), .Q(mem[935]) );
  DFFPOSX1 mem_reg_28__10_ ( .D(n2472), .CLK(clk), .Q(mem[934]) );
  DFFPOSX1 mem_reg_28__9_ ( .D(n2471), .CLK(clk), .Q(mem[933]) );
  DFFPOSX1 mem_reg_28__8_ ( .D(n2470), .CLK(clk), .Q(mem[932]) );
  DFFPOSX1 mem_reg_28__7_ ( .D(n2469), .CLK(clk), .Q(mem[931]) );
  DFFPOSX1 mem_reg_28__6_ ( .D(n2468), .CLK(clk), .Q(mem[930]) );
  DFFPOSX1 mem_reg_28__5_ ( .D(n2467), .CLK(clk), .Q(mem[929]) );
  DFFPOSX1 mem_reg_28__4_ ( .D(n2466), .CLK(clk), .Q(mem[928]) );
  DFFPOSX1 mem_reg_28__3_ ( .D(n2465), .CLK(clk), .Q(mem[927]) );
  DFFPOSX1 mem_reg_28__2_ ( .D(n2464), .CLK(clk), .Q(mem[926]) );
  DFFPOSX1 mem_reg_28__1_ ( .D(n2463), .CLK(clk), .Q(mem[925]) );
  DFFPOSX1 mem_reg_28__0_ ( .D(n2462), .CLK(clk), .Q(mem[924]) );
  DFFPOSX1 mem_reg_27__32_ ( .D(n2461), .CLK(clk), .Q(mem[923]) );
  DFFPOSX1 mem_reg_27__31_ ( .D(n2460), .CLK(clk), .Q(mem[922]) );
  DFFPOSX1 mem_reg_27__30_ ( .D(n2459), .CLK(clk), .Q(mem[921]) );
  DFFPOSX1 mem_reg_27__29_ ( .D(n2458), .CLK(clk), .Q(mem[920]) );
  DFFPOSX1 mem_reg_27__28_ ( .D(n2457), .CLK(clk), .Q(mem[919]) );
  DFFPOSX1 mem_reg_27__27_ ( .D(n2456), .CLK(clk), .Q(mem[918]) );
  DFFPOSX1 mem_reg_27__26_ ( .D(n2455), .CLK(clk), .Q(mem[917]) );
  DFFPOSX1 mem_reg_27__25_ ( .D(n2454), .CLK(clk), .Q(mem[916]) );
  DFFPOSX1 mem_reg_27__24_ ( .D(n2453), .CLK(clk), .Q(mem[915]) );
  DFFPOSX1 mem_reg_27__23_ ( .D(n2452), .CLK(clk), .Q(mem[914]) );
  DFFPOSX1 mem_reg_27__22_ ( .D(n2451), .CLK(clk), .Q(mem[913]) );
  DFFPOSX1 mem_reg_27__21_ ( .D(n2450), .CLK(clk), .Q(mem[912]) );
  DFFPOSX1 mem_reg_27__20_ ( .D(n2449), .CLK(clk), .Q(mem[911]) );
  DFFPOSX1 mem_reg_27__19_ ( .D(n2448), .CLK(clk), .Q(mem[910]) );
  DFFPOSX1 mem_reg_27__18_ ( .D(n2447), .CLK(clk), .Q(mem[909]) );
  DFFPOSX1 mem_reg_27__17_ ( .D(n2446), .CLK(clk), .Q(mem[908]) );
  DFFPOSX1 mem_reg_27__16_ ( .D(n2445), .CLK(clk), .Q(mem[907]) );
  DFFPOSX1 mem_reg_27__15_ ( .D(n2444), .CLK(clk), .Q(mem[906]) );
  DFFPOSX1 mem_reg_27__14_ ( .D(n2443), .CLK(clk), .Q(mem[905]) );
  DFFPOSX1 mem_reg_27__13_ ( .D(n2442), .CLK(clk), .Q(mem[904]) );
  DFFPOSX1 mem_reg_27__12_ ( .D(n2441), .CLK(clk), .Q(mem[903]) );
  DFFPOSX1 mem_reg_27__11_ ( .D(n2440), .CLK(clk), .Q(mem[902]) );
  DFFPOSX1 mem_reg_27__10_ ( .D(n2439), .CLK(clk), .Q(mem[901]) );
  DFFPOSX1 mem_reg_27__9_ ( .D(n2438), .CLK(clk), .Q(mem[900]) );
  DFFPOSX1 mem_reg_27__8_ ( .D(n2437), .CLK(clk), .Q(mem[899]) );
  DFFPOSX1 mem_reg_27__7_ ( .D(n2436), .CLK(clk), .Q(mem[898]) );
  DFFPOSX1 mem_reg_27__6_ ( .D(n2435), .CLK(clk), .Q(mem[897]) );
  DFFPOSX1 mem_reg_27__5_ ( .D(n2434), .CLK(clk), .Q(mem[896]) );
  DFFPOSX1 mem_reg_27__4_ ( .D(n2433), .CLK(clk), .Q(mem[895]) );
  DFFPOSX1 mem_reg_27__3_ ( .D(n2432), .CLK(clk), .Q(mem[894]) );
  DFFPOSX1 mem_reg_27__2_ ( .D(n2431), .CLK(clk), .Q(mem[893]) );
  DFFPOSX1 mem_reg_27__1_ ( .D(n2430), .CLK(clk), .Q(mem[892]) );
  DFFPOSX1 mem_reg_27__0_ ( .D(n2429), .CLK(clk), .Q(mem[891]) );
  DFFPOSX1 mem_reg_26__32_ ( .D(n2428), .CLK(clk), .Q(mem[890]) );
  DFFPOSX1 mem_reg_26__31_ ( .D(n2427), .CLK(clk), .Q(mem[889]) );
  DFFPOSX1 mem_reg_26__30_ ( .D(n2426), .CLK(clk), .Q(mem[888]) );
  DFFPOSX1 mem_reg_26__29_ ( .D(n2425), .CLK(clk), .Q(mem[887]) );
  DFFPOSX1 mem_reg_26__28_ ( .D(n2424), .CLK(clk), .Q(mem[886]) );
  DFFPOSX1 mem_reg_26__27_ ( .D(n2423), .CLK(clk), .Q(mem[885]) );
  DFFPOSX1 mem_reg_26__26_ ( .D(n2422), .CLK(clk), .Q(mem[884]) );
  DFFPOSX1 mem_reg_26__25_ ( .D(n2421), .CLK(clk), .Q(mem[883]) );
  DFFPOSX1 mem_reg_26__24_ ( .D(n2420), .CLK(clk), .Q(mem[882]) );
  DFFPOSX1 mem_reg_26__23_ ( .D(n2419), .CLK(clk), .Q(mem[881]) );
  DFFPOSX1 mem_reg_26__22_ ( .D(n2418), .CLK(clk), .Q(mem[880]) );
  DFFPOSX1 mem_reg_26__21_ ( .D(n2417), .CLK(clk), .Q(mem[879]) );
  DFFPOSX1 mem_reg_26__20_ ( .D(n2416), .CLK(clk), .Q(mem[878]) );
  DFFPOSX1 mem_reg_26__19_ ( .D(n2415), .CLK(clk), .Q(mem[877]) );
  DFFPOSX1 mem_reg_26__18_ ( .D(n2414), .CLK(clk), .Q(mem[876]) );
  DFFPOSX1 mem_reg_26__17_ ( .D(n2413), .CLK(clk), .Q(mem[875]) );
  DFFPOSX1 mem_reg_26__16_ ( .D(n2412), .CLK(clk), .Q(mem[874]) );
  DFFPOSX1 mem_reg_26__15_ ( .D(n2411), .CLK(clk), .Q(mem[873]) );
  DFFPOSX1 mem_reg_26__14_ ( .D(n2410), .CLK(clk), .Q(mem[872]) );
  DFFPOSX1 mem_reg_26__13_ ( .D(n2409), .CLK(clk), .Q(mem[871]) );
  DFFPOSX1 mem_reg_26__12_ ( .D(n2408), .CLK(clk), .Q(mem[870]) );
  DFFPOSX1 mem_reg_26__11_ ( .D(n2407), .CLK(clk), .Q(mem[869]) );
  DFFPOSX1 mem_reg_26__10_ ( .D(n2406), .CLK(clk), .Q(mem[868]) );
  DFFPOSX1 mem_reg_26__9_ ( .D(n2405), .CLK(clk), .Q(mem[867]) );
  DFFPOSX1 mem_reg_26__8_ ( .D(n2404), .CLK(clk), .Q(mem[866]) );
  DFFPOSX1 mem_reg_26__7_ ( .D(n2403), .CLK(clk), .Q(mem[865]) );
  DFFPOSX1 mem_reg_26__6_ ( .D(n2402), .CLK(clk), .Q(mem[864]) );
  DFFPOSX1 mem_reg_26__5_ ( .D(n2401), .CLK(clk), .Q(mem[863]) );
  DFFPOSX1 mem_reg_26__4_ ( .D(n2400), .CLK(clk), .Q(mem[862]) );
  DFFPOSX1 mem_reg_26__3_ ( .D(n2399), .CLK(clk), .Q(mem[861]) );
  DFFPOSX1 mem_reg_26__2_ ( .D(n2398), .CLK(clk), .Q(mem[860]) );
  DFFPOSX1 mem_reg_26__1_ ( .D(n2397), .CLK(clk), .Q(mem[859]) );
  DFFPOSX1 mem_reg_26__0_ ( .D(n2396), .CLK(clk), .Q(mem[858]) );
  DFFPOSX1 mem_reg_25__32_ ( .D(n2395), .CLK(clk), .Q(mem[857]) );
  DFFPOSX1 mem_reg_25__31_ ( .D(n2394), .CLK(clk), .Q(mem[856]) );
  DFFPOSX1 mem_reg_25__30_ ( .D(n2393), .CLK(clk), .Q(mem[855]) );
  DFFPOSX1 mem_reg_25__29_ ( .D(n2392), .CLK(clk), .Q(mem[854]) );
  DFFPOSX1 mem_reg_25__28_ ( .D(n2391), .CLK(clk), .Q(mem[853]) );
  DFFPOSX1 mem_reg_25__27_ ( .D(n2390), .CLK(clk), .Q(mem[852]) );
  DFFPOSX1 mem_reg_25__26_ ( .D(n2389), .CLK(clk), .Q(mem[851]) );
  DFFPOSX1 mem_reg_25__25_ ( .D(n2388), .CLK(clk), .Q(mem[850]) );
  DFFPOSX1 mem_reg_25__24_ ( .D(n2387), .CLK(clk), .Q(mem[849]) );
  DFFPOSX1 mem_reg_25__23_ ( .D(n2386), .CLK(clk), .Q(mem[848]) );
  DFFPOSX1 mem_reg_25__22_ ( .D(n2385), .CLK(clk), .Q(mem[847]) );
  DFFPOSX1 mem_reg_25__21_ ( .D(n2384), .CLK(clk), .Q(mem[846]) );
  DFFPOSX1 mem_reg_25__20_ ( .D(n2383), .CLK(clk), .Q(mem[845]) );
  DFFPOSX1 mem_reg_25__19_ ( .D(n2382), .CLK(clk), .Q(mem[844]) );
  DFFPOSX1 mem_reg_25__18_ ( .D(n2381), .CLK(clk), .Q(mem[843]) );
  DFFPOSX1 mem_reg_25__17_ ( .D(n2380), .CLK(clk), .Q(mem[842]) );
  DFFPOSX1 mem_reg_25__16_ ( .D(n2379), .CLK(clk), .Q(mem[841]) );
  DFFPOSX1 mem_reg_25__15_ ( .D(n2378), .CLK(clk), .Q(mem[840]) );
  DFFPOSX1 mem_reg_25__14_ ( .D(n2377), .CLK(clk), .Q(mem[839]) );
  DFFPOSX1 mem_reg_25__13_ ( .D(n2376), .CLK(clk), .Q(mem[838]) );
  DFFPOSX1 mem_reg_25__12_ ( .D(n2375), .CLK(clk), .Q(mem[837]) );
  DFFPOSX1 mem_reg_25__11_ ( .D(n2374), .CLK(clk), .Q(mem[836]) );
  DFFPOSX1 mem_reg_25__10_ ( .D(n2373), .CLK(clk), .Q(mem[835]) );
  DFFPOSX1 mem_reg_25__9_ ( .D(n2372), .CLK(clk), .Q(mem[834]) );
  DFFPOSX1 mem_reg_25__8_ ( .D(n2371), .CLK(clk), .Q(mem[833]) );
  DFFPOSX1 mem_reg_25__7_ ( .D(n2370), .CLK(clk), .Q(mem[832]) );
  DFFPOSX1 mem_reg_25__6_ ( .D(n2369), .CLK(clk), .Q(mem[831]) );
  DFFPOSX1 mem_reg_25__5_ ( .D(n2368), .CLK(clk), .Q(mem[830]) );
  DFFPOSX1 mem_reg_25__4_ ( .D(n2367), .CLK(clk), .Q(mem[829]) );
  DFFPOSX1 mem_reg_25__3_ ( .D(n2366), .CLK(clk), .Q(mem[828]) );
  DFFPOSX1 mem_reg_25__2_ ( .D(n2365), .CLK(clk), .Q(mem[827]) );
  DFFPOSX1 mem_reg_25__1_ ( .D(n2364), .CLK(clk), .Q(mem[826]) );
  DFFPOSX1 mem_reg_25__0_ ( .D(n2363), .CLK(clk), .Q(mem[825]) );
  DFFPOSX1 mem_reg_24__32_ ( .D(n2362), .CLK(clk), .Q(mem[824]) );
  DFFPOSX1 mem_reg_24__31_ ( .D(n2361), .CLK(clk), .Q(mem[823]) );
  DFFPOSX1 mem_reg_24__30_ ( .D(n2360), .CLK(clk), .Q(mem[822]) );
  DFFPOSX1 mem_reg_24__29_ ( .D(n2359), .CLK(clk), .Q(mem[821]) );
  DFFPOSX1 mem_reg_24__28_ ( .D(n2358), .CLK(clk), .Q(mem[820]) );
  DFFPOSX1 mem_reg_24__27_ ( .D(n2357), .CLK(clk), .Q(mem[819]) );
  DFFPOSX1 mem_reg_24__26_ ( .D(n2356), .CLK(clk), .Q(mem[818]) );
  DFFPOSX1 mem_reg_24__25_ ( .D(n2355), .CLK(clk), .Q(mem[817]) );
  DFFPOSX1 mem_reg_24__24_ ( .D(n2354), .CLK(clk), .Q(mem[816]) );
  DFFPOSX1 mem_reg_24__23_ ( .D(n2353), .CLK(clk), .Q(mem[815]) );
  DFFPOSX1 mem_reg_24__22_ ( .D(n2352), .CLK(clk), .Q(mem[814]) );
  DFFPOSX1 mem_reg_24__21_ ( .D(n2351), .CLK(clk), .Q(mem[813]) );
  DFFPOSX1 mem_reg_24__20_ ( .D(n2350), .CLK(clk), .Q(mem[812]) );
  DFFPOSX1 mem_reg_24__19_ ( .D(n2349), .CLK(clk), .Q(mem[811]) );
  DFFPOSX1 mem_reg_24__18_ ( .D(n2348), .CLK(clk), .Q(mem[810]) );
  DFFPOSX1 mem_reg_24__17_ ( .D(n2347), .CLK(clk), .Q(mem[809]) );
  DFFPOSX1 mem_reg_24__16_ ( .D(n2346), .CLK(clk), .Q(mem[808]) );
  DFFPOSX1 mem_reg_24__15_ ( .D(n2345), .CLK(clk), .Q(mem[807]) );
  DFFPOSX1 mem_reg_24__14_ ( .D(n2344), .CLK(clk), .Q(mem[806]) );
  DFFPOSX1 mem_reg_24__13_ ( .D(n2343), .CLK(clk), .Q(mem[805]) );
  DFFPOSX1 mem_reg_24__12_ ( .D(n2342), .CLK(clk), .Q(mem[804]) );
  DFFPOSX1 mem_reg_24__11_ ( .D(n2341), .CLK(clk), .Q(mem[803]) );
  DFFPOSX1 mem_reg_24__10_ ( .D(n2340), .CLK(clk), .Q(mem[802]) );
  DFFPOSX1 mem_reg_24__9_ ( .D(n2339), .CLK(clk), .Q(mem[801]) );
  DFFPOSX1 mem_reg_24__8_ ( .D(n2338), .CLK(clk), .Q(mem[800]) );
  DFFPOSX1 mem_reg_24__7_ ( .D(n2337), .CLK(clk), .Q(mem[799]) );
  DFFPOSX1 mem_reg_24__6_ ( .D(n2336), .CLK(clk), .Q(mem[798]) );
  DFFPOSX1 mem_reg_24__5_ ( .D(n2335), .CLK(clk), .Q(mem[797]) );
  DFFPOSX1 mem_reg_24__4_ ( .D(n2334), .CLK(clk), .Q(mem[796]) );
  DFFPOSX1 mem_reg_24__3_ ( .D(n2333), .CLK(clk), .Q(mem[795]) );
  DFFPOSX1 mem_reg_24__2_ ( .D(n2332), .CLK(clk), .Q(mem[794]) );
  DFFPOSX1 mem_reg_24__1_ ( .D(n2331), .CLK(clk), .Q(mem[793]) );
  DFFPOSX1 mem_reg_24__0_ ( .D(n2330), .CLK(clk), .Q(mem[792]) );
  DFFPOSX1 mem_reg_23__32_ ( .D(n2329), .CLK(clk), .Q(mem[791]) );
  DFFPOSX1 mem_reg_23__31_ ( .D(n2328), .CLK(clk), .Q(mem[790]) );
  DFFPOSX1 mem_reg_23__30_ ( .D(n2327), .CLK(clk), .Q(mem[789]) );
  DFFPOSX1 mem_reg_23__29_ ( .D(n2326), .CLK(clk), .Q(mem[788]) );
  DFFPOSX1 mem_reg_23__28_ ( .D(n2325), .CLK(clk), .Q(mem[787]) );
  DFFPOSX1 mem_reg_23__27_ ( .D(n2324), .CLK(clk), .Q(mem[786]) );
  DFFPOSX1 mem_reg_23__26_ ( .D(n2323), .CLK(clk), .Q(mem[785]) );
  DFFPOSX1 mem_reg_23__25_ ( .D(n2322), .CLK(clk), .Q(mem[784]) );
  DFFPOSX1 mem_reg_23__24_ ( .D(n2321), .CLK(clk), .Q(mem[783]) );
  DFFPOSX1 mem_reg_23__23_ ( .D(n2320), .CLK(clk), .Q(mem[782]) );
  DFFPOSX1 mem_reg_23__22_ ( .D(n2319), .CLK(clk), .Q(mem[781]) );
  DFFPOSX1 mem_reg_23__21_ ( .D(n2318), .CLK(clk), .Q(mem[780]) );
  DFFPOSX1 mem_reg_23__20_ ( .D(n2317), .CLK(clk), .Q(mem[779]) );
  DFFPOSX1 mem_reg_23__19_ ( .D(n2316), .CLK(clk), .Q(mem[778]) );
  DFFPOSX1 mem_reg_23__18_ ( .D(n2315), .CLK(clk), .Q(mem[777]) );
  DFFPOSX1 mem_reg_23__17_ ( .D(n2314), .CLK(clk), .Q(mem[776]) );
  DFFPOSX1 mem_reg_23__16_ ( .D(n2313), .CLK(clk), .Q(mem[775]) );
  DFFPOSX1 mem_reg_23__15_ ( .D(n2312), .CLK(clk), .Q(mem[774]) );
  DFFPOSX1 mem_reg_23__14_ ( .D(n2311), .CLK(clk), .Q(mem[773]) );
  DFFPOSX1 mem_reg_23__13_ ( .D(n2310), .CLK(clk), .Q(mem[772]) );
  DFFPOSX1 mem_reg_23__12_ ( .D(n2309), .CLK(clk), .Q(mem[771]) );
  DFFPOSX1 mem_reg_23__11_ ( .D(n2308), .CLK(clk), .Q(mem[770]) );
  DFFPOSX1 mem_reg_23__10_ ( .D(n2307), .CLK(clk), .Q(mem[769]) );
  DFFPOSX1 mem_reg_23__9_ ( .D(n2306), .CLK(clk), .Q(mem[768]) );
  DFFPOSX1 mem_reg_23__8_ ( .D(n2305), .CLK(clk), .Q(mem[767]) );
  DFFPOSX1 mem_reg_23__7_ ( .D(n2304), .CLK(clk), .Q(mem[766]) );
  DFFPOSX1 mem_reg_23__6_ ( .D(n2303), .CLK(clk), .Q(mem[765]) );
  DFFPOSX1 mem_reg_23__5_ ( .D(n2302), .CLK(clk), .Q(mem[764]) );
  DFFPOSX1 mem_reg_23__4_ ( .D(n2301), .CLK(clk), .Q(mem[763]) );
  DFFPOSX1 mem_reg_23__3_ ( .D(n2300), .CLK(clk), .Q(mem[762]) );
  DFFPOSX1 mem_reg_23__2_ ( .D(n2299), .CLK(clk), .Q(mem[761]) );
  DFFPOSX1 mem_reg_23__1_ ( .D(n2298), .CLK(clk), .Q(mem[760]) );
  DFFPOSX1 mem_reg_23__0_ ( .D(n2297), .CLK(clk), .Q(mem[759]) );
  DFFPOSX1 mem_reg_22__32_ ( .D(n2296), .CLK(clk), .Q(mem[758]) );
  DFFPOSX1 mem_reg_22__31_ ( .D(n2295), .CLK(clk), .Q(mem[757]) );
  DFFPOSX1 mem_reg_22__30_ ( .D(n2294), .CLK(clk), .Q(mem[756]) );
  DFFPOSX1 mem_reg_22__29_ ( .D(n2293), .CLK(clk), .Q(mem[755]) );
  DFFPOSX1 mem_reg_22__28_ ( .D(n2292), .CLK(clk), .Q(mem[754]) );
  DFFPOSX1 mem_reg_22__27_ ( .D(n2291), .CLK(clk), .Q(mem[753]) );
  DFFPOSX1 mem_reg_22__26_ ( .D(n2290), .CLK(clk), .Q(mem[752]) );
  DFFPOSX1 mem_reg_22__25_ ( .D(n2289), .CLK(clk), .Q(mem[751]) );
  DFFPOSX1 mem_reg_22__24_ ( .D(n2288), .CLK(clk), .Q(mem[750]) );
  DFFPOSX1 mem_reg_22__23_ ( .D(n2287), .CLK(clk), .Q(mem[749]) );
  DFFPOSX1 mem_reg_22__22_ ( .D(n2286), .CLK(clk), .Q(mem[748]) );
  DFFPOSX1 mem_reg_22__21_ ( .D(n2285), .CLK(clk), .Q(mem[747]) );
  DFFPOSX1 mem_reg_22__20_ ( .D(n2284), .CLK(clk), .Q(mem[746]) );
  DFFPOSX1 mem_reg_22__19_ ( .D(n2283), .CLK(clk), .Q(mem[745]) );
  DFFPOSX1 mem_reg_22__18_ ( .D(n2282), .CLK(clk), .Q(mem[744]) );
  DFFPOSX1 mem_reg_22__17_ ( .D(n2281), .CLK(clk), .Q(mem[743]) );
  DFFPOSX1 mem_reg_22__16_ ( .D(n2280), .CLK(clk), .Q(mem[742]) );
  DFFPOSX1 mem_reg_22__15_ ( .D(n2279), .CLK(clk), .Q(mem[741]) );
  DFFPOSX1 mem_reg_22__14_ ( .D(n2278), .CLK(clk), .Q(mem[740]) );
  DFFPOSX1 mem_reg_22__13_ ( .D(n2277), .CLK(clk), .Q(mem[739]) );
  DFFPOSX1 mem_reg_22__12_ ( .D(n2276), .CLK(clk), .Q(mem[738]) );
  DFFPOSX1 mem_reg_22__11_ ( .D(n2275), .CLK(clk), .Q(mem[737]) );
  DFFPOSX1 mem_reg_22__10_ ( .D(n2274), .CLK(clk), .Q(mem[736]) );
  DFFPOSX1 mem_reg_22__9_ ( .D(n2273), .CLK(clk), .Q(mem[735]) );
  DFFPOSX1 mem_reg_22__8_ ( .D(n2272), .CLK(clk), .Q(mem[734]) );
  DFFPOSX1 mem_reg_22__7_ ( .D(n2271), .CLK(clk), .Q(mem[733]) );
  DFFPOSX1 mem_reg_22__6_ ( .D(n2270), .CLK(clk), .Q(mem[732]) );
  DFFPOSX1 mem_reg_22__5_ ( .D(n2269), .CLK(clk), .Q(mem[731]) );
  DFFPOSX1 mem_reg_22__4_ ( .D(n2268), .CLK(clk), .Q(mem[730]) );
  DFFPOSX1 mem_reg_22__3_ ( .D(n2267), .CLK(clk), .Q(mem[729]) );
  DFFPOSX1 mem_reg_22__2_ ( .D(n2266), .CLK(clk), .Q(mem[728]) );
  DFFPOSX1 mem_reg_22__1_ ( .D(n2265), .CLK(clk), .Q(mem[727]) );
  DFFPOSX1 mem_reg_22__0_ ( .D(n2264), .CLK(clk), .Q(mem[726]) );
  DFFPOSX1 mem_reg_21__32_ ( .D(n2263), .CLK(clk), .Q(mem[725]) );
  DFFPOSX1 mem_reg_21__31_ ( .D(n2262), .CLK(clk), .Q(mem[724]) );
  DFFPOSX1 mem_reg_21__30_ ( .D(n2261), .CLK(clk), .Q(mem[723]) );
  DFFPOSX1 mem_reg_21__29_ ( .D(n2260), .CLK(clk), .Q(mem[722]) );
  DFFPOSX1 mem_reg_21__28_ ( .D(n2259), .CLK(clk), .Q(mem[721]) );
  DFFPOSX1 mem_reg_21__27_ ( .D(n2258), .CLK(clk), .Q(mem[720]) );
  DFFPOSX1 mem_reg_21__26_ ( .D(n2257), .CLK(clk), .Q(mem[719]) );
  DFFPOSX1 mem_reg_21__25_ ( .D(n2256), .CLK(clk), .Q(mem[718]) );
  DFFPOSX1 mem_reg_21__24_ ( .D(n2255), .CLK(clk), .Q(mem[717]) );
  DFFPOSX1 mem_reg_21__23_ ( .D(n2254), .CLK(clk), .Q(mem[716]) );
  DFFPOSX1 mem_reg_21__22_ ( .D(n2253), .CLK(clk), .Q(mem[715]) );
  DFFPOSX1 mem_reg_21__21_ ( .D(n2252), .CLK(clk), .Q(mem[714]) );
  DFFPOSX1 mem_reg_21__20_ ( .D(n2251), .CLK(clk), .Q(mem[713]) );
  DFFPOSX1 mem_reg_21__19_ ( .D(n2250), .CLK(clk), .Q(mem[712]) );
  DFFPOSX1 mem_reg_21__18_ ( .D(n2249), .CLK(clk), .Q(mem[711]) );
  DFFPOSX1 mem_reg_21__17_ ( .D(n2248), .CLK(clk), .Q(mem[710]) );
  DFFPOSX1 mem_reg_21__16_ ( .D(n2247), .CLK(clk), .Q(mem[709]) );
  DFFPOSX1 mem_reg_21__15_ ( .D(n2246), .CLK(clk), .Q(mem[708]) );
  DFFPOSX1 mem_reg_21__14_ ( .D(n2245), .CLK(clk), .Q(mem[707]) );
  DFFPOSX1 mem_reg_21__13_ ( .D(n2244), .CLK(clk), .Q(mem[706]) );
  DFFPOSX1 mem_reg_21__12_ ( .D(n2243), .CLK(clk), .Q(mem[705]) );
  DFFPOSX1 mem_reg_21__11_ ( .D(n2242), .CLK(clk), .Q(mem[704]) );
  DFFPOSX1 mem_reg_21__10_ ( .D(n2241), .CLK(clk), .Q(mem[703]) );
  DFFPOSX1 mem_reg_21__9_ ( .D(n2240), .CLK(clk), .Q(mem[702]) );
  DFFPOSX1 mem_reg_21__8_ ( .D(n2239), .CLK(clk), .Q(mem[701]) );
  DFFPOSX1 mem_reg_21__7_ ( .D(n2238), .CLK(clk), .Q(mem[700]) );
  DFFPOSX1 mem_reg_21__6_ ( .D(n2237), .CLK(clk), .Q(mem[699]) );
  DFFPOSX1 mem_reg_21__5_ ( .D(n2236), .CLK(clk), .Q(mem[698]) );
  DFFPOSX1 mem_reg_21__4_ ( .D(n2235), .CLK(clk), .Q(mem[697]) );
  DFFPOSX1 mem_reg_21__3_ ( .D(n2234), .CLK(clk), .Q(mem[696]) );
  DFFPOSX1 mem_reg_21__2_ ( .D(n2233), .CLK(clk), .Q(mem[695]) );
  DFFPOSX1 mem_reg_21__1_ ( .D(n2232), .CLK(clk), .Q(mem[694]) );
  DFFPOSX1 mem_reg_21__0_ ( .D(n2231), .CLK(clk), .Q(mem[693]) );
  DFFPOSX1 mem_reg_20__32_ ( .D(n2230), .CLK(clk), .Q(mem[692]) );
  DFFPOSX1 mem_reg_20__31_ ( .D(n2229), .CLK(clk), .Q(mem[691]) );
  DFFPOSX1 mem_reg_20__30_ ( .D(n2228), .CLK(clk), .Q(mem[690]) );
  DFFPOSX1 mem_reg_20__29_ ( .D(n2227), .CLK(clk), .Q(mem[689]) );
  DFFPOSX1 mem_reg_20__28_ ( .D(n2226), .CLK(clk), .Q(mem[688]) );
  DFFPOSX1 mem_reg_20__27_ ( .D(n2225), .CLK(clk), .Q(mem[687]) );
  DFFPOSX1 mem_reg_20__26_ ( .D(n2224), .CLK(clk), .Q(mem[686]) );
  DFFPOSX1 mem_reg_20__25_ ( .D(n2223), .CLK(clk), .Q(mem[685]) );
  DFFPOSX1 mem_reg_20__24_ ( .D(n2222), .CLK(clk), .Q(mem[684]) );
  DFFPOSX1 mem_reg_20__23_ ( .D(n2221), .CLK(clk), .Q(mem[683]) );
  DFFPOSX1 mem_reg_20__22_ ( .D(n2220), .CLK(clk), .Q(mem[682]) );
  DFFPOSX1 mem_reg_20__21_ ( .D(n2219), .CLK(clk), .Q(mem[681]) );
  DFFPOSX1 mem_reg_20__20_ ( .D(n2218), .CLK(clk), .Q(mem[680]) );
  DFFPOSX1 mem_reg_20__19_ ( .D(n2217), .CLK(clk), .Q(mem[679]) );
  DFFPOSX1 mem_reg_20__18_ ( .D(n2216), .CLK(clk), .Q(mem[678]) );
  DFFPOSX1 mem_reg_20__17_ ( .D(n2215), .CLK(clk), .Q(mem[677]) );
  DFFPOSX1 mem_reg_20__16_ ( .D(n2214), .CLK(clk), .Q(mem[676]) );
  DFFPOSX1 mem_reg_20__15_ ( .D(n2213), .CLK(clk), .Q(mem[675]) );
  DFFPOSX1 mem_reg_20__14_ ( .D(n2212), .CLK(clk), .Q(mem[674]) );
  DFFPOSX1 mem_reg_20__13_ ( .D(n2211), .CLK(clk), .Q(mem[673]) );
  DFFPOSX1 mem_reg_20__12_ ( .D(n2210), .CLK(clk), .Q(mem[672]) );
  DFFPOSX1 mem_reg_20__11_ ( .D(n2209), .CLK(clk), .Q(mem[671]) );
  DFFPOSX1 mem_reg_20__10_ ( .D(n2208), .CLK(clk), .Q(mem[670]) );
  DFFPOSX1 mem_reg_20__9_ ( .D(n2207), .CLK(clk), .Q(mem[669]) );
  DFFPOSX1 mem_reg_20__8_ ( .D(n2206), .CLK(clk), .Q(mem[668]) );
  DFFPOSX1 mem_reg_20__7_ ( .D(n2205), .CLK(clk), .Q(mem[667]) );
  DFFPOSX1 mem_reg_20__6_ ( .D(n2204), .CLK(clk), .Q(mem[666]) );
  DFFPOSX1 mem_reg_20__5_ ( .D(n2203), .CLK(clk), .Q(mem[665]) );
  DFFPOSX1 mem_reg_20__4_ ( .D(n2202), .CLK(clk), .Q(mem[664]) );
  DFFPOSX1 mem_reg_20__3_ ( .D(n2201), .CLK(clk), .Q(mem[663]) );
  DFFPOSX1 mem_reg_20__2_ ( .D(n2200), .CLK(clk), .Q(mem[662]) );
  DFFPOSX1 mem_reg_20__1_ ( .D(n2199), .CLK(clk), .Q(mem[661]) );
  DFFPOSX1 mem_reg_20__0_ ( .D(n2198), .CLK(clk), .Q(mem[660]) );
  DFFPOSX1 mem_reg_19__32_ ( .D(n2197), .CLK(clk), .Q(mem[659]) );
  DFFPOSX1 mem_reg_19__31_ ( .D(n2196), .CLK(clk), .Q(mem[658]) );
  DFFPOSX1 mem_reg_19__30_ ( .D(n2195), .CLK(clk), .Q(mem[657]) );
  DFFPOSX1 mem_reg_19__29_ ( .D(n2194), .CLK(clk), .Q(mem[656]) );
  DFFPOSX1 mem_reg_19__28_ ( .D(n2193), .CLK(clk), .Q(mem[655]) );
  DFFPOSX1 mem_reg_19__27_ ( .D(n2192), .CLK(clk), .Q(mem[654]) );
  DFFPOSX1 mem_reg_19__26_ ( .D(n2191), .CLK(clk), .Q(mem[653]) );
  DFFPOSX1 mem_reg_19__25_ ( .D(n2190), .CLK(clk), .Q(mem[652]) );
  DFFPOSX1 mem_reg_19__24_ ( .D(n2189), .CLK(clk), .Q(mem[651]) );
  DFFPOSX1 mem_reg_19__23_ ( .D(n2188), .CLK(clk), .Q(mem[650]) );
  DFFPOSX1 mem_reg_19__22_ ( .D(n2187), .CLK(clk), .Q(mem[649]) );
  DFFPOSX1 mem_reg_19__21_ ( .D(n2186), .CLK(clk), .Q(mem[648]) );
  DFFPOSX1 mem_reg_19__20_ ( .D(n2185), .CLK(clk), .Q(mem[647]) );
  DFFPOSX1 mem_reg_19__19_ ( .D(n2184), .CLK(clk), .Q(mem[646]) );
  DFFPOSX1 mem_reg_19__18_ ( .D(n2183), .CLK(clk), .Q(mem[645]) );
  DFFPOSX1 mem_reg_19__17_ ( .D(n2182), .CLK(clk), .Q(mem[644]) );
  DFFPOSX1 mem_reg_19__16_ ( .D(n2181), .CLK(clk), .Q(mem[643]) );
  DFFPOSX1 mem_reg_19__15_ ( .D(n2180), .CLK(clk), .Q(mem[642]) );
  DFFPOSX1 mem_reg_19__14_ ( .D(n2179), .CLK(clk), .Q(mem[641]) );
  DFFPOSX1 mem_reg_19__13_ ( .D(n2178), .CLK(clk), .Q(mem[640]) );
  DFFPOSX1 mem_reg_19__12_ ( .D(n2177), .CLK(clk), .Q(mem[639]) );
  DFFPOSX1 mem_reg_19__11_ ( .D(n2176), .CLK(clk), .Q(mem[638]) );
  DFFPOSX1 mem_reg_19__10_ ( .D(n2175), .CLK(clk), .Q(mem[637]) );
  DFFPOSX1 mem_reg_19__9_ ( .D(n2174), .CLK(clk), .Q(mem[636]) );
  DFFPOSX1 mem_reg_19__8_ ( .D(n2173), .CLK(clk), .Q(mem[635]) );
  DFFPOSX1 mem_reg_19__7_ ( .D(n2172), .CLK(clk), .Q(mem[634]) );
  DFFPOSX1 mem_reg_19__6_ ( .D(n2171), .CLK(clk), .Q(mem[633]) );
  DFFPOSX1 mem_reg_19__5_ ( .D(n2170), .CLK(clk), .Q(mem[632]) );
  DFFPOSX1 mem_reg_19__4_ ( .D(n2169), .CLK(clk), .Q(mem[631]) );
  DFFPOSX1 mem_reg_19__3_ ( .D(n2168), .CLK(clk), .Q(mem[630]) );
  DFFPOSX1 mem_reg_19__2_ ( .D(n2167), .CLK(clk), .Q(mem[629]) );
  DFFPOSX1 mem_reg_19__1_ ( .D(n2166), .CLK(clk), .Q(mem[628]) );
  DFFPOSX1 mem_reg_19__0_ ( .D(n2165), .CLK(clk), .Q(mem[627]) );
  DFFPOSX1 mem_reg_18__32_ ( .D(n2164), .CLK(clk), .Q(mem[626]) );
  DFFPOSX1 mem_reg_18__31_ ( .D(n2163), .CLK(clk), .Q(mem[625]) );
  DFFPOSX1 mem_reg_18__30_ ( .D(n2162), .CLK(clk), .Q(mem[624]) );
  DFFPOSX1 mem_reg_18__29_ ( .D(n2161), .CLK(clk), .Q(mem[623]) );
  DFFPOSX1 mem_reg_18__28_ ( .D(n2160), .CLK(clk), .Q(mem[622]) );
  DFFPOSX1 mem_reg_18__27_ ( .D(n2159), .CLK(clk), .Q(mem[621]) );
  DFFPOSX1 mem_reg_18__26_ ( .D(n2158), .CLK(clk), .Q(mem[620]) );
  DFFPOSX1 mem_reg_18__25_ ( .D(n2157), .CLK(clk), .Q(mem[619]) );
  DFFPOSX1 mem_reg_18__24_ ( .D(n2156), .CLK(clk), .Q(mem[618]) );
  DFFPOSX1 mem_reg_18__23_ ( .D(n2155), .CLK(clk), .Q(mem[617]) );
  DFFPOSX1 mem_reg_18__22_ ( .D(n2154), .CLK(clk), .Q(mem[616]) );
  DFFPOSX1 mem_reg_18__21_ ( .D(n2153), .CLK(clk), .Q(mem[615]) );
  DFFPOSX1 mem_reg_18__20_ ( .D(n2152), .CLK(clk), .Q(mem[614]) );
  DFFPOSX1 mem_reg_18__19_ ( .D(n2151), .CLK(clk), .Q(mem[613]) );
  DFFPOSX1 mem_reg_18__18_ ( .D(n2150), .CLK(clk), .Q(mem[612]) );
  DFFPOSX1 mem_reg_18__17_ ( .D(n2149), .CLK(clk), .Q(mem[611]) );
  DFFPOSX1 mem_reg_18__16_ ( .D(n2148), .CLK(clk), .Q(mem[610]) );
  DFFPOSX1 mem_reg_18__15_ ( .D(n2147), .CLK(clk), .Q(mem[609]) );
  DFFPOSX1 mem_reg_18__14_ ( .D(n2146), .CLK(clk), .Q(mem[608]) );
  DFFPOSX1 mem_reg_18__13_ ( .D(n2145), .CLK(clk), .Q(mem[607]) );
  DFFPOSX1 mem_reg_18__12_ ( .D(n2144), .CLK(clk), .Q(mem[606]) );
  DFFPOSX1 mem_reg_18__11_ ( .D(n2143), .CLK(clk), .Q(mem[605]) );
  DFFPOSX1 mem_reg_18__10_ ( .D(n2142), .CLK(clk), .Q(mem[604]) );
  DFFPOSX1 mem_reg_18__9_ ( .D(n2141), .CLK(clk), .Q(mem[603]) );
  DFFPOSX1 mem_reg_18__8_ ( .D(n2140), .CLK(clk), .Q(mem[602]) );
  DFFPOSX1 mem_reg_18__7_ ( .D(n2139), .CLK(clk), .Q(mem[601]) );
  DFFPOSX1 mem_reg_18__6_ ( .D(n2138), .CLK(clk), .Q(mem[600]) );
  DFFPOSX1 mem_reg_18__5_ ( .D(n2137), .CLK(clk), .Q(mem[599]) );
  DFFPOSX1 mem_reg_18__4_ ( .D(n2136), .CLK(clk), .Q(mem[598]) );
  DFFPOSX1 mem_reg_18__3_ ( .D(n2135), .CLK(clk), .Q(mem[597]) );
  DFFPOSX1 mem_reg_18__2_ ( .D(n2134), .CLK(clk), .Q(mem[596]) );
  DFFPOSX1 mem_reg_18__1_ ( .D(n2133), .CLK(clk), .Q(mem[595]) );
  DFFPOSX1 mem_reg_18__0_ ( .D(n2132), .CLK(clk), .Q(mem[594]) );
  DFFPOSX1 mem_reg_17__32_ ( .D(n2131), .CLK(clk), .Q(mem[593]) );
  DFFPOSX1 mem_reg_17__31_ ( .D(n2130), .CLK(clk), .Q(mem[592]) );
  DFFPOSX1 mem_reg_17__30_ ( .D(n2129), .CLK(clk), .Q(mem[591]) );
  DFFPOSX1 mem_reg_17__29_ ( .D(n2128), .CLK(clk), .Q(mem[590]) );
  DFFPOSX1 mem_reg_17__28_ ( .D(n2127), .CLK(clk), .Q(mem[589]) );
  DFFPOSX1 mem_reg_17__27_ ( .D(n2126), .CLK(clk), .Q(mem[588]) );
  DFFPOSX1 mem_reg_17__26_ ( .D(n2125), .CLK(clk), .Q(mem[587]) );
  DFFPOSX1 mem_reg_17__25_ ( .D(n2124), .CLK(clk), .Q(mem[586]) );
  DFFPOSX1 mem_reg_17__24_ ( .D(n2123), .CLK(clk), .Q(mem[585]) );
  DFFPOSX1 mem_reg_17__23_ ( .D(n2122), .CLK(clk), .Q(mem[584]) );
  DFFPOSX1 mem_reg_17__22_ ( .D(n2121), .CLK(clk), .Q(mem[583]) );
  DFFPOSX1 mem_reg_17__21_ ( .D(n2120), .CLK(clk), .Q(mem[582]) );
  DFFPOSX1 mem_reg_17__20_ ( .D(n2119), .CLK(clk), .Q(mem[581]) );
  DFFPOSX1 mem_reg_17__19_ ( .D(n2118), .CLK(clk), .Q(mem[580]) );
  DFFPOSX1 mem_reg_17__18_ ( .D(n2117), .CLK(clk), .Q(mem[579]) );
  DFFPOSX1 mem_reg_17__17_ ( .D(n2116), .CLK(clk), .Q(mem[578]) );
  DFFPOSX1 mem_reg_17__16_ ( .D(n2115), .CLK(clk), .Q(mem[577]) );
  DFFPOSX1 mem_reg_17__15_ ( .D(n2114), .CLK(clk), .Q(mem[576]) );
  DFFPOSX1 mem_reg_17__14_ ( .D(n2113), .CLK(clk), .Q(mem[575]) );
  DFFPOSX1 mem_reg_17__13_ ( .D(n2112), .CLK(clk), .Q(mem[574]) );
  DFFPOSX1 mem_reg_17__12_ ( .D(n2111), .CLK(clk), .Q(mem[573]) );
  DFFPOSX1 mem_reg_17__11_ ( .D(n2110), .CLK(clk), .Q(mem[572]) );
  DFFPOSX1 mem_reg_17__10_ ( .D(n2109), .CLK(clk), .Q(mem[571]) );
  DFFPOSX1 mem_reg_17__9_ ( .D(n2108), .CLK(clk), .Q(mem[570]) );
  DFFPOSX1 mem_reg_17__8_ ( .D(n2107), .CLK(clk), .Q(mem[569]) );
  DFFPOSX1 mem_reg_17__7_ ( .D(n2106), .CLK(clk), .Q(mem[568]) );
  DFFPOSX1 mem_reg_17__6_ ( .D(n2105), .CLK(clk), .Q(mem[567]) );
  DFFPOSX1 mem_reg_17__5_ ( .D(n2104), .CLK(clk), .Q(mem[566]) );
  DFFPOSX1 mem_reg_17__4_ ( .D(n2103), .CLK(clk), .Q(mem[565]) );
  DFFPOSX1 mem_reg_17__3_ ( .D(n2102), .CLK(clk), .Q(mem[564]) );
  DFFPOSX1 mem_reg_17__2_ ( .D(n2101), .CLK(clk), .Q(mem[563]) );
  DFFPOSX1 mem_reg_17__1_ ( .D(n2100), .CLK(clk), .Q(mem[562]) );
  DFFPOSX1 mem_reg_17__0_ ( .D(n2099), .CLK(clk), .Q(mem[561]) );
  DFFPOSX1 mem_reg_16__32_ ( .D(n2098), .CLK(clk), .Q(mem[560]) );
  DFFPOSX1 mem_reg_16__31_ ( .D(n2097), .CLK(clk), .Q(mem[559]) );
  DFFPOSX1 mem_reg_16__30_ ( .D(n2096), .CLK(clk), .Q(mem[558]) );
  DFFPOSX1 mem_reg_16__29_ ( .D(n2095), .CLK(clk), .Q(mem[557]) );
  DFFPOSX1 mem_reg_16__28_ ( .D(n2094), .CLK(clk), .Q(mem[556]) );
  DFFPOSX1 mem_reg_16__27_ ( .D(n2093), .CLK(clk), .Q(mem[555]) );
  DFFPOSX1 mem_reg_16__26_ ( .D(n2092), .CLK(clk), .Q(mem[554]) );
  DFFPOSX1 mem_reg_16__25_ ( .D(n2091), .CLK(clk), .Q(mem[553]) );
  DFFPOSX1 mem_reg_16__24_ ( .D(n2090), .CLK(clk), .Q(mem[552]) );
  DFFPOSX1 mem_reg_16__23_ ( .D(n2089), .CLK(clk), .Q(mem[551]) );
  DFFPOSX1 mem_reg_16__22_ ( .D(n2088), .CLK(clk), .Q(mem[550]) );
  DFFPOSX1 mem_reg_16__21_ ( .D(n2087), .CLK(clk), .Q(mem[549]) );
  DFFPOSX1 mem_reg_16__20_ ( .D(n2086), .CLK(clk), .Q(mem[548]) );
  DFFPOSX1 mem_reg_16__19_ ( .D(n2085), .CLK(clk), .Q(mem[547]) );
  DFFPOSX1 mem_reg_16__18_ ( .D(n2084), .CLK(clk), .Q(mem[546]) );
  DFFPOSX1 mem_reg_16__17_ ( .D(n2083), .CLK(clk), .Q(mem[545]) );
  DFFPOSX1 mem_reg_16__16_ ( .D(n2082), .CLK(clk), .Q(mem[544]) );
  DFFPOSX1 mem_reg_16__15_ ( .D(n2081), .CLK(clk), .Q(mem[543]) );
  DFFPOSX1 mem_reg_16__14_ ( .D(n2080), .CLK(clk), .Q(mem[542]) );
  DFFPOSX1 mem_reg_16__13_ ( .D(n2079), .CLK(clk), .Q(mem[541]) );
  DFFPOSX1 mem_reg_16__12_ ( .D(n2078), .CLK(clk), .Q(mem[540]) );
  DFFPOSX1 mem_reg_16__11_ ( .D(n2077), .CLK(clk), .Q(mem[539]) );
  DFFPOSX1 mem_reg_16__10_ ( .D(n2076), .CLK(clk), .Q(mem[538]) );
  DFFPOSX1 mem_reg_16__9_ ( .D(n2075), .CLK(clk), .Q(mem[537]) );
  DFFPOSX1 mem_reg_16__8_ ( .D(n2074), .CLK(clk), .Q(mem[536]) );
  DFFPOSX1 mem_reg_16__7_ ( .D(n2073), .CLK(clk), .Q(mem[535]) );
  DFFPOSX1 mem_reg_16__6_ ( .D(n2072), .CLK(clk), .Q(mem[534]) );
  DFFPOSX1 mem_reg_16__5_ ( .D(n2071), .CLK(clk), .Q(mem[533]) );
  DFFPOSX1 mem_reg_16__4_ ( .D(n2070), .CLK(clk), .Q(mem[532]) );
  DFFPOSX1 mem_reg_16__3_ ( .D(n2069), .CLK(clk), .Q(mem[531]) );
  DFFPOSX1 mem_reg_16__2_ ( .D(n2068), .CLK(clk), .Q(mem[530]) );
  DFFPOSX1 mem_reg_16__1_ ( .D(n2067), .CLK(clk), .Q(mem[529]) );
  DFFPOSX1 mem_reg_16__0_ ( .D(n2066), .CLK(clk), .Q(mem[528]) );
  DFFPOSX1 mem_reg_15__32_ ( .D(n2065), .CLK(clk), .Q(mem[527]) );
  DFFPOSX1 mem_reg_15__31_ ( .D(n2064), .CLK(clk), .Q(mem[526]) );
  DFFPOSX1 mem_reg_15__30_ ( .D(n2063), .CLK(clk), .Q(mem[525]) );
  DFFPOSX1 mem_reg_15__29_ ( .D(n2062), .CLK(clk), .Q(mem[524]) );
  DFFPOSX1 mem_reg_15__28_ ( .D(n2061), .CLK(clk), .Q(mem[523]) );
  DFFPOSX1 mem_reg_15__27_ ( .D(n2060), .CLK(clk), .Q(mem[522]) );
  DFFPOSX1 mem_reg_15__26_ ( .D(n2059), .CLK(clk), .Q(mem[521]) );
  DFFPOSX1 mem_reg_15__25_ ( .D(n2058), .CLK(clk), .Q(mem[520]) );
  DFFPOSX1 mem_reg_15__24_ ( .D(n2057), .CLK(clk), .Q(mem[519]) );
  DFFPOSX1 mem_reg_15__23_ ( .D(n2056), .CLK(clk), .Q(mem[518]) );
  DFFPOSX1 mem_reg_15__22_ ( .D(n2055), .CLK(clk), .Q(mem[517]) );
  DFFPOSX1 mem_reg_15__21_ ( .D(n2054), .CLK(clk), .Q(mem[516]) );
  DFFPOSX1 mem_reg_15__20_ ( .D(n2053), .CLK(clk), .Q(mem[515]) );
  DFFPOSX1 mem_reg_15__19_ ( .D(n2052), .CLK(clk), .Q(mem[514]) );
  DFFPOSX1 mem_reg_15__18_ ( .D(n2051), .CLK(clk), .Q(mem[513]) );
  DFFPOSX1 mem_reg_15__17_ ( .D(n2050), .CLK(clk), .Q(mem[512]) );
  DFFPOSX1 mem_reg_15__16_ ( .D(n2049), .CLK(clk), .Q(mem[511]) );
  DFFPOSX1 mem_reg_15__15_ ( .D(n2048), .CLK(clk), .Q(mem[510]) );
  DFFPOSX1 mem_reg_15__14_ ( .D(n2047), .CLK(clk), .Q(mem[509]) );
  DFFPOSX1 mem_reg_15__13_ ( .D(n2046), .CLK(clk), .Q(mem[508]) );
  DFFPOSX1 mem_reg_15__12_ ( .D(n2045), .CLK(clk), .Q(mem[507]) );
  DFFPOSX1 mem_reg_15__11_ ( .D(n2044), .CLK(clk), .Q(mem[506]) );
  DFFPOSX1 mem_reg_15__10_ ( .D(n2043), .CLK(clk), .Q(mem[505]) );
  DFFPOSX1 mem_reg_15__9_ ( .D(n2042), .CLK(clk), .Q(mem[504]) );
  DFFPOSX1 mem_reg_15__8_ ( .D(n2041), .CLK(clk), .Q(mem[503]) );
  DFFPOSX1 mem_reg_15__7_ ( .D(n2040), .CLK(clk), .Q(mem[502]) );
  DFFPOSX1 mem_reg_15__6_ ( .D(n2039), .CLK(clk), .Q(mem[501]) );
  DFFPOSX1 mem_reg_15__5_ ( .D(n2038), .CLK(clk), .Q(mem[500]) );
  DFFPOSX1 mem_reg_15__4_ ( .D(n2037), .CLK(clk), .Q(mem[499]) );
  DFFPOSX1 mem_reg_15__3_ ( .D(n2036), .CLK(clk), .Q(mem[498]) );
  DFFPOSX1 mem_reg_15__2_ ( .D(n2035), .CLK(clk), .Q(mem[497]) );
  DFFPOSX1 mem_reg_15__1_ ( .D(n2034), .CLK(clk), .Q(mem[496]) );
  DFFPOSX1 mem_reg_15__0_ ( .D(n2033), .CLK(clk), .Q(mem[495]) );
  DFFPOSX1 mem_reg_14__32_ ( .D(n2032), .CLK(clk), .Q(mem[494]) );
  DFFPOSX1 mem_reg_14__31_ ( .D(n2031), .CLK(clk), .Q(mem[493]) );
  DFFPOSX1 mem_reg_14__30_ ( .D(n2030), .CLK(clk), .Q(mem[492]) );
  DFFPOSX1 mem_reg_14__29_ ( .D(n2029), .CLK(clk), .Q(mem[491]) );
  DFFPOSX1 mem_reg_14__28_ ( .D(n2028), .CLK(clk), .Q(mem[490]) );
  DFFPOSX1 mem_reg_14__27_ ( .D(n2027), .CLK(clk), .Q(mem[489]) );
  DFFPOSX1 mem_reg_14__26_ ( .D(n2026), .CLK(clk), .Q(mem[488]) );
  DFFPOSX1 mem_reg_14__25_ ( .D(n2025), .CLK(clk), .Q(mem[487]) );
  DFFPOSX1 mem_reg_14__24_ ( .D(n2024), .CLK(clk), .Q(mem[486]) );
  DFFPOSX1 mem_reg_14__23_ ( .D(n2023), .CLK(clk), .Q(mem[485]) );
  DFFPOSX1 mem_reg_14__22_ ( .D(n2022), .CLK(clk), .Q(mem[484]) );
  DFFPOSX1 mem_reg_14__21_ ( .D(n2021), .CLK(clk), .Q(mem[483]) );
  DFFPOSX1 mem_reg_14__20_ ( .D(n2020), .CLK(clk), .Q(mem[482]) );
  DFFPOSX1 mem_reg_14__19_ ( .D(n2019), .CLK(clk), .Q(mem[481]) );
  DFFPOSX1 mem_reg_14__18_ ( .D(n2018), .CLK(clk), .Q(mem[480]) );
  DFFPOSX1 mem_reg_14__17_ ( .D(n2017), .CLK(clk), .Q(mem[479]) );
  DFFPOSX1 mem_reg_14__16_ ( .D(n2016), .CLK(clk), .Q(mem[478]) );
  DFFPOSX1 mem_reg_14__15_ ( .D(n2015), .CLK(clk), .Q(mem[477]) );
  DFFPOSX1 mem_reg_14__14_ ( .D(n2014), .CLK(clk), .Q(mem[476]) );
  DFFPOSX1 mem_reg_14__13_ ( .D(n2013), .CLK(clk), .Q(mem[475]) );
  DFFPOSX1 mem_reg_14__12_ ( .D(n2012), .CLK(clk), .Q(mem[474]) );
  DFFPOSX1 mem_reg_14__11_ ( .D(n2011), .CLK(clk), .Q(mem[473]) );
  DFFPOSX1 mem_reg_14__10_ ( .D(n2010), .CLK(clk), .Q(mem[472]) );
  DFFPOSX1 mem_reg_14__9_ ( .D(n2009), .CLK(clk), .Q(mem[471]) );
  DFFPOSX1 mem_reg_14__8_ ( .D(n2008), .CLK(clk), .Q(mem[470]) );
  DFFPOSX1 mem_reg_14__7_ ( .D(n2007), .CLK(clk), .Q(mem[469]) );
  DFFPOSX1 mem_reg_14__6_ ( .D(n2006), .CLK(clk), .Q(mem[468]) );
  DFFPOSX1 mem_reg_14__5_ ( .D(n2005), .CLK(clk), .Q(mem[467]) );
  DFFPOSX1 mem_reg_14__4_ ( .D(n2004), .CLK(clk), .Q(mem[466]) );
  DFFPOSX1 mem_reg_14__3_ ( .D(n2003), .CLK(clk), .Q(mem[465]) );
  DFFPOSX1 mem_reg_14__2_ ( .D(n2002), .CLK(clk), .Q(mem[464]) );
  DFFPOSX1 mem_reg_14__1_ ( .D(n2001), .CLK(clk), .Q(mem[463]) );
  DFFPOSX1 mem_reg_14__0_ ( .D(n2000), .CLK(clk), .Q(mem[462]) );
  DFFPOSX1 mem_reg_13__32_ ( .D(n1999), .CLK(clk), .Q(mem[461]) );
  DFFPOSX1 mem_reg_13__31_ ( .D(n1998), .CLK(clk), .Q(mem[460]) );
  DFFPOSX1 mem_reg_13__30_ ( .D(n1997), .CLK(clk), .Q(mem[459]) );
  DFFPOSX1 mem_reg_13__29_ ( .D(n1996), .CLK(clk), .Q(mem[458]) );
  DFFPOSX1 mem_reg_13__28_ ( .D(n1995), .CLK(clk), .Q(mem[457]) );
  DFFPOSX1 mem_reg_13__27_ ( .D(n1994), .CLK(clk), .Q(mem[456]) );
  DFFPOSX1 mem_reg_13__26_ ( .D(n1993), .CLK(clk), .Q(mem[455]) );
  DFFPOSX1 mem_reg_13__25_ ( .D(n1992), .CLK(clk), .Q(mem[454]) );
  DFFPOSX1 mem_reg_13__24_ ( .D(n1991), .CLK(clk), .Q(mem[453]) );
  DFFPOSX1 mem_reg_13__23_ ( .D(n1990), .CLK(clk), .Q(mem[452]) );
  DFFPOSX1 mem_reg_13__22_ ( .D(n1989), .CLK(clk), .Q(mem[451]) );
  DFFPOSX1 mem_reg_13__21_ ( .D(n1988), .CLK(clk), .Q(mem[450]) );
  DFFPOSX1 mem_reg_13__20_ ( .D(n1987), .CLK(clk), .Q(mem[449]) );
  DFFPOSX1 mem_reg_13__19_ ( .D(n1986), .CLK(clk), .Q(mem[448]) );
  DFFPOSX1 mem_reg_13__18_ ( .D(n1985), .CLK(clk), .Q(mem[447]) );
  DFFPOSX1 mem_reg_13__17_ ( .D(n1984), .CLK(clk), .Q(mem[446]) );
  DFFPOSX1 mem_reg_13__16_ ( .D(n1983), .CLK(clk), .Q(mem[445]) );
  DFFPOSX1 mem_reg_13__15_ ( .D(n1982), .CLK(clk), .Q(mem[444]) );
  DFFPOSX1 mem_reg_13__14_ ( .D(n1981), .CLK(clk), .Q(mem[443]) );
  DFFPOSX1 mem_reg_13__13_ ( .D(n1980), .CLK(clk), .Q(mem[442]) );
  DFFPOSX1 mem_reg_13__12_ ( .D(n1979), .CLK(clk), .Q(mem[441]) );
  DFFPOSX1 mem_reg_13__11_ ( .D(n1978), .CLK(clk), .Q(mem[440]) );
  DFFPOSX1 mem_reg_13__10_ ( .D(n1977), .CLK(clk), .Q(mem[439]) );
  DFFPOSX1 mem_reg_13__9_ ( .D(n1976), .CLK(clk), .Q(mem[438]) );
  DFFPOSX1 mem_reg_13__8_ ( .D(n1975), .CLK(clk), .Q(mem[437]) );
  DFFPOSX1 mem_reg_13__7_ ( .D(n1974), .CLK(clk), .Q(mem[436]) );
  DFFPOSX1 mem_reg_13__6_ ( .D(n1973), .CLK(clk), .Q(mem[435]) );
  DFFPOSX1 mem_reg_13__5_ ( .D(n1972), .CLK(clk), .Q(mem[434]) );
  DFFPOSX1 mem_reg_13__4_ ( .D(n1971), .CLK(clk), .Q(mem[433]) );
  DFFPOSX1 mem_reg_13__3_ ( .D(n1970), .CLK(clk), .Q(mem[432]) );
  DFFPOSX1 mem_reg_13__2_ ( .D(n1969), .CLK(clk), .Q(mem[431]) );
  DFFPOSX1 mem_reg_13__1_ ( .D(n1968), .CLK(clk), .Q(mem[430]) );
  DFFPOSX1 mem_reg_13__0_ ( .D(n1967), .CLK(clk), .Q(mem[429]) );
  DFFPOSX1 mem_reg_12__32_ ( .D(n1966), .CLK(clk), .Q(mem[428]) );
  DFFPOSX1 mem_reg_12__31_ ( .D(n1965), .CLK(clk), .Q(mem[427]) );
  DFFPOSX1 mem_reg_12__30_ ( .D(n1964), .CLK(clk), .Q(mem[426]) );
  DFFPOSX1 mem_reg_12__29_ ( .D(n1963), .CLK(clk), .Q(mem[425]) );
  DFFPOSX1 mem_reg_12__28_ ( .D(n1962), .CLK(clk), .Q(mem[424]) );
  DFFPOSX1 mem_reg_12__27_ ( .D(n1961), .CLK(clk), .Q(mem[423]) );
  DFFPOSX1 mem_reg_12__26_ ( .D(n1960), .CLK(clk), .Q(mem[422]) );
  DFFPOSX1 mem_reg_12__25_ ( .D(n1959), .CLK(clk), .Q(mem[421]) );
  DFFPOSX1 mem_reg_12__24_ ( .D(n1958), .CLK(clk), .Q(mem[420]) );
  DFFPOSX1 mem_reg_12__23_ ( .D(n1957), .CLK(clk), .Q(mem[419]) );
  DFFPOSX1 mem_reg_12__22_ ( .D(n1956), .CLK(clk), .Q(mem[418]) );
  DFFPOSX1 mem_reg_12__21_ ( .D(n1955), .CLK(clk), .Q(mem[417]) );
  DFFPOSX1 mem_reg_12__20_ ( .D(n1954), .CLK(clk), .Q(mem[416]) );
  DFFPOSX1 mem_reg_12__19_ ( .D(n1953), .CLK(clk), .Q(mem[415]) );
  DFFPOSX1 mem_reg_12__18_ ( .D(n1952), .CLK(clk), .Q(mem[414]) );
  DFFPOSX1 mem_reg_12__17_ ( .D(n1951), .CLK(clk), .Q(mem[413]) );
  DFFPOSX1 mem_reg_12__16_ ( .D(n1950), .CLK(clk), .Q(mem[412]) );
  DFFPOSX1 mem_reg_12__15_ ( .D(n1949), .CLK(clk), .Q(mem[411]) );
  DFFPOSX1 mem_reg_12__14_ ( .D(n1948), .CLK(clk), .Q(mem[410]) );
  DFFPOSX1 mem_reg_12__13_ ( .D(n1947), .CLK(clk), .Q(mem[409]) );
  DFFPOSX1 mem_reg_12__12_ ( .D(n1946), .CLK(clk), .Q(mem[408]) );
  DFFPOSX1 mem_reg_12__11_ ( .D(n1945), .CLK(clk), .Q(mem[407]) );
  DFFPOSX1 mem_reg_12__10_ ( .D(n1944), .CLK(clk), .Q(mem[406]) );
  DFFPOSX1 mem_reg_12__9_ ( .D(n1943), .CLK(clk), .Q(mem[405]) );
  DFFPOSX1 mem_reg_12__8_ ( .D(n1942), .CLK(clk), .Q(mem[404]) );
  DFFPOSX1 mem_reg_12__7_ ( .D(n1941), .CLK(clk), .Q(mem[403]) );
  DFFPOSX1 mem_reg_12__6_ ( .D(n1940), .CLK(clk), .Q(mem[402]) );
  DFFPOSX1 mem_reg_12__5_ ( .D(n1939), .CLK(clk), .Q(mem[401]) );
  DFFPOSX1 mem_reg_12__4_ ( .D(n1938), .CLK(clk), .Q(mem[400]) );
  DFFPOSX1 mem_reg_12__3_ ( .D(n1937), .CLK(clk), .Q(mem[399]) );
  DFFPOSX1 mem_reg_12__2_ ( .D(n1936), .CLK(clk), .Q(mem[398]) );
  DFFPOSX1 mem_reg_12__1_ ( .D(n1935), .CLK(clk), .Q(mem[397]) );
  DFFPOSX1 mem_reg_12__0_ ( .D(n1934), .CLK(clk), .Q(mem[396]) );
  DFFPOSX1 mem_reg_11__32_ ( .D(n1933), .CLK(clk), .Q(mem[395]) );
  DFFPOSX1 mem_reg_11__31_ ( .D(n1932), .CLK(clk), .Q(mem[394]) );
  DFFPOSX1 mem_reg_11__30_ ( .D(n1931), .CLK(clk), .Q(mem[393]) );
  DFFPOSX1 mem_reg_11__29_ ( .D(n1930), .CLK(clk), .Q(mem[392]) );
  DFFPOSX1 mem_reg_11__28_ ( .D(n1929), .CLK(clk), .Q(mem[391]) );
  DFFPOSX1 mem_reg_11__27_ ( .D(n1928), .CLK(clk), .Q(mem[390]) );
  DFFPOSX1 mem_reg_11__26_ ( .D(n1927), .CLK(clk), .Q(mem[389]) );
  DFFPOSX1 mem_reg_11__25_ ( .D(n1926), .CLK(clk), .Q(mem[388]) );
  DFFPOSX1 mem_reg_11__24_ ( .D(n1925), .CLK(clk), .Q(mem[387]) );
  DFFPOSX1 mem_reg_11__23_ ( .D(n1924), .CLK(clk), .Q(mem[386]) );
  DFFPOSX1 mem_reg_11__22_ ( .D(n1923), .CLK(clk), .Q(mem[385]) );
  DFFPOSX1 mem_reg_11__21_ ( .D(n1922), .CLK(clk), .Q(mem[384]) );
  DFFPOSX1 mem_reg_11__20_ ( .D(n1921), .CLK(clk), .Q(mem[383]) );
  DFFPOSX1 mem_reg_11__19_ ( .D(n1920), .CLK(clk), .Q(mem[382]) );
  DFFPOSX1 mem_reg_11__18_ ( .D(n1919), .CLK(clk), .Q(mem[381]) );
  DFFPOSX1 mem_reg_11__17_ ( .D(n1918), .CLK(clk), .Q(mem[380]) );
  DFFPOSX1 mem_reg_11__16_ ( .D(n1917), .CLK(clk), .Q(mem[379]) );
  DFFPOSX1 mem_reg_11__15_ ( .D(n1916), .CLK(clk), .Q(mem[378]) );
  DFFPOSX1 mem_reg_11__14_ ( .D(n1915), .CLK(clk), .Q(mem[377]) );
  DFFPOSX1 mem_reg_11__13_ ( .D(n1914), .CLK(clk), .Q(mem[376]) );
  DFFPOSX1 mem_reg_11__12_ ( .D(n1913), .CLK(clk), .Q(mem[375]) );
  DFFPOSX1 mem_reg_11__11_ ( .D(n1912), .CLK(clk), .Q(mem[374]) );
  DFFPOSX1 mem_reg_11__10_ ( .D(n1911), .CLK(clk), .Q(mem[373]) );
  DFFPOSX1 mem_reg_11__9_ ( .D(n1910), .CLK(clk), .Q(mem[372]) );
  DFFPOSX1 mem_reg_11__8_ ( .D(n1909), .CLK(clk), .Q(mem[371]) );
  DFFPOSX1 mem_reg_11__7_ ( .D(n1908), .CLK(clk), .Q(mem[370]) );
  DFFPOSX1 mem_reg_11__6_ ( .D(n1907), .CLK(clk), .Q(mem[369]) );
  DFFPOSX1 mem_reg_11__5_ ( .D(n1906), .CLK(clk), .Q(mem[368]) );
  DFFPOSX1 mem_reg_11__4_ ( .D(n1905), .CLK(clk), .Q(mem[367]) );
  DFFPOSX1 mem_reg_11__3_ ( .D(n1904), .CLK(clk), .Q(mem[366]) );
  DFFPOSX1 mem_reg_11__2_ ( .D(n1903), .CLK(clk), .Q(mem[365]) );
  DFFPOSX1 mem_reg_11__1_ ( .D(n1902), .CLK(clk), .Q(mem[364]) );
  DFFPOSX1 mem_reg_11__0_ ( .D(n1901), .CLK(clk), .Q(mem[363]) );
  DFFPOSX1 mem_reg_10__32_ ( .D(n1900), .CLK(clk), .Q(mem[362]) );
  DFFPOSX1 mem_reg_10__31_ ( .D(n1899), .CLK(clk), .Q(mem[361]) );
  DFFPOSX1 mem_reg_10__30_ ( .D(n1898), .CLK(clk), .Q(mem[360]) );
  DFFPOSX1 mem_reg_10__29_ ( .D(n1897), .CLK(clk), .Q(mem[359]) );
  DFFPOSX1 mem_reg_10__28_ ( .D(n1896), .CLK(clk), .Q(mem[358]) );
  DFFPOSX1 mem_reg_10__27_ ( .D(n1895), .CLK(clk), .Q(mem[357]) );
  DFFPOSX1 mem_reg_10__26_ ( .D(n1894), .CLK(clk), .Q(mem[356]) );
  DFFPOSX1 mem_reg_10__25_ ( .D(n1893), .CLK(clk), .Q(mem[355]) );
  DFFPOSX1 mem_reg_10__24_ ( .D(n1892), .CLK(clk), .Q(mem[354]) );
  DFFPOSX1 mem_reg_10__23_ ( .D(n1891), .CLK(clk), .Q(mem[353]) );
  DFFPOSX1 mem_reg_10__22_ ( .D(n1890), .CLK(clk), .Q(mem[352]) );
  DFFPOSX1 mem_reg_10__21_ ( .D(n1889), .CLK(clk), .Q(mem[351]) );
  DFFPOSX1 mem_reg_10__20_ ( .D(n1888), .CLK(clk), .Q(mem[350]) );
  DFFPOSX1 mem_reg_10__19_ ( .D(n1887), .CLK(clk), .Q(mem[349]) );
  DFFPOSX1 mem_reg_10__18_ ( .D(n1886), .CLK(clk), .Q(mem[348]) );
  DFFPOSX1 mem_reg_10__17_ ( .D(n1885), .CLK(clk), .Q(mem[347]) );
  DFFPOSX1 mem_reg_10__16_ ( .D(n1884), .CLK(clk), .Q(mem[346]) );
  DFFPOSX1 mem_reg_10__15_ ( .D(n1883), .CLK(clk), .Q(mem[345]) );
  DFFPOSX1 mem_reg_10__14_ ( .D(n1882), .CLK(clk), .Q(mem[344]) );
  DFFPOSX1 mem_reg_10__13_ ( .D(n1881), .CLK(clk), .Q(mem[343]) );
  DFFPOSX1 mem_reg_10__12_ ( .D(n1880), .CLK(clk), .Q(mem[342]) );
  DFFPOSX1 mem_reg_10__11_ ( .D(n1879), .CLK(clk), .Q(mem[341]) );
  DFFPOSX1 mem_reg_10__10_ ( .D(n1878), .CLK(clk), .Q(mem[340]) );
  DFFPOSX1 mem_reg_10__9_ ( .D(n1877), .CLK(clk), .Q(mem[339]) );
  DFFPOSX1 mem_reg_10__8_ ( .D(n1876), .CLK(clk), .Q(mem[338]) );
  DFFPOSX1 mem_reg_10__7_ ( .D(n1875), .CLK(clk), .Q(mem[337]) );
  DFFPOSX1 mem_reg_10__6_ ( .D(n1874), .CLK(clk), .Q(mem[336]) );
  DFFPOSX1 mem_reg_10__5_ ( .D(n1873), .CLK(clk), .Q(mem[335]) );
  DFFPOSX1 mem_reg_10__4_ ( .D(n1872), .CLK(clk), .Q(mem[334]) );
  DFFPOSX1 mem_reg_10__3_ ( .D(n1871), .CLK(clk), .Q(mem[333]) );
  DFFPOSX1 mem_reg_10__2_ ( .D(n1870), .CLK(clk), .Q(mem[332]) );
  DFFPOSX1 mem_reg_10__1_ ( .D(n1869), .CLK(clk), .Q(mem[331]) );
  DFFPOSX1 mem_reg_10__0_ ( .D(n1868), .CLK(clk), .Q(mem[330]) );
  DFFPOSX1 mem_reg_9__32_ ( .D(n1867), .CLK(clk), .Q(mem[329]) );
  DFFPOSX1 mem_reg_9__31_ ( .D(n1866), .CLK(clk), .Q(mem[328]) );
  DFFPOSX1 mem_reg_9__30_ ( .D(n1865), .CLK(clk), .Q(mem[327]) );
  DFFPOSX1 mem_reg_9__29_ ( .D(n1864), .CLK(clk), .Q(mem[326]) );
  DFFPOSX1 mem_reg_9__28_ ( .D(n1863), .CLK(clk), .Q(mem[325]) );
  DFFPOSX1 mem_reg_9__27_ ( .D(n1862), .CLK(clk), .Q(mem[324]) );
  DFFPOSX1 mem_reg_9__26_ ( .D(n1861), .CLK(clk), .Q(mem[323]) );
  DFFPOSX1 mem_reg_9__25_ ( .D(n1860), .CLK(clk), .Q(mem[322]) );
  DFFPOSX1 mem_reg_9__24_ ( .D(n1859), .CLK(clk), .Q(mem[321]) );
  DFFPOSX1 mem_reg_9__23_ ( .D(n1858), .CLK(clk), .Q(mem[320]) );
  DFFPOSX1 mem_reg_9__22_ ( .D(n1857), .CLK(clk), .Q(mem[319]) );
  DFFPOSX1 mem_reg_9__21_ ( .D(n1856), .CLK(clk), .Q(mem[318]) );
  DFFPOSX1 mem_reg_9__20_ ( .D(n1855), .CLK(clk), .Q(mem[317]) );
  DFFPOSX1 mem_reg_9__19_ ( .D(n1854), .CLK(clk), .Q(mem[316]) );
  DFFPOSX1 mem_reg_9__18_ ( .D(n1853), .CLK(clk), .Q(mem[315]) );
  DFFPOSX1 mem_reg_9__17_ ( .D(n1852), .CLK(clk), .Q(mem[314]) );
  DFFPOSX1 mem_reg_9__16_ ( .D(n1851), .CLK(clk), .Q(mem[313]) );
  DFFPOSX1 mem_reg_9__15_ ( .D(n1850), .CLK(clk), .Q(mem[312]) );
  DFFPOSX1 mem_reg_9__14_ ( .D(n1849), .CLK(clk), .Q(mem[311]) );
  DFFPOSX1 mem_reg_9__13_ ( .D(n1848), .CLK(clk), .Q(mem[310]) );
  DFFPOSX1 mem_reg_9__12_ ( .D(n1847), .CLK(clk), .Q(mem[309]) );
  DFFPOSX1 mem_reg_9__11_ ( .D(n1846), .CLK(clk), .Q(mem[308]) );
  DFFPOSX1 mem_reg_9__10_ ( .D(n1845), .CLK(clk), .Q(mem[307]) );
  DFFPOSX1 mem_reg_9__9_ ( .D(n1844), .CLK(clk), .Q(mem[306]) );
  DFFPOSX1 mem_reg_9__8_ ( .D(n1843), .CLK(clk), .Q(mem[305]) );
  DFFPOSX1 mem_reg_9__7_ ( .D(n1842), .CLK(clk), .Q(mem[304]) );
  DFFPOSX1 mem_reg_9__6_ ( .D(n1841), .CLK(clk), .Q(mem[303]) );
  DFFPOSX1 mem_reg_9__5_ ( .D(n1840), .CLK(clk), .Q(mem[302]) );
  DFFPOSX1 mem_reg_9__4_ ( .D(n1839), .CLK(clk), .Q(mem[301]) );
  DFFPOSX1 mem_reg_9__3_ ( .D(n1838), .CLK(clk), .Q(mem[300]) );
  DFFPOSX1 mem_reg_9__2_ ( .D(n1837), .CLK(clk), .Q(mem[299]) );
  DFFPOSX1 mem_reg_9__1_ ( .D(n1836), .CLK(clk), .Q(mem[298]) );
  DFFPOSX1 mem_reg_9__0_ ( .D(n1835), .CLK(clk), .Q(mem[297]) );
  DFFPOSX1 mem_reg_8__32_ ( .D(n1834), .CLK(clk), .Q(mem[296]) );
  DFFPOSX1 mem_reg_8__31_ ( .D(n1833), .CLK(clk), .Q(mem[295]) );
  DFFPOSX1 mem_reg_8__30_ ( .D(n1832), .CLK(clk), .Q(mem[294]) );
  DFFPOSX1 mem_reg_8__29_ ( .D(n1831), .CLK(clk), .Q(mem[293]) );
  DFFPOSX1 mem_reg_8__28_ ( .D(n1830), .CLK(clk), .Q(mem[292]) );
  DFFPOSX1 mem_reg_8__27_ ( .D(n1829), .CLK(clk), .Q(mem[291]) );
  DFFPOSX1 mem_reg_8__26_ ( .D(n1828), .CLK(clk), .Q(mem[290]) );
  DFFPOSX1 mem_reg_8__25_ ( .D(n1827), .CLK(clk), .Q(mem[289]) );
  DFFPOSX1 mem_reg_8__24_ ( .D(n1826), .CLK(clk), .Q(mem[288]) );
  DFFPOSX1 mem_reg_8__23_ ( .D(n1825), .CLK(clk), .Q(mem[287]) );
  DFFPOSX1 mem_reg_8__22_ ( .D(n1824), .CLK(clk), .Q(mem[286]) );
  DFFPOSX1 mem_reg_8__21_ ( .D(n1823), .CLK(clk), .Q(mem[285]) );
  DFFPOSX1 mem_reg_8__20_ ( .D(n1822), .CLK(clk), .Q(mem[284]) );
  DFFPOSX1 mem_reg_8__19_ ( .D(n1821), .CLK(clk), .Q(mem[283]) );
  DFFPOSX1 mem_reg_8__18_ ( .D(n1820), .CLK(clk), .Q(mem[282]) );
  DFFPOSX1 mem_reg_8__17_ ( .D(n1819), .CLK(clk), .Q(mem[281]) );
  DFFPOSX1 mem_reg_8__16_ ( .D(n1818), .CLK(clk), .Q(mem[280]) );
  DFFPOSX1 mem_reg_8__15_ ( .D(n1817), .CLK(clk), .Q(mem[279]) );
  DFFPOSX1 mem_reg_8__14_ ( .D(n1816), .CLK(clk), .Q(mem[278]) );
  DFFPOSX1 mem_reg_8__13_ ( .D(n1815), .CLK(clk), .Q(mem[277]) );
  DFFPOSX1 mem_reg_8__12_ ( .D(n1814), .CLK(clk), .Q(mem[276]) );
  DFFPOSX1 mem_reg_8__11_ ( .D(n1813), .CLK(clk), .Q(mem[275]) );
  DFFPOSX1 mem_reg_8__10_ ( .D(n1812), .CLK(clk), .Q(mem[274]) );
  DFFPOSX1 mem_reg_8__9_ ( .D(n1811), .CLK(clk), .Q(mem[273]) );
  DFFPOSX1 mem_reg_8__8_ ( .D(n1810), .CLK(clk), .Q(mem[272]) );
  DFFPOSX1 mem_reg_8__7_ ( .D(n1809), .CLK(clk), .Q(mem[271]) );
  DFFPOSX1 mem_reg_8__6_ ( .D(n1808), .CLK(clk), .Q(mem[270]) );
  DFFPOSX1 mem_reg_8__5_ ( .D(n1807), .CLK(clk), .Q(mem[269]) );
  DFFPOSX1 mem_reg_8__4_ ( .D(n1806), .CLK(clk), .Q(mem[268]) );
  DFFPOSX1 mem_reg_8__3_ ( .D(n1805), .CLK(clk), .Q(mem[267]) );
  DFFPOSX1 mem_reg_8__2_ ( .D(n1804), .CLK(clk), .Q(mem[266]) );
  DFFPOSX1 mem_reg_8__1_ ( .D(n1803), .CLK(clk), .Q(mem[265]) );
  DFFPOSX1 mem_reg_8__0_ ( .D(n1802), .CLK(clk), .Q(mem[264]) );
  DFFPOSX1 mem_reg_7__32_ ( .D(n1801), .CLK(clk), .Q(mem[263]) );
  DFFPOSX1 mem_reg_7__31_ ( .D(n1800), .CLK(clk), .Q(mem[262]) );
  DFFPOSX1 mem_reg_7__30_ ( .D(n1799), .CLK(clk), .Q(mem[261]) );
  DFFPOSX1 mem_reg_7__29_ ( .D(n1798), .CLK(clk), .Q(mem[260]) );
  DFFPOSX1 mem_reg_7__28_ ( .D(n1797), .CLK(clk), .Q(mem[259]) );
  DFFPOSX1 mem_reg_7__27_ ( .D(n1796), .CLK(clk), .Q(mem[258]) );
  DFFPOSX1 mem_reg_7__26_ ( .D(n1795), .CLK(clk), .Q(mem[257]) );
  DFFPOSX1 mem_reg_7__25_ ( .D(n1794), .CLK(clk), .Q(mem[256]) );
  DFFPOSX1 mem_reg_7__24_ ( .D(n1793), .CLK(clk), .Q(mem[255]) );
  DFFPOSX1 mem_reg_7__23_ ( .D(n1792), .CLK(clk), .Q(mem[254]) );
  DFFPOSX1 mem_reg_7__22_ ( .D(n1791), .CLK(clk), .Q(mem[253]) );
  DFFPOSX1 mem_reg_7__21_ ( .D(n1790), .CLK(clk), .Q(mem[252]) );
  DFFPOSX1 mem_reg_7__20_ ( .D(n1789), .CLK(clk), .Q(mem[251]) );
  DFFPOSX1 mem_reg_7__19_ ( .D(n1788), .CLK(clk), .Q(mem[250]) );
  DFFPOSX1 mem_reg_7__18_ ( .D(n1787), .CLK(clk), .Q(mem[249]) );
  DFFPOSX1 mem_reg_7__17_ ( .D(n1786), .CLK(clk), .Q(mem[248]) );
  DFFPOSX1 mem_reg_7__16_ ( .D(n1785), .CLK(clk), .Q(mem[247]) );
  DFFPOSX1 mem_reg_7__15_ ( .D(n1784), .CLK(clk), .Q(mem[246]) );
  DFFPOSX1 mem_reg_7__14_ ( .D(n1783), .CLK(clk), .Q(mem[245]) );
  DFFPOSX1 mem_reg_7__13_ ( .D(n1782), .CLK(clk), .Q(mem[244]) );
  DFFPOSX1 mem_reg_7__12_ ( .D(n1781), .CLK(clk), .Q(mem[243]) );
  DFFPOSX1 mem_reg_7__11_ ( .D(n1780), .CLK(clk), .Q(mem[242]) );
  DFFPOSX1 mem_reg_7__10_ ( .D(n1779), .CLK(clk), .Q(mem[241]) );
  DFFPOSX1 mem_reg_7__9_ ( .D(n1778), .CLK(clk), .Q(mem[240]) );
  DFFPOSX1 mem_reg_7__8_ ( .D(n1777), .CLK(clk), .Q(mem[239]) );
  DFFPOSX1 mem_reg_7__7_ ( .D(n1776), .CLK(clk), .Q(mem[238]) );
  DFFPOSX1 mem_reg_7__6_ ( .D(n1775), .CLK(clk), .Q(mem[237]) );
  DFFPOSX1 mem_reg_7__5_ ( .D(n1774), .CLK(clk), .Q(mem[236]) );
  DFFPOSX1 mem_reg_7__4_ ( .D(n1773), .CLK(clk), .Q(mem[235]) );
  DFFPOSX1 mem_reg_7__3_ ( .D(n1772), .CLK(clk), .Q(mem[234]) );
  DFFPOSX1 mem_reg_7__2_ ( .D(n1771), .CLK(clk), .Q(mem[233]) );
  DFFPOSX1 mem_reg_7__1_ ( .D(n1770), .CLK(clk), .Q(mem[232]) );
  DFFPOSX1 mem_reg_7__0_ ( .D(n1769), .CLK(clk), .Q(mem[231]) );
  DFFPOSX1 mem_reg_6__32_ ( .D(n1768), .CLK(clk), .Q(mem[230]) );
  DFFPOSX1 mem_reg_6__31_ ( .D(n1767), .CLK(clk), .Q(mem[229]) );
  DFFPOSX1 mem_reg_6__30_ ( .D(n1766), .CLK(clk), .Q(mem[228]) );
  DFFPOSX1 mem_reg_6__29_ ( .D(n1765), .CLK(clk), .Q(mem[227]) );
  DFFPOSX1 mem_reg_6__28_ ( .D(n1764), .CLK(clk), .Q(mem[226]) );
  DFFPOSX1 mem_reg_6__27_ ( .D(n1763), .CLK(clk), .Q(mem[225]) );
  DFFPOSX1 mem_reg_6__26_ ( .D(n1762), .CLK(clk), .Q(mem[224]) );
  DFFPOSX1 mem_reg_6__25_ ( .D(n1761), .CLK(clk), .Q(mem[223]) );
  DFFPOSX1 mem_reg_6__24_ ( .D(n1760), .CLK(clk), .Q(mem[222]) );
  DFFPOSX1 mem_reg_6__23_ ( .D(n1759), .CLK(clk), .Q(mem[221]) );
  DFFPOSX1 mem_reg_6__22_ ( .D(n1758), .CLK(clk), .Q(mem[220]) );
  DFFPOSX1 mem_reg_6__21_ ( .D(n1757), .CLK(clk), .Q(mem[219]) );
  DFFPOSX1 mem_reg_6__20_ ( .D(n1756), .CLK(clk), .Q(mem[218]) );
  DFFPOSX1 mem_reg_6__19_ ( .D(n1755), .CLK(clk), .Q(mem[217]) );
  DFFPOSX1 mem_reg_6__18_ ( .D(n1754), .CLK(clk), .Q(mem[216]) );
  DFFPOSX1 mem_reg_6__17_ ( .D(n1753), .CLK(clk), .Q(mem[215]) );
  DFFPOSX1 mem_reg_6__16_ ( .D(n1752), .CLK(clk), .Q(mem[214]) );
  DFFPOSX1 mem_reg_6__15_ ( .D(n1751), .CLK(clk), .Q(mem[213]) );
  DFFPOSX1 mem_reg_6__14_ ( .D(n1750), .CLK(clk), .Q(mem[212]) );
  DFFPOSX1 mem_reg_6__13_ ( .D(n1749), .CLK(clk), .Q(mem[211]) );
  DFFPOSX1 mem_reg_6__12_ ( .D(n1748), .CLK(clk), .Q(mem[210]) );
  DFFPOSX1 mem_reg_6__11_ ( .D(n1747), .CLK(clk), .Q(mem[209]) );
  DFFPOSX1 mem_reg_6__10_ ( .D(n1746), .CLK(clk), .Q(mem[208]) );
  DFFPOSX1 mem_reg_6__9_ ( .D(n1745), .CLK(clk), .Q(mem[207]) );
  DFFPOSX1 mem_reg_6__8_ ( .D(n1744), .CLK(clk), .Q(mem[206]) );
  DFFPOSX1 mem_reg_6__7_ ( .D(n1743), .CLK(clk), .Q(mem[205]) );
  DFFPOSX1 mem_reg_6__6_ ( .D(n1742), .CLK(clk), .Q(mem[204]) );
  DFFPOSX1 mem_reg_6__5_ ( .D(n1741), .CLK(clk), .Q(mem[203]) );
  DFFPOSX1 mem_reg_6__4_ ( .D(n1740), .CLK(clk), .Q(mem[202]) );
  DFFPOSX1 mem_reg_6__3_ ( .D(n1739), .CLK(clk), .Q(mem[201]) );
  DFFPOSX1 mem_reg_6__2_ ( .D(n1738), .CLK(clk), .Q(mem[200]) );
  DFFPOSX1 mem_reg_6__1_ ( .D(n1737), .CLK(clk), .Q(mem[199]) );
  DFFPOSX1 mem_reg_6__0_ ( .D(n1736), .CLK(clk), .Q(mem[198]) );
  DFFPOSX1 mem_reg_5__32_ ( .D(n1735), .CLK(clk), .Q(mem[197]) );
  DFFPOSX1 mem_reg_5__31_ ( .D(n1734), .CLK(clk), .Q(mem[196]) );
  DFFPOSX1 mem_reg_5__30_ ( .D(n1733), .CLK(clk), .Q(mem[195]) );
  DFFPOSX1 mem_reg_5__29_ ( .D(n1732), .CLK(clk), .Q(mem[194]) );
  DFFPOSX1 mem_reg_5__28_ ( .D(n1731), .CLK(clk), .Q(mem[193]) );
  DFFPOSX1 mem_reg_5__27_ ( .D(n1730), .CLK(clk), .Q(mem[192]) );
  DFFPOSX1 mem_reg_5__26_ ( .D(n1729), .CLK(clk), .Q(mem[191]) );
  DFFPOSX1 mem_reg_5__25_ ( .D(n1728), .CLK(clk), .Q(mem[190]) );
  DFFPOSX1 mem_reg_5__24_ ( .D(n1727), .CLK(clk), .Q(mem[189]) );
  DFFPOSX1 mem_reg_5__23_ ( .D(n1726), .CLK(clk), .Q(mem[188]) );
  DFFPOSX1 mem_reg_5__22_ ( .D(n1725), .CLK(clk), .Q(mem[187]) );
  DFFPOSX1 mem_reg_5__21_ ( .D(n1724), .CLK(clk), .Q(mem[186]) );
  DFFPOSX1 mem_reg_5__20_ ( .D(n1723), .CLK(clk), .Q(mem[185]) );
  DFFPOSX1 mem_reg_5__19_ ( .D(n1722), .CLK(clk), .Q(mem[184]) );
  DFFPOSX1 mem_reg_5__18_ ( .D(n1721), .CLK(clk), .Q(mem[183]) );
  DFFPOSX1 mem_reg_5__17_ ( .D(n1720), .CLK(clk), .Q(mem[182]) );
  DFFPOSX1 mem_reg_5__16_ ( .D(n1719), .CLK(clk), .Q(mem[181]) );
  DFFPOSX1 mem_reg_5__15_ ( .D(n1718), .CLK(clk), .Q(mem[180]) );
  DFFPOSX1 mem_reg_5__14_ ( .D(n1717), .CLK(clk), .Q(mem[179]) );
  DFFPOSX1 mem_reg_5__13_ ( .D(n1716), .CLK(clk), .Q(mem[178]) );
  DFFPOSX1 mem_reg_5__12_ ( .D(n1715), .CLK(clk), .Q(mem[177]) );
  DFFPOSX1 mem_reg_5__11_ ( .D(n1714), .CLK(clk), .Q(mem[176]) );
  DFFPOSX1 mem_reg_5__10_ ( .D(n1713), .CLK(clk), .Q(mem[175]) );
  DFFPOSX1 mem_reg_5__9_ ( .D(n1712), .CLK(clk), .Q(mem[174]) );
  DFFPOSX1 mem_reg_5__8_ ( .D(n1711), .CLK(clk), .Q(mem[173]) );
  DFFPOSX1 mem_reg_5__7_ ( .D(n1710), .CLK(clk), .Q(mem[172]) );
  DFFPOSX1 mem_reg_5__6_ ( .D(n1709), .CLK(clk), .Q(mem[171]) );
  DFFPOSX1 mem_reg_5__5_ ( .D(n1708), .CLK(clk), .Q(mem[170]) );
  DFFPOSX1 mem_reg_5__4_ ( .D(n1707), .CLK(clk), .Q(mem[169]) );
  DFFPOSX1 mem_reg_5__3_ ( .D(n1706), .CLK(clk), .Q(mem[168]) );
  DFFPOSX1 mem_reg_5__2_ ( .D(n1705), .CLK(clk), .Q(mem[167]) );
  DFFPOSX1 mem_reg_5__1_ ( .D(n1704), .CLK(clk), .Q(mem[166]) );
  DFFPOSX1 mem_reg_5__0_ ( .D(n1703), .CLK(clk), .Q(mem[165]) );
  DFFPOSX1 mem_reg_4__32_ ( .D(n1702), .CLK(clk), .Q(mem[164]) );
  DFFPOSX1 mem_reg_4__31_ ( .D(n1701), .CLK(clk), .Q(mem[163]) );
  DFFPOSX1 mem_reg_4__30_ ( .D(n1700), .CLK(clk), .Q(mem[162]) );
  DFFPOSX1 mem_reg_4__29_ ( .D(n1699), .CLK(clk), .Q(mem[161]) );
  DFFPOSX1 mem_reg_4__28_ ( .D(n1698), .CLK(clk), .Q(mem[160]) );
  DFFPOSX1 mem_reg_4__27_ ( .D(n1697), .CLK(clk), .Q(mem[159]) );
  DFFPOSX1 mem_reg_4__26_ ( .D(n1696), .CLK(clk), .Q(mem[158]) );
  DFFPOSX1 mem_reg_4__25_ ( .D(n1695), .CLK(clk), .Q(mem[157]) );
  DFFPOSX1 mem_reg_4__24_ ( .D(n1694), .CLK(clk), .Q(mem[156]) );
  DFFPOSX1 mem_reg_4__23_ ( .D(n1693), .CLK(clk), .Q(mem[155]) );
  DFFPOSX1 mem_reg_4__22_ ( .D(n1692), .CLK(clk), .Q(mem[154]) );
  DFFPOSX1 mem_reg_4__21_ ( .D(n1691), .CLK(clk), .Q(mem[153]) );
  DFFPOSX1 mem_reg_4__20_ ( .D(n1690), .CLK(clk), .Q(mem[152]) );
  DFFPOSX1 mem_reg_4__19_ ( .D(n1689), .CLK(clk), .Q(mem[151]) );
  DFFPOSX1 mem_reg_4__18_ ( .D(n1688), .CLK(clk), .Q(mem[150]) );
  DFFPOSX1 mem_reg_4__17_ ( .D(n1687), .CLK(clk), .Q(mem[149]) );
  DFFPOSX1 mem_reg_4__16_ ( .D(n1686), .CLK(clk), .Q(mem[148]) );
  DFFPOSX1 mem_reg_4__15_ ( .D(n1685), .CLK(clk), .Q(mem[147]) );
  DFFPOSX1 mem_reg_4__14_ ( .D(n1684), .CLK(clk), .Q(mem[146]) );
  DFFPOSX1 mem_reg_4__13_ ( .D(n1683), .CLK(clk), .Q(mem[145]) );
  DFFPOSX1 mem_reg_4__12_ ( .D(n1682), .CLK(clk), .Q(mem[144]) );
  DFFPOSX1 mem_reg_4__11_ ( .D(n1681), .CLK(clk), .Q(mem[143]) );
  DFFPOSX1 mem_reg_4__10_ ( .D(n1680), .CLK(clk), .Q(mem[142]) );
  DFFPOSX1 mem_reg_4__9_ ( .D(n1679), .CLK(clk), .Q(mem[141]) );
  DFFPOSX1 mem_reg_4__8_ ( .D(n1678), .CLK(clk), .Q(mem[140]) );
  DFFPOSX1 mem_reg_4__7_ ( .D(n1677), .CLK(clk), .Q(mem[139]) );
  DFFPOSX1 mem_reg_4__6_ ( .D(n1676), .CLK(clk), .Q(mem[138]) );
  DFFPOSX1 mem_reg_4__5_ ( .D(n1675), .CLK(clk), .Q(mem[137]) );
  DFFPOSX1 mem_reg_4__4_ ( .D(n1674), .CLK(clk), .Q(mem[136]) );
  DFFPOSX1 mem_reg_4__3_ ( .D(n1673), .CLK(clk), .Q(mem[135]) );
  DFFPOSX1 mem_reg_4__2_ ( .D(n1672), .CLK(clk), .Q(mem[134]) );
  DFFPOSX1 mem_reg_4__1_ ( .D(n1671), .CLK(clk), .Q(mem[133]) );
  DFFPOSX1 mem_reg_4__0_ ( .D(n1670), .CLK(clk), .Q(mem[132]) );
  DFFPOSX1 mem_reg_3__32_ ( .D(n1669), .CLK(clk), .Q(mem[131]) );
  DFFPOSX1 mem_reg_3__31_ ( .D(n1668), .CLK(clk), .Q(mem[130]) );
  DFFPOSX1 mem_reg_3__30_ ( .D(n1667), .CLK(clk), .Q(mem[129]) );
  DFFPOSX1 mem_reg_3__29_ ( .D(n1666), .CLK(clk), .Q(mem[128]) );
  DFFPOSX1 mem_reg_3__28_ ( .D(n1665), .CLK(clk), .Q(mem[127]) );
  DFFPOSX1 mem_reg_3__27_ ( .D(n1664), .CLK(clk), .Q(mem[126]) );
  DFFPOSX1 mem_reg_3__26_ ( .D(n1663), .CLK(clk), .Q(mem[125]) );
  DFFPOSX1 mem_reg_3__25_ ( .D(n1662), .CLK(clk), .Q(mem[124]) );
  DFFPOSX1 mem_reg_3__24_ ( .D(n1661), .CLK(clk), .Q(mem[123]) );
  DFFPOSX1 mem_reg_3__23_ ( .D(n1660), .CLK(clk), .Q(mem[122]) );
  DFFPOSX1 mem_reg_3__22_ ( .D(n1659), .CLK(clk), .Q(mem[121]) );
  DFFPOSX1 mem_reg_3__21_ ( .D(n1658), .CLK(clk), .Q(mem[120]) );
  DFFPOSX1 mem_reg_3__20_ ( .D(n1657), .CLK(clk), .Q(mem[119]) );
  DFFPOSX1 mem_reg_3__19_ ( .D(n1656), .CLK(clk), .Q(mem[118]) );
  DFFPOSX1 mem_reg_3__18_ ( .D(n1655), .CLK(clk), .Q(mem[117]) );
  DFFPOSX1 mem_reg_3__17_ ( .D(n1654), .CLK(clk), .Q(mem[116]) );
  DFFPOSX1 mem_reg_3__16_ ( .D(n1653), .CLK(clk), .Q(mem[115]) );
  DFFPOSX1 mem_reg_3__15_ ( .D(n1652), .CLK(clk), .Q(mem[114]) );
  DFFPOSX1 mem_reg_3__14_ ( .D(n1651), .CLK(clk), .Q(mem[113]) );
  DFFPOSX1 mem_reg_3__13_ ( .D(n1650), .CLK(clk), .Q(mem[112]) );
  DFFPOSX1 mem_reg_3__12_ ( .D(n1649), .CLK(clk), .Q(mem[111]) );
  DFFPOSX1 mem_reg_3__11_ ( .D(n1648), .CLK(clk), .Q(mem[110]) );
  DFFPOSX1 mem_reg_3__10_ ( .D(n1647), .CLK(clk), .Q(mem[109]) );
  DFFPOSX1 mem_reg_3__9_ ( .D(n1646), .CLK(clk), .Q(mem[108]) );
  DFFPOSX1 mem_reg_3__8_ ( .D(n1645), .CLK(clk), .Q(mem[107]) );
  DFFPOSX1 mem_reg_3__7_ ( .D(n1644), .CLK(clk), .Q(mem[106]) );
  DFFPOSX1 mem_reg_3__6_ ( .D(n1643), .CLK(clk), .Q(mem[105]) );
  DFFPOSX1 mem_reg_3__5_ ( .D(n1642), .CLK(clk), .Q(mem[104]) );
  DFFPOSX1 mem_reg_3__4_ ( .D(n1641), .CLK(clk), .Q(mem[103]) );
  DFFPOSX1 mem_reg_3__3_ ( .D(n1640), .CLK(clk), .Q(mem[102]) );
  DFFPOSX1 mem_reg_3__2_ ( .D(n1639), .CLK(clk), .Q(mem[101]) );
  DFFPOSX1 mem_reg_3__1_ ( .D(n1638), .CLK(clk), .Q(mem[100]) );
  DFFPOSX1 mem_reg_3__0_ ( .D(n1637), .CLK(clk), .Q(mem[99]) );
  DFFPOSX1 mem_reg_2__32_ ( .D(n1636), .CLK(clk), .Q(mem[98]) );
  DFFPOSX1 mem_reg_2__31_ ( .D(n1635), .CLK(clk), .Q(mem[97]) );
  DFFPOSX1 mem_reg_2__30_ ( .D(n1634), .CLK(clk), .Q(mem[96]) );
  DFFPOSX1 mem_reg_2__29_ ( .D(n1633), .CLK(clk), .Q(mem[95]) );
  DFFPOSX1 mem_reg_2__28_ ( .D(n1632), .CLK(clk), .Q(mem[94]) );
  DFFPOSX1 mem_reg_2__27_ ( .D(n1631), .CLK(clk), .Q(mem[93]) );
  DFFPOSX1 mem_reg_2__26_ ( .D(n1630), .CLK(clk), .Q(mem[92]) );
  DFFPOSX1 mem_reg_2__25_ ( .D(n1629), .CLK(clk), .Q(mem[91]) );
  DFFPOSX1 mem_reg_2__24_ ( .D(n1628), .CLK(clk), .Q(mem[90]) );
  DFFPOSX1 mem_reg_2__23_ ( .D(n1627), .CLK(clk), .Q(mem[89]) );
  DFFPOSX1 mem_reg_2__22_ ( .D(n1626), .CLK(clk), .Q(mem[88]) );
  DFFPOSX1 mem_reg_2__21_ ( .D(n1625), .CLK(clk), .Q(mem[87]) );
  DFFPOSX1 mem_reg_2__20_ ( .D(n1624), .CLK(clk), .Q(mem[86]) );
  DFFPOSX1 mem_reg_2__19_ ( .D(n1623), .CLK(clk), .Q(mem[85]) );
  DFFPOSX1 mem_reg_2__18_ ( .D(n1622), .CLK(clk), .Q(mem[84]) );
  DFFPOSX1 mem_reg_2__17_ ( .D(n1621), .CLK(clk), .Q(mem[83]) );
  DFFPOSX1 mem_reg_2__16_ ( .D(n1620), .CLK(clk), .Q(mem[82]) );
  DFFPOSX1 mem_reg_2__15_ ( .D(n1619), .CLK(clk), .Q(mem[81]) );
  DFFPOSX1 mem_reg_2__14_ ( .D(n1618), .CLK(clk), .Q(mem[80]) );
  DFFPOSX1 mem_reg_2__13_ ( .D(n1617), .CLK(clk), .Q(mem[79]) );
  DFFPOSX1 mem_reg_2__12_ ( .D(n1616), .CLK(clk), .Q(mem[78]) );
  DFFPOSX1 mem_reg_2__11_ ( .D(n1615), .CLK(clk), .Q(mem[77]) );
  DFFPOSX1 mem_reg_2__10_ ( .D(n1614), .CLK(clk), .Q(mem[76]) );
  DFFPOSX1 mem_reg_2__9_ ( .D(n1613), .CLK(clk), .Q(mem[75]) );
  DFFPOSX1 mem_reg_2__8_ ( .D(n1612), .CLK(clk), .Q(mem[74]) );
  DFFPOSX1 mem_reg_2__7_ ( .D(n1611), .CLK(clk), .Q(mem[73]) );
  DFFPOSX1 mem_reg_2__6_ ( .D(n1610), .CLK(clk), .Q(mem[72]) );
  DFFPOSX1 mem_reg_2__5_ ( .D(n1609), .CLK(clk), .Q(mem[71]) );
  DFFPOSX1 mem_reg_2__4_ ( .D(n1608), .CLK(clk), .Q(mem[70]) );
  DFFPOSX1 mem_reg_2__3_ ( .D(n1607), .CLK(clk), .Q(mem[69]) );
  DFFPOSX1 mem_reg_2__2_ ( .D(n1606), .CLK(clk), .Q(mem[68]) );
  DFFPOSX1 mem_reg_2__1_ ( .D(n1605), .CLK(clk), .Q(mem[67]) );
  DFFPOSX1 mem_reg_2__0_ ( .D(n1604), .CLK(clk), .Q(mem[66]) );
  DFFPOSX1 mem_reg_1__32_ ( .D(n1603), .CLK(clk), .Q(mem[65]) );
  DFFPOSX1 mem_reg_1__31_ ( .D(n1602), .CLK(clk), .Q(mem[64]) );
  DFFPOSX1 mem_reg_1__30_ ( .D(n1601), .CLK(clk), .Q(mem[63]) );
  DFFPOSX1 mem_reg_1__29_ ( .D(n1600), .CLK(clk), .Q(mem[62]) );
  DFFPOSX1 mem_reg_1__28_ ( .D(n1599), .CLK(clk), .Q(mem[61]) );
  DFFPOSX1 mem_reg_1__27_ ( .D(n1598), .CLK(clk), .Q(mem[60]) );
  DFFPOSX1 mem_reg_1__26_ ( .D(n1597), .CLK(clk), .Q(mem[59]) );
  DFFPOSX1 mem_reg_1__25_ ( .D(n1596), .CLK(clk), .Q(mem[58]) );
  DFFPOSX1 mem_reg_1__24_ ( .D(n1595), .CLK(clk), .Q(mem[57]) );
  DFFPOSX1 mem_reg_1__23_ ( .D(n1594), .CLK(clk), .Q(mem[56]) );
  DFFPOSX1 mem_reg_1__22_ ( .D(n1593), .CLK(clk), .Q(mem[55]) );
  DFFPOSX1 mem_reg_1__21_ ( .D(n1592), .CLK(clk), .Q(mem[54]) );
  DFFPOSX1 mem_reg_1__20_ ( .D(n1591), .CLK(clk), .Q(mem[53]) );
  DFFPOSX1 mem_reg_1__19_ ( .D(n1590), .CLK(clk), .Q(mem[52]) );
  DFFPOSX1 mem_reg_1__18_ ( .D(n1589), .CLK(clk), .Q(mem[51]) );
  DFFPOSX1 mem_reg_1__17_ ( .D(n1588), .CLK(clk), .Q(mem[50]) );
  DFFPOSX1 mem_reg_1__16_ ( .D(n1587), .CLK(clk), .Q(mem[49]) );
  DFFPOSX1 mem_reg_1__15_ ( .D(n1586), .CLK(clk), .Q(mem[48]) );
  DFFPOSX1 mem_reg_1__14_ ( .D(n1585), .CLK(clk), .Q(mem[47]) );
  DFFPOSX1 mem_reg_1__13_ ( .D(n1584), .CLK(clk), .Q(mem[46]) );
  DFFPOSX1 mem_reg_1__12_ ( .D(n1583), .CLK(clk), .Q(mem[45]) );
  DFFPOSX1 mem_reg_1__11_ ( .D(n1582), .CLK(clk), .Q(mem[44]) );
  DFFPOSX1 mem_reg_1__10_ ( .D(n1581), .CLK(clk), .Q(mem[43]) );
  DFFPOSX1 mem_reg_1__9_ ( .D(n1580), .CLK(clk), .Q(mem[42]) );
  DFFPOSX1 mem_reg_1__8_ ( .D(n1579), .CLK(clk), .Q(mem[41]) );
  DFFPOSX1 mem_reg_1__7_ ( .D(n1578), .CLK(clk), .Q(mem[40]) );
  DFFPOSX1 mem_reg_1__6_ ( .D(n1577), .CLK(clk), .Q(mem[39]) );
  DFFPOSX1 mem_reg_1__5_ ( .D(n1576), .CLK(clk), .Q(mem[38]) );
  DFFPOSX1 mem_reg_1__4_ ( .D(n1575), .CLK(clk), .Q(mem[37]) );
  DFFPOSX1 mem_reg_1__3_ ( .D(n1574), .CLK(clk), .Q(mem[36]) );
  DFFPOSX1 mem_reg_1__2_ ( .D(n1573), .CLK(clk), .Q(mem[35]) );
  DFFPOSX1 mem_reg_1__1_ ( .D(n1572), .CLK(clk), .Q(mem[34]) );
  DFFPOSX1 mem_reg_1__0_ ( .D(n1571), .CLK(clk), .Q(mem[33]) );
  DFFPOSX1 mem_reg_0__32_ ( .D(n1570), .CLK(clk), .Q(mem[32]) );
  DFFPOSX1 mem_reg_0__31_ ( .D(n1569), .CLK(clk), .Q(mem[31]) );
  DFFPOSX1 mem_reg_0__30_ ( .D(n1568), .CLK(clk), .Q(mem[30]) );
  DFFPOSX1 mem_reg_0__29_ ( .D(n1567), .CLK(clk), .Q(mem[29]) );
  DFFPOSX1 mem_reg_0__28_ ( .D(n1566), .CLK(clk), .Q(mem[28]) );
  DFFPOSX1 mem_reg_0__27_ ( .D(n1565), .CLK(clk), .Q(mem[27]) );
  DFFPOSX1 mem_reg_0__26_ ( .D(n1564), .CLK(clk), .Q(mem[26]) );
  DFFPOSX1 mem_reg_0__25_ ( .D(n1563), .CLK(clk), .Q(mem[25]) );
  DFFPOSX1 mem_reg_0__24_ ( .D(n1562), .CLK(clk), .Q(mem[24]) );
  DFFPOSX1 mem_reg_0__23_ ( .D(n1561), .CLK(clk), .Q(mem[23]) );
  DFFPOSX1 mem_reg_0__22_ ( .D(n1560), .CLK(clk), .Q(mem[22]) );
  DFFPOSX1 mem_reg_0__21_ ( .D(n1559), .CLK(clk), .Q(mem[21]) );
  DFFPOSX1 mem_reg_0__20_ ( .D(n1558), .CLK(clk), .Q(mem[20]) );
  DFFPOSX1 mem_reg_0__19_ ( .D(n1557), .CLK(clk), .Q(mem[19]) );
  DFFPOSX1 mem_reg_0__18_ ( .D(n1556), .CLK(clk), .Q(mem[18]) );
  DFFPOSX1 mem_reg_0__17_ ( .D(n1555), .CLK(clk), .Q(mem[17]) );
  DFFPOSX1 mem_reg_0__16_ ( .D(n1554), .CLK(clk), .Q(mem[16]) );
  DFFPOSX1 mem_reg_0__15_ ( .D(n1553), .CLK(clk), .Q(mem[15]) );
  DFFPOSX1 mem_reg_0__14_ ( .D(n1552), .CLK(clk), .Q(mem[14]) );
  DFFPOSX1 mem_reg_0__13_ ( .D(n1551), .CLK(clk), .Q(mem[13]) );
  DFFPOSX1 mem_reg_0__12_ ( .D(n1550), .CLK(clk), .Q(mem[12]) );
  DFFPOSX1 mem_reg_0__11_ ( .D(n1549), .CLK(clk), .Q(mem[11]) );
  DFFPOSX1 mem_reg_0__10_ ( .D(n1548), .CLK(clk), .Q(mem[10]) );
  DFFPOSX1 mem_reg_0__9_ ( .D(n1547), .CLK(clk), .Q(mem[9]) );
  DFFPOSX1 mem_reg_0__8_ ( .D(n1546), .CLK(clk), .Q(mem[8]) );
  DFFPOSX1 mem_reg_0__7_ ( .D(n1545), .CLK(clk), .Q(mem[7]) );
  DFFPOSX1 mem_reg_0__6_ ( .D(n1544), .CLK(clk), .Q(mem[6]) );
  DFFPOSX1 mem_reg_0__5_ ( .D(n1543), .CLK(clk), .Q(mem[5]) );
  DFFPOSX1 mem_reg_0__4_ ( .D(n1542), .CLK(clk), .Q(mem[4]) );
  DFFPOSX1 mem_reg_0__3_ ( .D(n1541), .CLK(clk), .Q(mem[3]) );
  DFFPOSX1 mem_reg_0__2_ ( .D(n1540), .CLK(clk), .Q(mem[2]) );
  DFFPOSX1 mem_reg_0__1_ ( .D(n1539), .CLK(clk), .Q(mem[1]) );
  DFFPOSX1 mem_reg_0__0_ ( .D(n1538), .CLK(clk), .Q(mem[0]) );
  NAND3X1 U1161 ( .A(n5187), .B(n1087), .C(n1088), .Y(n4460) );
  NOR3X1 U1162 ( .A(n5750), .B(n5783), .C(n5816), .Y(n1088) );
  NAND3X1 U1164 ( .A(n3260), .B(n5452), .C(n5717), .Y(n1093) );
  AOI22X1 U1165 ( .A(n6837), .B(n7258), .C(n6836), .D(n7159), .Y(n1095) );
  NAND3X1 U1167 ( .A(n5153), .B(n5451), .C(n5716), .Y(n1092) );
  AOI22X1 U1168 ( .A(n1101), .B(n7324), .C(n1102), .D(n7192), .Y(n1100) );
  AOI22X1 U1170 ( .A(n1104), .B(n7357), .C(n1105), .D(n7291), .Y(n1098) );
  NAND3X1 U1172 ( .A(n1108), .B(n5450), .C(n5715), .Y(n1107) );
  AOI22X1 U1173 ( .A(n6837), .B(n6994), .C(n6836), .D(n6895), .Y(n1110) );
  NAND3X1 U1175 ( .A(n5152), .B(n5449), .C(n5714), .Y(n1106) );
  AOI22X1 U1176 ( .A(n1101), .B(n7060), .C(n1102), .D(n6928), .Y(n1113) );
  AOI22X1 U1178 ( .A(n1104), .B(n7093), .C(n1105), .D(n7027), .Y(n1111) );
  NAND3X1 U1180 ( .A(n1116), .B(n5448), .C(n5713), .Y(n1115) );
  AOI22X1 U1181 ( .A(n6837), .B(n7786), .C(n6835), .D(n7687), .Y(n1118) );
  NAND3X1 U1183 ( .A(n5151), .B(n5447), .C(n5712), .Y(n1114) );
  AOI22X1 U1184 ( .A(n6830), .B(n7852), .C(n1102), .D(n7720), .Y(n1121) );
  AOI22X1 U1186 ( .A(n6817), .B(n7885), .C(n1105), .D(n7819), .Y(n1119) );
  NAND3X1 U1187 ( .A(n1124), .B(n5446), .C(n5711), .Y(n1123) );
  AOI22X1 U1188 ( .A(n6837), .B(n7522), .C(n1097), .D(n7423), .Y(n1126) );
  NAND3X1 U1190 ( .A(n5150), .B(n5445), .C(n5710), .Y(n1122) );
  AOI22X1 U1191 ( .A(n1101), .B(n7588), .C(n1102), .D(n7456), .Y(n1129) );
  AOI22X1 U1193 ( .A(n1104), .B(n7621), .C(n1105), .D(n7555), .Y(n1127) );
  NAND3X1 U1195 ( .A(n5186), .B(n1131), .C(n1132), .Y(n4461) );
  NOR3X1 U1196 ( .A(n5749), .B(n5782), .C(n5815), .Y(n1132) );
  NAND3X1 U1198 ( .A(n3260), .B(n5444), .C(n5709), .Y(n1137) );
  AOI22X1 U1199 ( .A(n6837), .B(n7260), .C(n1097), .D(n7161), .Y(n1139) );
  NAND3X1 U1201 ( .A(n5149), .B(n5443), .C(n5708), .Y(n1136) );
  AOI22X1 U1202 ( .A(n1101), .B(n7326), .C(n1102), .D(n7194), .Y(n1142) );
  AOI22X1 U1204 ( .A(n1104), .B(n7359), .C(n1105), .D(n7293), .Y(n1140) );
  NAND3X1 U1206 ( .A(n1108), .B(n5442), .C(n5707), .Y(n1144) );
  AOI22X1 U1207 ( .A(n6837), .B(n6996), .C(n6835), .D(n6897), .Y(n1146) );
  NAND3X1 U1209 ( .A(n5148), .B(n5441), .C(n5706), .Y(n1143) );
  AOI22X1 U1210 ( .A(n1101), .B(n7062), .C(n1102), .D(n6930), .Y(n1149) );
  AOI22X1 U1212 ( .A(n1104), .B(n7095), .C(n1105), .D(n7029), .Y(n1147) );
  NAND3X1 U1214 ( .A(n1116), .B(n5440), .C(n5705), .Y(n1151) );
  AOI22X1 U1215 ( .A(n6837), .B(n7788), .C(n6833), .D(n7689), .Y(n1153) );
  NAND3X1 U1217 ( .A(n5147), .B(n5439), .C(n5704), .Y(n1150) );
  AOI22X1 U1218 ( .A(n6829), .B(n7854), .C(n1102), .D(n7722), .Y(n1156) );
  AOI22X1 U1220 ( .A(n6818), .B(n7887), .C(n1105), .D(n7821), .Y(n1154) );
  NAND3X1 U1221 ( .A(n1124), .B(n5438), .C(n5703), .Y(n1158) );
  AOI22X1 U1222 ( .A(n6837), .B(n7524), .C(n1097), .D(n7425), .Y(n1160) );
  NAND3X1 U1224 ( .A(n5146), .B(n5437), .C(n5702), .Y(n1157) );
  AOI22X1 U1225 ( .A(n1101), .B(n7590), .C(n1102), .D(n7458), .Y(n1163) );
  AOI22X1 U1227 ( .A(n1104), .B(n7623), .C(n1105), .D(n7557), .Y(n1161) );
  NAND3X1 U1229 ( .A(n5185), .B(n1165), .C(n1166), .Y(n4462) );
  NOR3X1 U1230 ( .A(n5748), .B(n5781), .C(n5814), .Y(n1166) );
  NAND3X1 U1232 ( .A(n3260), .B(n5436), .C(n5701), .Y(n1171) );
  AOI22X1 U1233 ( .A(n6837), .B(n7262), .C(n6833), .D(n7163), .Y(n1173) );
  NAND3X1 U1235 ( .A(n5145), .B(n5435), .C(n5700), .Y(n1170) );
  AOI22X1 U1236 ( .A(n1101), .B(n7328), .C(n1102), .D(n7196), .Y(n1176) );
  AOI22X1 U1238 ( .A(n1104), .B(n7361), .C(n1105), .D(n7295), .Y(n1174) );
  NAND3X1 U1240 ( .A(n1108), .B(n5434), .C(n5699), .Y(n1178) );
  AOI22X1 U1241 ( .A(n6837), .B(n6998), .C(n6836), .D(n6899), .Y(n1180) );
  NAND3X1 U1243 ( .A(n5144), .B(n5433), .C(n5698), .Y(n1177) );
  AOI22X1 U1244 ( .A(n1101), .B(n7064), .C(n1102), .D(n6932), .Y(n1183) );
  AOI22X1 U1246 ( .A(n1104), .B(n7097), .C(n1105), .D(n7031), .Y(n1181) );
  NAND3X1 U1248 ( .A(n1116), .B(n5432), .C(n5697), .Y(n1185) );
  AOI22X1 U1249 ( .A(n6837), .B(n7790), .C(n6834), .D(n7691), .Y(n1187) );
  NAND3X1 U1251 ( .A(n5143), .B(n5431), .C(n5696), .Y(n1184) );
  AOI22X1 U1252 ( .A(n6830), .B(n7856), .C(n1102), .D(n7724), .Y(n1190) );
  AOI22X1 U1254 ( .A(n6818), .B(n7889), .C(n1105), .D(n7823), .Y(n1188) );
  NAND3X1 U1255 ( .A(n1124), .B(n5430), .C(n5695), .Y(n1192) );
  AOI22X1 U1256 ( .A(n6837), .B(n7526), .C(n1097), .D(n7427), .Y(n1194) );
  NAND3X1 U1258 ( .A(n5142), .B(n5429), .C(n5694), .Y(n1191) );
  AOI22X1 U1259 ( .A(n1101), .B(n7592), .C(n1102), .D(n7460), .Y(n1197) );
  AOI22X1 U1261 ( .A(n1104), .B(n7625), .C(n1105), .D(n7559), .Y(n1195) );
  NAND3X1 U1263 ( .A(n5184), .B(n1199), .C(n1200), .Y(n4463) );
  NOR3X1 U1264 ( .A(n5747), .B(n5780), .C(n5813), .Y(n1200) );
  NAND3X1 U1266 ( .A(n3260), .B(n5428), .C(n5693), .Y(n1205) );
  AOI22X1 U1267 ( .A(n6837), .B(n7264), .C(n6833), .D(n7165), .Y(n1207) );
  NAND3X1 U1269 ( .A(n5141), .B(n5427), .C(n5692), .Y(n1204) );
  AOI22X1 U1270 ( .A(n1101), .B(n7330), .C(n1102), .D(n7198), .Y(n1210) );
  AOI22X1 U1272 ( .A(n1104), .B(n7363), .C(n1105), .D(n7297), .Y(n1208) );
  NAND3X1 U1274 ( .A(n1108), .B(n5426), .C(n5691), .Y(n1212) );
  AOI22X1 U1275 ( .A(n6840), .B(n7000), .C(n6836), .D(n6901), .Y(n1214) );
  NAND3X1 U1277 ( .A(n5140), .B(n5425), .C(n5690), .Y(n1211) );
  AOI22X1 U1278 ( .A(n6830), .B(n7066), .C(n1102), .D(n6934), .Y(n1217) );
  AOI22X1 U1280 ( .A(n6817), .B(n7099), .C(n1105), .D(n7033), .Y(n1215) );
  NAND3X1 U1282 ( .A(n1116), .B(n5424), .C(n5689), .Y(n1219) );
  AOI22X1 U1283 ( .A(n6838), .B(n7792), .C(n6833), .D(n7693), .Y(n1221) );
  NAND3X1 U1285 ( .A(n5139), .B(n5423), .C(n5688), .Y(n1218) );
  AOI22X1 U1286 ( .A(n6828), .B(n7858), .C(n1102), .D(n7726), .Y(n1224) );
  AOI22X1 U1288 ( .A(n6818), .B(n7891), .C(n1105), .D(n7825), .Y(n1222) );
  NAND3X1 U1289 ( .A(n1124), .B(n5422), .C(n5687), .Y(n1226) );
  AOI22X1 U1290 ( .A(n1096), .B(n7528), .C(n1097), .D(n7429), .Y(n1228) );
  NAND3X1 U1292 ( .A(n5138), .B(n5421), .C(n5686), .Y(n1225) );
  AOI22X1 U1293 ( .A(n6828), .B(n7594), .C(n1102), .D(n7462), .Y(n1231) );
  AOI22X1 U1295 ( .A(n1104), .B(n7627), .C(n1105), .D(n7561), .Y(n1229) );
  NAND3X1 U1297 ( .A(n5183), .B(n1233), .C(n1234), .Y(n4464) );
  NOR3X1 U1298 ( .A(n5746), .B(n5779), .C(n5812), .Y(n1234) );
  NAND3X1 U1300 ( .A(n3260), .B(n5420), .C(n5685), .Y(n1239) );
  AOI22X1 U1301 ( .A(n6838), .B(n7266), .C(n6834), .D(n7167), .Y(n1241) );
  NAND3X1 U1303 ( .A(n5137), .B(n5419), .C(n5684), .Y(n1238) );
  AOI22X1 U1304 ( .A(n6829), .B(n7332), .C(n1102), .D(n7200), .Y(n1244) );
  AOI22X1 U1306 ( .A(n1104), .B(n7365), .C(n1105), .D(n7299), .Y(n1242) );
  NAND3X1 U1308 ( .A(n1108), .B(n5418), .C(n5683), .Y(n1246) );
  AOI22X1 U1309 ( .A(n1096), .B(n7002), .C(n6833), .D(n6903), .Y(n1248) );
  NAND3X1 U1311 ( .A(n5136), .B(n5417), .C(n5682), .Y(n1245) );
  AOI22X1 U1312 ( .A(n6830), .B(n7068), .C(n1102), .D(n6936), .Y(n1251) );
  AOI22X1 U1314 ( .A(n6816), .B(n7101), .C(n1105), .D(n7035), .Y(n1249) );
  NAND3X1 U1316 ( .A(n1116), .B(n5416), .C(n5681), .Y(n1253) );
  AOI22X1 U1317 ( .A(n6838), .B(n7794), .C(n6835), .D(n7695), .Y(n1255) );
  NAND3X1 U1319 ( .A(n5135), .B(n5415), .C(n5680), .Y(n1252) );
  AOI22X1 U1320 ( .A(n6829), .B(n7860), .C(n1102), .D(n7728), .Y(n1258) );
  AOI22X1 U1322 ( .A(n6816), .B(n7893), .C(n1105), .D(n7827), .Y(n1256) );
  NAND3X1 U1323 ( .A(n1124), .B(n5414), .C(n5679), .Y(n1260) );
  AOI22X1 U1324 ( .A(n6839), .B(n7530), .C(n1097), .D(n7431), .Y(n1262) );
  NAND3X1 U1326 ( .A(n5134), .B(n5413), .C(n5678), .Y(n1259) );
  AOI22X1 U1327 ( .A(n1101), .B(n7596), .C(n1102), .D(n7464), .Y(n1265) );
  AOI22X1 U1329 ( .A(n1104), .B(n7629), .C(n1105), .D(n7563), .Y(n1263) );
  NAND3X1 U1331 ( .A(n5182), .B(n1267), .C(n1268), .Y(n4465) );
  NOR3X1 U1332 ( .A(n5745), .B(n5778), .C(n5811), .Y(n1268) );
  NAND3X1 U1334 ( .A(n3260), .B(n5412), .C(n5677), .Y(n1273) );
  AOI22X1 U1335 ( .A(n6839), .B(n7267), .C(n1097), .D(n7168), .Y(n1275) );
  NAND3X1 U1337 ( .A(n5133), .B(n5411), .C(n5676), .Y(n1272) );
  AOI22X1 U1338 ( .A(n1101), .B(n7333), .C(n1102), .D(n7201), .Y(n1278) );
  AOI22X1 U1340 ( .A(n1104), .B(n7366), .C(n1105), .D(n7300), .Y(n1276) );
  NAND3X1 U1342 ( .A(n1108), .B(n5410), .C(n5675), .Y(n1280) );
  AOI22X1 U1343 ( .A(n1096), .B(n7003), .C(n6835), .D(n6904), .Y(n1282) );
  NAND3X1 U1345 ( .A(n5132), .B(n5409), .C(n5674), .Y(n1279) );
  AOI22X1 U1346 ( .A(n6828), .B(n7069), .C(n1102), .D(n6937), .Y(n1285) );
  AOI22X1 U1348 ( .A(n6818), .B(n7102), .C(n1105), .D(n7036), .Y(n1283) );
  NAND3X1 U1350 ( .A(n1116), .B(n5408), .C(n5673), .Y(n1287) );
  AOI22X1 U1351 ( .A(n1096), .B(n7795), .C(n6835), .D(n7696), .Y(n1289) );
  NAND3X1 U1353 ( .A(n5131), .B(n5407), .C(n5672), .Y(n1286) );
  AOI22X1 U1354 ( .A(n6828), .B(n7861), .C(n1102), .D(n7729), .Y(n1292) );
  AOI22X1 U1356 ( .A(n6816), .B(n7894), .C(n1105), .D(n7828), .Y(n1290) );
  NAND3X1 U1357 ( .A(n1124), .B(n5406), .C(n5671), .Y(n1294) );
  AOI22X1 U1358 ( .A(n1096), .B(n7531), .C(n1097), .D(n7432), .Y(n1296) );
  NAND3X1 U1360 ( .A(n5130), .B(n5405), .C(n5670), .Y(n1293) );
  AOI22X1 U1361 ( .A(n6828), .B(n7597), .C(n1102), .D(n7465), .Y(n1299) );
  AOI22X1 U1363 ( .A(n1104), .B(n7630), .C(n1105), .D(n7564), .Y(n1297) );
  NAND3X1 U1365 ( .A(n5181), .B(n1301), .C(n1302), .Y(n4466) );
  NOR3X1 U1366 ( .A(n5744), .B(n5777), .C(n5810), .Y(n1302) );
  NAND3X1 U1368 ( .A(n3260), .B(n5404), .C(n5669), .Y(n1307) );
  AOI22X1 U1369 ( .A(n1096), .B(n7268), .C(n1097), .D(n7169), .Y(n1309) );
  NAND3X1 U1371 ( .A(n5129), .B(n5403), .C(n5668), .Y(n1306) );
  AOI22X1 U1372 ( .A(n1101), .B(n7334), .C(n1102), .D(n7202), .Y(n1312) );
  AOI22X1 U1374 ( .A(n1104), .B(n7367), .C(n6812), .D(n7301), .Y(n1310) );
  NAND3X1 U1376 ( .A(n1108), .B(n5402), .C(n5667), .Y(n1314) );
  AOI22X1 U1377 ( .A(n6839), .B(n7004), .C(n6836), .D(n6905), .Y(n1316) );
  NAND3X1 U1379 ( .A(n5128), .B(n5401), .C(n5666), .Y(n1313) );
  AOI22X1 U1380 ( .A(n6830), .B(n7070), .C(n1102), .D(n6938), .Y(n1319) );
  AOI22X1 U1382 ( .A(n6816), .B(n7103), .C(n6813), .D(n7037), .Y(n1317) );
  NAND3X1 U1384 ( .A(n1116), .B(n5400), .C(n5665), .Y(n1321) );
  AOI22X1 U1385 ( .A(n6838), .B(n7796), .C(n6833), .D(n7697), .Y(n1323) );
  NAND3X1 U1387 ( .A(n5127), .B(n5399), .C(n5664), .Y(n1320) );
  AOI22X1 U1388 ( .A(n6828), .B(n7862), .C(n1102), .D(n7730), .Y(n1326) );
  AOI22X1 U1390 ( .A(n6816), .B(n7895), .C(n6814), .D(n7829), .Y(n1324) );
  NAND3X1 U1391 ( .A(n1124), .B(n5398), .C(n5663), .Y(n1328) );
  AOI22X1 U1392 ( .A(n6838), .B(n7532), .C(n1097), .D(n7433), .Y(n1330) );
  NAND3X1 U1394 ( .A(n5126), .B(n5397), .C(n5662), .Y(n1327) );
  AOI22X1 U1395 ( .A(n1101), .B(n7598), .C(n6826), .D(n7466), .Y(n1333) );
  AOI22X1 U1397 ( .A(n1104), .B(n7631), .C(n6813), .D(n7565), .Y(n1331) );
  NAND3X1 U1399 ( .A(n5180), .B(n1335), .C(n1336), .Y(n4467) );
  NOR3X1 U1400 ( .A(n5743), .B(n5776), .C(n5809), .Y(n1336) );
  NAND3X1 U1402 ( .A(n3260), .B(n5396), .C(n5661), .Y(n1341) );
  AOI22X1 U1403 ( .A(n6838), .B(n7269), .C(n1097), .D(n7170), .Y(n1343) );
  NAND3X1 U1405 ( .A(n5125), .B(n5395), .C(n5660), .Y(n1340) );
  AOI22X1 U1406 ( .A(n1101), .B(n7335), .C(n1102), .D(n7203), .Y(n1346) );
  AOI22X1 U1408 ( .A(n6817), .B(n7368), .C(n6814), .D(n7302), .Y(n1344) );
  NAND3X1 U1410 ( .A(n1108), .B(n5394), .C(n5659), .Y(n1348) );
  AOI22X1 U1411 ( .A(n6838), .B(n7005), .C(n6833), .D(n6906), .Y(n1350) );
  NAND3X1 U1413 ( .A(n5124), .B(n5393), .C(n5658), .Y(n1347) );
  AOI22X1 U1414 ( .A(n6829), .B(n7071), .C(n1102), .D(n6939), .Y(n1353) );
  AOI22X1 U1416 ( .A(n6817), .B(n7104), .C(n6813), .D(n7038), .Y(n1351) );
  NAND3X1 U1418 ( .A(n1116), .B(n5392), .C(n5657), .Y(n1355) );
  AOI22X1 U1419 ( .A(n6838), .B(n7797), .C(n6836), .D(n7698), .Y(n1357) );
  NAND3X1 U1421 ( .A(n5123), .B(n5391), .C(n5656), .Y(n1354) );
  AOI22X1 U1422 ( .A(n6829), .B(n7863), .C(n1102), .D(n7731), .Y(n1360) );
  AOI22X1 U1424 ( .A(n6817), .B(n7896), .C(n6812), .D(n7830), .Y(n1358) );
  NAND3X1 U1425 ( .A(n1124), .B(n5390), .C(n5655), .Y(n1362) );
  AOI22X1 U1426 ( .A(n6838), .B(n7533), .C(n1097), .D(n7434), .Y(n1364) );
  NAND3X1 U1428 ( .A(n5122), .B(n5389), .C(n5654), .Y(n1361) );
  AOI22X1 U1429 ( .A(n1101), .B(n7599), .C(n1102), .D(n7467), .Y(n1367) );
  AOI22X1 U1431 ( .A(n6818), .B(n7632), .C(n6812), .D(n7566), .Y(n1365) );
  NAND3X1 U1433 ( .A(n5179), .B(n1369), .C(n1370), .Y(n4468) );
  NOR3X1 U1434 ( .A(n5742), .B(n5775), .C(n5808), .Y(n1370) );
  NAND3X1 U1436 ( .A(n3260), .B(n5388), .C(n5653), .Y(n1375) );
  AOI22X1 U1437 ( .A(n6838), .B(n7270), .C(n1097), .D(n7171), .Y(n1377) );
  NAND3X1 U1439 ( .A(n5121), .B(n5387), .C(n5652), .Y(n1374) );
  AOI22X1 U1440 ( .A(n6828), .B(n7336), .C(n1102), .D(n7204), .Y(n1380) );
  AOI22X1 U1442 ( .A(n1104), .B(n7369), .C(n6814), .D(n7303), .Y(n1378) );
  NAND3X1 U1444 ( .A(n1108), .B(n5386), .C(n5651), .Y(n1382) );
  AOI22X1 U1445 ( .A(n6838), .B(n7006), .C(n6834), .D(n6907), .Y(n1384) );
  NAND3X1 U1447 ( .A(n5120), .B(n5385), .C(n5650), .Y(n1381) );
  AOI22X1 U1448 ( .A(n6829), .B(n7072), .C(n1102), .D(n6940), .Y(n1387) );
  AOI22X1 U1450 ( .A(n1104), .B(n7105), .C(n6812), .D(n7039), .Y(n1385) );
  NAND3X1 U1452 ( .A(n1116), .B(n5384), .C(n5649), .Y(n1389) );
  AOI22X1 U1453 ( .A(n6838), .B(n7798), .C(n1097), .D(n7699), .Y(n1391) );
  NAND3X1 U1455 ( .A(n5119), .B(n5383), .C(n5648), .Y(n1388) );
  AOI22X1 U1456 ( .A(n6829), .B(n7864), .C(n1102), .D(n7732), .Y(n1394) );
  AOI22X1 U1458 ( .A(n6818), .B(n7897), .C(n6813), .D(n7831), .Y(n1392) );
  NAND3X1 U1459 ( .A(n1124), .B(n5382), .C(n5647), .Y(n1396) );
  AOI22X1 U1460 ( .A(n6838), .B(n7534), .C(n1097), .D(n7435), .Y(n1398) );
  NAND3X1 U1462 ( .A(n5118), .B(n5381), .C(n5646), .Y(n1395) );
  AOI22X1 U1463 ( .A(n1101), .B(n7600), .C(n1102), .D(n7468), .Y(n1401) );
  AOI22X1 U1465 ( .A(n6816), .B(n7633), .C(n6813), .D(n7567), .Y(n1399) );
  NAND3X1 U1467 ( .A(n5178), .B(n1403), .C(n1404), .Y(n4469) );
  NOR3X1 U1468 ( .A(n5741), .B(n5774), .C(n5807), .Y(n1404) );
  NAND3X1 U1470 ( .A(n3260), .B(n5380), .C(n5645), .Y(n1409) );
  AOI22X1 U1471 ( .A(n6838), .B(n7271), .C(n1097), .D(n7172), .Y(n1411) );
  NAND3X1 U1473 ( .A(n5117), .B(n5379), .C(n5644), .Y(n1408) );
  AOI22X1 U1474 ( .A(n6829), .B(n7337), .C(n6826), .D(n7205), .Y(n1414) );
  AOI22X1 U1476 ( .A(n1104), .B(n7370), .C(n1105), .D(n7304), .Y(n1412) );
  NAND3X1 U1478 ( .A(n1108), .B(n5378), .C(n5643), .Y(n1416) );
  AOI22X1 U1479 ( .A(n6838), .B(n7007), .C(n6835), .D(n6908), .Y(n1418) );
  NAND3X1 U1481 ( .A(n5116), .B(n5377), .C(n5642), .Y(n1415) );
  AOI22X1 U1482 ( .A(n6830), .B(n7073), .C(n6824), .D(n6941), .Y(n1421) );
  AOI22X1 U1484 ( .A(n6818), .B(n7106), .C(n1105), .D(n7040), .Y(n1419) );
  NAND3X1 U1486 ( .A(n1116), .B(n5376), .C(n5641), .Y(n1423) );
  AOI22X1 U1487 ( .A(n6838), .B(n7799), .C(n6835), .D(n7700), .Y(n1425) );
  NAND3X1 U1489 ( .A(n5115), .B(n5375), .C(n5640), .Y(n1422) );
  AOI22X1 U1490 ( .A(n6828), .B(n7865), .C(n6825), .D(n7733), .Y(n1428) );
  AOI22X1 U1492 ( .A(n6816), .B(n7898), .C(n1105), .D(n7832), .Y(n1426) );
  NAND3X1 U1493 ( .A(n1124), .B(n5374), .C(n5639), .Y(n1430) );
  AOI22X1 U1494 ( .A(n6839), .B(n7535), .C(n1097), .D(n7436), .Y(n1432) );
  NAND3X1 U1496 ( .A(n5114), .B(n5373), .C(n5638), .Y(n1429) );
  AOI22X1 U1497 ( .A(n6828), .B(n7601), .C(n6824), .D(n7469), .Y(n1435) );
  AOI22X1 U1499 ( .A(n1104), .B(n7634), .C(n1105), .D(n7568), .Y(n1433) );
  NAND3X1 U1501 ( .A(n5177), .B(n1437), .C(n1438), .Y(n4470) );
  NOR3X1 U1502 ( .A(n5740), .B(n5773), .C(n5806), .Y(n1438) );
  NAND3X1 U1504 ( .A(n3260), .B(n5372), .C(n5637), .Y(n1443) );
  AOI22X1 U1505 ( .A(n6839), .B(n7272), .C(n1097), .D(n7173), .Y(n1445) );
  NAND3X1 U1507 ( .A(n5113), .B(n5371), .C(n5636), .Y(n1442) );
  AOI22X1 U1508 ( .A(n6828), .B(n7338), .C(n6825), .D(n7206), .Y(n1448) );
  AOI22X1 U1510 ( .A(n1104), .B(n7371), .C(n1105), .D(n7305), .Y(n1446) );
  NAND3X1 U1512 ( .A(n1108), .B(n5370), .C(n5635), .Y(n1450) );
  AOI22X1 U1513 ( .A(n6839), .B(n7008), .C(n1097), .D(n6909), .Y(n1452) );
  NAND3X1 U1515 ( .A(n5112), .B(n5369), .C(n5634), .Y(n1449) );
  AOI22X1 U1516 ( .A(n6828), .B(n7074), .C(n6826), .D(n6942), .Y(n1455) );
  AOI22X1 U1518 ( .A(n1104), .B(n7107), .C(n1105), .D(n7041), .Y(n1453) );
  NAND3X1 U1520 ( .A(n1116), .B(n5368), .C(n5633), .Y(n1457) );
  AOI22X1 U1521 ( .A(n6839), .B(n7800), .C(n6833), .D(n7701), .Y(n1459) );
  NAND3X1 U1523 ( .A(n5111), .B(n5367), .C(n5632), .Y(n1456) );
  AOI22X1 U1524 ( .A(n6828), .B(n7866), .C(n6825), .D(n7734), .Y(n1462) );
  AOI22X1 U1526 ( .A(n6817), .B(n7899), .C(n1105), .D(n7833), .Y(n1460) );
  NAND3X1 U1527 ( .A(n1124), .B(n5366), .C(n5631), .Y(n1464) );
  AOI22X1 U1528 ( .A(n6839), .B(n7536), .C(n1097), .D(n7437), .Y(n1466) );
  NAND3X1 U1530 ( .A(n5110), .B(n5365), .C(n5630), .Y(n1463) );
  AOI22X1 U1531 ( .A(n6828), .B(n7602), .C(n6826), .D(n7470), .Y(n1469) );
  AOI22X1 U1533 ( .A(n1104), .B(n7635), .C(n1105), .D(n7569), .Y(n1467) );
  NAND3X1 U1535 ( .A(n5176), .B(n1471), .C(n1472), .Y(n4471) );
  NOR3X1 U1536 ( .A(n5739), .B(n5772), .C(n5805), .Y(n1472) );
  NAND3X1 U1538 ( .A(n3260), .B(n5364), .C(n5629), .Y(n1477) );
  AOI22X1 U1539 ( .A(n6839), .B(n7273), .C(n1097), .D(n7174), .Y(n1479) );
  NAND3X1 U1541 ( .A(n5109), .B(n5363), .C(n5628), .Y(n1476) );
  AOI22X1 U1542 ( .A(n6828), .B(n7339), .C(n6825), .D(n7207), .Y(n1482) );
  AOI22X1 U1544 ( .A(n1104), .B(n7372), .C(n1105), .D(n7306), .Y(n1480) );
  NAND3X1 U1546 ( .A(n1108), .B(n5362), .C(n5627), .Y(n1484) );
  AOI22X1 U1547 ( .A(n6839), .B(n7009), .C(n1097), .D(n6910), .Y(n1486) );
  NAND3X1 U1549 ( .A(n5108), .B(n5361), .C(n5626), .Y(n1483) );
  AOI22X1 U1550 ( .A(n6828), .B(n7075), .C(n6824), .D(n6943), .Y(n1489) );
  AOI22X1 U1552 ( .A(n6816), .B(n7108), .C(n1105), .D(n7042), .Y(n1487) );
  NAND3X1 U1554 ( .A(n1116), .B(n5360), .C(n5625), .Y(n1491) );
  AOI22X1 U1555 ( .A(n6839), .B(n7801), .C(n6834), .D(n7702), .Y(n1493) );
  NAND3X1 U1557 ( .A(n5107), .B(n5359), .C(n5624), .Y(n1490) );
  AOI22X1 U1558 ( .A(n6828), .B(n7867), .C(n6826), .D(n7735), .Y(n1496) );
  AOI22X1 U1560 ( .A(n6818), .B(n7900), .C(n1105), .D(n7834), .Y(n1494) );
  NAND3X1 U1561 ( .A(n1124), .B(n5358), .C(n5623), .Y(n1498) );
  AOI22X1 U1562 ( .A(n6839), .B(n7537), .C(n1097), .D(n7438), .Y(n1500) );
  NAND3X1 U1564 ( .A(n5106), .B(n5357), .C(n5622), .Y(n1497) );
  AOI22X1 U1565 ( .A(n6828), .B(n7603), .C(n6824), .D(n7471), .Y(n1503) );
  AOI22X1 U1567 ( .A(n1104), .B(n7636), .C(n1105), .D(n7570), .Y(n1501) );
  NAND3X1 U1569 ( .A(n5175), .B(n1505), .C(n1506), .Y(n4472) );
  NOR3X1 U1570 ( .A(n5738), .B(n5771), .C(n5804), .Y(n1506) );
  NAND3X1 U1572 ( .A(n3260), .B(n5356), .C(n5621), .Y(n1511) );
  AOI22X1 U1573 ( .A(n6839), .B(n7274), .C(n1097), .D(n7175), .Y(n1513) );
  NAND3X1 U1575 ( .A(n5105), .B(n5355), .C(n5620), .Y(n1510) );
  AOI22X1 U1576 ( .A(n6828), .B(n7340), .C(n1102), .D(n7208), .Y(n1516) );
  AOI22X1 U1578 ( .A(n1104), .B(n7373), .C(n1105), .D(n7307), .Y(n1514) );
  NAND3X1 U1580 ( .A(n1108), .B(n5354), .C(n5619), .Y(n1518) );
  AOI22X1 U1581 ( .A(n6839), .B(n7010), .C(n6835), .D(n6911), .Y(n1520) );
  NAND3X1 U1583 ( .A(n5104), .B(n5353), .C(n5618), .Y(n1517) );
  AOI22X1 U1584 ( .A(n6828), .B(n7076), .C(n1102), .D(n6944), .Y(n1523) );
  AOI22X1 U1586 ( .A(n6816), .B(n7109), .C(n1105), .D(n7043), .Y(n1521) );
  NAND3X1 U1588 ( .A(n1116), .B(n5352), .C(n5617), .Y(n1525) );
  AOI22X1 U1589 ( .A(n6839), .B(n7802), .C(n6833), .D(n7703), .Y(n1527) );
  NAND3X1 U1591 ( .A(n5103), .B(n5351), .C(n5616), .Y(n1524) );
  AOI22X1 U1592 ( .A(n6828), .B(n7868), .C(n1102), .D(n7736), .Y(n1530) );
  AOI22X1 U1594 ( .A(n6816), .B(n7901), .C(n1105), .D(n7835), .Y(n1528) );
  NAND3X1 U1595 ( .A(n1124), .B(n5350), .C(n5615), .Y(n1532) );
  AOI22X1 U1596 ( .A(n6839), .B(n7538), .C(n1097), .D(n7439), .Y(n1534) );
  NAND3X1 U1598 ( .A(n5102), .B(n5349), .C(n5614), .Y(n1531) );
  AOI22X1 U1599 ( .A(n6828), .B(n7604), .C(n1102), .D(n7472), .Y(n1537) );
  AOI22X1 U1601 ( .A(n1104), .B(n7637), .C(n6812), .D(n7571), .Y(n1535) );
  NAND3X1 U1603 ( .A(n5174), .B(n2605), .C(n2606), .Y(n4473) );
  NOR3X1 U1604 ( .A(n5737), .B(n5770), .C(n5803), .Y(n2606) );
  NAND3X1 U1606 ( .A(n3260), .B(n5348), .C(n5613), .Y(n2611) );
  AOI22X1 U1607 ( .A(n1096), .B(n7275), .C(n6834), .D(n7176), .Y(n2613) );
  NAND3X1 U1609 ( .A(n5101), .B(n5347), .C(n5612), .Y(n2610) );
  AOI22X1 U1610 ( .A(n6829), .B(n7341), .C(n1102), .D(n7209), .Y(n2616) );
  AOI22X1 U1612 ( .A(n6816), .B(n7374), .C(n1105), .D(n7308), .Y(n2614) );
  NAND3X1 U1614 ( .A(n1108), .B(n5346), .C(n5611), .Y(n2618) );
  AOI22X1 U1615 ( .A(n6839), .B(n7011), .C(n6834), .D(n6912), .Y(n2620) );
  NAND3X1 U1617 ( .A(n5100), .B(n5345), .C(n5610), .Y(n2617) );
  AOI22X1 U1618 ( .A(n6829), .B(n7077), .C(n1102), .D(n6945), .Y(n2623) );
  AOI22X1 U1620 ( .A(n6816), .B(n7110), .C(n1105), .D(n7044), .Y(n2621) );
  NAND3X1 U1622 ( .A(n1116), .B(n5344), .C(n5609), .Y(n2625) );
  AOI22X1 U1623 ( .A(n6840), .B(n7803), .C(n1097), .D(n7704), .Y(n2627) );
  NAND3X1 U1625 ( .A(n5099), .B(n5343), .C(n5608), .Y(n2624) );
  AOI22X1 U1626 ( .A(n6829), .B(n7869), .C(n1102), .D(n7737), .Y(n2630) );
  AOI22X1 U1628 ( .A(n6816), .B(n7902), .C(n1105), .D(n7836), .Y(n2628) );
  NAND3X1 U1629 ( .A(n1124), .B(n5342), .C(n5607), .Y(n2632) );
  AOI22X1 U1630 ( .A(n1096), .B(n7539), .C(n1097), .D(n7440), .Y(n2634) );
  NAND3X1 U1632 ( .A(n5098), .B(n5341), .C(n5606), .Y(n2631) );
  AOI22X1 U1633 ( .A(n6829), .B(n7605), .C(n1102), .D(n7473), .Y(n2637) );
  AOI22X1 U1635 ( .A(n6816), .B(n7638), .C(n1105), .D(n7572), .Y(n2635) );
  NAND3X1 U1637 ( .A(n5173), .B(n2639), .C(n2640), .Y(n4474) );
  NOR3X1 U1638 ( .A(n5736), .B(n5769), .C(n5802), .Y(n2640) );
  NAND3X1 U1640 ( .A(n3260), .B(n5340), .C(n5605), .Y(n2645) );
  AOI22X1 U1641 ( .A(n1096), .B(n7276), .C(n6833), .D(n7177), .Y(n2647) );
  NAND3X1 U1643 ( .A(n5097), .B(n5339), .C(n5604), .Y(n2644) );
  AOI22X1 U1644 ( .A(n6829), .B(n7342), .C(n1102), .D(n7210), .Y(n2650) );
  AOI22X1 U1646 ( .A(n6816), .B(n7375), .C(n1105), .D(n7309), .Y(n2648) );
  NAND3X1 U1648 ( .A(n1108), .B(n5338), .C(n5603), .Y(n2652) );
  AOI22X1 U1649 ( .A(n6838), .B(n7012), .C(n6836), .D(n6913), .Y(n2654) );
  NAND3X1 U1651 ( .A(n5096), .B(n5337), .C(n5602), .Y(n2651) );
  AOI22X1 U1652 ( .A(n6829), .B(n7078), .C(n1102), .D(n6946), .Y(n2657) );
  AOI22X1 U1654 ( .A(n6816), .B(n7111), .C(n1105), .D(n7045), .Y(n2655) );
  NAND3X1 U1656 ( .A(n1116), .B(n5336), .C(n5601), .Y(n2659) );
  AOI22X1 U1657 ( .A(n6837), .B(n7804), .C(n6835), .D(n7705), .Y(n2661) );
  NAND3X1 U1659 ( .A(n5095), .B(n5335), .C(n5600), .Y(n2658) );
  AOI22X1 U1660 ( .A(n6829), .B(n7870), .C(n1102), .D(n7738), .Y(n2664) );
  AOI22X1 U1662 ( .A(n6816), .B(n7903), .C(n1105), .D(n7837), .Y(n2662) );
  NAND3X1 U1663 ( .A(n1124), .B(n5334), .C(n5599), .Y(n2666) );
  AOI22X1 U1664 ( .A(n1096), .B(n7540), .C(n1097), .D(n7441), .Y(n2668) );
  NAND3X1 U1666 ( .A(n5094), .B(n5333), .C(n5598), .Y(n2665) );
  AOI22X1 U1667 ( .A(n6829), .B(n7606), .C(n1102), .D(n7474), .Y(n2671) );
  AOI22X1 U1669 ( .A(n6816), .B(n7639), .C(n1105), .D(n7573), .Y(n2669) );
  NAND3X1 U1671 ( .A(n5172), .B(n2673), .C(n2674), .Y(n4475) );
  NOR3X1 U1672 ( .A(n5735), .B(n5768), .C(n5801), .Y(n2674) );
  NAND3X1 U1674 ( .A(n3260), .B(n5332), .C(n5597), .Y(n2679) );
  AOI22X1 U1675 ( .A(n6840), .B(n7277), .C(n6836), .D(n7178), .Y(n2681) );
  NAND3X1 U1677 ( .A(n5093), .B(n5331), .C(n5596), .Y(n2678) );
  AOI22X1 U1678 ( .A(n6829), .B(n7343), .C(n6824), .D(n7211), .Y(n2684) );
  AOI22X1 U1680 ( .A(n6816), .B(n7376), .C(n6813), .D(n7310), .Y(n2682) );
  NAND3X1 U1682 ( .A(n1108), .B(n5330), .C(n5595), .Y(n2686) );
  AOI22X1 U1683 ( .A(n6838), .B(n7013), .C(n6836), .D(n6914), .Y(n2688) );
  NAND3X1 U1685 ( .A(n5092), .B(n5329), .C(n5594), .Y(n2685) );
  AOI22X1 U1686 ( .A(n6829), .B(n7079), .C(n6825), .D(n6947), .Y(n2691) );
  AOI22X1 U1688 ( .A(n6816), .B(n7112), .C(n6812), .D(n7046), .Y(n2689) );
  NAND3X1 U1690 ( .A(n1116), .B(n5328), .C(n5593), .Y(n2693) );
  AOI22X1 U1691 ( .A(n6839), .B(n7805), .C(n6835), .D(n7706), .Y(n2695) );
  NAND3X1 U1693 ( .A(n5091), .B(n5327), .C(n5592), .Y(n2692) );
  AOI22X1 U1694 ( .A(n6829), .B(n7871), .C(n6824), .D(n7739), .Y(n2698) );
  AOI22X1 U1696 ( .A(n6816), .B(n7904), .C(n6813), .D(n7838), .Y(n2696) );
  NAND3X1 U1697 ( .A(n1124), .B(n5326), .C(n5591), .Y(n2700) );
  AOI22X1 U1698 ( .A(n1096), .B(n7541), .C(n6833), .D(n7442), .Y(n2702) );
  NAND3X1 U1700 ( .A(n5090), .B(n5325), .C(n5590), .Y(n2699) );
  AOI22X1 U1701 ( .A(n6829), .B(n7607), .C(n6826), .D(n7475), .Y(n2705) );
  AOI22X1 U1703 ( .A(n6816), .B(n7640), .C(n6813), .D(n7574), .Y(n2703) );
  NAND3X1 U1705 ( .A(n5171), .B(n2707), .C(n2708), .Y(n4476) );
  NOR3X1 U1706 ( .A(n5734), .B(n5767), .C(n5800), .Y(n2708) );
  NAND3X1 U1708 ( .A(n3260), .B(n5324), .C(n5589), .Y(n2713) );
  AOI22X1 U1709 ( .A(n6837), .B(n7257), .C(n6835), .D(n7158), .Y(n2715) );
  NAND3X1 U1711 ( .A(n5089), .B(n5323), .C(n5588), .Y(n2712) );
  AOI22X1 U1712 ( .A(n6829), .B(n7323), .C(n6824), .D(n7191), .Y(n2718) );
  AOI22X1 U1714 ( .A(n6816), .B(n7356), .C(n6814), .D(n7290), .Y(n2716) );
  NAND3X1 U1716 ( .A(n1108), .B(n5322), .C(n5587), .Y(n2720) );
  AOI22X1 U1717 ( .A(n6838), .B(n6993), .C(n6834), .D(n6894), .Y(n2722) );
  NAND3X1 U1719 ( .A(n5088), .B(n5321), .C(n5586), .Y(n2719) );
  AOI22X1 U1720 ( .A(n6830), .B(n7059), .C(n6824), .D(n6927), .Y(n2725) );
  AOI22X1 U1722 ( .A(n6817), .B(n7092), .C(n6812), .D(n7026), .Y(n2723) );
  NAND3X1 U1724 ( .A(n1116), .B(n5320), .C(n5585), .Y(n2727) );
  AOI22X1 U1725 ( .A(n6837), .B(n7785), .C(n6834), .D(n7686), .Y(n2729) );
  NAND3X1 U1727 ( .A(n5087), .B(n5319), .C(n5584), .Y(n2726) );
  AOI22X1 U1728 ( .A(n6830), .B(n7851), .C(n6825), .D(n7719), .Y(n2732) );
  AOI22X1 U1730 ( .A(n6817), .B(n7884), .C(n6814), .D(n7818), .Y(n2730) );
  NAND3X1 U1731 ( .A(n1124), .B(n5318), .C(n5583), .Y(n2734) );
  AOI22X1 U1732 ( .A(n6837), .B(n7521), .C(n6835), .D(n7422), .Y(n2736) );
  NAND3X1 U1734 ( .A(n5086), .B(n5317), .C(n5582), .Y(n2733) );
  AOI22X1 U1735 ( .A(n6830), .B(n7587), .C(n6824), .D(n7455), .Y(n2739) );
  AOI22X1 U1737 ( .A(n6817), .B(n7620), .C(n6812), .D(n7554), .Y(n2737) );
  NAND3X1 U1739 ( .A(n5170), .B(n2741), .C(n2742), .Y(n4477) );
  NOR3X1 U1740 ( .A(n5733), .B(n5766), .C(n5799), .Y(n2742) );
  NAND3X1 U1742 ( .A(n3260), .B(n5316), .C(n5581), .Y(n2747) );
  AOI22X1 U1743 ( .A(n6838), .B(n7259), .C(n6834), .D(n7160), .Y(n2749) );
  NAND3X1 U1745 ( .A(n5085), .B(n5315), .C(n5580), .Y(n2746) );
  AOI22X1 U1746 ( .A(n6830), .B(n7325), .C(n6826), .D(n7193), .Y(n2752) );
  AOI22X1 U1748 ( .A(n6817), .B(n7358), .C(n6813), .D(n7292), .Y(n2750) );
  NAND3X1 U1750 ( .A(n1108), .B(n5314), .C(n5579), .Y(n2754) );
  AOI22X1 U1751 ( .A(n6837), .B(n6995), .C(n6834), .D(n6896), .Y(n2756) );
  NAND3X1 U1753 ( .A(n5084), .B(n5313), .C(n5578), .Y(n2753) );
  AOI22X1 U1754 ( .A(n6830), .B(n7061), .C(n6826), .D(n6929), .Y(n2759) );
  AOI22X1 U1756 ( .A(n6817), .B(n7094), .C(n6814), .D(n7028), .Y(n2757) );
  NAND3X1 U1758 ( .A(n1116), .B(n5312), .C(n5577), .Y(n2761) );
  AOI22X1 U1759 ( .A(n1096), .B(n7787), .C(n6836), .D(n7688), .Y(n2763) );
  NAND3X1 U1761 ( .A(n5083), .B(n5311), .C(n5576), .Y(n2760) );
  AOI22X1 U1762 ( .A(n6830), .B(n7853), .C(n6825), .D(n7721), .Y(n2766) );
  AOI22X1 U1764 ( .A(n6817), .B(n7886), .C(n6814), .D(n7820), .Y(n2764) );
  NAND3X1 U1765 ( .A(n1124), .B(n5310), .C(n5575), .Y(n2768) );
  AOI22X1 U1766 ( .A(n6840), .B(n7523), .C(n6836), .D(n7424), .Y(n2770) );
  NAND3X1 U1768 ( .A(n5082), .B(n5309), .C(n5574), .Y(n2767) );
  AOI22X1 U1769 ( .A(n6830), .B(n7589), .C(n6825), .D(n7457), .Y(n2773) );
  AOI22X1 U1771 ( .A(n6817), .B(n7622), .C(n6814), .D(n7556), .Y(n2771) );
  NAND3X1 U1773 ( .A(n5169), .B(n2775), .C(n2776), .Y(n4478) );
  NOR3X1 U1774 ( .A(n5732), .B(n5765), .C(n5798), .Y(n2776) );
  NAND3X1 U1776 ( .A(n3260), .B(n5308), .C(n5573), .Y(n2781) );
  AOI22X1 U1777 ( .A(n6837), .B(n7261), .C(n1097), .D(n7162), .Y(n2783) );
  NAND3X1 U1779 ( .A(n5081), .B(n5307), .C(n5572), .Y(n2780) );
  AOI22X1 U1780 ( .A(n6830), .B(n7327), .C(n6825), .D(n7195), .Y(n2786) );
  AOI22X1 U1782 ( .A(n6817), .B(n7360), .C(n6813), .D(n7294), .Y(n2784) );
  NAND3X1 U1784 ( .A(n1108), .B(n5306), .C(n5571), .Y(n2788) );
  AOI22X1 U1785 ( .A(n6840), .B(n6997), .C(n6834), .D(n6898), .Y(n2790) );
  NAND3X1 U1787 ( .A(n5080), .B(n5305), .C(n5570), .Y(n2787) );
  AOI22X1 U1788 ( .A(n6830), .B(n7063), .C(n6826), .D(n6931), .Y(n2793) );
  AOI22X1 U1790 ( .A(n6817), .B(n7096), .C(n6814), .D(n7030), .Y(n2791) );
  NAND3X1 U1792 ( .A(n1116), .B(n5304), .C(n5569), .Y(n2795) );
  AOI22X1 U1793 ( .A(n1096), .B(n7789), .C(n6836), .D(n7690), .Y(n2797) );
  NAND3X1 U1795 ( .A(n5079), .B(n5303), .C(n5568), .Y(n2794) );
  AOI22X1 U1796 ( .A(n6830), .B(n7855), .C(n6825), .D(n7723), .Y(n2800) );
  AOI22X1 U1798 ( .A(n6817), .B(n7888), .C(n6813), .D(n7822), .Y(n2798) );
  NAND3X1 U1799 ( .A(n1124), .B(n5302), .C(n5567), .Y(n2802) );
  AOI22X1 U1800 ( .A(n6839), .B(n7525), .C(n1097), .D(n7426), .Y(n2804) );
  NAND3X1 U1802 ( .A(n5078), .B(n5301), .C(n5566), .Y(n2801) );
  AOI22X1 U1803 ( .A(n6830), .B(n7591), .C(n6825), .D(n7459), .Y(n2807) );
  AOI22X1 U1805 ( .A(n6817), .B(n7624), .C(n6812), .D(n7558), .Y(n2805) );
  NAND3X1 U1807 ( .A(n5168), .B(n2809), .C(n2810), .Y(n4479) );
  NOR3X1 U1808 ( .A(n5731), .B(n5764), .C(n5797), .Y(n2810) );
  NAND3X1 U1810 ( .A(n3260), .B(n5300), .C(n5565), .Y(n2815) );
  AOI22X1 U1811 ( .A(n6840), .B(n7263), .C(n1097), .D(n7164), .Y(n2817) );
  NAND3X1 U1813 ( .A(n5077), .B(n5299), .C(n5564), .Y(n2814) );
  AOI22X1 U1814 ( .A(n6830), .B(n7329), .C(n6824), .D(n7197), .Y(n2820) );
  AOI22X1 U1816 ( .A(n6817), .B(n7362), .C(n6814), .D(n7296), .Y(n2818) );
  NAND3X1 U1818 ( .A(n1108), .B(n5298), .C(n5563), .Y(n2822) );
  AOI22X1 U1819 ( .A(n6839), .B(n6999), .C(n6833), .D(n6900), .Y(n2824) );
  NAND3X1 U1821 ( .A(n5076), .B(n5297), .C(n5562), .Y(n2821) );
  AOI22X1 U1822 ( .A(n6830), .B(n7065), .C(n6825), .D(n6933), .Y(n2827) );
  AOI22X1 U1824 ( .A(n6817), .B(n7098), .C(n6812), .D(n7032), .Y(n2825) );
  NAND3X1 U1826 ( .A(n1116), .B(n5296), .C(n5561), .Y(n2829) );
  AOI22X1 U1827 ( .A(n1096), .B(n7791), .C(n6835), .D(n7692), .Y(n2831) );
  NAND3X1 U1829 ( .A(n5075), .B(n5295), .C(n5560), .Y(n2828) );
  AOI22X1 U1830 ( .A(n1101), .B(n7857), .C(n6824), .D(n7725), .Y(n2834) );
  AOI22X1 U1832 ( .A(n1104), .B(n7890), .C(n6814), .D(n7824), .Y(n2832) );
  NAND3X1 U1833 ( .A(n1124), .B(n5294), .C(n5559), .Y(n2836) );
  AOI22X1 U1834 ( .A(n1096), .B(n7527), .C(n1097), .D(n7428), .Y(n2838) );
  NAND3X1 U1836 ( .A(n5074), .B(n5293), .C(n5558), .Y(n2835) );
  AOI22X1 U1837 ( .A(n1101), .B(n7593), .C(n6825), .D(n7461), .Y(n2841) );
  AOI22X1 U1839 ( .A(n1104), .B(n7626), .C(n6812), .D(n7560), .Y(n2839) );
  NAND3X1 U1841 ( .A(n5167), .B(n2843), .C(n2844), .Y(n4480) );
  NOR3X1 U1842 ( .A(n5730), .B(n5763), .C(n5796), .Y(n2844) );
  NAND3X1 U1844 ( .A(n3260), .B(n5292), .C(n5557), .Y(n2849) );
  AOI22X1 U1845 ( .A(n1096), .B(n7265), .C(n6833), .D(n7166), .Y(n2851) );
  NAND3X1 U1847 ( .A(n5073), .B(n5291), .C(n5556), .Y(n2848) );
  AOI22X1 U1848 ( .A(n1101), .B(n7331), .C(n6824), .D(n7199), .Y(n2854) );
  AOI22X1 U1850 ( .A(n1104), .B(n7364), .C(n6813), .D(n7298), .Y(n2852) );
  NAND3X1 U1852 ( .A(n1108), .B(n5290), .C(n5555), .Y(n2856) );
  AOI22X1 U1853 ( .A(n1096), .B(n7001), .C(n6834), .D(n6902), .Y(n2858) );
  NAND3X1 U1855 ( .A(n5072), .B(n5289), .C(n5554), .Y(n2855) );
  AOI22X1 U1856 ( .A(n1101), .B(n7067), .C(n6826), .D(n6935), .Y(n2861) );
  AOI22X1 U1858 ( .A(n1104), .B(n7100), .C(n6812), .D(n7034), .Y(n2859) );
  NAND3X1 U1860 ( .A(n1116), .B(n5288), .C(n5553), .Y(n2863) );
  AOI22X1 U1861 ( .A(n1096), .B(n7793), .C(n6836), .D(n7694), .Y(n2865) );
  NAND3X1 U1863 ( .A(n5071), .B(n5287), .C(n5552), .Y(n2862) );
  AOI22X1 U1864 ( .A(n1101), .B(n7859), .C(n6826), .D(n7727), .Y(n2868) );
  AOI22X1 U1866 ( .A(n1104), .B(n7892), .C(n6814), .D(n7826), .Y(n2866) );
  NAND3X1 U1867 ( .A(n1124), .B(n5286), .C(n5551), .Y(n2870) );
  AOI22X1 U1868 ( .A(n1096), .B(n7529), .C(n1097), .D(n7430), .Y(n2872) );
  NAND3X1 U1870 ( .A(n5070), .B(n5285), .C(n5550), .Y(n2869) );
  AOI22X1 U1871 ( .A(n1101), .B(n7595), .C(n6824), .D(n7463), .Y(n2875) );
  AOI22X1 U1873 ( .A(n1104), .B(n7628), .C(n6812), .D(n7562), .Y(n2873) );
  NAND3X1 U1875 ( .A(n5166), .B(n2877), .C(n2878), .Y(n4481) );
  NOR3X1 U1876 ( .A(n5729), .B(n5762), .C(n5795), .Y(n2878) );
  NAND3X1 U1878 ( .A(n3260), .B(n5284), .C(n5549), .Y(n2883) );
  AOI22X1 U1879 ( .A(n1096), .B(n7278), .C(n6836), .D(n7179), .Y(n2885) );
  NAND3X1 U1881 ( .A(n5069), .B(n5283), .C(n5548), .Y(n2882) );
  AOI22X1 U1882 ( .A(n1101), .B(n7344), .C(n6826), .D(n7212), .Y(n2888) );
  AOI22X1 U1884 ( .A(n1104), .B(n7377), .C(n6813), .D(n7311), .Y(n2886) );
  NAND3X1 U1886 ( .A(n1108), .B(n5282), .C(n5547), .Y(n2890) );
  AOI22X1 U1887 ( .A(n1096), .B(n7014), .C(n6836), .D(n6915), .Y(n2892) );
  NAND3X1 U1889 ( .A(n5068), .B(n5281), .C(n5546), .Y(n2889) );
  AOI22X1 U1890 ( .A(n1101), .B(n7080), .C(n6825), .D(n6948), .Y(n2895) );
  AOI22X1 U1892 ( .A(n1104), .B(n7113), .C(n6813), .D(n7047), .Y(n2893) );
  NAND3X1 U1894 ( .A(n1116), .B(n5280), .C(n5545), .Y(n2897) );
  AOI22X1 U1895 ( .A(n1096), .B(n7806), .C(n6836), .D(n7707), .Y(n2899) );
  NAND3X1 U1897 ( .A(n5067), .B(n5279), .C(n5544), .Y(n2896) );
  AOI22X1 U1898 ( .A(n1101), .B(n7872), .C(n6824), .D(n7740), .Y(n2902) );
  AOI22X1 U1900 ( .A(n1104), .B(n7905), .C(n6814), .D(n7839), .Y(n2900) );
  NAND3X1 U1901 ( .A(n1124), .B(n5278), .C(n5543), .Y(n2904) );
  AOI22X1 U1902 ( .A(n1096), .B(n7542), .C(n6836), .D(n7443), .Y(n2906) );
  NAND3X1 U1904 ( .A(n5066), .B(n5277), .C(n5542), .Y(n2903) );
  AOI22X1 U1905 ( .A(n1101), .B(n7608), .C(n6825), .D(n7476), .Y(n2909) );
  AOI22X1 U1907 ( .A(n1104), .B(n7641), .C(n6813), .D(n7575), .Y(n2907) );
  NAND3X1 U1909 ( .A(n5165), .B(n2911), .C(n2912), .Y(n4482) );
  NOR3X1 U1910 ( .A(n5728), .B(n5761), .C(n5794), .Y(n2912) );
  NAND3X1 U1912 ( .A(n3260), .B(n5276), .C(n5541), .Y(n2917) );
  AOI22X1 U1913 ( .A(n1096), .B(n7279), .C(n6836), .D(n7180), .Y(n2919) );
  NAND3X1 U1915 ( .A(n5065), .B(n5275), .C(n5540), .Y(n2916) );
  AOI22X1 U1916 ( .A(n1101), .B(n7345), .C(n6824), .D(n7213), .Y(n2922) );
  AOI22X1 U1918 ( .A(n1104), .B(n7378), .C(n6812), .D(n7312), .Y(n2920) );
  NAND3X1 U1920 ( .A(n1108), .B(n5274), .C(n5539), .Y(n2924) );
  AOI22X1 U1921 ( .A(n1096), .B(n7015), .C(n6836), .D(n6916), .Y(n2926) );
  NAND3X1 U1923 ( .A(n5064), .B(n5273), .C(n5538), .Y(n2923) );
  AOI22X1 U1924 ( .A(n1101), .B(n7081), .C(n6826), .D(n6949), .Y(n2929) );
  AOI22X1 U1926 ( .A(n1104), .B(n7114), .C(n6812), .D(n7048), .Y(n2927) );
  NAND3X1 U1928 ( .A(n1116), .B(n5272), .C(n5537), .Y(n2931) );
  AOI22X1 U1929 ( .A(n1096), .B(n7807), .C(n6836), .D(n7708), .Y(n2933) );
  NAND3X1 U1931 ( .A(n5063), .B(n5271), .C(n5536), .Y(n2930) );
  AOI22X1 U1932 ( .A(n6828), .B(n7873), .C(n6825), .D(n7741), .Y(n2936) );
  AOI22X1 U1934 ( .A(n6817), .B(n7906), .C(n6813), .D(n7840), .Y(n2934) );
  NAND3X1 U1935 ( .A(n1124), .B(n5270), .C(n5535), .Y(n2938) );
  AOI22X1 U1936 ( .A(n1096), .B(n7543), .C(n6836), .D(n7444), .Y(n2940) );
  NAND3X1 U1938 ( .A(n5062), .B(n5269), .C(n5534), .Y(n2937) );
  AOI22X1 U1939 ( .A(n6828), .B(n7609), .C(n6826), .D(n7477), .Y(n2943) );
  AOI22X1 U1941 ( .A(n6817), .B(n7642), .C(n6812), .D(n7576), .Y(n2941) );
  NAND3X1 U1943 ( .A(n5164), .B(n2945), .C(n2946), .Y(n4483) );
  NOR3X1 U1944 ( .A(n5727), .B(n5760), .C(n5793), .Y(n2946) );
  NAND3X1 U1946 ( .A(n3260), .B(n5268), .C(n5533), .Y(n2951) );
  AOI22X1 U1947 ( .A(n1096), .B(n7280), .C(n6836), .D(n7181), .Y(n2953) );
  NAND3X1 U1949 ( .A(n5061), .B(n5267), .C(n5532), .Y(n2950) );
  AOI22X1 U1950 ( .A(n6829), .B(n7346), .C(n6826), .D(n7214), .Y(n2956) );
  AOI22X1 U1952 ( .A(n6817), .B(n7379), .C(n6814), .D(n7313), .Y(n2954) );
  NAND3X1 U1954 ( .A(n1108), .B(n5266), .C(n5531), .Y(n2958) );
  AOI22X1 U1955 ( .A(n1096), .B(n7016), .C(n6836), .D(n6917), .Y(n2960) );
  NAND3X1 U1957 ( .A(n5060), .B(n5265), .C(n5530), .Y(n2957) );
  AOI22X1 U1958 ( .A(n1101), .B(n7082), .C(n6825), .D(n6950), .Y(n2963) );
  AOI22X1 U1960 ( .A(n1104), .B(n7115), .C(n6813), .D(n7049), .Y(n2961) );
  NAND3X1 U1962 ( .A(n1116), .B(n5264), .C(n5529), .Y(n2965) );
  AOI22X1 U1963 ( .A(n1096), .B(n7808), .C(n6836), .D(n7709), .Y(n2967) );
  NAND3X1 U1965 ( .A(n5059), .B(n5263), .C(n5528), .Y(n2964) );
  AOI22X1 U1966 ( .A(n1101), .B(n7874), .C(n6824), .D(n7742), .Y(n2970) );
  AOI22X1 U1968 ( .A(n1104), .B(n7907), .C(n6814), .D(n7841), .Y(n2968) );
  NAND3X1 U1969 ( .A(n1124), .B(n5262), .C(n5527), .Y(n2972) );
  AOI22X1 U1970 ( .A(n1096), .B(n7544), .C(n6836), .D(n7445), .Y(n2974) );
  NAND3X1 U1972 ( .A(n5058), .B(n5261), .C(n5526), .Y(n2971) );
  AOI22X1 U1973 ( .A(n6829), .B(n7610), .C(n6826), .D(n7478), .Y(n2977) );
  AOI22X1 U1975 ( .A(n6818), .B(n7643), .C(n6814), .D(n7577), .Y(n2975) );
  NAND3X1 U1977 ( .A(n5163), .B(n2979), .C(n2980), .Y(n4484) );
  NOR3X1 U1978 ( .A(n5726), .B(n5759), .C(n5792), .Y(n2980) );
  NAND3X1 U1980 ( .A(n3260), .B(n5260), .C(n5525), .Y(n2985) );
  AOI22X1 U1981 ( .A(n1096), .B(n7281), .C(n6835), .D(n7182), .Y(n2987) );
  NAND3X1 U1983 ( .A(n5057), .B(n5259), .C(n5524), .Y(n2984) );
  AOI22X1 U1984 ( .A(n1101), .B(n7347), .C(n6824), .D(n7215), .Y(n2990) );
  AOI22X1 U1986 ( .A(n6818), .B(n7380), .C(n6812), .D(n7314), .Y(n2988) );
  NAND3X1 U1988 ( .A(n1108), .B(n5258), .C(n5523), .Y(n2992) );
  AOI22X1 U1989 ( .A(n6840), .B(n7017), .C(n6835), .D(n6918), .Y(n2994) );
  NAND3X1 U1991 ( .A(n5056), .B(n5257), .C(n5522), .Y(n2991) );
  AOI22X1 U1992 ( .A(n1101), .B(n7083), .C(n6824), .D(n6951), .Y(n2997) );
  AOI22X1 U1994 ( .A(n1104), .B(n7116), .C(n6812), .D(n7050), .Y(n2995) );
  NAND3X1 U1996 ( .A(n1116), .B(n5256), .C(n5521), .Y(n2999) );
  AOI22X1 U1997 ( .A(n6840), .B(n7809), .C(n6835), .D(n7710), .Y(n3001) );
  NAND3X1 U1999 ( .A(n5055), .B(n5255), .C(n5520), .Y(n2998) );
  AOI22X1 U2000 ( .A(n1101), .B(n7875), .C(n6824), .D(n7743), .Y(n3004) );
  AOI22X1 U2002 ( .A(n1104), .B(n7908), .C(n6812), .D(n7842), .Y(n3002) );
  NAND3X1 U2003 ( .A(n1124), .B(n5254), .C(n5519), .Y(n3006) );
  AOI22X1 U2004 ( .A(n1096), .B(n7545), .C(n6835), .D(n7446), .Y(n3008) );
  NAND3X1 U2006 ( .A(n5054), .B(n5253), .C(n5518), .Y(n3005) );
  AOI22X1 U2007 ( .A(n6830), .B(n7611), .C(n6824), .D(n7479), .Y(n3011) );
  AOI22X1 U2009 ( .A(n6816), .B(n7644), .C(n6812), .D(n7578), .Y(n3009) );
  NAND3X1 U2011 ( .A(n5162), .B(n3013), .C(n3014), .Y(n4485) );
  NOR3X1 U2012 ( .A(n5725), .B(n5758), .C(n5791), .Y(n3014) );
  NAND3X1 U2014 ( .A(n3260), .B(n5252), .C(n5517), .Y(n3019) );
  AOI22X1 U2015 ( .A(n1096), .B(n7282), .C(n6835), .D(n7183), .Y(n3021) );
  NAND3X1 U2017 ( .A(n5053), .B(n5251), .C(n5516), .Y(n3018) );
  AOI22X1 U2018 ( .A(n1101), .B(n7348), .C(n6824), .D(n7216), .Y(n3024) );
  AOI22X1 U2020 ( .A(n1104), .B(n7381), .C(n6812), .D(n7315), .Y(n3022) );
  NAND3X1 U2022 ( .A(n1108), .B(n5250), .C(n5515), .Y(n3026) );
  AOI22X1 U2023 ( .A(n6837), .B(n7018), .C(n6835), .D(n6919), .Y(n3028) );
  NAND3X1 U2025 ( .A(n5052), .B(n5249), .C(n5514), .Y(n3025) );
  AOI22X1 U2026 ( .A(n1101), .B(n7084), .C(n6824), .D(n6952), .Y(n3031) );
  AOI22X1 U2028 ( .A(n1104), .B(n7117), .C(n6812), .D(n7051), .Y(n3029) );
  NAND3X1 U2030 ( .A(n1116), .B(n5248), .C(n5513), .Y(n3033) );
  AOI22X1 U2031 ( .A(n6837), .B(n7810), .C(n6835), .D(n7711), .Y(n3035) );
  NAND3X1 U2033 ( .A(n5051), .B(n5247), .C(n5512), .Y(n3032) );
  AOI22X1 U2034 ( .A(n1101), .B(n7876), .C(n6824), .D(n7744), .Y(n3038) );
  AOI22X1 U2036 ( .A(n1104), .B(n7909), .C(n6812), .D(n7843), .Y(n3036) );
  NAND3X1 U2037 ( .A(n1124), .B(n5246), .C(n5511), .Y(n3040) );
  AOI22X1 U2038 ( .A(n1096), .B(n7546), .C(n6835), .D(n7447), .Y(n3042) );
  NAND3X1 U2040 ( .A(n5050), .B(n5245), .C(n5510), .Y(n3039) );
  AOI22X1 U2041 ( .A(n6830), .B(n7612), .C(n6824), .D(n7480), .Y(n3045) );
  AOI22X1 U2043 ( .A(n6816), .B(n7645), .C(n6812), .D(n7579), .Y(n3043) );
  NAND3X1 U2045 ( .A(n5161), .B(n3047), .C(n3048), .Y(n4486) );
  NOR3X1 U2046 ( .A(n5724), .B(n5757), .C(n5790), .Y(n3048) );
  NAND3X1 U2048 ( .A(n3260), .B(n5244), .C(n5509), .Y(n3053) );
  AOI22X1 U2049 ( .A(n1096), .B(n7283), .C(n6835), .D(n7184), .Y(n3055) );
  NAND3X1 U2051 ( .A(n5049), .B(n5243), .C(n5508), .Y(n3052) );
  AOI22X1 U2052 ( .A(n1101), .B(n7349), .C(n6824), .D(n7217), .Y(n3058) );
  AOI22X1 U2054 ( .A(n6818), .B(n7382), .C(n6812), .D(n7316), .Y(n3056) );
  NAND3X1 U2056 ( .A(n1108), .B(n5242), .C(n5507), .Y(n3060) );
  AOI22X1 U2057 ( .A(n1096), .B(n7019), .C(n6835), .D(n6920), .Y(n3062) );
  NAND3X1 U2059 ( .A(n5048), .B(n5241), .C(n5506), .Y(n3059) );
  AOI22X1 U2060 ( .A(n1101), .B(n7085), .C(n6824), .D(n6953), .Y(n3065) );
  AOI22X1 U2062 ( .A(n6817), .B(n7118), .C(n6812), .D(n7052), .Y(n3063) );
  NAND3X1 U2064 ( .A(n1116), .B(n5240), .C(n5505), .Y(n3067) );
  AOI22X1 U2065 ( .A(n6839), .B(n7811), .C(n6835), .D(n7712), .Y(n3069) );
  NAND3X1 U2067 ( .A(n5047), .B(n5239), .C(n5504), .Y(n3066) );
  AOI22X1 U2068 ( .A(n1101), .B(n7877), .C(n6824), .D(n7745), .Y(n3072) );
  AOI22X1 U2070 ( .A(n6817), .B(n7910), .C(n6812), .D(n7844), .Y(n3070) );
  NAND3X1 U2071 ( .A(n1124), .B(n5238), .C(n5503), .Y(n3074) );
  AOI22X1 U2072 ( .A(n1096), .B(n7547), .C(n6835), .D(n7448), .Y(n3076) );
  NAND3X1 U2074 ( .A(n5046), .B(n5237), .C(n5502), .Y(n3073) );
  AOI22X1 U2075 ( .A(n1101), .B(n7613), .C(n6824), .D(n7481), .Y(n3079) );
  AOI22X1 U2077 ( .A(n6817), .B(n7646), .C(n6812), .D(n7580), .Y(n3077) );
  NAND3X1 U2079 ( .A(n5160), .B(n3081), .C(n3082), .Y(n4487) );
  NOR3X1 U2080 ( .A(n5723), .B(n5756), .C(n5789), .Y(n3082) );
  NAND3X1 U2082 ( .A(n3260), .B(n5236), .C(n5501), .Y(n3087) );
  AOI22X1 U2083 ( .A(n1096), .B(n7284), .C(n6834), .D(n7185), .Y(n3089) );
  NAND3X1 U2085 ( .A(n5045), .B(n5235), .C(n5500), .Y(n3086) );
  AOI22X1 U2086 ( .A(n1101), .B(n7350), .C(n6825), .D(n7218), .Y(n3092) );
  AOI22X1 U2088 ( .A(n6817), .B(n7383), .C(n6813), .D(n7317), .Y(n3090) );
  NAND3X1 U2090 ( .A(n1108), .B(n5234), .C(n5499), .Y(n3094) );
  AOI22X1 U2091 ( .A(n1096), .B(n7020), .C(n6834), .D(n6921), .Y(n3096) );
  NAND3X1 U2093 ( .A(n5044), .B(n5233), .C(n5498), .Y(n3093) );
  AOI22X1 U2094 ( .A(n6829), .B(n7086), .C(n6825), .D(n6954), .Y(n3099) );
  AOI22X1 U2096 ( .A(n6816), .B(n7119), .C(n6813), .D(n7053), .Y(n3097) );
  NAND3X1 U2098 ( .A(n1116), .B(n5232), .C(n5497), .Y(n3101) );
  AOI22X1 U2099 ( .A(n1096), .B(n7812), .C(n6834), .D(n7713), .Y(n3103) );
  NAND3X1 U2101 ( .A(n5043), .B(n5231), .C(n5496), .Y(n3100) );
  AOI22X1 U2102 ( .A(n6830), .B(n7878), .C(n6825), .D(n7746), .Y(n3106) );
  AOI22X1 U2104 ( .A(n6818), .B(n7911), .C(n6813), .D(n7845), .Y(n3104) );
  NAND3X1 U2105 ( .A(n1124), .B(n5230), .C(n5495), .Y(n3108) );
  AOI22X1 U2106 ( .A(n1096), .B(n7548), .C(n6834), .D(n7449), .Y(n3110) );
  NAND3X1 U2108 ( .A(n5042), .B(n5229), .C(n5494), .Y(n3107) );
  AOI22X1 U2109 ( .A(n1101), .B(n7614), .C(n6825), .D(n7482), .Y(n3113) );
  AOI22X1 U2111 ( .A(n6818), .B(n7647), .C(n6813), .D(n7581), .Y(n3111) );
  NAND3X1 U2113 ( .A(n5159), .B(n3115), .C(n3116), .Y(n4488) );
  NOR3X1 U2114 ( .A(n5722), .B(n5755), .C(n5788), .Y(n3116) );
  NAND3X1 U2116 ( .A(n3260), .B(n5228), .C(n5493), .Y(n3121) );
  AOI22X1 U2117 ( .A(n1096), .B(n7285), .C(n6834), .D(n7186), .Y(n3123) );
  NAND3X1 U2119 ( .A(n5041), .B(n5227), .C(n5492), .Y(n3120) );
  AOI22X1 U2120 ( .A(n1101), .B(n7351), .C(n6825), .D(n7219), .Y(n3126) );
  AOI22X1 U2122 ( .A(n6816), .B(n7384), .C(n6813), .D(n7318), .Y(n3124) );
  NAND3X1 U2124 ( .A(n1108), .B(n5226), .C(n5491), .Y(n3128) );
  AOI22X1 U2125 ( .A(n1096), .B(n7021), .C(n6834), .D(n6922), .Y(n3130) );
  NAND3X1 U2127 ( .A(n5040), .B(n5225), .C(n5490), .Y(n3127) );
  AOI22X1 U2128 ( .A(n6830), .B(n7087), .C(n6825), .D(n6955), .Y(n3133) );
  AOI22X1 U2130 ( .A(n6818), .B(n7120), .C(n6813), .D(n7054), .Y(n3131) );
  NAND3X1 U2132 ( .A(n1116), .B(n5224), .C(n5489), .Y(n3135) );
  AOI22X1 U2133 ( .A(n6838), .B(n7813), .C(n6834), .D(n7714), .Y(n3137) );
  NAND3X1 U2135 ( .A(n5039), .B(n5223), .C(n5488), .Y(n3134) );
  AOI22X1 U2136 ( .A(n6830), .B(n7879), .C(n6825), .D(n7747), .Y(n3140) );
  AOI22X1 U2138 ( .A(n6817), .B(n7912), .C(n6813), .D(n7846), .Y(n3138) );
  NAND3X1 U2139 ( .A(n1124), .B(n5222), .C(n5487), .Y(n3142) );
  AOI22X1 U2140 ( .A(n1096), .B(n7549), .C(n6834), .D(n7450), .Y(n3144) );
  NAND3X1 U2142 ( .A(n5038), .B(n5221), .C(n5486), .Y(n3141) );
  AOI22X1 U2143 ( .A(n1101), .B(n7615), .C(n6825), .D(n7483), .Y(n3147) );
  AOI22X1 U2145 ( .A(n6817), .B(n7648), .C(n6813), .D(n7582), .Y(n3145) );
  NAND3X1 U2147 ( .A(n5158), .B(n3149), .C(n3150), .Y(n4489) );
  NOR3X1 U2148 ( .A(n5721), .B(n5754), .C(n5787), .Y(n3150) );
  NAND3X1 U2150 ( .A(n3260), .B(n5220), .C(n5485), .Y(n3155) );
  AOI22X1 U2151 ( .A(n1096), .B(n7286), .C(n6834), .D(n7187), .Y(n3157) );
  NAND3X1 U2153 ( .A(n5037), .B(n5219), .C(n5484), .Y(n3154) );
  AOI22X1 U2154 ( .A(n1101), .B(n7352), .C(n6825), .D(n7220), .Y(n3160) );
  AOI22X1 U2156 ( .A(n6818), .B(n7385), .C(n6813), .D(n7319), .Y(n3158) );
  NAND3X1 U2158 ( .A(n1108), .B(n5218), .C(n5483), .Y(n3162) );
  AOI22X1 U2159 ( .A(n6840), .B(n7022), .C(n6834), .D(n6923), .Y(n3164) );
  NAND3X1 U2161 ( .A(n5036), .B(n5217), .C(n5482), .Y(n3161) );
  AOI22X1 U2162 ( .A(n6828), .B(n7088), .C(n6825), .D(n6956), .Y(n3167) );
  AOI22X1 U2164 ( .A(n6818), .B(n7121), .C(n6813), .D(n7055), .Y(n3165) );
  NAND3X1 U2166 ( .A(n1116), .B(n5216), .C(n5481), .Y(n3169) );
  AOI22X1 U2167 ( .A(n6840), .B(n7814), .C(n6834), .D(n7715), .Y(n3171) );
  NAND3X1 U2169 ( .A(n5035), .B(n5215), .C(n5480), .Y(n3168) );
  AOI22X1 U2170 ( .A(n6830), .B(n7880), .C(n6825), .D(n7748), .Y(n3174) );
  AOI22X1 U2172 ( .A(n6818), .B(n7913), .C(n6813), .D(n7847), .Y(n3172) );
  NAND3X1 U2173 ( .A(n1124), .B(n5214), .C(n5479), .Y(n3176) );
  AOI22X1 U2174 ( .A(n6840), .B(n7550), .C(n6834), .D(n7451), .Y(n3178) );
  NAND3X1 U2176 ( .A(n5034), .B(n5213), .C(n5478), .Y(n3175) );
  AOI22X1 U2177 ( .A(n6830), .B(n7616), .C(n6825), .D(n7484), .Y(n3181) );
  AOI22X1 U2179 ( .A(n6818), .B(n7649), .C(n6813), .D(n7583), .Y(n3179) );
  NAND3X1 U2181 ( .A(n5157), .B(n3183), .C(n3184), .Y(n4490) );
  NOR3X1 U2182 ( .A(n5720), .B(n5753), .C(n5786), .Y(n3184) );
  NAND3X1 U2184 ( .A(n3260), .B(n5212), .C(n5477), .Y(n3189) );
  AOI22X1 U2185 ( .A(n6840), .B(n7287), .C(n6833), .D(n7188), .Y(n3191) );
  NAND3X1 U2187 ( .A(n5033), .B(n5211), .C(n5476), .Y(n3188) );
  AOI22X1 U2188 ( .A(n6828), .B(n7353), .C(n6826), .D(n7221), .Y(n3194) );
  AOI22X1 U2190 ( .A(n6818), .B(n7386), .C(n6814), .D(n7320), .Y(n3192) );
  NAND3X1 U2192 ( .A(n1108), .B(n5210), .C(n5475), .Y(n3196) );
  AOI22X1 U2193 ( .A(n6840), .B(n7023), .C(n6833), .D(n6924), .Y(n3198) );
  NAND3X1 U2195 ( .A(n5032), .B(n5209), .C(n5474), .Y(n3195) );
  AOI22X1 U2196 ( .A(n6829), .B(n7089), .C(n6826), .D(n6957), .Y(n3201) );
  AOI22X1 U2198 ( .A(n6818), .B(n7122), .C(n6814), .D(n7056), .Y(n3199) );
  NAND3X1 U2200 ( .A(n1116), .B(n5208), .C(n5473), .Y(n3203) );
  AOI22X1 U2201 ( .A(n6840), .B(n7815), .C(n6833), .D(n7716), .Y(n3205) );
  NAND3X1 U2203 ( .A(n5031), .B(n5207), .C(n5472), .Y(n3202) );
  AOI22X1 U2204 ( .A(n6828), .B(n7881), .C(n6826), .D(n7749), .Y(n3208) );
  AOI22X1 U2206 ( .A(n6818), .B(n7914), .C(n6814), .D(n7848), .Y(n3206) );
  NAND3X1 U2207 ( .A(n1124), .B(n5206), .C(n5471), .Y(n3210) );
  AOI22X1 U2208 ( .A(n6840), .B(n7551), .C(n6833), .D(n7452), .Y(n3212) );
  NAND3X1 U2210 ( .A(n5030), .B(n5205), .C(n5470), .Y(n3209) );
  AOI22X1 U2211 ( .A(n6828), .B(n7617), .C(n6826), .D(n7485), .Y(n3215) );
  AOI22X1 U2213 ( .A(n6818), .B(n7650), .C(n6814), .D(n7584), .Y(n3213) );
  NAND3X1 U2215 ( .A(n5156), .B(n3217), .C(n3218), .Y(n4491) );
  NOR3X1 U2216 ( .A(n5719), .B(n5752), .C(n5785), .Y(n3218) );
  NAND3X1 U2218 ( .A(n3260), .B(n5204), .C(n5469), .Y(n3223) );
  AOI22X1 U2219 ( .A(n6840), .B(n7288), .C(n6833), .D(n7189), .Y(n3225) );
  NAND3X1 U2221 ( .A(n5029), .B(n5203), .C(n5468), .Y(n3222) );
  AOI22X1 U2222 ( .A(n6829), .B(n7354), .C(n6826), .D(n7222), .Y(n3228) );
  AOI22X1 U2224 ( .A(n6818), .B(n7387), .C(n6814), .D(n7321), .Y(n3226) );
  NAND3X1 U2226 ( .A(n1108), .B(n5202), .C(n5467), .Y(n3230) );
  AOI22X1 U2227 ( .A(n6840), .B(n7024), .C(n6833), .D(n6925), .Y(n3232) );
  NAND3X1 U2229 ( .A(n5028), .B(n5201), .C(n5466), .Y(n3229) );
  AOI22X1 U2230 ( .A(n6830), .B(n7090), .C(n6826), .D(n6958), .Y(n3235) );
  AOI22X1 U2232 ( .A(n6818), .B(n7123), .C(n6814), .D(n7057), .Y(n3233) );
  NAND3X1 U2234 ( .A(n1116), .B(n5200), .C(n5465), .Y(n3237) );
  AOI22X1 U2235 ( .A(n6840), .B(n7816), .C(n6833), .D(n7717), .Y(n3239) );
  NAND3X1 U2237 ( .A(n5027), .B(n5199), .C(n5464), .Y(n3236) );
  AOI22X1 U2238 ( .A(n6829), .B(n7882), .C(n6826), .D(n7750), .Y(n3242) );
  AOI22X1 U2240 ( .A(n6818), .B(n7915), .C(n6814), .D(n7849), .Y(n3240) );
  NAND3X1 U2241 ( .A(n1124), .B(n5198), .C(n5463), .Y(n3244) );
  AOI22X1 U2242 ( .A(n6840), .B(n7552), .C(n6833), .D(n7453), .Y(n3246) );
  NAND3X1 U2244 ( .A(n5026), .B(n5197), .C(n5462), .Y(n3243) );
  AOI22X1 U2245 ( .A(n6829), .B(n7618), .C(n6826), .D(n7486), .Y(n3249) );
  AOI22X1 U2247 ( .A(n6818), .B(n7651), .C(n6814), .D(n7585), .Y(n3247) );
  NAND3X1 U2249 ( .A(n5155), .B(n3251), .C(n3252), .Y(n4492) );
  NOR3X1 U2250 ( .A(n5718), .B(n5751), .C(n5784), .Y(n3252) );
  NAND3X1 U2252 ( .A(n3260), .B(n5196), .C(n5461), .Y(n3257) );
  AOI22X1 U2253 ( .A(n6840), .B(n7289), .C(n6833), .D(n7190), .Y(n3259) );
  NAND3X1 U2255 ( .A(n5025), .B(n5195), .C(n5460), .Y(n3256) );
  AOI22X1 U2256 ( .A(n6830), .B(n7355), .C(n6826), .D(n7223), .Y(n3263) );
  AOI22X1 U2258 ( .A(n6818), .B(n7388), .C(n6814), .D(n7322), .Y(n3261) );
  NAND3X1 U2260 ( .A(n1108), .B(n5194), .C(n5459), .Y(n3265) );
  AOI22X1 U2261 ( .A(n6840), .B(n7025), .C(n6833), .D(n6926), .Y(n3267) );
  NAND3X1 U2263 ( .A(n5024), .B(n5193), .C(n5458), .Y(n3264) );
  AOI22X1 U2264 ( .A(n6828), .B(n7091), .C(n6826), .D(n6959), .Y(n3271) );
  AOI22X1 U2266 ( .A(n6818), .B(n7124), .C(n6814), .D(n7058), .Y(n3269) );
  NAND3X1 U2268 ( .A(n1116), .B(n5192), .C(n5457), .Y(n3273) );
  AOI22X1 U2269 ( .A(n6837), .B(n7817), .C(n6833), .D(n7718), .Y(n3275) );
  NOR3X1 U2271 ( .A(n15), .B(n16), .C(n6662), .Y(n1116) );
  NAND3X1 U2272 ( .A(n5023), .B(n5191), .C(n5456), .Y(n3272) );
  AOI22X1 U2273 ( .A(n1101), .B(n7883), .C(n6826), .D(n7751), .Y(n3279) );
  AOI22X1 U2275 ( .A(n6816), .B(n7916), .C(n6814), .D(n7850), .Y(n3277) );
  NAND3X1 U2276 ( .A(n1124), .B(n5190), .C(n5455), .Y(n3281) );
  AOI22X1 U2277 ( .A(n1096), .B(n7553), .C(n6833), .D(n7454), .Y(n3283) );
  NOR3X1 U2278 ( .A(n6855), .B(n12), .C(n6854), .Y(n1097) );
  NAND3X1 U2280 ( .A(n5022), .B(n5189), .C(n5454), .Y(n3280) );
  AOI22X1 U2281 ( .A(n1101), .B(n7619), .C(n6826), .D(n7487), .Y(n3286) );
  AOI22X1 U2283 ( .A(n1104), .B(n7652), .C(n6814), .D(n7586), .Y(n3284) );
  AOI21X1 U2285 ( .A(n16), .B(n6663), .C(n6846), .Y(n3290) );
  OAI21X1 U2286 ( .A(n6663), .B(n16), .C(n6857), .Y(n3292) );
  OAI21X1 U2288 ( .A(wr_ptr[0]), .B(n6807), .C(n3294), .Y(n2603) );
  NAND3X1 U2289 ( .A(n5154), .B(n6805), .C(n5453), .Y(n2602) );
  AOI22X1 U2290 ( .A(n3268), .B(n6734), .C(n3299), .D(n16), .Y(n3297) );
  NOR3X1 U2293 ( .A(n6856), .B(n16), .C(n6662), .Y(n1124) );
  OAI21X1 U2294 ( .A(n6853), .B(n6590), .C(n6456), .Y(n2601) );
  OAI21X1 U2296 ( .A(n5817), .B(n6854), .C(n4661), .Y(n2600) );
  NAND3X1 U2297 ( .A(n12), .B(n6854), .C(n3276), .Y(n3302) );
  OAI21X1 U2298 ( .A(n5817), .B(n6855), .C(n3303), .Y(n2599) );
  OAI21X1 U2299 ( .A(n1096), .B(n3287), .C(n3276), .Y(n3303) );
  AOI21X1 U2300 ( .A(n6853), .B(n3276), .C(n3299), .Y(n3301) );
  OAI21X1 U2301 ( .A(n5188), .B(n6856), .C(n4660), .Y(n2598) );
  NAND3X1 U2302 ( .A(n3276), .B(n6856), .C(n6810), .Y(n3305) );
  AOI21X1 U2303 ( .A(n3276), .B(n6734), .C(n3299), .Y(n3304) );
  NAND3X1 U2304 ( .A(n14), .B(n12), .C(n13), .Y(n3298) );
  NAND3X1 U2308 ( .A(n3307), .B(n3308), .C(n3309), .Y(n4624) );
  NOR3X1 U2309 ( .A(n3310), .B(fillcount[0]), .C(n3311), .Y(n3309) );
  OAI21X1 U2310 ( .A(n6519), .B(n6857), .C(n6518), .Y(n2597) );
  NAND3X1 U2311 ( .A(n6852), .B(n3293), .C(n6520), .Y(n3313) );
  AOI21X1 U2313 ( .A(n3293), .B(n6860), .C(n3315), .Y(n3312) );
  OAI21X1 U2314 ( .A(n6850), .B(n6858), .C(n6266), .Y(n2596) );
  NAND3X1 U2315 ( .A(wr_ptr[0]), .B(n6858), .C(n3293), .Y(n3316) );
  OAI21X1 U2316 ( .A(n6328), .B(n6859), .C(n3319), .Y(n2595) );
  AOI21X1 U2317 ( .A(n3293), .B(n6858), .C(n3317), .Y(n3318) );
  OAI21X1 U2318 ( .A(wr_ptr[0]), .B(n6807), .C(n6735), .Y(n3317) );
  OAI21X1 U2319 ( .A(n6851), .B(n6860), .C(n6453), .Y(n2594) );
  NAND3X1 U2320 ( .A(n3293), .B(n6860), .C(n6852), .Y(n3321) );
  OAI21X1 U2321 ( .A(n6852), .B(n6807), .C(n6735), .Y(n3315) );
  OAI21X1 U2324 ( .A(n3323), .B(n6861), .C(n6329), .Y(n2593) );
  OAI21X1 U2326 ( .A(n3323), .B(n6862), .C(n6738), .Y(n2592) );
  OAI21X1 U2328 ( .A(n3323), .B(n6863), .C(n6667), .Y(n2591) );
  OAI21X1 U2330 ( .A(n3323), .B(n6864), .C(n4757), .Y(n2590) );
  OAI21X1 U2332 ( .A(n3323), .B(n6865), .C(n4756), .Y(n2589) );
  OAI21X1 U2334 ( .A(n3323), .B(n6866), .C(n4755), .Y(n2588) );
  OAI21X1 U2336 ( .A(n3323), .B(n6867), .C(n6457), .Y(n2587) );
  OAI21X1 U2338 ( .A(n3323), .B(n6868), .C(n6392), .Y(n2586) );
  OAI21X1 U2340 ( .A(n3323), .B(n6869), .C(n6330), .Y(n2585) );
  OAI21X1 U2342 ( .A(n3323), .B(n6870), .C(n6038), .Y(n2584) );
  OAI21X1 U2344 ( .A(n3323), .B(n6871), .C(n6523), .Y(n2583) );
  OAI21X1 U2346 ( .A(n3323), .B(n6872), .C(n6267), .Y(n2582) );
  OAI21X1 U2348 ( .A(n3323), .B(n6873), .C(n5983), .Y(n2581) );
  OAI21X1 U2350 ( .A(n3323), .B(n6874), .C(n6595), .Y(n2580) );
  OAI21X1 U2352 ( .A(n3323), .B(n6875), .C(n5928), .Y(n2579) );
  OAI21X1 U2354 ( .A(n3323), .B(n6876), .C(n5873), .Y(n2578) );
  OAI21X1 U2356 ( .A(n3323), .B(n6877), .C(n5818), .Y(n2577) );
  OAI21X1 U2358 ( .A(n3323), .B(n6878), .C(n6209), .Y(n2576) );
  OAI21X1 U2360 ( .A(n3323), .B(n6879), .C(n6152), .Y(n2575) );
  OAI21X1 U2362 ( .A(n3323), .B(n6880), .C(n6095), .Y(n2574) );
  OAI21X1 U2364 ( .A(n3323), .B(n6881), .C(n6039), .Y(n2573) );
  OAI21X1 U2366 ( .A(n3323), .B(n6882), .C(n6739), .Y(n2572) );
  OAI21X1 U2368 ( .A(n3323), .B(n6883), .C(n6668), .Y(n2571) );
  OAI21X1 U2370 ( .A(n3323), .B(n6884), .C(n6596), .Y(n2570) );
  OAI21X1 U2372 ( .A(n3323), .B(n6885), .C(n6524), .Y(n2569) );
  OAI21X1 U2374 ( .A(n3323), .B(n6886), .C(n5984), .Y(n2568) );
  OAI21X1 U2376 ( .A(n3323), .B(n6887), .C(n5929), .Y(n2567) );
  OAI21X1 U2378 ( .A(n3323), .B(n6888), .C(n5874), .Y(n2566) );
  OAI21X1 U2380 ( .A(n3323), .B(n6889), .C(n5819), .Y(n2565) );
  OAI21X1 U2382 ( .A(n3323), .B(n6890), .C(n6210), .Y(n2564) );
  OAI21X1 U2384 ( .A(n3323), .B(n6891), .C(n6153), .Y(n2563) );
  OAI21X1 U2386 ( .A(n3323), .B(n6892), .C(n6096), .Y(n2562) );
  OAI21X1 U2388 ( .A(n3323), .B(n6893), .C(n6040), .Y(n2561) );
  OAI21X1 U2390 ( .A(n6594), .B(n6808), .C(n6842), .Y(n3323) );
  OAI21X1 U2391 ( .A(n3391), .B(n6894), .C(n6268), .Y(n2560) );
  OAI21X1 U2393 ( .A(n3391), .B(n6895), .C(n6669), .Y(n2559) );
  OAI21X1 U2395 ( .A(n3391), .B(n6896), .C(n6740), .Y(n2558) );
  OAI21X1 U2397 ( .A(n3391), .B(n6897), .C(n4754), .Y(n2557) );
  OAI21X1 U2399 ( .A(n3391), .B(n6898), .C(n4753), .Y(n2556) );
  OAI21X1 U2401 ( .A(n3391), .B(n6899), .C(n4752), .Y(n2555) );
  OAI21X1 U2403 ( .A(n3391), .B(n6900), .C(n6393), .Y(n2554) );
  OAI21X1 U2405 ( .A(n3391), .B(n6901), .C(n6458), .Y(n2553) );
  OAI21X1 U2407 ( .A(n3391), .B(n6902), .C(n6269), .Y(n2552) );
  OAI21X1 U2409 ( .A(n3391), .B(n6903), .C(n6097), .Y(n2551) );
  OAI21X1 U2411 ( .A(n3391), .B(n6904), .C(n6597), .Y(n2550) );
  OAI21X1 U2413 ( .A(n3391), .B(n6905), .C(n6331), .Y(n2549) );
  OAI21X1 U2415 ( .A(n3391), .B(n6906), .C(n5930), .Y(n2548) );
  OAI21X1 U2417 ( .A(n3391), .B(n6907), .C(n6525), .Y(n2547) );
  OAI21X1 U2419 ( .A(n3391), .B(n6908), .C(n5985), .Y(n2546) );
  OAI21X1 U2421 ( .A(n3391), .B(n6909), .C(n5820), .Y(n2545) );
  OAI21X1 U2423 ( .A(n3391), .B(n6910), .C(n5875), .Y(n2544) );
  OAI21X1 U2425 ( .A(n3391), .B(n6911), .C(n6154), .Y(n2543) );
  OAI21X1 U2427 ( .A(n3391), .B(n6912), .C(n6211), .Y(n2542) );
  OAI21X1 U2429 ( .A(n3391), .B(n6913), .C(n6041), .Y(n2541) );
  OAI21X1 U2431 ( .A(n3391), .B(n6914), .C(n6098), .Y(n2540) );
  OAI21X1 U2433 ( .A(n3391), .B(n6915), .C(n6670), .Y(n2539) );
  OAI21X1 U2435 ( .A(n3391), .B(n6916), .C(n6741), .Y(n2538) );
  OAI21X1 U2437 ( .A(n3391), .B(n6917), .C(n6526), .Y(n2537) );
  OAI21X1 U2439 ( .A(n3391), .B(n6918), .C(n6598), .Y(n2536) );
  OAI21X1 U2441 ( .A(n3391), .B(n6919), .C(n5931), .Y(n2535) );
  OAI21X1 U2443 ( .A(n3391), .B(n6920), .C(n5986), .Y(n2534) );
  OAI21X1 U2445 ( .A(n3391), .B(n6921), .C(n5821), .Y(n2533) );
  OAI21X1 U2447 ( .A(n3391), .B(n6922), .C(n5876), .Y(n2532) );
  OAI21X1 U2449 ( .A(n3391), .B(n6923), .C(n6155), .Y(n2531) );
  OAI21X1 U2451 ( .A(n3391), .B(n6924), .C(n6212), .Y(n2530) );
  OAI21X1 U2453 ( .A(n3391), .B(n6925), .C(n6042), .Y(n2529) );
  OAI21X1 U2455 ( .A(n3391), .B(n6926), .C(n6099), .Y(n2528) );
  OAI21X1 U2457 ( .A(n6808), .B(n6521), .C(n6842), .Y(n3391) );
  OAI21X1 U2458 ( .A(n3426), .B(n6927), .C(n6459), .Y(n2527) );
  OAI21X1 U2460 ( .A(n3426), .B(n6928), .C(n6599), .Y(n2526) );
  OAI21X1 U2462 ( .A(n3426), .B(n6929), .C(n6527), .Y(n2525) );
  OAI21X1 U2464 ( .A(n3426), .B(n6930), .C(n4751), .Y(n2524) );
  OAI21X1 U2466 ( .A(n3426), .B(n6931), .C(n4750), .Y(n2523) );
  OAI21X1 U2468 ( .A(n3426), .B(n6932), .C(n4749), .Y(n2522) );
  OAI21X1 U2470 ( .A(n3426), .B(n6933), .C(n6332), .Y(n2521) );
  OAI21X1 U2472 ( .A(n3426), .B(n6934), .C(n6270), .Y(n2520) );
  OAI21X1 U2474 ( .A(n3426), .B(n6935), .C(n6460), .Y(n2519) );
  OAI21X1 U2476 ( .A(n3426), .B(n6936), .C(n6156), .Y(n2518) );
  OAI21X1 U2478 ( .A(n3426), .B(n6937), .C(n6671), .Y(n2517) );
  OAI21X1 U2480 ( .A(n3426), .B(n6938), .C(n6394), .Y(n2516) );
  OAI21X1 U2482 ( .A(n3426), .B(n6939), .C(n5877), .Y(n2515) );
  OAI21X1 U2484 ( .A(n3426), .B(n6940), .C(n6742), .Y(n2514) );
  OAI21X1 U2486 ( .A(n3426), .B(n6941), .C(n5822), .Y(n2513) );
  OAI21X1 U2488 ( .A(n3426), .B(n6942), .C(n5987), .Y(n2512) );
  OAI21X1 U2490 ( .A(n3426), .B(n6943), .C(n5932), .Y(n2511) );
  OAI21X1 U2492 ( .A(n3426), .B(n6944), .C(n6100), .Y(n2510) );
  OAI21X1 U2494 ( .A(n3426), .B(n6945), .C(n6043), .Y(n2509) );
  OAI21X1 U2496 ( .A(n3426), .B(n6946), .C(n6213), .Y(n2508) );
  OAI21X1 U2498 ( .A(n3426), .B(n6947), .C(n6157), .Y(n2507) );
  OAI21X1 U2500 ( .A(n3426), .B(n6948), .C(n6600), .Y(n2506) );
  OAI21X1 U2502 ( .A(n3426), .B(n6949), .C(n6528), .Y(n2505) );
  OAI21X1 U2504 ( .A(n3426), .B(n6950), .C(n6743), .Y(n2504) );
  OAI21X1 U2506 ( .A(n3426), .B(n6951), .C(n6672), .Y(n2503) );
  OAI21X1 U2508 ( .A(n3426), .B(n6952), .C(n5878), .Y(n2502) );
  OAI21X1 U2510 ( .A(n3426), .B(n6953), .C(n5823), .Y(n2501) );
  OAI21X1 U2512 ( .A(n3426), .B(n6954), .C(n5988), .Y(n2500) );
  OAI21X1 U2514 ( .A(n3426), .B(n6955), .C(n5933), .Y(n2499) );
  OAI21X1 U2516 ( .A(n3426), .B(n6956), .C(n6101), .Y(n2498) );
  OAI21X1 U2518 ( .A(n3426), .B(n6957), .C(n6044), .Y(n2497) );
  OAI21X1 U2520 ( .A(n3426), .B(n6958), .C(n6214), .Y(n2496) );
  OAI21X1 U2522 ( .A(n3426), .B(n6959), .C(n6158), .Y(n2495) );
  OAI21X1 U2524 ( .A(n6808), .B(n6454), .C(n6842), .Y(n3426) );
  OAI21X1 U2525 ( .A(n3461), .B(n6960), .C(n6395), .Y(n2494) );
  OAI21X1 U2527 ( .A(n3461), .B(n6961), .C(n6529), .Y(n2493) );
  OAI21X1 U2529 ( .A(n3461), .B(n6962), .C(n6601), .Y(n2492) );
  OAI21X1 U2531 ( .A(n3461), .B(n6963), .C(n4748), .Y(n2491) );
  OAI21X1 U2533 ( .A(n3461), .B(n6964), .C(n4747), .Y(n2490) );
  OAI21X1 U2535 ( .A(n3461), .B(n6965), .C(n4746), .Y(n2489) );
  OAI21X1 U2537 ( .A(n3461), .B(n6966), .C(n6271), .Y(n2488) );
  OAI21X1 U2539 ( .A(n3461), .B(n6967), .C(n6333), .Y(n2487) );
  OAI21X1 U2541 ( .A(n3461), .B(n6968), .C(n6396), .Y(n2486) );
  OAI21X1 U2543 ( .A(n3461), .B(n6969), .C(n6215), .Y(n2485) );
  OAI21X1 U2545 ( .A(n3461), .B(n6970), .C(n6744), .Y(n2484) );
  OAI21X1 U2547 ( .A(n3461), .B(n6971), .C(n6461), .Y(n2483) );
  OAI21X1 U2549 ( .A(n3461), .B(n6972), .C(n5824), .Y(n2482) );
  OAI21X1 U2551 ( .A(n3461), .B(n6973), .C(n6673), .Y(n2481) );
  OAI21X1 U2553 ( .A(n3461), .B(n6974), .C(n5879), .Y(n2480) );
  OAI21X1 U2555 ( .A(n3461), .B(n6975), .C(n5934), .Y(n2479) );
  OAI21X1 U2557 ( .A(n3461), .B(n6976), .C(n5989), .Y(n2478) );
  OAI21X1 U2559 ( .A(n3461), .B(n6977), .C(n6045), .Y(n2477) );
  OAI21X1 U2561 ( .A(n3461), .B(n6978), .C(n6102), .Y(n2476) );
  OAI21X1 U2563 ( .A(n3461), .B(n6979), .C(n6159), .Y(n2475) );
  OAI21X1 U2565 ( .A(n3461), .B(n6980), .C(n6216), .Y(n2474) );
  OAI21X1 U2567 ( .A(n3461), .B(n6981), .C(n6530), .Y(n2473) );
  OAI21X1 U2569 ( .A(n3461), .B(n6982), .C(n6602), .Y(n2472) );
  OAI21X1 U2571 ( .A(n3461), .B(n6983), .C(n6674), .Y(n2471) );
  OAI21X1 U2573 ( .A(n3461), .B(n6984), .C(n6745), .Y(n2470) );
  OAI21X1 U2575 ( .A(n3461), .B(n6985), .C(n5825), .Y(n2469) );
  OAI21X1 U2577 ( .A(n3461), .B(n6986), .C(n5880), .Y(n2468) );
  OAI21X1 U2579 ( .A(n3461), .B(n6987), .C(n5935), .Y(n2467) );
  OAI21X1 U2581 ( .A(n3461), .B(n6988), .C(n5990), .Y(n2466) );
  OAI21X1 U2583 ( .A(n3461), .B(n6989), .C(n6046), .Y(n2465) );
  OAI21X1 U2585 ( .A(n3461), .B(n6990), .C(n6103), .Y(n2464) );
  OAI21X1 U2587 ( .A(n3461), .B(n6991), .C(n6160), .Y(n2463) );
  OAI21X1 U2589 ( .A(n3461), .B(n6992), .C(n6217), .Y(n2462) );
  OAI21X1 U2591 ( .A(n6808), .B(n6665), .C(n6842), .Y(n3461) );
  OAI21X1 U2592 ( .A(n3496), .B(n6993), .C(n6104), .Y(n2461) );
  OAI21X1 U2594 ( .A(n3496), .B(n6994), .C(n5991), .Y(n2460) );
  OAI21X1 U2596 ( .A(n3496), .B(n6995), .C(n5936), .Y(n2459) );
  OAI21X1 U2598 ( .A(n3496), .B(n6996), .C(n4745), .Y(n2458) );
  OAI21X1 U2600 ( .A(n3496), .B(n6997), .C(n4744), .Y(n2457) );
  OAI21X1 U2602 ( .A(n3496), .B(n6998), .C(n4743), .Y(n2456) );
  OAI21X1 U2604 ( .A(n3496), .B(n6999), .C(n6218), .Y(n2455) );
  OAI21X1 U2606 ( .A(n3496), .B(n7000), .C(n6161), .Y(n2454) );
  OAI21X1 U2608 ( .A(n3496), .B(n7001), .C(n6105), .Y(n2453) );
  OAI21X1 U2610 ( .A(n3496), .B(n7002), .C(n6272), .Y(n2452) );
  OAI21X1 U2612 ( .A(n3496), .B(n7003), .C(n5826), .Y(n2451) );
  OAI21X1 U2614 ( .A(n3496), .B(n7004), .C(n6047), .Y(n2450) );
  OAI21X1 U2616 ( .A(n3496), .B(n7005), .C(n6746), .Y(n2449) );
  OAI21X1 U2618 ( .A(n3496), .B(n7006), .C(n5881), .Y(n2448) );
  OAI21X1 U2620 ( .A(n3496), .B(n7007), .C(n6675), .Y(n2447) );
  OAI21X1 U2622 ( .A(n3496), .B(n7008), .C(n6603), .Y(n2446) );
  OAI21X1 U2624 ( .A(n3496), .B(n7009), .C(n6531), .Y(n2445) );
  OAI21X1 U2626 ( .A(n3496), .B(n7010), .C(n6462), .Y(n2444) );
  OAI21X1 U2628 ( .A(n3496), .B(n7011), .C(n6397), .Y(n2443) );
  OAI21X1 U2630 ( .A(n3496), .B(n7012), .C(n6334), .Y(n2442) );
  OAI21X1 U2632 ( .A(n3496), .B(n7013), .C(n6273), .Y(n2441) );
  OAI21X1 U2634 ( .A(n3496), .B(n7014), .C(n5992), .Y(n2440) );
  OAI21X1 U2636 ( .A(n3496), .B(n7015), .C(n5937), .Y(n2439) );
  OAI21X1 U2638 ( .A(n3496), .B(n7016), .C(n5882), .Y(n2438) );
  OAI21X1 U2640 ( .A(n3496), .B(n7017), .C(n5827), .Y(n2437) );
  OAI21X1 U2642 ( .A(n3496), .B(n7018), .C(n6747), .Y(n2436) );
  OAI21X1 U2644 ( .A(n3496), .B(n7019), .C(n6676), .Y(n2435) );
  OAI21X1 U2646 ( .A(n3496), .B(n7020), .C(n6604), .Y(n2434) );
  OAI21X1 U2648 ( .A(n3496), .B(n7021), .C(n6532), .Y(n2433) );
  OAI21X1 U2650 ( .A(n3496), .B(n7022), .C(n6463), .Y(n2432) );
  OAI21X1 U2652 ( .A(n3496), .B(n7023), .C(n6398), .Y(n2431) );
  OAI21X1 U2654 ( .A(n3496), .B(n7024), .C(n6335), .Y(n2430) );
  OAI21X1 U2656 ( .A(n3496), .B(n7025), .C(n6274), .Y(n2429) );
  OAI21X1 U2658 ( .A(n6666), .B(n6808), .C(n6842), .Y(n3496) );
  OAI21X1 U2659 ( .A(n3530), .B(n7026), .C(n6048), .Y(n2428) );
  OAI21X1 U2661 ( .A(n3530), .B(n7027), .C(n5938), .Y(n2427) );
  OAI21X1 U2663 ( .A(n3530), .B(n7028), .C(n5993), .Y(n2426) );
  OAI21X1 U2665 ( .A(n3530), .B(n7029), .C(n4742), .Y(n2425) );
  OAI21X1 U2667 ( .A(n3530), .B(n7030), .C(n4741), .Y(n2424) );
  OAI21X1 U2669 ( .A(n3530), .B(n7031), .C(n4740), .Y(n2423) );
  OAI21X1 U2671 ( .A(n3530), .B(n7032), .C(n6162), .Y(n2422) );
  OAI21X1 U2673 ( .A(n3530), .B(n7033), .C(n6219), .Y(n2421) );
  OAI21X1 U2675 ( .A(n3530), .B(n7034), .C(n6049), .Y(n2420) );
  OAI21X1 U2677 ( .A(n3530), .B(n7035), .C(n6336), .Y(n2419) );
  OAI21X1 U2679 ( .A(n3530), .B(n7036), .C(n5883), .Y(n2418) );
  OAI21X1 U2681 ( .A(n3530), .B(n7037), .C(n6106), .Y(n2417) );
  OAI21X1 U2683 ( .A(n3530), .B(n7038), .C(n6677), .Y(n2416) );
  OAI21X1 U2685 ( .A(n3530), .B(n7039), .C(n5828), .Y(n2415) );
  OAI21X1 U2687 ( .A(n3530), .B(n7040), .C(n6748), .Y(n2414) );
  OAI21X1 U2689 ( .A(n3530), .B(n7041), .C(n6533), .Y(n2413) );
  OAI21X1 U2691 ( .A(n3530), .B(n7042), .C(n6605), .Y(n2412) );
  OAI21X1 U2693 ( .A(n3530), .B(n7043), .C(n6399), .Y(n2411) );
  OAI21X1 U2695 ( .A(n3530), .B(n7044), .C(n6464), .Y(n2410) );
  OAI21X1 U2697 ( .A(n3530), .B(n7045), .C(n6275), .Y(n2409) );
  OAI21X1 U2699 ( .A(n3530), .B(n7046), .C(n6337), .Y(n2408) );
  OAI21X1 U2701 ( .A(n3530), .B(n7047), .C(n5939), .Y(n2407) );
  OAI21X1 U2703 ( .A(n3530), .B(n7048), .C(n5994), .Y(n2406) );
  OAI21X1 U2705 ( .A(n3530), .B(n7049), .C(n5829), .Y(n2405) );
  OAI21X1 U2707 ( .A(n3530), .B(n7050), .C(n5884), .Y(n2404) );
  OAI21X1 U2709 ( .A(n3530), .B(n7051), .C(n6678), .Y(n2403) );
  OAI21X1 U2711 ( .A(n3530), .B(n7052), .C(n6749), .Y(n2402) );
  OAI21X1 U2713 ( .A(n3530), .B(n7053), .C(n6534), .Y(n2401) );
  OAI21X1 U2715 ( .A(n3530), .B(n7054), .C(n6606), .Y(n2400) );
  OAI21X1 U2717 ( .A(n3530), .B(n7055), .C(n6400), .Y(n2399) );
  OAI21X1 U2719 ( .A(n3530), .B(n7056), .C(n6465), .Y(n2398) );
  OAI21X1 U2721 ( .A(n3530), .B(n7057), .C(n6276), .Y(n2397) );
  OAI21X1 U2723 ( .A(n3530), .B(n7058), .C(n6338), .Y(n2396) );
  OAI21X1 U2725 ( .A(n6808), .B(n6455), .C(n6842), .Y(n3530) );
  OAI21X1 U2726 ( .A(n3565), .B(n7059), .C(n6220), .Y(n2395) );
  OAI21X1 U2728 ( .A(n3565), .B(n7060), .C(n5885), .Y(n2394) );
  OAI21X1 U2730 ( .A(n3565), .B(n7061), .C(n5830), .Y(n2393) );
  OAI21X1 U2732 ( .A(n3565), .B(n7062), .C(n4739), .Y(n2392) );
  OAI21X1 U2734 ( .A(n3565), .B(n7063), .C(n4738), .Y(n2391) );
  OAI21X1 U2736 ( .A(n3565), .B(n7064), .C(n4737), .Y(n2390) );
  OAI21X1 U2738 ( .A(n3565), .B(n7065), .C(n6107), .Y(n2389) );
  OAI21X1 U2740 ( .A(n3565), .B(n7066), .C(n6050), .Y(n2388) );
  OAI21X1 U2742 ( .A(n3565), .B(n7067), .C(n6221), .Y(n2387) );
  OAI21X1 U2744 ( .A(n3565), .B(n7068), .C(n6401), .Y(n2386) );
  OAI21X1 U2746 ( .A(n3565), .B(n7069), .C(n5940), .Y(n2385) );
  OAI21X1 U2748 ( .A(n3565), .B(n7070), .C(n6163), .Y(n2384) );
  OAI21X1 U2750 ( .A(n3565), .B(n7071), .C(n6607), .Y(n2383) );
  OAI21X1 U2752 ( .A(n3565), .B(n7072), .C(n5995), .Y(n2382) );
  OAI21X1 U2754 ( .A(n3565), .B(n7073), .C(n6535), .Y(n2381) );
  OAI21X1 U2756 ( .A(n3565), .B(n7074), .C(n6750), .Y(n2380) );
  OAI21X1 U2758 ( .A(n3565), .B(n7075), .C(n6679), .Y(n2379) );
  OAI21X1 U2760 ( .A(n3565), .B(n7076), .C(n6339), .Y(n2378) );
  OAI21X1 U2762 ( .A(n3565), .B(n7077), .C(n6277), .Y(n2377) );
  OAI21X1 U2764 ( .A(n3565), .B(n7078), .C(n6466), .Y(n2376) );
  OAI21X1 U2766 ( .A(n3565), .B(n7079), .C(n6402), .Y(n2375) );
  OAI21X1 U2768 ( .A(n3565), .B(n7080), .C(n5886), .Y(n2374) );
  OAI21X1 U2770 ( .A(n3565), .B(n7081), .C(n5831), .Y(n2373) );
  OAI21X1 U2772 ( .A(n3565), .B(n7082), .C(n5996), .Y(n2372) );
  OAI21X1 U2774 ( .A(n3565), .B(n7083), .C(n5941), .Y(n2371) );
  OAI21X1 U2776 ( .A(n3565), .B(n7084), .C(n6608), .Y(n2370) );
  OAI21X1 U2778 ( .A(n3565), .B(n7085), .C(n6536), .Y(n2369) );
  OAI21X1 U2780 ( .A(n3565), .B(n7086), .C(n6751), .Y(n2368) );
  OAI21X1 U2782 ( .A(n3565), .B(n7087), .C(n6680), .Y(n2367) );
  OAI21X1 U2784 ( .A(n3565), .B(n7088), .C(n6340), .Y(n2366) );
  OAI21X1 U2786 ( .A(n3565), .B(n7089), .C(n6278), .Y(n2365) );
  OAI21X1 U2788 ( .A(n3565), .B(n7090), .C(n6467), .Y(n2364) );
  OAI21X1 U2790 ( .A(n3565), .B(n7091), .C(n6403), .Y(n2363) );
  OAI21X1 U2792 ( .A(n6808), .B(n6522), .C(n6842), .Y(n3565) );
  OAI21X1 U2793 ( .A(n3600), .B(n7092), .C(n6164), .Y(n2362) );
  OAI21X1 U2795 ( .A(n3600), .B(n7093), .C(n5832), .Y(n2361) );
  OAI21X1 U2797 ( .A(n3600), .B(n7094), .C(n5887), .Y(n2360) );
  OAI21X1 U2799 ( .A(n3600), .B(n7095), .C(n4736), .Y(n2359) );
  OAI21X1 U2801 ( .A(n3600), .B(n7096), .C(n4735), .Y(n2358) );
  OAI21X1 U2803 ( .A(n3600), .B(n7097), .C(n4734), .Y(n2357) );
  OAI21X1 U2805 ( .A(n3600), .B(n7098), .C(n6051), .Y(n2356) );
  OAI21X1 U2807 ( .A(n3600), .B(n7099), .C(n6108), .Y(n2355) );
  OAI21X1 U2809 ( .A(n3600), .B(n7100), .C(n6165), .Y(n2354) );
  OAI21X1 U2811 ( .A(n3600), .B(n7101), .C(n6468), .Y(n2353) );
  OAI21X1 U2813 ( .A(n3600), .B(n7102), .C(n5997), .Y(n2352) );
  OAI21X1 U2815 ( .A(n3600), .B(n7103), .C(n6222), .Y(n2351) );
  OAI21X1 U2817 ( .A(n3600), .B(n7104), .C(n6537), .Y(n2350) );
  OAI21X1 U2819 ( .A(n3600), .B(n7105), .C(n5942), .Y(n2349) );
  OAI21X1 U2821 ( .A(n3600), .B(n7106), .C(n6609), .Y(n2348) );
  OAI21X1 U2823 ( .A(n3600), .B(n7107), .C(n6681), .Y(n2347) );
  OAI21X1 U2825 ( .A(n3600), .B(n7108), .C(n6752), .Y(n2346) );
  OAI21X1 U2827 ( .A(n3600), .B(n7109), .C(n6279), .Y(n2345) );
  OAI21X1 U2829 ( .A(n3600), .B(n7110), .C(n6341), .Y(n2344) );
  OAI21X1 U2831 ( .A(n3600), .B(n7111), .C(n6404), .Y(n2343) );
  OAI21X1 U2833 ( .A(n3600), .B(n7112), .C(n6469), .Y(n2342) );
  OAI21X1 U2835 ( .A(n3600), .B(n7113), .C(n5833), .Y(n2341) );
  OAI21X1 U2837 ( .A(n3600), .B(n7114), .C(n5888), .Y(n2340) );
  OAI21X1 U2839 ( .A(n3600), .B(n7115), .C(n5943), .Y(n2339) );
  OAI21X1 U2841 ( .A(n3600), .B(n7116), .C(n5998), .Y(n2338) );
  OAI21X1 U2843 ( .A(n3600), .B(n7117), .C(n6538), .Y(n2337) );
  OAI21X1 U2845 ( .A(n3600), .B(n7118), .C(n6610), .Y(n2336) );
  OAI21X1 U2847 ( .A(n3600), .B(n7119), .C(n6682), .Y(n2335) );
  OAI21X1 U2849 ( .A(n3600), .B(n7120), .C(n6753), .Y(n2334) );
  OAI21X1 U2851 ( .A(n3600), .B(n7121), .C(n6280), .Y(n2333) );
  OAI21X1 U2853 ( .A(n3600), .B(n7122), .C(n6342), .Y(n2332) );
  OAI21X1 U2855 ( .A(n3600), .B(n7123), .C(n6405), .Y(n2331) );
  OAI21X1 U2857 ( .A(n3600), .B(n7124), .C(n6470), .Y(n2330) );
  OAI21X1 U2859 ( .A(n6808), .B(n6593), .C(n6842), .Y(n3600) );
  NAND3X1 U2860 ( .A(wr_ptr[4]), .B(wr_ptr[3]), .C(put), .Y(n3390) );
  OAI21X1 U2861 ( .A(n3635), .B(n7125), .C(n5889), .Y(n2329) );
  OAI21X1 U2863 ( .A(n3635), .B(n7126), .C(n6223), .Y(n2328) );
  OAI21X1 U2865 ( .A(n3635), .B(n7127), .C(n6166), .Y(n2327) );
  OAI21X1 U2867 ( .A(n3635), .B(n7128), .C(n4733), .Y(n2326) );
  OAI21X1 U2869 ( .A(n3635), .B(n7129), .C(n4732), .Y(n2325) );
  OAI21X1 U2871 ( .A(n3635), .B(n7130), .C(n4731), .Y(n2324) );
  OAI21X1 U2873 ( .A(n3635), .B(n7131), .C(n5999), .Y(n2323) );
  OAI21X1 U2875 ( .A(n3635), .B(n7132), .C(n5944), .Y(n2322) );
  OAI21X1 U2877 ( .A(n3635), .B(n7133), .C(n5890), .Y(n2321) );
  OAI21X1 U2879 ( .A(n3635), .B(n7134), .C(n6539), .Y(n2320) );
  OAI21X1 U2881 ( .A(n3635), .B(n7135), .C(n6052), .Y(n2319) );
  OAI21X1 U2883 ( .A(n3635), .B(n7136), .C(n5834), .Y(n2318) );
  OAI21X1 U2885 ( .A(n3635), .B(n7137), .C(n6471), .Y(n2317) );
  OAI21X1 U2887 ( .A(n3635), .B(n7138), .C(n6109), .Y(n2316) );
  OAI21X1 U2889 ( .A(n3635), .B(n7139), .C(n6406), .Y(n2315) );
  OAI21X1 U2891 ( .A(n3635), .B(n7140), .C(n6343), .Y(n2314) );
  OAI21X1 U2893 ( .A(n3635), .B(n7141), .C(n6281), .Y(n2313) );
  OAI21X1 U2895 ( .A(n3635), .B(n7142), .C(n6754), .Y(n2312) );
  OAI21X1 U2897 ( .A(n3635), .B(n7143), .C(n6683), .Y(n2311) );
  OAI21X1 U2899 ( .A(n3635), .B(n7144), .C(n6611), .Y(n2310) );
  OAI21X1 U2901 ( .A(n3635), .B(n7145), .C(n6540), .Y(n2309) );
  OAI21X1 U2903 ( .A(n3635), .B(n7146), .C(n6224), .Y(n2308) );
  OAI21X1 U2905 ( .A(n3635), .B(n7147), .C(n6167), .Y(n2307) );
  OAI21X1 U2907 ( .A(n3635), .B(n7148), .C(n6110), .Y(n2306) );
  OAI21X1 U2909 ( .A(n3635), .B(n7149), .C(n6053), .Y(n2305) );
  OAI21X1 U2911 ( .A(n3635), .B(n7150), .C(n6472), .Y(n2304) );
  OAI21X1 U2913 ( .A(n3635), .B(n7151), .C(n6407), .Y(n2303) );
  OAI21X1 U2915 ( .A(n3635), .B(n7152), .C(n6344), .Y(n2302) );
  OAI21X1 U2917 ( .A(n3635), .B(n7153), .C(n6282), .Y(n2301) );
  OAI21X1 U2919 ( .A(n3635), .B(n7154), .C(n6755), .Y(n2300) );
  OAI21X1 U2921 ( .A(n3635), .B(n7155), .C(n6684), .Y(n2299) );
  OAI21X1 U2923 ( .A(n3635), .B(n7156), .C(n6612), .Y(n2298) );
  OAI21X1 U2925 ( .A(n3635), .B(n7157), .C(n6541), .Y(n2297) );
  OAI21X1 U2927 ( .A(n6594), .B(n6736), .C(n6842), .Y(n3635) );
  OAI21X1 U2928 ( .A(n3670), .B(n7158), .C(n5835), .Y(n2296) );
  OAI21X1 U2930 ( .A(n3670), .B(n7159), .C(n6168), .Y(n2295) );
  OAI21X1 U2932 ( .A(n3670), .B(n7160), .C(n6225), .Y(n2294) );
  OAI21X1 U2934 ( .A(n3670), .B(n7161), .C(n4730), .Y(n2293) );
  OAI21X1 U2936 ( .A(n3670), .B(n7162), .C(n4729), .Y(n2292) );
  OAI21X1 U2938 ( .A(n3670), .B(n7163), .C(n4728), .Y(n2291) );
  OAI21X1 U2940 ( .A(n3670), .B(n7164), .C(n5945), .Y(n2290) );
  OAI21X1 U2942 ( .A(n3670), .B(n7165), .C(n6000), .Y(n2289) );
  OAI21X1 U2944 ( .A(n3670), .B(n7166), .C(n5836), .Y(n2288) );
  OAI21X1 U2946 ( .A(n3670), .B(n7167), .C(n6613), .Y(n2287) );
  OAI21X1 U2948 ( .A(n3670), .B(n7168), .C(n6111), .Y(n2286) );
  OAI21X1 U2950 ( .A(n3670), .B(n7169), .C(n5891), .Y(n2285) );
  OAI21X1 U2952 ( .A(n3670), .B(n7170), .C(n6408), .Y(n2284) );
  OAI21X1 U2954 ( .A(n3670), .B(n7171), .C(n6054), .Y(n2283) );
  OAI21X1 U2956 ( .A(n3670), .B(n7172), .C(n6473), .Y(n2282) );
  OAI21X1 U2958 ( .A(n3670), .B(n7173), .C(n6283), .Y(n2281) );
  OAI21X1 U2960 ( .A(n3670), .B(n7174), .C(n6345), .Y(n2280) );
  OAI21X1 U2962 ( .A(n3670), .B(n7175), .C(n6685), .Y(n2279) );
  OAI21X1 U2964 ( .A(n3670), .B(n7176), .C(n6756), .Y(n2278) );
  OAI21X1 U2966 ( .A(n3670), .B(n7177), .C(n6542), .Y(n2277) );
  OAI21X1 U2968 ( .A(n3670), .B(n7178), .C(n6614), .Y(n2276) );
  OAI21X1 U2970 ( .A(n3670), .B(n7179), .C(n6169), .Y(n2275) );
  OAI21X1 U2972 ( .A(n3670), .B(n7180), .C(n6226), .Y(n2274) );
  OAI21X1 U2974 ( .A(n3670), .B(n7181), .C(n6055), .Y(n2273) );
  OAI21X1 U2976 ( .A(n3670), .B(n7182), .C(n6112), .Y(n2272) );
  OAI21X1 U2978 ( .A(n3670), .B(n7183), .C(n6409), .Y(n2271) );
  OAI21X1 U2980 ( .A(n3670), .B(n7184), .C(n6474), .Y(n2270) );
  OAI21X1 U2982 ( .A(n3670), .B(n7185), .C(n6284), .Y(n2269) );
  OAI21X1 U2984 ( .A(n3670), .B(n7186), .C(n6346), .Y(n2268) );
  OAI21X1 U2986 ( .A(n3670), .B(n7187), .C(n6686), .Y(n2267) );
  OAI21X1 U2988 ( .A(n3670), .B(n7188), .C(n6757), .Y(n2266) );
  OAI21X1 U2990 ( .A(n3670), .B(n7189), .C(n6543), .Y(n2265) );
  OAI21X1 U2992 ( .A(n3670), .B(n7190), .C(n6615), .Y(n2264) );
  OAI21X1 U2994 ( .A(n6521), .B(n6736), .C(n6843), .Y(n3670) );
  OAI21X1 U2995 ( .A(n3704), .B(n7191), .C(n6001), .Y(n2263) );
  OAI21X1 U2997 ( .A(n3704), .B(n7192), .C(n6113), .Y(n2262) );
  OAI21X1 U2999 ( .A(n3704), .B(n7193), .C(n6056), .Y(n2261) );
  OAI21X1 U3001 ( .A(n3704), .B(n7194), .C(n4727), .Y(n2260) );
  OAI21X1 U3003 ( .A(n3704), .B(n7195), .C(n4726), .Y(n2259) );
  OAI21X1 U3005 ( .A(n3704), .B(n7196), .C(n4725), .Y(n2258) );
  OAI21X1 U3007 ( .A(n3704), .B(n7197), .C(n5892), .Y(n2257) );
  OAI21X1 U3009 ( .A(n3704), .B(n7198), .C(n5837), .Y(n2256) );
  OAI21X1 U3011 ( .A(n3704), .B(n7199), .C(n6002), .Y(n2255) );
  OAI21X1 U3013 ( .A(n3704), .B(n7200), .C(n6687), .Y(n2254) );
  OAI21X1 U3015 ( .A(n3704), .B(n7201), .C(n6170), .Y(n2253) );
  OAI21X1 U3017 ( .A(n3704), .B(n7202), .C(n5946), .Y(n2252) );
  OAI21X1 U3019 ( .A(n3704), .B(n7203), .C(n6347), .Y(n2251) );
  OAI21X1 U3021 ( .A(n3704), .B(n7204), .C(n6227), .Y(n2250) );
  OAI21X1 U3023 ( .A(n3704), .B(n7205), .C(n6285), .Y(n2249) );
  OAI21X1 U3025 ( .A(n3704), .B(n7206), .C(n6475), .Y(n2248) );
  OAI21X1 U3027 ( .A(n3704), .B(n7207), .C(n6410), .Y(n2247) );
  OAI21X1 U3029 ( .A(n3704), .B(n7208), .C(n6616), .Y(n2246) );
  OAI21X1 U3031 ( .A(n3704), .B(n7209), .C(n6544), .Y(n2245) );
  OAI21X1 U3033 ( .A(n3704), .B(n7210), .C(n6758), .Y(n2244) );
  OAI21X1 U3035 ( .A(n3704), .B(n7211), .C(n6688), .Y(n2243) );
  OAI21X1 U3037 ( .A(n3704), .B(n7212), .C(n6114), .Y(n2242) );
  OAI21X1 U3039 ( .A(n3704), .B(n7213), .C(n6057), .Y(n2241) );
  OAI21X1 U3041 ( .A(n3704), .B(n7214), .C(n6228), .Y(n2240) );
  OAI21X1 U3043 ( .A(n3704), .B(n7215), .C(n6171), .Y(n2239) );
  OAI21X1 U3045 ( .A(n3704), .B(n7216), .C(n6348), .Y(n2238) );
  OAI21X1 U3047 ( .A(n3704), .B(n7217), .C(n6286), .Y(n2237) );
  OAI21X1 U3049 ( .A(n3704), .B(n7218), .C(n6476), .Y(n2236) );
  OAI21X1 U3051 ( .A(n3704), .B(n7219), .C(n6411), .Y(n2235) );
  OAI21X1 U3053 ( .A(n3704), .B(n7220), .C(n6617), .Y(n2234) );
  OAI21X1 U3055 ( .A(n3704), .B(n7221), .C(n6545), .Y(n2233) );
  OAI21X1 U3057 ( .A(n3704), .B(n7222), .C(n6759), .Y(n2232) );
  OAI21X1 U3059 ( .A(n3704), .B(n7223), .C(n6689), .Y(n2231) );
  OAI21X1 U3061 ( .A(n6454), .B(n6736), .C(n6843), .Y(n3704) );
  OAI21X1 U3062 ( .A(n3738), .B(n7224), .C(n5947), .Y(n2230) );
  OAI21X1 U3064 ( .A(n3738), .B(n7225), .C(n6058), .Y(n2229) );
  OAI21X1 U3066 ( .A(n3738), .B(n7226), .C(n6115), .Y(n2228) );
  OAI21X1 U3068 ( .A(n3738), .B(n7227), .C(n4724), .Y(n2227) );
  OAI21X1 U3070 ( .A(n3738), .B(n7228), .C(n4723), .Y(n2226) );
  OAI21X1 U3072 ( .A(n3738), .B(n7229), .C(n4722), .Y(n2225) );
  OAI21X1 U3074 ( .A(n3738), .B(n7230), .C(n5838), .Y(n2224) );
  OAI21X1 U3076 ( .A(n3738), .B(n7231), .C(n5893), .Y(n2223) );
  OAI21X1 U3078 ( .A(n3738), .B(n7232), .C(n5948), .Y(n2222) );
  OAI21X1 U3080 ( .A(n3738), .B(n7233), .C(n6760), .Y(n2221) );
  OAI21X1 U3082 ( .A(n3738), .B(n7234), .C(n6229), .Y(n2220) );
  OAI21X1 U3084 ( .A(n3738), .B(n7235), .C(n6003), .Y(n2219) );
  OAI21X1 U3086 ( .A(n3738), .B(n7236), .C(n6287), .Y(n2218) );
  OAI21X1 U3088 ( .A(n3738), .B(n7237), .C(n6172), .Y(n2217) );
  OAI21X1 U3090 ( .A(n3738), .B(n7238), .C(n6349), .Y(n2216) );
  OAI21X1 U3092 ( .A(n3738), .B(n7239), .C(n6412), .Y(n2215) );
  OAI21X1 U3094 ( .A(n3738), .B(n7240), .C(n6477), .Y(n2214) );
  OAI21X1 U3096 ( .A(n3738), .B(n7241), .C(n6546), .Y(n2213) );
  OAI21X1 U3098 ( .A(n3738), .B(n7242), .C(n6618), .Y(n2212) );
  OAI21X1 U3100 ( .A(n3738), .B(n7243), .C(n6690), .Y(n2211) );
  OAI21X1 U3102 ( .A(n3738), .B(n7244), .C(n6761), .Y(n2210) );
  OAI21X1 U3104 ( .A(n3738), .B(n7245), .C(n6059), .Y(n2209) );
  OAI21X1 U3106 ( .A(n3738), .B(n7246), .C(n6116), .Y(n2208) );
  OAI21X1 U3108 ( .A(n3738), .B(n7247), .C(n6173), .Y(n2207) );
  OAI21X1 U3110 ( .A(n3738), .B(n7248), .C(n6230), .Y(n2206) );
  OAI21X1 U3112 ( .A(n3738), .B(n7249), .C(n6288), .Y(n2205) );
  OAI21X1 U3114 ( .A(n3738), .B(n7250), .C(n6350), .Y(n2204) );
  OAI21X1 U3116 ( .A(n3738), .B(n7251), .C(n6413), .Y(n2203) );
  OAI21X1 U3118 ( .A(n3738), .B(n7252), .C(n6478), .Y(n2202) );
  OAI21X1 U3120 ( .A(n3738), .B(n7253), .C(n6547), .Y(n2201) );
  OAI21X1 U3122 ( .A(n3738), .B(n7254), .C(n6619), .Y(n2200) );
  OAI21X1 U3124 ( .A(n3738), .B(n7255), .C(n6691), .Y(n2199) );
  OAI21X1 U3126 ( .A(n3738), .B(n7256), .C(n6762), .Y(n2198) );
  OAI21X1 U3128 ( .A(n6665), .B(n6736), .C(n6843), .Y(n3738) );
  OAI21X1 U3129 ( .A(n3772), .B(n7257), .C(n6351), .Y(n2197) );
  OAI21X1 U3131 ( .A(n3772), .B(n7258), .C(n6763), .Y(n2196) );
  OAI21X1 U3133 ( .A(n3772), .B(n7259), .C(n6692), .Y(n2195) );
  OAI21X1 U3135 ( .A(n3772), .B(n7260), .C(n4721), .Y(n2194) );
  OAI21X1 U3137 ( .A(n3772), .B(n7261), .C(n4720), .Y(n2193) );
  OAI21X1 U3139 ( .A(n3772), .B(n7262), .C(n4719), .Y(n2192) );
  OAI21X1 U3141 ( .A(n3772), .B(n7263), .C(n6479), .Y(n2191) );
  OAI21X1 U3143 ( .A(n3772), .B(n7264), .C(n6414), .Y(n2190) );
  OAI21X1 U3145 ( .A(n3772), .B(n7265), .C(n6352), .Y(n2189) );
  OAI21X1 U3147 ( .A(n3772), .B(n7266), .C(n6060), .Y(n2188) );
  OAI21X1 U3149 ( .A(n3772), .B(n7267), .C(n6548), .Y(n2187) );
  OAI21X1 U3151 ( .A(n3772), .B(n7268), .C(n6289), .Y(n2186) );
  OAI21X1 U3153 ( .A(n3772), .B(n7269), .C(n6004), .Y(n2185) );
  OAI21X1 U3155 ( .A(n3772), .B(n7270), .C(n6620), .Y(n2184) );
  OAI21X1 U3157 ( .A(n3772), .B(n7271), .C(n5949), .Y(n2183) );
  OAI21X1 U3159 ( .A(n3772), .B(n7272), .C(n5894), .Y(n2182) );
  OAI21X1 U3161 ( .A(n3772), .B(n7273), .C(n5839), .Y(n2181) );
  OAI21X1 U3163 ( .A(n3772), .B(n7274), .C(n6231), .Y(n2180) );
  OAI21X1 U3165 ( .A(n3772), .B(n7275), .C(n6174), .Y(n2179) );
  OAI21X1 U3167 ( .A(n3772), .B(n7276), .C(n6117), .Y(n2178) );
  OAI21X1 U3169 ( .A(n3772), .B(n7277), .C(n6061), .Y(n2177) );
  OAI21X1 U3171 ( .A(n3772), .B(n7278), .C(n6764), .Y(n2176) );
  OAI21X1 U3173 ( .A(n3772), .B(n7279), .C(n6693), .Y(n2175) );
  OAI21X1 U3175 ( .A(n3772), .B(n7280), .C(n6621), .Y(n2174) );
  OAI21X1 U3177 ( .A(n3772), .B(n7281), .C(n6549), .Y(n2173) );
  OAI21X1 U3179 ( .A(n3772), .B(n7282), .C(n6005), .Y(n2172) );
  OAI21X1 U3181 ( .A(n3772), .B(n7283), .C(n5950), .Y(n2171) );
  OAI21X1 U3183 ( .A(n3772), .B(n7284), .C(n5895), .Y(n2170) );
  OAI21X1 U3185 ( .A(n3772), .B(n7285), .C(n5840), .Y(n2169) );
  OAI21X1 U3187 ( .A(n3772), .B(n7286), .C(n6232), .Y(n2168) );
  OAI21X1 U3189 ( .A(n3772), .B(n7287), .C(n6175), .Y(n2167) );
  OAI21X1 U3191 ( .A(n3772), .B(n7288), .C(n6118), .Y(n2166) );
  OAI21X1 U3193 ( .A(n3772), .B(n7289), .C(n6062), .Y(n2165) );
  OAI21X1 U3195 ( .A(n6666), .B(n6736), .C(n6843), .Y(n3772) );
  OAI21X1 U3196 ( .A(n3806), .B(n7290), .C(n6290), .Y(n2164) );
  OAI21X1 U3198 ( .A(n3806), .B(n7291), .C(n6694), .Y(n2163) );
  OAI21X1 U3200 ( .A(n3806), .B(n7292), .C(n6765), .Y(n2162) );
  OAI21X1 U3202 ( .A(n3806), .B(n7293), .C(n4718), .Y(n2161) );
  OAI21X1 U3204 ( .A(n3806), .B(n7294), .C(n4717), .Y(n2160) );
  OAI21X1 U3206 ( .A(n3806), .B(n7295), .C(n4716), .Y(n2159) );
  OAI21X1 U3208 ( .A(n3806), .B(n7296), .C(n6415), .Y(n2158) );
  OAI21X1 U3210 ( .A(n3806), .B(n7297), .C(n6480), .Y(n2157) );
  OAI21X1 U3212 ( .A(n3806), .B(n7298), .C(n6291), .Y(n2156) );
  OAI21X1 U3214 ( .A(n3806), .B(n7299), .C(n6119), .Y(n2155) );
  OAI21X1 U3216 ( .A(n3806), .B(n7300), .C(n6622), .Y(n2154) );
  OAI21X1 U3218 ( .A(n3806), .B(n7301), .C(n6353), .Y(n2153) );
  OAI21X1 U3220 ( .A(n3806), .B(n7302), .C(n5951), .Y(n2152) );
  OAI21X1 U3222 ( .A(n3806), .B(n7303), .C(n6550), .Y(n2151) );
  OAI21X1 U3224 ( .A(n3806), .B(n7304), .C(n6006), .Y(n2150) );
  OAI21X1 U3226 ( .A(n3806), .B(n7305), .C(n5841), .Y(n2149) );
  OAI21X1 U3228 ( .A(n3806), .B(n7306), .C(n5896), .Y(n2148) );
  OAI21X1 U3230 ( .A(n3806), .B(n7307), .C(n6176), .Y(n2147) );
  OAI21X1 U3232 ( .A(n3806), .B(n7308), .C(n6233), .Y(n2146) );
  OAI21X1 U3234 ( .A(n3806), .B(n7309), .C(n6063), .Y(n2145) );
  OAI21X1 U3236 ( .A(n3806), .B(n7310), .C(n6120), .Y(n2144) );
  OAI21X1 U3238 ( .A(n3806), .B(n7311), .C(n6695), .Y(n2143) );
  OAI21X1 U3240 ( .A(n3806), .B(n7312), .C(n6766), .Y(n2142) );
  OAI21X1 U3242 ( .A(n3806), .B(n7313), .C(n6551), .Y(n2141) );
  OAI21X1 U3244 ( .A(n3806), .B(n7314), .C(n6623), .Y(n2140) );
  OAI21X1 U3246 ( .A(n3806), .B(n7315), .C(n5952), .Y(n2139) );
  OAI21X1 U3248 ( .A(n3806), .B(n7316), .C(n6007), .Y(n2138) );
  OAI21X1 U3250 ( .A(n3806), .B(n7317), .C(n5842), .Y(n2137) );
  OAI21X1 U3252 ( .A(n3806), .B(n7318), .C(n5897), .Y(n2136) );
  OAI21X1 U3254 ( .A(n3806), .B(n7319), .C(n6177), .Y(n2135) );
  OAI21X1 U3256 ( .A(n3806), .B(n7320), .C(n6234), .Y(n2134) );
  OAI21X1 U3258 ( .A(n3806), .B(n7321), .C(n6064), .Y(n2133) );
  OAI21X1 U3260 ( .A(n3806), .B(n7322), .C(n6121), .Y(n2132) );
  OAI21X1 U3262 ( .A(n6455), .B(n6736), .C(n6843), .Y(n3806) );
  OAI21X1 U3263 ( .A(n3840), .B(n7323), .C(n6481), .Y(n2131) );
  OAI21X1 U3265 ( .A(n3840), .B(n7324), .C(n6624), .Y(n2130) );
  OAI21X1 U3267 ( .A(n3840), .B(n7325), .C(n6552), .Y(n2129) );
  OAI21X1 U3269 ( .A(n3840), .B(n7326), .C(n4715), .Y(n2128) );
  OAI21X1 U3271 ( .A(n3840), .B(n7327), .C(n4714), .Y(n2127) );
  OAI21X1 U3273 ( .A(n3840), .B(n7328), .C(n4713), .Y(n2126) );
  OAI21X1 U3275 ( .A(n3840), .B(n7329), .C(n6354), .Y(n2125) );
  OAI21X1 U3277 ( .A(n3840), .B(n7330), .C(n6292), .Y(n2124) );
  OAI21X1 U3279 ( .A(n3840), .B(n7331), .C(n6482), .Y(n2123) );
  OAI21X1 U3281 ( .A(n3840), .B(n7332), .C(n6178), .Y(n2122) );
  OAI21X1 U3283 ( .A(n3840), .B(n7333), .C(n6696), .Y(n2121) );
  OAI21X1 U3285 ( .A(n3840), .B(n7334), .C(n6416), .Y(n2120) );
  OAI21X1 U3287 ( .A(n3840), .B(n7335), .C(n5898), .Y(n2119) );
  OAI21X1 U3289 ( .A(n3840), .B(n7336), .C(n6767), .Y(n2118) );
  OAI21X1 U3291 ( .A(n3840), .B(n7337), .C(n5843), .Y(n2117) );
  OAI21X1 U3293 ( .A(n3840), .B(n7338), .C(n6008), .Y(n2116) );
  OAI21X1 U3295 ( .A(n3840), .B(n7339), .C(n5953), .Y(n2115) );
  OAI21X1 U3297 ( .A(n3840), .B(n7340), .C(n6122), .Y(n2114) );
  OAI21X1 U3299 ( .A(n3840), .B(n7341), .C(n6065), .Y(n2113) );
  OAI21X1 U3301 ( .A(n3840), .B(n7342), .C(n6235), .Y(n2112) );
  OAI21X1 U3303 ( .A(n3840), .B(n7343), .C(n6179), .Y(n2111) );
  OAI21X1 U3305 ( .A(n3840), .B(n7344), .C(n6625), .Y(n2110) );
  OAI21X1 U3307 ( .A(n3840), .B(n7345), .C(n6553), .Y(n2109) );
  OAI21X1 U3309 ( .A(n3840), .B(n7346), .C(n6768), .Y(n2108) );
  OAI21X1 U3311 ( .A(n3840), .B(n7347), .C(n6697), .Y(n2107) );
  OAI21X1 U3313 ( .A(n3840), .B(n7348), .C(n5899), .Y(n2106) );
  OAI21X1 U3315 ( .A(n3840), .B(n7349), .C(n5844), .Y(n2105) );
  OAI21X1 U3317 ( .A(n3840), .B(n7350), .C(n6009), .Y(n2104) );
  OAI21X1 U3319 ( .A(n3840), .B(n7351), .C(n5954), .Y(n2103) );
  OAI21X1 U3321 ( .A(n3840), .B(n7352), .C(n6123), .Y(n2102) );
  OAI21X1 U3323 ( .A(n3840), .B(n7353), .C(n6066), .Y(n2101) );
  OAI21X1 U3325 ( .A(n3840), .B(n7354), .C(n6236), .Y(n2100) );
  OAI21X1 U3327 ( .A(n3840), .B(n7355), .C(n6180), .Y(n2099) );
  OAI21X1 U3329 ( .A(n6522), .B(n6736), .C(n6843), .Y(n3840) );
  OAI21X1 U3330 ( .A(n3874), .B(n7356), .C(n6417), .Y(n2098) );
  OAI21X1 U3332 ( .A(n3874), .B(n7357), .C(n6554), .Y(n2097) );
  OAI21X1 U3334 ( .A(n3874), .B(n7358), .C(n6626), .Y(n2096) );
  OAI21X1 U3336 ( .A(n3874), .B(n7359), .C(n4712), .Y(n2095) );
  OAI21X1 U3338 ( .A(n3874), .B(n7360), .C(n4711), .Y(n2094) );
  OAI21X1 U3340 ( .A(n3874), .B(n7361), .C(n4710), .Y(n2093) );
  OAI21X1 U3342 ( .A(n3874), .B(n7362), .C(n6293), .Y(n2092) );
  OAI21X1 U3344 ( .A(n3874), .B(n7363), .C(n6355), .Y(n2091) );
  OAI21X1 U3346 ( .A(n3874), .B(n7364), .C(n6418), .Y(n2090) );
  OAI21X1 U3348 ( .A(n3874), .B(n7365), .C(n6237), .Y(n2089) );
  OAI21X1 U3350 ( .A(n3874), .B(n7366), .C(n6769), .Y(n2088) );
  OAI21X1 U3352 ( .A(n3874), .B(n7367), .C(n6483), .Y(n2087) );
  OAI21X1 U3354 ( .A(n3874), .B(n7368), .C(n5845), .Y(n2086) );
  OAI21X1 U3356 ( .A(n3874), .B(n7369), .C(n6698), .Y(n2085) );
  OAI21X1 U3358 ( .A(n3874), .B(n7370), .C(n5900), .Y(n2084) );
  OAI21X1 U3360 ( .A(n3874), .B(n7371), .C(n5955), .Y(n2083) );
  OAI21X1 U3362 ( .A(n3874), .B(n7372), .C(n6010), .Y(n2082) );
  OAI21X1 U3364 ( .A(n3874), .B(n7373), .C(n6067), .Y(n2081) );
  OAI21X1 U3366 ( .A(n3874), .B(n7374), .C(n6124), .Y(n2080) );
  OAI21X1 U3368 ( .A(n3874), .B(n7375), .C(n6181), .Y(n2079) );
  OAI21X1 U3370 ( .A(n3874), .B(n7376), .C(n6238), .Y(n2078) );
  OAI21X1 U3372 ( .A(n3874), .B(n7377), .C(n6555), .Y(n2077) );
  OAI21X1 U3374 ( .A(n3874), .B(n7378), .C(n6627), .Y(n2076) );
  OAI21X1 U3376 ( .A(n3874), .B(n7379), .C(n6699), .Y(n2075) );
  OAI21X1 U3378 ( .A(n3874), .B(n7380), .C(n6770), .Y(n2074) );
  OAI21X1 U3380 ( .A(n3874), .B(n7381), .C(n5846), .Y(n2073) );
  OAI21X1 U3382 ( .A(n3874), .B(n7382), .C(n5901), .Y(n2072) );
  OAI21X1 U3384 ( .A(n3874), .B(n7383), .C(n5956), .Y(n2071) );
  OAI21X1 U3386 ( .A(n3874), .B(n7384), .C(n6011), .Y(n2070) );
  OAI21X1 U3388 ( .A(n3874), .B(n7385), .C(n6068), .Y(n2069) );
  OAI21X1 U3390 ( .A(n3874), .B(n7386), .C(n6125), .Y(n2068) );
  OAI21X1 U3392 ( .A(n3874), .B(n7387), .C(n6182), .Y(n2067) );
  OAI21X1 U3394 ( .A(n3874), .B(n7388), .C(n6239), .Y(n2066) );
  OAI21X1 U3396 ( .A(n6593), .B(n6736), .C(n6843), .Y(n3874) );
  NAND3X1 U3397 ( .A(wr_ptr[4]), .B(n6860), .C(put), .Y(n3669) );
  OAI21X1 U3398 ( .A(n3908), .B(n7389), .C(n6126), .Y(n2065) );
  OAI21X1 U3400 ( .A(n3908), .B(n7390), .C(n6012), .Y(n2064) );
  OAI21X1 U3402 ( .A(n3908), .B(n7391), .C(n5957), .Y(n2063) );
  OAI21X1 U3404 ( .A(n3908), .B(n7392), .C(n4709), .Y(n2062) );
  OAI21X1 U3406 ( .A(n3908), .B(n7393), .C(n4708), .Y(n2061) );
  OAI21X1 U3408 ( .A(n3908), .B(n7394), .C(n4707), .Y(n2060) );
  OAI21X1 U3410 ( .A(n3908), .B(n7395), .C(n6240), .Y(n2059) );
  OAI21X1 U3412 ( .A(n3908), .B(n7396), .C(n6183), .Y(n2058) );
  OAI21X1 U3414 ( .A(n3908), .B(n7397), .C(n6127), .Y(n2057) );
  OAI21X1 U3416 ( .A(n3908), .B(n7398), .C(n6294), .Y(n2056) );
  OAI21X1 U3418 ( .A(n3908), .B(n7399), .C(n5847), .Y(n2055) );
  OAI21X1 U3420 ( .A(n3908), .B(n7400), .C(n6069), .Y(n2054) );
  OAI21X1 U3422 ( .A(n3908), .B(n7401), .C(n6771), .Y(n2053) );
  OAI21X1 U3424 ( .A(n3908), .B(n7402), .C(n5902), .Y(n2052) );
  OAI21X1 U3426 ( .A(n3908), .B(n7403), .C(n6700), .Y(n2051) );
  OAI21X1 U3428 ( .A(n3908), .B(n7404), .C(n6628), .Y(n2050) );
  OAI21X1 U3430 ( .A(n3908), .B(n7405), .C(n6556), .Y(n2049) );
  OAI21X1 U3432 ( .A(n3908), .B(n7406), .C(n6484), .Y(n2048) );
  OAI21X1 U3434 ( .A(n3908), .B(n7407), .C(n6419), .Y(n2047) );
  OAI21X1 U3436 ( .A(n3908), .B(n7408), .C(n6356), .Y(n2046) );
  OAI21X1 U3438 ( .A(n3908), .B(n7409), .C(n6295), .Y(n2045) );
  OAI21X1 U3440 ( .A(n3908), .B(n7410), .C(n6013), .Y(n2044) );
  OAI21X1 U3442 ( .A(n3908), .B(n7411), .C(n5958), .Y(n2043) );
  OAI21X1 U3444 ( .A(n3908), .B(n7412), .C(n5903), .Y(n2042) );
  OAI21X1 U3446 ( .A(n3908), .B(n7413), .C(n5848), .Y(n2041) );
  OAI21X1 U3448 ( .A(n3908), .B(n7414), .C(n6772), .Y(n2040) );
  OAI21X1 U3450 ( .A(n3908), .B(n7415), .C(n6701), .Y(n2039) );
  OAI21X1 U3452 ( .A(n3908), .B(n7416), .C(n6629), .Y(n2038) );
  OAI21X1 U3454 ( .A(n3908), .B(n7417), .C(n6557), .Y(n2037) );
  OAI21X1 U3456 ( .A(n3908), .B(n7418), .C(n6485), .Y(n2036) );
  OAI21X1 U3458 ( .A(n3908), .B(n7419), .C(n6420), .Y(n2035) );
  OAI21X1 U3460 ( .A(n3908), .B(n7420), .C(n6357), .Y(n2034) );
  OAI21X1 U3462 ( .A(n3908), .B(n7421), .C(n6296), .Y(n2033) );
  OAI21X1 U3464 ( .A(n6594), .B(n6737), .C(n6843), .Y(n3908) );
  OAI21X1 U3465 ( .A(n3943), .B(n7422), .C(n6070), .Y(n2032) );
  OAI21X1 U3467 ( .A(n3943), .B(n7423), .C(n5959), .Y(n2031) );
  OAI21X1 U3469 ( .A(n3943), .B(n7424), .C(n6014), .Y(n2030) );
  OAI21X1 U3471 ( .A(n3943), .B(n7425), .C(n4706), .Y(n2029) );
  OAI21X1 U3473 ( .A(n3943), .B(n7426), .C(n4705), .Y(n2028) );
  OAI21X1 U3475 ( .A(n3943), .B(n7427), .C(n4704), .Y(n2027) );
  OAI21X1 U3477 ( .A(n3943), .B(n7428), .C(n6184), .Y(n2026) );
  OAI21X1 U3479 ( .A(n3943), .B(n7429), .C(n6241), .Y(n2025) );
  OAI21X1 U3481 ( .A(n3943), .B(n7430), .C(n6071), .Y(n2024) );
  OAI21X1 U3483 ( .A(n3943), .B(n7431), .C(n6358), .Y(n2023) );
  OAI21X1 U3485 ( .A(n3943), .B(n7432), .C(n5904), .Y(n2022) );
  OAI21X1 U3487 ( .A(n3943), .B(n7433), .C(n6128), .Y(n2021) );
  OAI21X1 U3489 ( .A(n3943), .B(n7434), .C(n6702), .Y(n2020) );
  OAI21X1 U3491 ( .A(n3943), .B(n7435), .C(n5849), .Y(n2019) );
  OAI21X1 U3493 ( .A(n3943), .B(n7436), .C(n6773), .Y(n2018) );
  OAI21X1 U3495 ( .A(n3943), .B(n7437), .C(n6558), .Y(n2017) );
  OAI21X1 U3497 ( .A(n3943), .B(n7438), .C(n6630), .Y(n2016) );
  OAI21X1 U3499 ( .A(n3943), .B(n7439), .C(n6421), .Y(n2015) );
  OAI21X1 U3501 ( .A(n3943), .B(n7440), .C(n6486), .Y(n2014) );
  OAI21X1 U3503 ( .A(n3943), .B(n7441), .C(n6297), .Y(n2013) );
  OAI21X1 U3505 ( .A(n3943), .B(n7442), .C(n6359), .Y(n2012) );
  OAI21X1 U3507 ( .A(n3943), .B(n7443), .C(n5960), .Y(n2011) );
  OAI21X1 U3509 ( .A(n3943), .B(n7444), .C(n6015), .Y(n2010) );
  OAI21X1 U3511 ( .A(n3943), .B(n7445), .C(n5850), .Y(n2009) );
  OAI21X1 U3513 ( .A(n3943), .B(n7446), .C(n5905), .Y(n2008) );
  OAI21X1 U3515 ( .A(n3943), .B(n7447), .C(n6703), .Y(n2007) );
  OAI21X1 U3517 ( .A(n3943), .B(n7448), .C(n6774), .Y(n2006) );
  OAI21X1 U3519 ( .A(n3943), .B(n7449), .C(n6559), .Y(n2005) );
  OAI21X1 U3521 ( .A(n3943), .B(n7450), .C(n6631), .Y(n2004) );
  OAI21X1 U3523 ( .A(n3943), .B(n7451), .C(n6422), .Y(n2003) );
  OAI21X1 U3525 ( .A(n3943), .B(n7452), .C(n6487), .Y(n2002) );
  OAI21X1 U3527 ( .A(n3943), .B(n7453), .C(n6298), .Y(n2001) );
  OAI21X1 U3529 ( .A(n3943), .B(n7454), .C(n6360), .Y(n2000) );
  OAI21X1 U3531 ( .A(n6521), .B(n6737), .C(n6843), .Y(n3943) );
  OAI21X1 U3532 ( .A(n3977), .B(n7455), .C(n6242), .Y(n1999) );
  OAI21X1 U3534 ( .A(n3977), .B(n7456), .C(n5906), .Y(n1998) );
  OAI21X1 U3536 ( .A(n3977), .B(n7457), .C(n5851), .Y(n1997) );
  OAI21X1 U3538 ( .A(n3977), .B(n7458), .C(n4703), .Y(n1996) );
  OAI21X1 U3540 ( .A(n3977), .B(n7459), .C(n4702), .Y(n1995) );
  OAI21X1 U3542 ( .A(n3977), .B(n7460), .C(n4701), .Y(n1994) );
  OAI21X1 U3544 ( .A(n3977), .B(n7461), .C(n6129), .Y(n1993) );
  OAI21X1 U3546 ( .A(n3977), .B(n7462), .C(n6072), .Y(n1992) );
  OAI21X1 U3548 ( .A(n3977), .B(n7463), .C(n6243), .Y(n1991) );
  OAI21X1 U3550 ( .A(n3977), .B(n7464), .C(n6423), .Y(n1990) );
  OAI21X1 U3552 ( .A(n3977), .B(n7465), .C(n5961), .Y(n1989) );
  OAI21X1 U3554 ( .A(n3977), .B(n7466), .C(n6185), .Y(n1988) );
  OAI21X1 U3556 ( .A(n3977), .B(n7467), .C(n6632), .Y(n1987) );
  OAI21X1 U3558 ( .A(n3977), .B(n7468), .C(n6016), .Y(n1986) );
  OAI21X1 U3560 ( .A(n3977), .B(n7469), .C(n6560), .Y(n1985) );
  OAI21X1 U3562 ( .A(n3977), .B(n7470), .C(n6775), .Y(n1984) );
  OAI21X1 U3564 ( .A(n3977), .B(n7471), .C(n6704), .Y(n1983) );
  OAI21X1 U3566 ( .A(n3977), .B(n7472), .C(n6361), .Y(n1982) );
  OAI21X1 U3568 ( .A(n3977), .B(n7473), .C(n6299), .Y(n1981) );
  OAI21X1 U3570 ( .A(n3977), .B(n7474), .C(n6488), .Y(n1980) );
  OAI21X1 U3572 ( .A(n3977), .B(n7475), .C(n6424), .Y(n1979) );
  OAI21X1 U3574 ( .A(n3977), .B(n7476), .C(n5907), .Y(n1978) );
  OAI21X1 U3576 ( .A(n3977), .B(n7477), .C(n5852), .Y(n1977) );
  OAI21X1 U3578 ( .A(n3977), .B(n7478), .C(n6017), .Y(n1976) );
  OAI21X1 U3580 ( .A(n3977), .B(n7479), .C(n5962), .Y(n1975) );
  OAI21X1 U3582 ( .A(n3977), .B(n7480), .C(n6633), .Y(n1974) );
  OAI21X1 U3584 ( .A(n3977), .B(n7481), .C(n6561), .Y(n1973) );
  OAI21X1 U3586 ( .A(n3977), .B(n7482), .C(n6776), .Y(n1972) );
  OAI21X1 U3588 ( .A(n3977), .B(n7483), .C(n6705), .Y(n1971) );
  OAI21X1 U3590 ( .A(n3977), .B(n7484), .C(n6362), .Y(n1970) );
  OAI21X1 U3592 ( .A(n3977), .B(n7485), .C(n6300), .Y(n1969) );
  OAI21X1 U3594 ( .A(n3977), .B(n7486), .C(n6489), .Y(n1968) );
  OAI21X1 U3596 ( .A(n3977), .B(n7487), .C(n6425), .Y(n1967) );
  OAI21X1 U3598 ( .A(n6454), .B(n6737), .C(n6843), .Y(n3977) );
  OAI21X1 U3599 ( .A(n4011), .B(n7488), .C(n6186), .Y(n1966) );
  OAI21X1 U3601 ( .A(n4011), .B(n7489), .C(n5853), .Y(n1965) );
  OAI21X1 U3603 ( .A(n4011), .B(n7490), .C(n5908), .Y(n1964) );
  OAI21X1 U3605 ( .A(n4011), .B(n7491), .C(n4700), .Y(n1963) );
  OAI21X1 U3607 ( .A(n4011), .B(n7492), .C(n4699), .Y(n1962) );
  OAI21X1 U3609 ( .A(n4011), .B(n7493), .C(n4698), .Y(n1961) );
  OAI21X1 U3611 ( .A(n4011), .B(n7494), .C(n6073), .Y(n1960) );
  OAI21X1 U3613 ( .A(n4011), .B(n7495), .C(n6130), .Y(n1959) );
  OAI21X1 U3615 ( .A(n4011), .B(n7496), .C(n6187), .Y(n1958) );
  OAI21X1 U3617 ( .A(n4011), .B(n7497), .C(n6490), .Y(n1957) );
  OAI21X1 U3619 ( .A(n4011), .B(n7498), .C(n6018), .Y(n1956) );
  OAI21X1 U3621 ( .A(n4011), .B(n7499), .C(n6244), .Y(n1955) );
  OAI21X1 U3623 ( .A(n4011), .B(n7500), .C(n6562), .Y(n1954) );
  OAI21X1 U3625 ( .A(n4011), .B(n7501), .C(n5963), .Y(n1953) );
  OAI21X1 U3627 ( .A(n4011), .B(n7502), .C(n6634), .Y(n1952) );
  OAI21X1 U3629 ( .A(n4011), .B(n7503), .C(n6706), .Y(n1951) );
  OAI21X1 U3631 ( .A(n4011), .B(n7504), .C(n6777), .Y(n1950) );
  OAI21X1 U3633 ( .A(n4011), .B(n7505), .C(n6301), .Y(n1949) );
  OAI21X1 U3635 ( .A(n4011), .B(n7506), .C(n6363), .Y(n1948) );
  OAI21X1 U3637 ( .A(n4011), .B(n7507), .C(n6426), .Y(n1947) );
  OAI21X1 U3639 ( .A(n4011), .B(n7508), .C(n6491), .Y(n1946) );
  OAI21X1 U3641 ( .A(n4011), .B(n7509), .C(n5854), .Y(n1945) );
  OAI21X1 U3643 ( .A(n4011), .B(n7510), .C(n5909), .Y(n1944) );
  OAI21X1 U3645 ( .A(n4011), .B(n7511), .C(n5964), .Y(n1943) );
  OAI21X1 U3647 ( .A(n4011), .B(n7512), .C(n6019), .Y(n1942) );
  OAI21X1 U3649 ( .A(n4011), .B(n7513), .C(n6563), .Y(n1941) );
  OAI21X1 U3651 ( .A(n4011), .B(n7514), .C(n6635), .Y(n1940) );
  OAI21X1 U3653 ( .A(n4011), .B(n7515), .C(n6707), .Y(n1939) );
  OAI21X1 U3655 ( .A(n4011), .B(n7516), .C(n6778), .Y(n1938) );
  OAI21X1 U3657 ( .A(n4011), .B(n7517), .C(n6302), .Y(n1937) );
  OAI21X1 U3659 ( .A(n4011), .B(n7518), .C(n6364), .Y(n1936) );
  OAI21X1 U3661 ( .A(n4011), .B(n7519), .C(n6427), .Y(n1935) );
  OAI21X1 U3663 ( .A(n4011), .B(n7520), .C(n6492), .Y(n1934) );
  OAI21X1 U3665 ( .A(n6665), .B(n6737), .C(n6843), .Y(n4011) );
  OAI21X1 U3666 ( .A(n4045), .B(n7521), .C(n5910), .Y(n1933) );
  OAI21X1 U3668 ( .A(n4045), .B(n7522), .C(n6245), .Y(n1932) );
  OAI21X1 U3670 ( .A(n4045), .B(n7523), .C(n6188), .Y(n1931) );
  OAI21X1 U3672 ( .A(n4045), .B(n7524), .C(n4697), .Y(n1930) );
  OAI21X1 U3674 ( .A(n4045), .B(n7525), .C(n4696), .Y(n1929) );
  OAI21X1 U3676 ( .A(n4045), .B(n7526), .C(n4695), .Y(n1928) );
  OAI21X1 U3678 ( .A(n4045), .B(n7527), .C(n6020), .Y(n1927) );
  OAI21X1 U3680 ( .A(n4045), .B(n7528), .C(n5965), .Y(n1926) );
  OAI21X1 U3682 ( .A(n4045), .B(n7529), .C(n5911), .Y(n1925) );
  OAI21X1 U3684 ( .A(n4045), .B(n7530), .C(n6564), .Y(n1924) );
  OAI21X1 U3686 ( .A(n4045), .B(n7531), .C(n6074), .Y(n1923) );
  OAI21X1 U3688 ( .A(n4045), .B(n7532), .C(n5855), .Y(n1922) );
  OAI21X1 U3690 ( .A(n4045), .B(n7533), .C(n6493), .Y(n1921) );
  OAI21X1 U3692 ( .A(n4045), .B(n7534), .C(n6131), .Y(n1920) );
  OAI21X1 U3694 ( .A(n4045), .B(n7535), .C(n6428), .Y(n1919) );
  OAI21X1 U3696 ( .A(n4045), .B(n7536), .C(n6365), .Y(n1918) );
  OAI21X1 U3698 ( .A(n4045), .B(n7537), .C(n6303), .Y(n1917) );
  OAI21X1 U3700 ( .A(n4045), .B(n7538), .C(n6779), .Y(n1916) );
  OAI21X1 U3702 ( .A(n4045), .B(n7539), .C(n6708), .Y(n1915) );
  OAI21X1 U3704 ( .A(n4045), .B(n7540), .C(n6636), .Y(n1914) );
  OAI21X1 U3706 ( .A(n4045), .B(n7541), .C(n6565), .Y(n1913) );
  OAI21X1 U3708 ( .A(n4045), .B(n7542), .C(n6246), .Y(n1912) );
  OAI21X1 U3710 ( .A(n4045), .B(n7543), .C(n6189), .Y(n1911) );
  OAI21X1 U3712 ( .A(n4045), .B(n7544), .C(n6132), .Y(n1910) );
  OAI21X1 U3714 ( .A(n4045), .B(n7545), .C(n6075), .Y(n1909) );
  OAI21X1 U3716 ( .A(n4045), .B(n7546), .C(n6494), .Y(n1908) );
  OAI21X1 U3718 ( .A(n4045), .B(n7547), .C(n6429), .Y(n1907) );
  OAI21X1 U3720 ( .A(n4045), .B(n7548), .C(n6366), .Y(n1906) );
  OAI21X1 U3722 ( .A(n4045), .B(n7549), .C(n6304), .Y(n1905) );
  OAI21X1 U3724 ( .A(n4045), .B(n7550), .C(n6780), .Y(n1904) );
  OAI21X1 U3726 ( .A(n4045), .B(n7551), .C(n6709), .Y(n1903) );
  OAI21X1 U3728 ( .A(n4045), .B(n7552), .C(n6637), .Y(n1902) );
  OAI21X1 U3730 ( .A(n4045), .B(n7553), .C(n6566), .Y(n1901) );
  OAI21X1 U3732 ( .A(n6666), .B(n6737), .C(n6843), .Y(n4045) );
  OAI21X1 U3733 ( .A(n4079), .B(n7554), .C(n5856), .Y(n1900) );
  OAI21X1 U3735 ( .A(n4079), .B(n7555), .C(n6190), .Y(n1899) );
  OAI21X1 U3737 ( .A(n4079), .B(n7556), .C(n6247), .Y(n1898) );
  OAI21X1 U3739 ( .A(n4079), .B(n7557), .C(n4694), .Y(n1897) );
  OAI21X1 U3741 ( .A(n4079), .B(n7558), .C(n4693), .Y(n1896) );
  OAI21X1 U3743 ( .A(n4079), .B(n7559), .C(n4692), .Y(n1895) );
  OAI21X1 U3745 ( .A(n4079), .B(n7560), .C(n5966), .Y(n1894) );
  OAI21X1 U3747 ( .A(n4079), .B(n7561), .C(n6021), .Y(n1893) );
  OAI21X1 U3749 ( .A(n4079), .B(n7562), .C(n5857), .Y(n1892) );
  OAI21X1 U3751 ( .A(n4079), .B(n7563), .C(n6638), .Y(n1891) );
  OAI21X1 U3753 ( .A(n4079), .B(n7564), .C(n6133), .Y(n1890) );
  OAI21X1 U3755 ( .A(n4079), .B(n7565), .C(n5912), .Y(n1889) );
  OAI21X1 U3757 ( .A(n4079), .B(n7566), .C(n6430), .Y(n1888) );
  OAI21X1 U3759 ( .A(n4079), .B(n7567), .C(n6076), .Y(n1887) );
  OAI21X1 U3761 ( .A(n4079), .B(n7568), .C(n6495), .Y(n1886) );
  OAI21X1 U3763 ( .A(n4079), .B(n7569), .C(n6305), .Y(n1885) );
  OAI21X1 U3765 ( .A(n4079), .B(n7570), .C(n6367), .Y(n1884) );
  OAI21X1 U3767 ( .A(n4079), .B(n7571), .C(n6710), .Y(n1883) );
  OAI21X1 U3769 ( .A(n4079), .B(n7572), .C(n6781), .Y(n1882) );
  OAI21X1 U3771 ( .A(n4079), .B(n7573), .C(n6567), .Y(n1881) );
  OAI21X1 U3773 ( .A(n4079), .B(n7574), .C(n6639), .Y(n1880) );
  OAI21X1 U3775 ( .A(n4079), .B(n7575), .C(n6191), .Y(n1879) );
  OAI21X1 U3777 ( .A(n4079), .B(n7576), .C(n6248), .Y(n1878) );
  OAI21X1 U3779 ( .A(n4079), .B(n7577), .C(n6077), .Y(n1877) );
  OAI21X1 U3781 ( .A(n4079), .B(n7578), .C(n6134), .Y(n1876) );
  OAI21X1 U3783 ( .A(n4079), .B(n7579), .C(n6431), .Y(n1875) );
  OAI21X1 U3785 ( .A(n4079), .B(n7580), .C(n6496), .Y(n1874) );
  OAI21X1 U3787 ( .A(n4079), .B(n7581), .C(n6306), .Y(n1873) );
  OAI21X1 U3789 ( .A(n4079), .B(n7582), .C(n6368), .Y(n1872) );
  OAI21X1 U3791 ( .A(n4079), .B(n7583), .C(n6711), .Y(n1871) );
  OAI21X1 U3793 ( .A(n4079), .B(n7584), .C(n6782), .Y(n1870) );
  OAI21X1 U3795 ( .A(n4079), .B(n7585), .C(n6568), .Y(n1869) );
  OAI21X1 U3797 ( .A(n4079), .B(n7586), .C(n6640), .Y(n1868) );
  OAI21X1 U3799 ( .A(n6455), .B(n6737), .C(n6843), .Y(n4079) );
  OAI21X1 U3800 ( .A(n4113), .B(n7587), .C(n6022), .Y(n1867) );
  OAI21X1 U3802 ( .A(n4113), .B(n7588), .C(n6135), .Y(n1866) );
  OAI21X1 U3804 ( .A(n4113), .B(n7589), .C(n6078), .Y(n1865) );
  OAI21X1 U3806 ( .A(n4113), .B(n7590), .C(n4691), .Y(n1864) );
  OAI21X1 U3808 ( .A(n4113), .B(n7591), .C(n4690), .Y(n1863) );
  OAI21X1 U3810 ( .A(n4113), .B(n7592), .C(n4689), .Y(n1862) );
  OAI21X1 U3812 ( .A(n4113), .B(n7593), .C(n5913), .Y(n1861) );
  OAI21X1 U3814 ( .A(n4113), .B(n7594), .C(n5858), .Y(n1860) );
  OAI21X1 U3816 ( .A(n4113), .B(n7595), .C(n6023), .Y(n1859) );
  OAI21X1 U3818 ( .A(n4113), .B(n7596), .C(n6712), .Y(n1858) );
  OAI21X1 U3820 ( .A(n4113), .B(n7597), .C(n6192), .Y(n1857) );
  OAI21X1 U3822 ( .A(n4113), .B(n7598), .C(n5967), .Y(n1856) );
  OAI21X1 U3824 ( .A(n4113), .B(n7599), .C(n6369), .Y(n1855) );
  OAI21X1 U3826 ( .A(n4113), .B(n7600), .C(n6249), .Y(n1854) );
  OAI21X1 U3828 ( .A(n4113), .B(n7601), .C(n6307), .Y(n1853) );
  OAI21X1 U3830 ( .A(n4113), .B(n7602), .C(n6497), .Y(n1852) );
  OAI21X1 U3832 ( .A(n4113), .B(n7603), .C(n6432), .Y(n1851) );
  OAI21X1 U3834 ( .A(n4113), .B(n7604), .C(n6641), .Y(n1850) );
  OAI21X1 U3836 ( .A(n4113), .B(n7605), .C(n6569), .Y(n1849) );
  OAI21X1 U3838 ( .A(n4113), .B(n7606), .C(n6783), .Y(n1848) );
  OAI21X1 U3840 ( .A(n4113), .B(n7607), .C(n6713), .Y(n1847) );
  OAI21X1 U3842 ( .A(n4113), .B(n7608), .C(n6136), .Y(n1846) );
  OAI21X1 U3844 ( .A(n4113), .B(n7609), .C(n6079), .Y(n1845) );
  OAI21X1 U3846 ( .A(n4113), .B(n7610), .C(n6250), .Y(n1844) );
  OAI21X1 U3848 ( .A(n4113), .B(n7611), .C(n6193), .Y(n1843) );
  OAI21X1 U3850 ( .A(n4113), .B(n7612), .C(n6370), .Y(n1842) );
  OAI21X1 U3852 ( .A(n4113), .B(n7613), .C(n6308), .Y(n1841) );
  OAI21X1 U3854 ( .A(n4113), .B(n7614), .C(n6498), .Y(n1840) );
  OAI21X1 U3856 ( .A(n4113), .B(n7615), .C(n6433), .Y(n1839) );
  OAI21X1 U3858 ( .A(n4113), .B(n7616), .C(n6642), .Y(n1838) );
  OAI21X1 U3860 ( .A(n4113), .B(n7617), .C(n6570), .Y(n1837) );
  OAI21X1 U3862 ( .A(n4113), .B(n7618), .C(n6784), .Y(n1836) );
  OAI21X1 U3864 ( .A(n4113), .B(n7619), .C(n6714), .Y(n1835) );
  OAI21X1 U3866 ( .A(n6522), .B(n6737), .C(n6843), .Y(n4113) );
  OAI21X1 U3867 ( .A(n4147), .B(n7620), .C(n5968), .Y(n1834) );
  OAI21X1 U3869 ( .A(n4147), .B(n7621), .C(n6080), .Y(n1833) );
  OAI21X1 U3871 ( .A(n4147), .B(n7622), .C(n6137), .Y(n1832) );
  OAI21X1 U3873 ( .A(n4147), .B(n7623), .C(n4688), .Y(n1831) );
  OAI21X1 U3875 ( .A(n4147), .B(n7624), .C(n4687), .Y(n1830) );
  OAI21X1 U3877 ( .A(n4147), .B(n7625), .C(n4686), .Y(n1829) );
  OAI21X1 U3879 ( .A(n4147), .B(n7626), .C(n5859), .Y(n1828) );
  OAI21X1 U3881 ( .A(n4147), .B(n7627), .C(n5914), .Y(n1827) );
  OAI21X1 U3883 ( .A(n4147), .B(n7628), .C(n5969), .Y(n1826) );
  OAI21X1 U3885 ( .A(n4147), .B(n7629), .C(n6785), .Y(n1825) );
  OAI21X1 U3887 ( .A(n4147), .B(n7630), .C(n6251), .Y(n1824) );
  OAI21X1 U3889 ( .A(n4147), .B(n7631), .C(n6024), .Y(n1823) );
  OAI21X1 U3891 ( .A(n4147), .B(n7632), .C(n6309), .Y(n1822) );
  OAI21X1 U3893 ( .A(n4147), .B(n7633), .C(n6194), .Y(n1821) );
  OAI21X1 U3895 ( .A(n4147), .B(n7634), .C(n6371), .Y(n1820) );
  OAI21X1 U3897 ( .A(n4147), .B(n7635), .C(n6434), .Y(n1819) );
  OAI21X1 U3899 ( .A(n4147), .B(n7636), .C(n6499), .Y(n1818) );
  OAI21X1 U3901 ( .A(n4147), .B(n7637), .C(n6571), .Y(n1817) );
  OAI21X1 U3903 ( .A(n4147), .B(n7638), .C(n6643), .Y(n1816) );
  OAI21X1 U3905 ( .A(n4147), .B(n7639), .C(n6715), .Y(n1815) );
  OAI21X1 U3907 ( .A(n4147), .B(n7640), .C(n6786), .Y(n1814) );
  OAI21X1 U3909 ( .A(n4147), .B(n7641), .C(n6081), .Y(n1813) );
  OAI21X1 U3911 ( .A(n4147), .B(n7642), .C(n6138), .Y(n1812) );
  OAI21X1 U3913 ( .A(n4147), .B(n7643), .C(n6195), .Y(n1811) );
  OAI21X1 U3915 ( .A(n4147), .B(n7644), .C(n6252), .Y(n1810) );
  OAI21X1 U3917 ( .A(n4147), .B(n7645), .C(n6310), .Y(n1809) );
  OAI21X1 U3919 ( .A(n4147), .B(n7646), .C(n6372), .Y(n1808) );
  OAI21X1 U3921 ( .A(n4147), .B(n7647), .C(n6435), .Y(n1807) );
  OAI21X1 U3923 ( .A(n4147), .B(n7648), .C(n6500), .Y(n1806) );
  OAI21X1 U3925 ( .A(n4147), .B(n7649), .C(n6572), .Y(n1805) );
  OAI21X1 U3927 ( .A(n4147), .B(n7650), .C(n6644), .Y(n1804) );
  OAI21X1 U3929 ( .A(n4147), .B(n7651), .C(n6716), .Y(n1803) );
  OAI21X1 U3931 ( .A(n4147), .B(n7652), .C(n6787), .Y(n1802) );
  OAI21X1 U3933 ( .A(n6593), .B(n6737), .C(n6843), .Y(n4147) );
  NAND3X1 U3934 ( .A(wr_ptr[3]), .B(n6857), .C(put), .Y(n3942) );
  OAI21X1 U3935 ( .A(n4181), .B(n7653), .C(n6139), .Y(n1801) );
  OAI21X1 U3937 ( .A(n4181), .B(n7654), .C(n6025), .Y(n1800) );
  OAI21X1 U3939 ( .A(n4181), .B(n7655), .C(n5970), .Y(n1799) );
  OAI21X1 U3941 ( .A(n4181), .B(n7656), .C(n4685), .Y(n1798) );
  OAI21X1 U3943 ( .A(n4181), .B(n7657), .C(n4684), .Y(n1797) );
  OAI21X1 U3945 ( .A(n4181), .B(n7658), .C(n4683), .Y(n1796) );
  OAI21X1 U3947 ( .A(n4181), .B(n7659), .C(n6253), .Y(n1795) );
  OAI21X1 U3949 ( .A(n4181), .B(n7660), .C(n6196), .Y(n1794) );
  OAI21X1 U3951 ( .A(n4181), .B(n7661), .C(n6140), .Y(n1793) );
  OAI21X1 U3953 ( .A(n4181), .B(n7662), .C(n6311), .Y(n1792) );
  OAI21X1 U3955 ( .A(n4181), .B(n7663), .C(n5860), .Y(n1791) );
  OAI21X1 U3957 ( .A(n4181), .B(n7664), .C(n6082), .Y(n1790) );
  OAI21X1 U3959 ( .A(n4181), .B(n7665), .C(n6788), .Y(n1789) );
  OAI21X1 U3961 ( .A(n4181), .B(n7666), .C(n5915), .Y(n1788) );
  OAI21X1 U3963 ( .A(n4181), .B(n7667), .C(n6717), .Y(n1787) );
  OAI21X1 U3965 ( .A(n4181), .B(n7668), .C(n6645), .Y(n1786) );
  OAI21X1 U3967 ( .A(n4181), .B(n7669), .C(n6573), .Y(n1785) );
  OAI21X1 U3969 ( .A(n4181), .B(n7670), .C(n6501), .Y(n1784) );
  OAI21X1 U3971 ( .A(n4181), .B(n7671), .C(n6436), .Y(n1783) );
  OAI21X1 U3973 ( .A(n4181), .B(n7672), .C(n6373), .Y(n1782) );
  OAI21X1 U3975 ( .A(n4181), .B(n7673), .C(n6312), .Y(n1781) );
  OAI21X1 U3977 ( .A(n4181), .B(n7674), .C(n6026), .Y(n1780) );
  OAI21X1 U3979 ( .A(n4181), .B(n7675), .C(n5971), .Y(n1779) );
  OAI21X1 U3981 ( .A(n4181), .B(n7676), .C(n5916), .Y(n1778) );
  OAI21X1 U3983 ( .A(n4181), .B(n7677), .C(n5861), .Y(n1777) );
  OAI21X1 U3985 ( .A(n4181), .B(n7678), .C(n6789), .Y(n1776) );
  OAI21X1 U3987 ( .A(n4181), .B(n7679), .C(n6718), .Y(n1775) );
  OAI21X1 U3989 ( .A(n4181), .B(n7680), .C(n6646), .Y(n1774) );
  OAI21X1 U3991 ( .A(n4181), .B(n7681), .C(n6574), .Y(n1773) );
  OAI21X1 U3993 ( .A(n4181), .B(n7682), .C(n6502), .Y(n1772) );
  OAI21X1 U3995 ( .A(n4181), .B(n7683), .C(n6437), .Y(n1771) );
  OAI21X1 U3997 ( .A(n4181), .B(n7684), .C(n6374), .Y(n1770) );
  OAI21X1 U3999 ( .A(n4181), .B(n7685), .C(n6313), .Y(n1769) );
  OAI21X1 U4001 ( .A(n6594), .B(n6809), .C(n6843), .Y(n4181) );
  NAND3X1 U4002 ( .A(wr_ptr[2]), .B(wr_ptr[0]), .C(wr_ptr[1]), .Y(n3322) );
  OAI21X1 U4003 ( .A(n4216), .B(n7686), .C(n6083), .Y(n1768) );
  OAI21X1 U4005 ( .A(n4216), .B(n7687), .C(n5972), .Y(n1767) );
  OAI21X1 U4007 ( .A(n4216), .B(n7688), .C(n6027), .Y(n1766) );
  OAI21X1 U4009 ( .A(n4216), .B(n7689), .C(n4682), .Y(n1765) );
  OAI21X1 U4011 ( .A(n4216), .B(n7690), .C(n4681), .Y(n1764) );
  OAI21X1 U4013 ( .A(n4216), .B(n7691), .C(n4680), .Y(n1763) );
  OAI21X1 U4015 ( .A(n4216), .B(n7692), .C(n6197), .Y(n1762) );
  OAI21X1 U4017 ( .A(n4216), .B(n7693), .C(n6254), .Y(n1761) );
  OAI21X1 U4019 ( .A(n4216), .B(n7694), .C(n6084), .Y(n1760) );
  OAI21X1 U4021 ( .A(n4216), .B(n7695), .C(n6375), .Y(n1759) );
  OAI21X1 U4023 ( .A(n4216), .B(n7696), .C(n5917), .Y(n1758) );
  OAI21X1 U4025 ( .A(n4216), .B(n7697), .C(n6141), .Y(n1757) );
  OAI21X1 U4027 ( .A(n4216), .B(n7698), .C(n6719), .Y(n1756) );
  OAI21X1 U4029 ( .A(n4216), .B(n7699), .C(n5862), .Y(n1755) );
  OAI21X1 U4031 ( .A(n4216), .B(n7700), .C(n6790), .Y(n1754) );
  OAI21X1 U4033 ( .A(n4216), .B(n7701), .C(n6575), .Y(n1753) );
  OAI21X1 U4035 ( .A(n4216), .B(n7702), .C(n6647), .Y(n1752) );
  OAI21X1 U4037 ( .A(n4216), .B(n7703), .C(n6438), .Y(n1751) );
  OAI21X1 U4039 ( .A(n4216), .B(n7704), .C(n6503), .Y(n1750) );
  OAI21X1 U4041 ( .A(n4216), .B(n7705), .C(n6314), .Y(n1749) );
  OAI21X1 U4043 ( .A(n4216), .B(n7706), .C(n6376), .Y(n1748) );
  OAI21X1 U4045 ( .A(n4216), .B(n7707), .C(n5973), .Y(n1747) );
  OAI21X1 U4047 ( .A(n4216), .B(n7708), .C(n6028), .Y(n1746) );
  OAI21X1 U4049 ( .A(n4216), .B(n7709), .C(n5863), .Y(n1745) );
  OAI21X1 U4051 ( .A(n4216), .B(n7710), .C(n5918), .Y(n1744) );
  OAI21X1 U4053 ( .A(n4216), .B(n7711), .C(n6720), .Y(n1743) );
  OAI21X1 U4055 ( .A(n4216), .B(n7712), .C(n6791), .Y(n1742) );
  OAI21X1 U4057 ( .A(n4216), .B(n7713), .C(n6576), .Y(n1741) );
  OAI21X1 U4059 ( .A(n4216), .B(n7714), .C(n6648), .Y(n1740) );
  OAI21X1 U4061 ( .A(n4216), .B(n7715), .C(n6439), .Y(n1739) );
  OAI21X1 U4063 ( .A(n4216), .B(n7716), .C(n6504), .Y(n1738) );
  OAI21X1 U4065 ( .A(n4216), .B(n7717), .C(n6315), .Y(n1737) );
  OAI21X1 U4067 ( .A(n4216), .B(n7718), .C(n6377), .Y(n1736) );
  OAI21X1 U4069 ( .A(n6521), .B(n6809), .C(n6843), .Y(n4216) );
  NAND3X1 U4070 ( .A(wr_ptr[2]), .B(n6849), .C(wr_ptr[1]), .Y(n3425) );
  OAI21X1 U4071 ( .A(n4250), .B(n7719), .C(n6255), .Y(n1735) );
  OAI21X1 U4073 ( .A(n4250), .B(n7720), .C(n5919), .Y(n1734) );
  OAI21X1 U4075 ( .A(n4250), .B(n7721), .C(n5864), .Y(n1733) );
  OAI21X1 U4077 ( .A(n4250), .B(n7722), .C(n4679), .Y(n1732) );
  OAI21X1 U4079 ( .A(n4250), .B(n7723), .C(n4678), .Y(n1731) );
  OAI21X1 U4081 ( .A(n4250), .B(n7724), .C(n4677), .Y(n1730) );
  OAI21X1 U4083 ( .A(n4250), .B(n7725), .C(n6142), .Y(n1729) );
  OAI21X1 U4085 ( .A(n4250), .B(n7726), .C(n6085), .Y(n1728) );
  OAI21X1 U4087 ( .A(n4250), .B(n7727), .C(n6256), .Y(n1727) );
  OAI21X1 U4089 ( .A(n4250), .B(n7728), .C(n6440), .Y(n1726) );
  OAI21X1 U4091 ( .A(n4250), .B(n7729), .C(n5974), .Y(n1725) );
  OAI21X1 U4093 ( .A(n4250), .B(n7730), .C(n6198), .Y(n1724) );
  OAI21X1 U4095 ( .A(n4250), .B(n7731), .C(n6649), .Y(n1723) );
  OAI21X1 U4097 ( .A(n4250), .B(n7732), .C(n6029), .Y(n1722) );
  OAI21X1 U4099 ( .A(n4250), .B(n7733), .C(n6577), .Y(n1721) );
  OAI21X1 U4101 ( .A(n4250), .B(n7734), .C(n6792), .Y(n1720) );
  OAI21X1 U4103 ( .A(n4250), .B(n7735), .C(n6721), .Y(n1719) );
  OAI21X1 U4105 ( .A(n4250), .B(n7736), .C(n6378), .Y(n1718) );
  OAI21X1 U4107 ( .A(n4250), .B(n7737), .C(n6316), .Y(n1717) );
  OAI21X1 U4109 ( .A(n4250), .B(n7738), .C(n6505), .Y(n1716) );
  OAI21X1 U4111 ( .A(n4250), .B(n7739), .C(n6441), .Y(n1715) );
  OAI21X1 U4113 ( .A(n4250), .B(n7740), .C(n5920), .Y(n1714) );
  OAI21X1 U4115 ( .A(n4250), .B(n7741), .C(n5865), .Y(n1713) );
  OAI21X1 U4117 ( .A(n4250), .B(n7742), .C(n6030), .Y(n1712) );
  OAI21X1 U4119 ( .A(n4250), .B(n7743), .C(n5975), .Y(n1711) );
  OAI21X1 U4121 ( .A(n4250), .B(n7744), .C(n6650), .Y(n1710) );
  OAI21X1 U4123 ( .A(n4250), .B(n7745), .C(n6578), .Y(n1709) );
  OAI21X1 U4125 ( .A(n4250), .B(n7746), .C(n6793), .Y(n1708) );
  OAI21X1 U4127 ( .A(n4250), .B(n7747), .C(n6722), .Y(n1707) );
  OAI21X1 U4129 ( .A(n4250), .B(n7748), .C(n6379), .Y(n1706) );
  OAI21X1 U4131 ( .A(n4250), .B(n7749), .C(n6317), .Y(n1705) );
  OAI21X1 U4133 ( .A(n4250), .B(n7750), .C(n6506), .Y(n1704) );
  OAI21X1 U4135 ( .A(n4250), .B(n7751), .C(n6442), .Y(n1703) );
  OAI21X1 U4137 ( .A(n6454), .B(n6809), .C(n6843), .Y(n4250) );
  NAND3X1 U4138 ( .A(wr_ptr[0]), .B(n6858), .C(wr_ptr[2]), .Y(n3460) );
  OAI21X1 U4139 ( .A(n4284), .B(n7752), .C(n6199), .Y(n1702) );
  OAI21X1 U4141 ( .A(n4284), .B(n7753), .C(n5866), .Y(n1701) );
  OAI21X1 U4143 ( .A(n4284), .B(n7754), .C(n5921), .Y(n1700) );
  OAI21X1 U4145 ( .A(n4284), .B(n7755), .C(n4676), .Y(n1699) );
  OAI21X1 U4147 ( .A(n4284), .B(n7756), .C(n4675), .Y(n1698) );
  OAI21X1 U4149 ( .A(n4284), .B(n7757), .C(n4674), .Y(n1697) );
  OAI21X1 U4151 ( .A(n4284), .B(n7758), .C(n6086), .Y(n1696) );
  OAI21X1 U4153 ( .A(n4284), .B(n7759), .C(n6143), .Y(n1695) );
  OAI21X1 U4155 ( .A(n4284), .B(n7760), .C(n6200), .Y(n1694) );
  OAI21X1 U4157 ( .A(n4284), .B(n7761), .C(n6507), .Y(n1693) );
  OAI21X1 U4159 ( .A(n4284), .B(n7762), .C(n6031), .Y(n1692) );
  OAI21X1 U4161 ( .A(n4284), .B(n7763), .C(n6257), .Y(n1691) );
  OAI21X1 U4163 ( .A(n4284), .B(n7764), .C(n6579), .Y(n1690) );
  OAI21X1 U4165 ( .A(n4284), .B(n7765), .C(n5976), .Y(n1689) );
  OAI21X1 U4167 ( .A(n4284), .B(n7766), .C(n6651), .Y(n1688) );
  OAI21X1 U4169 ( .A(n4284), .B(n7767), .C(n6723), .Y(n1687) );
  OAI21X1 U4171 ( .A(n4284), .B(n7768), .C(n6794), .Y(n1686) );
  OAI21X1 U4173 ( .A(n4284), .B(n7769), .C(n6318), .Y(n1685) );
  OAI21X1 U4175 ( .A(n4284), .B(n7770), .C(n6380), .Y(n1684) );
  OAI21X1 U4177 ( .A(n4284), .B(n7771), .C(n6443), .Y(n1683) );
  OAI21X1 U4179 ( .A(n4284), .B(n7772), .C(n6508), .Y(n1682) );
  OAI21X1 U4181 ( .A(n4284), .B(n7773), .C(n5867), .Y(n1681) );
  OAI21X1 U4183 ( .A(n4284), .B(n7774), .C(n5922), .Y(n1680) );
  OAI21X1 U4185 ( .A(n4284), .B(n7775), .C(n5977), .Y(n1679) );
  OAI21X1 U4187 ( .A(n4284), .B(n7776), .C(n6032), .Y(n1678) );
  OAI21X1 U4189 ( .A(n4284), .B(n7777), .C(n6580), .Y(n1677) );
  OAI21X1 U4191 ( .A(n4284), .B(n7778), .C(n6652), .Y(n1676) );
  OAI21X1 U4193 ( .A(n4284), .B(n7779), .C(n6724), .Y(n1675) );
  OAI21X1 U4195 ( .A(n4284), .B(n7780), .C(n6795), .Y(n1674) );
  OAI21X1 U4197 ( .A(n4284), .B(n7781), .C(n6319), .Y(n1673) );
  OAI21X1 U4199 ( .A(n4284), .B(n7782), .C(n6381), .Y(n1672) );
  OAI21X1 U4201 ( .A(n4284), .B(n7783), .C(n6444), .Y(n1671) );
  OAI21X1 U4203 ( .A(n4284), .B(n7784), .C(n6509), .Y(n1670) );
  OAI21X1 U4205 ( .A(n6665), .B(n6809), .C(n6843), .Y(n4284) );
  NAND3X1 U4206 ( .A(n6849), .B(n6858), .C(wr_ptr[2]), .Y(n3495) );
  OAI21X1 U4207 ( .A(n4318), .B(n7785), .C(n5923), .Y(n1669) );
  OAI21X1 U4209 ( .A(n4318), .B(n7786), .C(n6258), .Y(n1668) );
  OAI21X1 U4211 ( .A(n4318), .B(n7787), .C(n6201), .Y(n1667) );
  OAI21X1 U4213 ( .A(n4318), .B(n7788), .C(n4673), .Y(n1666) );
  OAI21X1 U4215 ( .A(n4318), .B(n7789), .C(n4672), .Y(n1665) );
  OAI21X1 U4217 ( .A(n4318), .B(n7790), .C(n4671), .Y(n1664) );
  OAI21X1 U4219 ( .A(n4318), .B(n7791), .C(n6033), .Y(n1663) );
  OAI21X1 U4221 ( .A(n4318), .B(n7792), .C(n5978), .Y(n1662) );
  OAI21X1 U4223 ( .A(n4318), .B(n7793), .C(n5924), .Y(n1661) );
  OAI21X1 U4225 ( .A(n4318), .B(n7794), .C(n6581), .Y(n1660) );
  OAI21X1 U4227 ( .A(n4318), .B(n7795), .C(n6087), .Y(n1659) );
  OAI21X1 U4229 ( .A(n4318), .B(n7796), .C(n5868), .Y(n1658) );
  OAI21X1 U4231 ( .A(n4318), .B(n7797), .C(n6510), .Y(n1657) );
  OAI21X1 U4233 ( .A(n4318), .B(n7798), .C(n6144), .Y(n1656) );
  OAI21X1 U4235 ( .A(n4318), .B(n7799), .C(n6445), .Y(n1655) );
  OAI21X1 U4237 ( .A(n4318), .B(n7800), .C(n6382), .Y(n1654) );
  OAI21X1 U4239 ( .A(n4318), .B(n7801), .C(n6320), .Y(n1653) );
  OAI21X1 U4241 ( .A(n4318), .B(n7802), .C(n6796), .Y(n1652) );
  OAI21X1 U4243 ( .A(n4318), .B(n7803), .C(n6725), .Y(n1651) );
  OAI21X1 U4245 ( .A(n4318), .B(n7804), .C(n6653), .Y(n1650) );
  OAI21X1 U4247 ( .A(n4318), .B(n7805), .C(n6582), .Y(n1649) );
  OAI21X1 U4249 ( .A(n4318), .B(n7806), .C(n6259), .Y(n1648) );
  OAI21X1 U4251 ( .A(n4318), .B(n7807), .C(n6202), .Y(n1647) );
  OAI21X1 U4253 ( .A(n4318), .B(n7808), .C(n6145), .Y(n1646) );
  OAI21X1 U4255 ( .A(n4318), .B(n7809), .C(n6088), .Y(n1645) );
  OAI21X1 U4257 ( .A(n4318), .B(n7810), .C(n6511), .Y(n1644) );
  OAI21X1 U4259 ( .A(n4318), .B(n7811), .C(n6446), .Y(n1643) );
  OAI21X1 U4261 ( .A(n4318), .B(n7812), .C(n6383), .Y(n1642) );
  OAI21X1 U4263 ( .A(n4318), .B(n7813), .C(n6321), .Y(n1641) );
  OAI21X1 U4265 ( .A(n4318), .B(n7814), .C(n6797), .Y(n1640) );
  OAI21X1 U4267 ( .A(n4318), .B(n7815), .C(n6726), .Y(n1639) );
  OAI21X1 U4269 ( .A(n4318), .B(n7816), .C(n6654), .Y(n1638) );
  OAI21X1 U4271 ( .A(n4318), .B(n7817), .C(n6583), .Y(n1637) );
  OAI21X1 U4273 ( .A(n6666), .B(n6809), .C(n6843), .Y(n4318) );
  NAND3X1 U4274 ( .A(wr_ptr[0]), .B(n6859), .C(wr_ptr[1]), .Y(n3320) );
  OAI21X1 U4275 ( .A(n4352), .B(n7818), .C(n5869), .Y(n1636) );
  OAI21X1 U4277 ( .A(n4352), .B(n7819), .C(n6203), .Y(n1635) );
  OAI21X1 U4279 ( .A(n4352), .B(n7820), .C(n6260), .Y(n1634) );
  OAI21X1 U4281 ( .A(n4352), .B(n7821), .C(n4670), .Y(n1633) );
  OAI21X1 U4283 ( .A(n4352), .B(n7822), .C(n4669), .Y(n1632) );
  OAI21X1 U4285 ( .A(n4352), .B(n7823), .C(n4668), .Y(n1631) );
  OAI21X1 U4287 ( .A(n4352), .B(n7824), .C(n5979), .Y(n1630) );
  OAI21X1 U4289 ( .A(n4352), .B(n7825), .C(n6034), .Y(n1629) );
  OAI21X1 U4291 ( .A(n4352), .B(n7826), .C(n5870), .Y(n1628) );
  OAI21X1 U4293 ( .A(n4352), .B(n7827), .C(n6655), .Y(n1627) );
  OAI21X1 U4295 ( .A(n4352), .B(n7828), .C(n6146), .Y(n1626) );
  OAI21X1 U4297 ( .A(n4352), .B(n7829), .C(n5925), .Y(n1625) );
  OAI21X1 U4299 ( .A(n4352), .B(n7830), .C(n6447), .Y(n1624) );
  OAI21X1 U4301 ( .A(n4352), .B(n7831), .C(n6089), .Y(n1623) );
  OAI21X1 U4303 ( .A(n4352), .B(n7832), .C(n6512), .Y(n1622) );
  OAI21X1 U4305 ( .A(n4352), .B(n7833), .C(n6322), .Y(n1621) );
  OAI21X1 U4307 ( .A(n4352), .B(n7834), .C(n6384), .Y(n1620) );
  OAI21X1 U4309 ( .A(n4352), .B(n7835), .C(n6727), .Y(n1619) );
  OAI21X1 U4311 ( .A(n4352), .B(n7836), .C(n6798), .Y(n1618) );
  OAI21X1 U4313 ( .A(n4352), .B(n7837), .C(n6584), .Y(n1617) );
  OAI21X1 U4315 ( .A(n4352), .B(n7838), .C(n6656), .Y(n1616) );
  OAI21X1 U4317 ( .A(n4352), .B(n7839), .C(n6204), .Y(n1615) );
  OAI21X1 U4319 ( .A(n4352), .B(n7840), .C(n6261), .Y(n1614) );
  OAI21X1 U4321 ( .A(n4352), .B(n7841), .C(n6090), .Y(n1613) );
  OAI21X1 U4323 ( .A(n4352), .B(n7842), .C(n6147), .Y(n1612) );
  OAI21X1 U4325 ( .A(n4352), .B(n7843), .C(n6448), .Y(n1611) );
  OAI21X1 U4327 ( .A(n4352), .B(n7844), .C(n6513), .Y(n1610) );
  OAI21X1 U4329 ( .A(n4352), .B(n7845), .C(n6323), .Y(n1609) );
  OAI21X1 U4331 ( .A(n4352), .B(n7846), .C(n6385), .Y(n1608) );
  OAI21X1 U4333 ( .A(n4352), .B(n7847), .C(n6728), .Y(n1607) );
  OAI21X1 U4335 ( .A(n4352), .B(n7848), .C(n6799), .Y(n1606) );
  OAI21X1 U4337 ( .A(n4352), .B(n7849), .C(n6585), .Y(n1605) );
  OAI21X1 U4339 ( .A(n4352), .B(n7850), .C(n6657), .Y(n1604) );
  OAI21X1 U4341 ( .A(n6455), .B(n6809), .C(n6843), .Y(n4352) );
  NAND3X1 U4342 ( .A(n6849), .B(n6859), .C(wr_ptr[1]), .Y(n3564) );
  OAI21X1 U4343 ( .A(n4386), .B(n7851), .C(n6035), .Y(n1603) );
  OAI21X1 U4345 ( .A(n4386), .B(n7852), .C(n6148), .Y(n1602) );
  OAI21X1 U4347 ( .A(n4386), .B(n7853), .C(n6091), .Y(n1601) );
  OAI21X1 U4349 ( .A(n4386), .B(n7854), .C(n4667), .Y(n1600) );
  OAI21X1 U4351 ( .A(n4386), .B(n7855), .C(n4666), .Y(n1599) );
  OAI21X1 U4353 ( .A(n4386), .B(n7856), .C(n4665), .Y(n1598) );
  OAI21X1 U4355 ( .A(n4386), .B(n7857), .C(n5926), .Y(n1597) );
  OAI21X1 U4357 ( .A(n4386), .B(n7858), .C(n5871), .Y(n1596) );
  OAI21X1 U4359 ( .A(n4386), .B(n7859), .C(n6036), .Y(n1595) );
  OAI21X1 U4361 ( .A(n4386), .B(n7860), .C(n6729), .Y(n1594) );
  OAI21X1 U4363 ( .A(n4386), .B(n7861), .C(n6205), .Y(n1593) );
  OAI21X1 U4365 ( .A(n4386), .B(n7862), .C(n5980), .Y(n1592) );
  OAI21X1 U4367 ( .A(n4386), .B(n7863), .C(n6386), .Y(n1591) );
  OAI21X1 U4369 ( .A(n4386), .B(n7864), .C(n6262), .Y(n1590) );
  OAI21X1 U4371 ( .A(n4386), .B(n7865), .C(n6324), .Y(n1589) );
  OAI21X1 U4373 ( .A(n4386), .B(n7866), .C(n6514), .Y(n1588) );
  OAI21X1 U4375 ( .A(n4386), .B(n7867), .C(n6449), .Y(n1587) );
  OAI21X1 U4377 ( .A(n4386), .B(n7868), .C(n6658), .Y(n1586) );
  OAI21X1 U4379 ( .A(n4386), .B(n7869), .C(n6586), .Y(n1585) );
  OAI21X1 U4381 ( .A(n4386), .B(n7870), .C(n6800), .Y(n1584) );
  OAI21X1 U4383 ( .A(n4386), .B(n7871), .C(n6730), .Y(n1583) );
  OAI21X1 U4385 ( .A(n4386), .B(n7872), .C(n6149), .Y(n1582) );
  OAI21X1 U4387 ( .A(n4386), .B(n7873), .C(n6092), .Y(n1581) );
  OAI21X1 U4389 ( .A(n4386), .B(n7874), .C(n6263), .Y(n1580) );
  OAI21X1 U4391 ( .A(n4386), .B(n7875), .C(n6206), .Y(n1579) );
  OAI21X1 U4393 ( .A(n4386), .B(n7876), .C(n6387), .Y(n1578) );
  OAI21X1 U4395 ( .A(n4386), .B(n7877), .C(n6325), .Y(n1577) );
  OAI21X1 U4397 ( .A(n4386), .B(n7878), .C(n6515), .Y(n1576) );
  OAI21X1 U4399 ( .A(n4386), .B(n7879), .C(n6450), .Y(n1575) );
  OAI21X1 U4401 ( .A(n4386), .B(n7880), .C(n6659), .Y(n1574) );
  OAI21X1 U4403 ( .A(n4386), .B(n7881), .C(n6587), .Y(n1573) );
  OAI21X1 U4405 ( .A(n4386), .B(n7882), .C(n6801), .Y(n1572) );
  OAI21X1 U4407 ( .A(n4386), .B(n7883), .C(n6731), .Y(n1571) );
  OAI21X1 U4409 ( .A(n6522), .B(n6809), .C(n6843), .Y(n4386) );
  NAND3X1 U4410 ( .A(n6858), .B(n6859), .C(wr_ptr[0]), .Y(n3599) );
  OAI21X1 U4411 ( .A(n4420), .B(n7884), .C(n5981), .Y(n1570) );
  OAI21X1 U4413 ( .A(n4420), .B(n7885), .C(n6093), .Y(n1569) );
  OAI21X1 U4415 ( .A(n4420), .B(n7886), .C(n6150), .Y(n1568) );
  OAI21X1 U4417 ( .A(n4420), .B(n7887), .C(n4664), .Y(n1567) );
  OAI21X1 U4419 ( .A(n4420), .B(n7888), .C(n4663), .Y(n1566) );
  OAI21X1 U4421 ( .A(n4420), .B(n7889), .C(n4662), .Y(n1565) );
  OAI21X1 U4423 ( .A(n4420), .B(n7890), .C(n5872), .Y(n1564) );
  OAI21X1 U4425 ( .A(n4420), .B(n7891), .C(n5927), .Y(n1563) );
  OAI21X1 U4427 ( .A(n4420), .B(n7892), .C(n5982), .Y(n1562) );
  OAI21X1 U4429 ( .A(n4420), .B(n7893), .C(n6802), .Y(n1561) );
  OAI21X1 U4431 ( .A(n4420), .B(n7894), .C(n6264), .Y(n1560) );
  OAI21X1 U4433 ( .A(n4420), .B(n7895), .C(n6037), .Y(n1559) );
  OAI21X1 U4435 ( .A(n4420), .B(n7896), .C(n6326), .Y(n1558) );
  OAI21X1 U4437 ( .A(n4420), .B(n7897), .C(n6207), .Y(n1557) );
  OAI21X1 U4439 ( .A(n4420), .B(n7898), .C(n6388), .Y(n1556) );
  OAI21X1 U4441 ( .A(n4420), .B(n7899), .C(n6451), .Y(n1555) );
  OAI21X1 U4443 ( .A(n4420), .B(n7900), .C(n6516), .Y(n1554) );
  OAI21X1 U4445 ( .A(n4420), .B(n7901), .C(n6588), .Y(n1553) );
  OAI21X1 U4447 ( .A(n4420), .B(n7902), .C(n6660), .Y(n1552) );
  OAI21X1 U4449 ( .A(n4420), .B(n7903), .C(n6732), .Y(n1551) );
  OAI21X1 U4451 ( .A(n4420), .B(n7904), .C(n6803), .Y(n1550) );
  OAI21X1 U4453 ( .A(n4420), .B(n7905), .C(n6094), .Y(n1549) );
  OAI21X1 U4455 ( .A(n4420), .B(n7906), .C(n6151), .Y(n1548) );
  OAI21X1 U4457 ( .A(n4420), .B(n7907), .C(n6208), .Y(n1547) );
  OAI21X1 U4459 ( .A(n4420), .B(n7908), .C(n6265), .Y(n1546) );
  OAI21X1 U4461 ( .A(n4420), .B(n7909), .C(n6327), .Y(n1545) );
  OAI21X1 U4463 ( .A(n4420), .B(n7910), .C(n6389), .Y(n1544) );
  OAI21X1 U4465 ( .A(n4420), .B(n7911), .C(n6452), .Y(n1543) );
  OAI21X1 U4467 ( .A(n4420), .B(n7912), .C(n6517), .Y(n1542) );
  OAI21X1 U4469 ( .A(n4420), .B(n7913), .C(n6589), .Y(n1541) );
  OAI21X1 U4471 ( .A(n4420), .B(n7914), .C(n6661), .Y(n1540) );
  OAI21X1 U4473 ( .A(n4420), .B(n7915), .C(n6733), .Y(n1539) );
  OAI21X1 U4475 ( .A(n4420), .B(n7916), .C(n6804), .Y(n1538) );
  OAI21X1 U4477 ( .A(n6593), .B(n6809), .C(n6843), .Y(n4420) );
  NAND3X1 U4478 ( .A(n6860), .B(n6857), .C(put), .Y(n4215) );
  NAND3X1 U4479 ( .A(n6858), .B(n6859), .C(n6849), .Y(n3634) );
  XOR2X1 U4480 ( .A(n6663), .B(n3311), .Y(fillcount[4]) );
  XNOR2X1 U4481 ( .A(n16), .B(n6857), .Y(n3311) );
  AOI21X1 U4482 ( .A(n6856), .B(n4454), .C(n6664), .Y(n3291) );
  AOI21X1 U4483 ( .A(n15), .B(n6847), .C(n6860), .Y(n4455) );
  XOR2X1 U4484 ( .A(n4454), .B(n3308), .Y(fillcount[3]) );
  XNOR2X1 U4485 ( .A(n15), .B(wr_ptr[3]), .Y(n3308) );
  OAI21X1 U4486 ( .A(n14), .B(n6390), .C(n4457), .Y(n4454) );
  OAI21X1 U4487 ( .A(n6855), .B(n6848), .C(wr_ptr[2]), .Y(n4457) );
  XOR2X1 U4488 ( .A(n6848), .B(n3307), .Y(fillcount[2]) );
  XNOR2X1 U4489 ( .A(n14), .B(wr_ptr[2]), .Y(n3307) );
  AOI21X1 U4490 ( .A(n6854), .B(n6806), .C(n6391), .Y(n4456) );
  AOI21X1 U4491 ( .A(n13), .B(n4458), .C(n6858), .Y(n4459) );
  XNOR2X1 U4492 ( .A(n6806), .B(n3310), .Y(fillcount[1]) );
  XNOR2X1 U4493 ( .A(n13), .B(n6858), .Y(n3310) );
  OAI21X1 U4494 ( .A(n12), .B(n6849), .C(n6806), .Y(fillcount[0]) );
  OR2X1 U3 ( .A(n4760), .B(n4892), .Y(n3254) );
  OR2X1 U4 ( .A(n4761), .B(n4893), .Y(n3255) );
  OR2X1 U5 ( .A(n4759), .B(n4891), .Y(n3253) );
  OR2X1 U6 ( .A(n4764), .B(n4896), .Y(n3220) );
  OR2X1 U7 ( .A(n4765), .B(n4897), .Y(n3221) );
  OR2X1 U8 ( .A(n4763), .B(n4895), .Y(n3219) );
  OR2X1 U9 ( .A(n4768), .B(n4900), .Y(n3186) );
  OR2X1 U10 ( .A(n4769), .B(n4901), .Y(n3187) );
  OR2X1 U11 ( .A(n4767), .B(n4899), .Y(n3185) );
  OR2X1 U12 ( .A(n4772), .B(n4904), .Y(n3152) );
  OR2X1 U13 ( .A(n4773), .B(n4905), .Y(n3153) );
  OR2X1 U14 ( .A(n4771), .B(n4903), .Y(n3151) );
  OR2X1 U15 ( .A(n4776), .B(n4908), .Y(n3118) );
  OR2X1 U16 ( .A(n4777), .B(n4909), .Y(n3119) );
  OR2X1 U17 ( .A(n4775), .B(n4907), .Y(n3117) );
  OR2X1 U18 ( .A(n4780), .B(n4912), .Y(n3084) );
  OR2X1 U19 ( .A(n4781), .B(n4913), .Y(n3085) );
  OR2X1 U20 ( .A(n4779), .B(n4911), .Y(n3083) );
  OR2X1 U21 ( .A(n4784), .B(n4916), .Y(n3050) );
  OR2X1 U22 ( .A(n4785), .B(n4917), .Y(n3051) );
  OR2X1 U23 ( .A(n4783), .B(n4915), .Y(n3049) );
  OR2X1 U24 ( .A(n4788), .B(n4920), .Y(n3016) );
  OR2X1 U25 ( .A(n4789), .B(n4921), .Y(n3017) );
  OR2X1 U26 ( .A(n4787), .B(n4919), .Y(n3015) );
  OR2X1 U27 ( .A(n4792), .B(n4924), .Y(n2982) );
  OR2X1 U28 ( .A(n4793), .B(n4925), .Y(n2983) );
  OR2X1 U29 ( .A(n4791), .B(n4923), .Y(n2981) );
  OR2X1 U30 ( .A(n4796), .B(n4928), .Y(n2948) );
  OR2X1 U31 ( .A(n4797), .B(n4929), .Y(n2949) );
  OR2X1 U32 ( .A(n4795), .B(n4927), .Y(n2947) );
  OR2X1 U33 ( .A(n4800), .B(n4932), .Y(n2914) );
  OR2X1 U34 ( .A(n4801), .B(n4933), .Y(n2915) );
  OR2X1 U35 ( .A(n4799), .B(n4931), .Y(n2913) );
  OR2X1 U36 ( .A(n4804), .B(n4936), .Y(n2880) );
  OR2X1 U37 ( .A(n4805), .B(n4937), .Y(n2881) );
  OR2X1 U38 ( .A(n4803), .B(n4935), .Y(n2879) );
  OR2X1 U39 ( .A(n4828), .B(n4960), .Y(n2676) );
  OR2X1 U40 ( .A(n4829), .B(n4961), .Y(n2677) );
  OR2X1 U41 ( .A(n4827), .B(n4959), .Y(n2675) );
  OR2X1 U42 ( .A(n4832), .B(n4964), .Y(n2642) );
  OR2X1 U43 ( .A(n4833), .B(n4965), .Y(n2643) );
  OR2X1 U44 ( .A(n4831), .B(n4963), .Y(n2641) );
  OR2X1 U45 ( .A(n4836), .B(n4968), .Y(n2608) );
  OR2X1 U46 ( .A(n4837), .B(n4969), .Y(n2609) );
  OR2X1 U47 ( .A(n4835), .B(n4967), .Y(n2607) );
  OR2X1 U48 ( .A(n4840), .B(n4972), .Y(n1508) );
  OR2X1 U49 ( .A(n4841), .B(n4973), .Y(n1509) );
  OR2X1 U50 ( .A(n4839), .B(n4971), .Y(n1507) );
  OR2X1 U51 ( .A(n4844), .B(n4976), .Y(n1474) );
  OR2X1 U52 ( .A(n4845), .B(n4977), .Y(n1475) );
  OR2X1 U53 ( .A(n4843), .B(n4975), .Y(n1473) );
  OR2X1 U54 ( .A(n4848), .B(n4980), .Y(n1440) );
  OR2X1 U55 ( .A(n4849), .B(n4981), .Y(n1441) );
  OR2X1 U56 ( .A(n4847), .B(n4979), .Y(n1439) );
  OR2X1 U57 ( .A(n4852), .B(n4984), .Y(n1406) );
  OR2X1 U58 ( .A(n4853), .B(n4985), .Y(n1407) );
  OR2X1 U59 ( .A(n4851), .B(n4983), .Y(n1405) );
  OR2X1 U60 ( .A(n4856), .B(n4988), .Y(n1372) );
  OR2X1 U61 ( .A(n4857), .B(n4989), .Y(n1373) );
  OR2X1 U62 ( .A(n4855), .B(n4987), .Y(n1371) );
  OR2X1 U63 ( .A(n4860), .B(n4992), .Y(n1338) );
  OR2X1 U64 ( .A(n4861), .B(n4993), .Y(n1339) );
  OR2X1 U65 ( .A(n4859), .B(n4991), .Y(n1337) );
  OR2X1 U66 ( .A(n4864), .B(n4996), .Y(n1304) );
  OR2X1 U67 ( .A(n4865), .B(n4997), .Y(n1305) );
  OR2X1 U68 ( .A(n4863), .B(n4995), .Y(n1303) );
  OR2X1 U69 ( .A(n4868), .B(n5000), .Y(n1270) );
  OR2X1 U70 ( .A(n4869), .B(n5001), .Y(n1271) );
  OR2X1 U71 ( .A(n4867), .B(n4999), .Y(n1269) );
  OR2X1 U72 ( .A(n4872), .B(n5004), .Y(n1236) );
  OR2X1 U73 ( .A(n4873), .B(n5005), .Y(n1237) );
  OR2X1 U74 ( .A(n4871), .B(n5003), .Y(n1235) );
  OR2X1 U75 ( .A(n4808), .B(n4940), .Y(n2846) );
  OR2X1 U76 ( .A(n4809), .B(n4941), .Y(n2847) );
  OR2X1 U77 ( .A(n4807), .B(n4939), .Y(n2845) );
  OR2X1 U78 ( .A(n4876), .B(n5008), .Y(n1202) );
  OR2X1 U79 ( .A(n4877), .B(n5009), .Y(n1203) );
  OR2X1 U80 ( .A(n4875), .B(n5007), .Y(n1201) );
  OR2X1 U81 ( .A(n4812), .B(n4944), .Y(n2812) );
  OR2X1 U82 ( .A(n4813), .B(n4945), .Y(n2813) );
  OR2X1 U83 ( .A(n4811), .B(n4943), .Y(n2811) );
  OR2X1 U84 ( .A(n4880), .B(n5012), .Y(n1168) );
  OR2X1 U85 ( .A(n4881), .B(n5013), .Y(n1169) );
  OR2X1 U86 ( .A(n4879), .B(n5011), .Y(n1167) );
  OR2X1 U87 ( .A(n4816), .B(n4948), .Y(n2778) );
  OR2X1 U88 ( .A(n4817), .B(n4949), .Y(n2779) );
  OR2X1 U89 ( .A(n4815), .B(n4947), .Y(n2777) );
  OR2X1 U90 ( .A(n4884), .B(n5016), .Y(n1134) );
  OR2X1 U91 ( .A(n4885), .B(n5017), .Y(n1135) );
  OR2X1 U92 ( .A(n4883), .B(n5015), .Y(n1133) );
  OR2X1 U93 ( .A(n4820), .B(n4952), .Y(n2744) );
  OR2X1 U94 ( .A(n4821), .B(n4953), .Y(n2745) );
  OR2X1 U95 ( .A(n4819), .B(n4951), .Y(n2743) );
  OR2X1 U96 ( .A(n4888), .B(n5020), .Y(n1090) );
  OR2X1 U97 ( .A(n4889), .B(n5021), .Y(n1091) );
  OR2X1 U98 ( .A(n4887), .B(n5019), .Y(n1089) );
  OR2X1 U99 ( .A(n4824), .B(n4956), .Y(n2710) );
  OR2X1 U100 ( .A(n4825), .B(n4957), .Y(n2711) );
  OR2X1 U101 ( .A(n4823), .B(n4955), .Y(n2709) );
  AND2X1 U102 ( .A(get), .B(empty_bar), .Y(n3306) );
  OR2X1 U103 ( .A(n4758), .B(n4890), .Y(n3251) );
  OR2X1 U104 ( .A(n4762), .B(n4894), .Y(n3217) );
  OR2X1 U105 ( .A(n4766), .B(n4898), .Y(n3183) );
  OR2X1 U106 ( .A(n4770), .B(n4902), .Y(n3149) );
  OR2X1 U107 ( .A(n4774), .B(n4906), .Y(n3115) );
  OR2X1 U108 ( .A(n4778), .B(n4910), .Y(n3081) );
  OR2X1 U109 ( .A(n4782), .B(n4914), .Y(n3047) );
  OR2X1 U110 ( .A(n4786), .B(n4918), .Y(n3013) );
  OR2X1 U111 ( .A(n4790), .B(n4922), .Y(n2979) );
  OR2X1 U112 ( .A(n4794), .B(n4926), .Y(n2945) );
  OR2X1 U113 ( .A(n4798), .B(n4930), .Y(n2911) );
  OR2X1 U114 ( .A(n4802), .B(n4934), .Y(n2877) );
  OR2X1 U115 ( .A(n4826), .B(n4958), .Y(n2673) );
  OR2X1 U116 ( .A(n4830), .B(n4962), .Y(n2639) );
  OR2X1 U117 ( .A(n4834), .B(n4966), .Y(n2605) );
  OR2X1 U118 ( .A(n4838), .B(n4970), .Y(n1505) );
  OR2X1 U119 ( .A(n4842), .B(n4974), .Y(n1471) );
  OR2X1 U120 ( .A(n4846), .B(n4978), .Y(n1437) );
  OR2X1 U121 ( .A(n4850), .B(n4982), .Y(n1403) );
  OR2X1 U122 ( .A(n4854), .B(n4986), .Y(n1369) );
  OR2X1 U123 ( .A(n4858), .B(n4990), .Y(n1335) );
  OR2X1 U124 ( .A(n4862), .B(n4994), .Y(n1301) );
  OR2X1 U125 ( .A(n4866), .B(n4998), .Y(n1267) );
  OR2X1 U126 ( .A(n4870), .B(n5002), .Y(n1233) );
  OR2X1 U127 ( .A(n4806), .B(n4938), .Y(n2843) );
  OR2X1 U128 ( .A(n4874), .B(n5006), .Y(n1199) );
  OR2X1 U129 ( .A(n4810), .B(n4942), .Y(n2809) );
  OR2X1 U130 ( .A(n4878), .B(n5010), .Y(n1165) );
  OR2X1 U131 ( .A(n4814), .B(n4946), .Y(n2775) );
  OR2X1 U132 ( .A(n4882), .B(n5014), .Y(n1131) );
  OR2X1 U133 ( .A(n4818), .B(n4950), .Y(n2741) );
  OR2X1 U134 ( .A(n4886), .B(n5018), .Y(n1087) );
  OR2X1 U135 ( .A(n4822), .B(n4954), .Y(n2707) );
  OR2X1 U136 ( .A(n6666), .B(n6807), .Y(n3319) );
  OR2X1 U137 ( .A(n6735), .B(n6849), .Y(n3294) );
  AND2X1 U138 ( .A(n6842), .B(n6591), .Y(n3299) );
  AND2X1 U139 ( .A(n6842), .B(n6590), .Y(n3276) );
  AND2X1 U140 ( .A(n6842), .B(n6735), .Y(n3293) );
  BUFX2 U141 ( .A(n2602), .Y(n4626) );
  BUFX2 U142 ( .A(n4492), .Y(n4627) );
  BUFX2 U143 ( .A(n4491), .Y(n4628) );
  BUFX2 U144 ( .A(n4490), .Y(n4629) );
  BUFX2 U145 ( .A(n4489), .Y(n4630) );
  BUFX2 U146 ( .A(n4488), .Y(n4631) );
  BUFX2 U147 ( .A(n4487), .Y(n4632) );
  BUFX2 U148 ( .A(n4486), .Y(n4633) );
  BUFX2 U149 ( .A(n4485), .Y(n4634) );
  BUFX2 U150 ( .A(n4484), .Y(n4635) );
  BUFX2 U151 ( .A(n4483), .Y(n4636) );
  BUFX2 U152 ( .A(n4482), .Y(n4637) );
  BUFX2 U153 ( .A(n4481), .Y(n4638) );
  BUFX2 U154 ( .A(n4480), .Y(n4639) );
  BUFX2 U155 ( .A(n4479), .Y(n4640) );
  BUFX2 U156 ( .A(n4478), .Y(n4641) );
  BUFX2 U157 ( .A(n4477), .Y(n4642) );
  BUFX2 U158 ( .A(n4476), .Y(n4643) );
  BUFX2 U159 ( .A(n4475), .Y(n4644) );
  BUFX2 U160 ( .A(n4474), .Y(n4645) );
  BUFX2 U161 ( .A(n4473), .Y(n4646) );
  BUFX2 U162 ( .A(n4472), .Y(n4647) );
  BUFX2 U163 ( .A(n4471), .Y(n4648) );
  BUFX2 U164 ( .A(n4470), .Y(n4649) );
  BUFX2 U165 ( .A(n4469), .Y(n4650) );
  BUFX2 U166 ( .A(n4468), .Y(n4651) );
  BUFX2 U167 ( .A(n4467), .Y(n4652) );
  BUFX2 U168 ( .A(n4466), .Y(n4653) );
  BUFX2 U169 ( .A(n4465), .Y(n4654) );
  BUFX2 U170 ( .A(n4464), .Y(n4655) );
  BUFX2 U171 ( .A(n4463), .Y(n4656) );
  BUFX2 U172 ( .A(n4462), .Y(n4657) );
  BUFX2 U173 ( .A(n4461), .Y(n4658) );
  BUFX2 U174 ( .A(n4460), .Y(n4659) );
  BUFX2 U175 ( .A(n3305), .Y(n4660) );
  BUFX2 U176 ( .A(n3302), .Y(n4661) );
  AND2X1 U177 ( .A(n3335), .B(n4420), .Y(n4426) );
  INVX1 U178 ( .A(n4426), .Y(n4662) );
  AND2X1 U179 ( .A(n3333), .B(n4420), .Y(n4425) );
  INVX1 U180 ( .A(n4425), .Y(n4663) );
  AND2X1 U181 ( .A(n3331), .B(n4420), .Y(n4424) );
  INVX1 U182 ( .A(n4424), .Y(n4664) );
  AND2X1 U183 ( .A(n3335), .B(n4386), .Y(n4392) );
  INVX1 U184 ( .A(n4392), .Y(n4665) );
  AND2X1 U185 ( .A(n3333), .B(n4386), .Y(n4391) );
  INVX1 U186 ( .A(n4391), .Y(n4666) );
  AND2X1 U187 ( .A(n3331), .B(n4386), .Y(n4390) );
  INVX1 U188 ( .A(n4390), .Y(n4667) );
  AND2X1 U189 ( .A(n3335), .B(n4352), .Y(n4358) );
  INVX1 U190 ( .A(n4358), .Y(n4668) );
  AND2X1 U191 ( .A(n3333), .B(n4352), .Y(n4357) );
  INVX1 U192 ( .A(n4357), .Y(n4669) );
  AND2X1 U193 ( .A(n3331), .B(n4352), .Y(n4356) );
  INVX1 U194 ( .A(n4356), .Y(n4670) );
  AND2X1 U195 ( .A(n3335), .B(n4318), .Y(n4324) );
  INVX1 U196 ( .A(n4324), .Y(n4671) );
  AND2X1 U197 ( .A(n3333), .B(n4318), .Y(n4323) );
  INVX1 U198 ( .A(n4323), .Y(n4672) );
  AND2X1 U199 ( .A(n3331), .B(n4318), .Y(n4322) );
  INVX1 U200 ( .A(n4322), .Y(n4673) );
  AND2X1 U201 ( .A(n3335), .B(n4284), .Y(n4290) );
  INVX1 U202 ( .A(n4290), .Y(n4674) );
  AND2X1 U203 ( .A(n3333), .B(n4284), .Y(n4289) );
  INVX1 U204 ( .A(n4289), .Y(n4675) );
  AND2X1 U205 ( .A(n3331), .B(n4284), .Y(n4288) );
  INVX1 U206 ( .A(n4288), .Y(n4676) );
  AND2X1 U207 ( .A(n3335), .B(n4250), .Y(n4256) );
  INVX1 U208 ( .A(n4256), .Y(n4677) );
  AND2X1 U209 ( .A(n3333), .B(n4250), .Y(n4255) );
  INVX1 U210 ( .A(n4255), .Y(n4678) );
  AND2X1 U211 ( .A(n3331), .B(n4250), .Y(n4254) );
  INVX1 U212 ( .A(n4254), .Y(n4679) );
  AND2X1 U213 ( .A(n3335), .B(n4216), .Y(n4222) );
  INVX1 U214 ( .A(n4222), .Y(n4680) );
  AND2X1 U215 ( .A(n3333), .B(n4216), .Y(n4221) );
  INVX1 U216 ( .A(n4221), .Y(n4681) );
  AND2X1 U217 ( .A(n3331), .B(n4216), .Y(n4220) );
  INVX1 U218 ( .A(n4220), .Y(n4682) );
  AND2X1 U219 ( .A(n3335), .B(n4181), .Y(n4187) );
  INVX1 U220 ( .A(n4187), .Y(n4683) );
  AND2X1 U221 ( .A(n3333), .B(n4181), .Y(n4186) );
  INVX1 U222 ( .A(n4186), .Y(n4684) );
  AND2X1 U223 ( .A(n3331), .B(n4181), .Y(n4185) );
  INVX1 U224 ( .A(n4185), .Y(n4685) );
  AND2X1 U225 ( .A(n3335), .B(n4147), .Y(n4153) );
  INVX1 U226 ( .A(n4153), .Y(n4686) );
  AND2X1 U227 ( .A(n3333), .B(n4147), .Y(n4152) );
  INVX1 U228 ( .A(n4152), .Y(n4687) );
  AND2X1 U229 ( .A(n3331), .B(n4147), .Y(n4151) );
  INVX1 U230 ( .A(n4151), .Y(n4688) );
  AND2X1 U231 ( .A(n3335), .B(n4113), .Y(n4119) );
  INVX1 U232 ( .A(n4119), .Y(n4689) );
  AND2X1 U233 ( .A(n3333), .B(n4113), .Y(n4118) );
  INVX1 U234 ( .A(n4118), .Y(n4690) );
  AND2X1 U235 ( .A(n3331), .B(n4113), .Y(n4117) );
  INVX1 U236 ( .A(n4117), .Y(n4691) );
  AND2X1 U237 ( .A(n3335), .B(n4079), .Y(n4085) );
  INVX1 U238 ( .A(n4085), .Y(n4692) );
  AND2X1 U239 ( .A(n3333), .B(n4079), .Y(n4084) );
  INVX1 U240 ( .A(n4084), .Y(n4693) );
  AND2X1 U241 ( .A(n3331), .B(n4079), .Y(n4083) );
  INVX1 U242 ( .A(n4083), .Y(n4694) );
  AND2X1 U243 ( .A(n3335), .B(n4045), .Y(n4051) );
  INVX1 U244 ( .A(n4051), .Y(n4695) );
  AND2X1 U245 ( .A(n3333), .B(n4045), .Y(n4050) );
  INVX1 U246 ( .A(n4050), .Y(n4696) );
  AND2X1 U247 ( .A(n3331), .B(n4045), .Y(n4049) );
  INVX1 U248 ( .A(n4049), .Y(n4697) );
  AND2X1 U249 ( .A(n3335), .B(n4011), .Y(n4017) );
  INVX1 U250 ( .A(n4017), .Y(n4698) );
  AND2X1 U251 ( .A(n3333), .B(n4011), .Y(n4016) );
  INVX1 U252 ( .A(n4016), .Y(n4699) );
  AND2X1 U253 ( .A(n3331), .B(n4011), .Y(n4015) );
  INVX1 U254 ( .A(n4015), .Y(n4700) );
  AND2X1 U255 ( .A(n3335), .B(n3977), .Y(n3983) );
  INVX1 U256 ( .A(n3983), .Y(n4701) );
  AND2X1 U257 ( .A(n3333), .B(n3977), .Y(n3982) );
  INVX1 U258 ( .A(n3982), .Y(n4702) );
  AND2X1 U259 ( .A(n3331), .B(n3977), .Y(n3981) );
  INVX1 U260 ( .A(n3981), .Y(n4703) );
  AND2X1 U261 ( .A(n3335), .B(n3943), .Y(n3949) );
  INVX1 U262 ( .A(n3949), .Y(n4704) );
  AND2X1 U263 ( .A(n3333), .B(n3943), .Y(n3948) );
  INVX1 U264 ( .A(n3948), .Y(n4705) );
  AND2X1 U265 ( .A(n3331), .B(n3943), .Y(n3947) );
  INVX1 U266 ( .A(n3947), .Y(n4706) );
  AND2X1 U267 ( .A(n3335), .B(n3908), .Y(n3914) );
  INVX1 U268 ( .A(n3914), .Y(n4707) );
  AND2X1 U269 ( .A(n3333), .B(n3908), .Y(n3913) );
  INVX1 U270 ( .A(n3913), .Y(n4708) );
  AND2X1 U271 ( .A(n3331), .B(n3908), .Y(n3912) );
  INVX1 U272 ( .A(n3912), .Y(n4709) );
  AND2X1 U273 ( .A(n3335), .B(n3874), .Y(n3880) );
  INVX1 U274 ( .A(n3880), .Y(n4710) );
  AND2X1 U275 ( .A(n3333), .B(n3874), .Y(n3879) );
  INVX1 U276 ( .A(n3879), .Y(n4711) );
  AND2X1 U277 ( .A(n3331), .B(n3874), .Y(n3878) );
  INVX1 U278 ( .A(n3878), .Y(n4712) );
  AND2X1 U279 ( .A(n3335), .B(n3840), .Y(n3846) );
  INVX1 U280 ( .A(n3846), .Y(n4713) );
  AND2X1 U281 ( .A(n3333), .B(n3840), .Y(n3845) );
  INVX1 U282 ( .A(n3845), .Y(n4714) );
  AND2X1 U283 ( .A(n3331), .B(n3840), .Y(n3844) );
  INVX1 U284 ( .A(n3844), .Y(n4715) );
  AND2X1 U285 ( .A(n3335), .B(n3806), .Y(n3812) );
  INVX1 U286 ( .A(n3812), .Y(n4716) );
  AND2X1 U287 ( .A(n3333), .B(n3806), .Y(n3811) );
  INVX1 U288 ( .A(n3811), .Y(n4717) );
  AND2X1 U289 ( .A(n3331), .B(n3806), .Y(n3810) );
  INVX1 U290 ( .A(n3810), .Y(n4718) );
  AND2X1 U291 ( .A(n3335), .B(n3772), .Y(n3778) );
  INVX1 U292 ( .A(n3778), .Y(n4719) );
  AND2X1 U293 ( .A(n3333), .B(n3772), .Y(n3777) );
  INVX1 U294 ( .A(n3777), .Y(n4720) );
  AND2X1 U295 ( .A(n3331), .B(n3772), .Y(n3776) );
  INVX1 U296 ( .A(n3776), .Y(n4721) );
  AND2X1 U297 ( .A(n3335), .B(n3738), .Y(n3744) );
  INVX1 U298 ( .A(n3744), .Y(n4722) );
  AND2X1 U299 ( .A(n3333), .B(n3738), .Y(n3743) );
  INVX1 U300 ( .A(n3743), .Y(n4723) );
  AND2X1 U301 ( .A(n3331), .B(n3738), .Y(n3742) );
  INVX1 U302 ( .A(n3742), .Y(n4724) );
  AND2X1 U303 ( .A(n3335), .B(n3704), .Y(n3710) );
  INVX1 U304 ( .A(n3710), .Y(n4725) );
  AND2X1 U305 ( .A(n3333), .B(n3704), .Y(n3709) );
  INVX1 U306 ( .A(n3709), .Y(n4726) );
  AND2X1 U307 ( .A(n3331), .B(n3704), .Y(n3708) );
  INVX1 U308 ( .A(n3708), .Y(n4727) );
  AND2X1 U309 ( .A(n3335), .B(n3670), .Y(n3676) );
  INVX1 U310 ( .A(n3676), .Y(n4728) );
  AND2X1 U311 ( .A(n3333), .B(n3670), .Y(n3675) );
  INVX1 U312 ( .A(n3675), .Y(n4729) );
  AND2X1 U313 ( .A(n3331), .B(n3670), .Y(n3674) );
  INVX1 U314 ( .A(n3674), .Y(n4730) );
  AND2X1 U315 ( .A(n3335), .B(n3635), .Y(n3641) );
  INVX1 U316 ( .A(n3641), .Y(n4731) );
  AND2X1 U317 ( .A(n3333), .B(n3635), .Y(n3640) );
  INVX1 U318 ( .A(n3640), .Y(n4732) );
  AND2X1 U319 ( .A(n3331), .B(n3635), .Y(n3639) );
  INVX1 U320 ( .A(n3639), .Y(n4733) );
  AND2X1 U321 ( .A(n3335), .B(n3600), .Y(n3606) );
  INVX1 U322 ( .A(n3606), .Y(n4734) );
  AND2X1 U323 ( .A(n3333), .B(n3600), .Y(n3605) );
  INVX1 U324 ( .A(n3605), .Y(n4735) );
  AND2X1 U325 ( .A(n3331), .B(n3600), .Y(n3604) );
  INVX1 U326 ( .A(n3604), .Y(n4736) );
  AND2X1 U327 ( .A(n3335), .B(n3565), .Y(n3571) );
  INVX1 U328 ( .A(n3571), .Y(n4737) );
  AND2X1 U329 ( .A(n3333), .B(n3565), .Y(n3570) );
  INVX1 U330 ( .A(n3570), .Y(n4738) );
  AND2X1 U331 ( .A(n3331), .B(n3565), .Y(n3569) );
  INVX1 U332 ( .A(n3569), .Y(n4739) );
  AND2X1 U333 ( .A(n3335), .B(n3530), .Y(n3536) );
  INVX1 U334 ( .A(n3536), .Y(n4740) );
  AND2X1 U335 ( .A(n3333), .B(n3530), .Y(n3535) );
  INVX1 U336 ( .A(n3535), .Y(n4741) );
  AND2X1 U337 ( .A(n3331), .B(n3530), .Y(n3534) );
  INVX1 U338 ( .A(n3534), .Y(n4742) );
  AND2X1 U339 ( .A(n3335), .B(n3496), .Y(n3502) );
  INVX1 U340 ( .A(n3502), .Y(n4743) );
  AND2X1 U341 ( .A(n3333), .B(n3496), .Y(n3501) );
  INVX1 U342 ( .A(n3501), .Y(n4744) );
  AND2X1 U343 ( .A(n3331), .B(n3496), .Y(n3500) );
  INVX1 U344 ( .A(n3500), .Y(n4745) );
  AND2X1 U345 ( .A(n3335), .B(n3461), .Y(n3467) );
  INVX1 U346 ( .A(n3467), .Y(n4746) );
  AND2X1 U347 ( .A(n3333), .B(n3461), .Y(n3466) );
  INVX1 U348 ( .A(n3466), .Y(n4747) );
  AND2X1 U349 ( .A(n3331), .B(n3461), .Y(n3465) );
  INVX1 U350 ( .A(n3465), .Y(n4748) );
  AND2X1 U351 ( .A(n3335), .B(n3426), .Y(n3432) );
  INVX1 U352 ( .A(n3432), .Y(n4749) );
  AND2X1 U353 ( .A(n3333), .B(n3426), .Y(n3431) );
  INVX1 U354 ( .A(n3431), .Y(n4750) );
  AND2X1 U355 ( .A(n3331), .B(n3426), .Y(n3430) );
  INVX1 U356 ( .A(n3430), .Y(n4751) );
  AND2X1 U357 ( .A(n3335), .B(n3391), .Y(n3397) );
  INVX1 U358 ( .A(n3397), .Y(n4752) );
  AND2X1 U359 ( .A(n3333), .B(n3391), .Y(n3396) );
  INVX1 U360 ( .A(n3396), .Y(n4753) );
  AND2X1 U361 ( .A(n3331), .B(n3391), .Y(n3395) );
  INVX1 U362 ( .A(n3395), .Y(n4754) );
  AND2X1 U363 ( .A(n3335), .B(n3323), .Y(n3334) );
  INVX1 U364 ( .A(n3334), .Y(n4755) );
  AND2X1 U365 ( .A(n3333), .B(n3323), .Y(n3332) );
  INVX1 U366 ( .A(n3332), .Y(n4756) );
  AND2X1 U367 ( .A(n3331), .B(n3323), .Y(n3330) );
  INVX1 U368 ( .A(n3330), .Y(n4757) );
  BUFX2 U369 ( .A(n3280), .Y(n4758) );
  BUFX2 U370 ( .A(n3272), .Y(n4759) );
  BUFX2 U371 ( .A(n3264), .Y(n4760) );
  BUFX2 U372 ( .A(n3256), .Y(n4761) );
  BUFX2 U373 ( .A(n3243), .Y(n4762) );
  BUFX2 U374 ( .A(n3236), .Y(n4763) );
  BUFX2 U375 ( .A(n3229), .Y(n4764) );
  BUFX2 U376 ( .A(n3222), .Y(n4765) );
  BUFX2 U377 ( .A(n3209), .Y(n4766) );
  BUFX2 U378 ( .A(n3202), .Y(n4767) );
  BUFX2 U379 ( .A(n3195), .Y(n4768) );
  BUFX2 U380 ( .A(n3188), .Y(n4769) );
  BUFX2 U381 ( .A(n3175), .Y(n4770) );
  BUFX2 U382 ( .A(n3168), .Y(n4771) );
  BUFX2 U383 ( .A(n3161), .Y(n4772) );
  BUFX2 U384 ( .A(n3154), .Y(n4773) );
  BUFX2 U385 ( .A(n3141), .Y(n4774) );
  BUFX2 U386 ( .A(n3134), .Y(n4775) );
  BUFX2 U387 ( .A(n3127), .Y(n4776) );
  BUFX2 U388 ( .A(n3120), .Y(n4777) );
  BUFX2 U389 ( .A(n3107), .Y(n4778) );
  BUFX2 U390 ( .A(n3100), .Y(n4779) );
  BUFX2 U391 ( .A(n3093), .Y(n4780) );
  BUFX2 U392 ( .A(n3086), .Y(n4781) );
  BUFX2 U393 ( .A(n3073), .Y(n4782) );
  BUFX2 U394 ( .A(n3066), .Y(n4783) );
  BUFX2 U395 ( .A(n3059), .Y(n4784) );
  BUFX2 U396 ( .A(n3052), .Y(n4785) );
  BUFX2 U397 ( .A(n3039), .Y(n4786) );
  BUFX2 U398 ( .A(n3032), .Y(n4787) );
  BUFX2 U399 ( .A(n3025), .Y(n4788) );
  BUFX2 U400 ( .A(n3018), .Y(n4789) );
  BUFX2 U401 ( .A(n3005), .Y(n4790) );
  BUFX2 U402 ( .A(n2998), .Y(n4791) );
  BUFX2 U403 ( .A(n2991), .Y(n4792) );
  BUFX2 U404 ( .A(n2984), .Y(n4793) );
  BUFX2 U405 ( .A(n2971), .Y(n4794) );
  BUFX2 U406 ( .A(n2964), .Y(n4795) );
  BUFX2 U407 ( .A(n2957), .Y(n4796) );
  BUFX2 U408 ( .A(n2950), .Y(n4797) );
  BUFX2 U409 ( .A(n2937), .Y(n4798) );
  BUFX2 U410 ( .A(n2930), .Y(n4799) );
  BUFX2 U411 ( .A(n2923), .Y(n4800) );
  BUFX2 U412 ( .A(n2916), .Y(n4801) );
  BUFX2 U413 ( .A(n2903), .Y(n4802) );
  BUFX2 U414 ( .A(n2896), .Y(n4803) );
  BUFX2 U415 ( .A(n2889), .Y(n4804) );
  BUFX2 U416 ( .A(n2882), .Y(n4805) );
  BUFX2 U417 ( .A(n2869), .Y(n4806) );
  BUFX2 U418 ( .A(n2862), .Y(n4807) );
  BUFX2 U419 ( .A(n2855), .Y(n4808) );
  BUFX2 U420 ( .A(n2848), .Y(n4809) );
  BUFX2 U421 ( .A(n2835), .Y(n4810) );
  BUFX2 U422 ( .A(n2828), .Y(n4811) );
  BUFX2 U423 ( .A(n2821), .Y(n4812) );
  BUFX2 U424 ( .A(n2814), .Y(n4813) );
  BUFX2 U425 ( .A(n2801), .Y(n4814) );
  BUFX2 U426 ( .A(n2794), .Y(n4815) );
  BUFX2 U427 ( .A(n2787), .Y(n4816) );
  BUFX2 U428 ( .A(n2780), .Y(n4817) );
  BUFX2 U429 ( .A(n2767), .Y(n4818) );
  BUFX2 U430 ( .A(n2760), .Y(n4819) );
  BUFX2 U431 ( .A(n2753), .Y(n4820) );
  BUFX2 U432 ( .A(n2746), .Y(n4821) );
  BUFX2 U433 ( .A(n2733), .Y(n4822) );
  BUFX2 U434 ( .A(n2726), .Y(n4823) );
  BUFX2 U435 ( .A(n2719), .Y(n4824) );
  BUFX2 U436 ( .A(n2712), .Y(n4825) );
  BUFX2 U437 ( .A(n2699), .Y(n4826) );
  BUFX2 U438 ( .A(n2692), .Y(n4827) );
  BUFX2 U439 ( .A(n2685), .Y(n4828) );
  BUFX2 U440 ( .A(n2678), .Y(n4829) );
  BUFX2 U441 ( .A(n2665), .Y(n4830) );
  BUFX2 U442 ( .A(n2658), .Y(n4831) );
  BUFX2 U443 ( .A(n2651), .Y(n4832) );
  BUFX2 U444 ( .A(n2644), .Y(n4833) );
  BUFX2 U445 ( .A(n2631), .Y(n4834) );
  BUFX2 U446 ( .A(n2624), .Y(n4835) );
  BUFX2 U447 ( .A(n2617), .Y(n4836) );
  BUFX2 U448 ( .A(n2610), .Y(n4837) );
  BUFX2 U449 ( .A(n1531), .Y(n4838) );
  BUFX2 U450 ( .A(n1524), .Y(n4839) );
  BUFX2 U451 ( .A(n1517), .Y(n4840) );
  BUFX2 U452 ( .A(n1510), .Y(n4841) );
  BUFX2 U453 ( .A(n1497), .Y(n4842) );
  BUFX2 U454 ( .A(n1490), .Y(n4843) );
  BUFX2 U455 ( .A(n1483), .Y(n4844) );
  BUFX2 U456 ( .A(n1476), .Y(n4845) );
  BUFX2 U457 ( .A(n1463), .Y(n4846) );
  BUFX2 U458 ( .A(n1456), .Y(n4847) );
  BUFX2 U459 ( .A(n1449), .Y(n4848) );
  BUFX2 U460 ( .A(n1442), .Y(n4849) );
  BUFX2 U461 ( .A(n1429), .Y(n4850) );
  BUFX2 U462 ( .A(n1422), .Y(n4851) );
  BUFX2 U463 ( .A(n1415), .Y(n4852) );
  BUFX2 U464 ( .A(n1408), .Y(n4853) );
  BUFX2 U465 ( .A(n1395), .Y(n4854) );
  BUFX2 U466 ( .A(n1388), .Y(n4855) );
  BUFX2 U467 ( .A(n1381), .Y(n4856) );
  BUFX2 U468 ( .A(n1374), .Y(n4857) );
  BUFX2 U469 ( .A(n1361), .Y(n4858) );
  BUFX2 U470 ( .A(n1354), .Y(n4859) );
  BUFX2 U471 ( .A(n1347), .Y(n4860) );
  BUFX2 U472 ( .A(n1340), .Y(n4861) );
  BUFX2 U473 ( .A(n1327), .Y(n4862) );
  BUFX2 U474 ( .A(n1320), .Y(n4863) );
  BUFX2 U475 ( .A(n1313), .Y(n4864) );
  BUFX2 U476 ( .A(n1306), .Y(n4865) );
  BUFX2 U477 ( .A(n1293), .Y(n4866) );
  BUFX2 U478 ( .A(n1286), .Y(n4867) );
  BUFX2 U479 ( .A(n1279), .Y(n4868) );
  BUFX2 U480 ( .A(n1272), .Y(n4869) );
  BUFX2 U481 ( .A(n1259), .Y(n4870) );
  BUFX2 U482 ( .A(n1252), .Y(n4871) );
  BUFX2 U483 ( .A(n1245), .Y(n4872) );
  BUFX2 U484 ( .A(n1238), .Y(n4873) );
  BUFX2 U485 ( .A(n1225), .Y(n4874) );
  BUFX2 U486 ( .A(n1218), .Y(n4875) );
  BUFX2 U487 ( .A(n1211), .Y(n4876) );
  BUFX2 U488 ( .A(n1204), .Y(n4877) );
  BUFX2 U489 ( .A(n1191), .Y(n4878) );
  BUFX2 U490 ( .A(n1184), .Y(n4879) );
  BUFX2 U491 ( .A(n1177), .Y(n4880) );
  BUFX2 U492 ( .A(n1170), .Y(n4881) );
  BUFX2 U493 ( .A(n1157), .Y(n4882) );
  BUFX2 U494 ( .A(n1150), .Y(n4883) );
  BUFX2 U495 ( .A(n1143), .Y(n4884) );
  BUFX2 U496 ( .A(n1136), .Y(n4885) );
  BUFX2 U497 ( .A(n1122), .Y(n4886) );
  BUFX2 U498 ( .A(n1114), .Y(n4887) );
  BUFX2 U499 ( .A(n1106), .Y(n4888) );
  BUFX2 U500 ( .A(n1092), .Y(n4889) );
  BUFX2 U501 ( .A(n3281), .Y(n4890) );
  BUFX2 U502 ( .A(n3273), .Y(n4891) );
  BUFX2 U503 ( .A(n3265), .Y(n4892) );
  BUFX2 U504 ( .A(n3257), .Y(n4893) );
  BUFX2 U505 ( .A(n3244), .Y(n4894) );
  BUFX2 U506 ( .A(n3237), .Y(n4895) );
  BUFX2 U507 ( .A(n3230), .Y(n4896) );
  BUFX2 U508 ( .A(n3223), .Y(n4897) );
  BUFX2 U509 ( .A(n3210), .Y(n4898) );
  BUFX2 U510 ( .A(n3203), .Y(n4899) );
  BUFX2 U511 ( .A(n3196), .Y(n4900) );
  BUFX2 U512 ( .A(n3189), .Y(n4901) );
  BUFX2 U513 ( .A(n3176), .Y(n4902) );
  BUFX2 U514 ( .A(n3169), .Y(n4903) );
  BUFX2 U515 ( .A(n3162), .Y(n4904) );
  BUFX2 U516 ( .A(n3155), .Y(n4905) );
  BUFX2 U517 ( .A(n3142), .Y(n4906) );
  BUFX2 U518 ( .A(n3135), .Y(n4907) );
  BUFX2 U519 ( .A(n3128), .Y(n4908) );
  BUFX2 U520 ( .A(n3121), .Y(n4909) );
  BUFX2 U521 ( .A(n3108), .Y(n4910) );
  BUFX2 U522 ( .A(n3101), .Y(n4911) );
  BUFX2 U523 ( .A(n3094), .Y(n4912) );
  BUFX2 U524 ( .A(n3087), .Y(n4913) );
  BUFX2 U525 ( .A(n3074), .Y(n4914) );
  BUFX2 U526 ( .A(n3067), .Y(n4915) );
  BUFX2 U527 ( .A(n3060), .Y(n4916) );
  BUFX2 U528 ( .A(n3053), .Y(n4917) );
  BUFX2 U529 ( .A(n3040), .Y(n4918) );
  BUFX2 U530 ( .A(n3033), .Y(n4919) );
  BUFX2 U531 ( .A(n3026), .Y(n4920) );
  BUFX2 U532 ( .A(n3019), .Y(n4921) );
  BUFX2 U533 ( .A(n3006), .Y(n4922) );
  BUFX2 U534 ( .A(n2999), .Y(n4923) );
  BUFX2 U535 ( .A(n2992), .Y(n4924) );
  BUFX2 U536 ( .A(n2985), .Y(n4925) );
  BUFX2 U537 ( .A(n2972), .Y(n4926) );
  BUFX2 U538 ( .A(n2965), .Y(n4927) );
  BUFX2 U539 ( .A(n2958), .Y(n4928) );
  BUFX2 U540 ( .A(n2951), .Y(n4929) );
  BUFX2 U541 ( .A(n2938), .Y(n4930) );
  BUFX2 U542 ( .A(n2931), .Y(n4931) );
  BUFX2 U543 ( .A(n2924), .Y(n4932) );
  BUFX2 U544 ( .A(n2917), .Y(n4933) );
  BUFX2 U545 ( .A(n2904), .Y(n4934) );
  BUFX2 U546 ( .A(n2897), .Y(n4935) );
  BUFX2 U547 ( .A(n2890), .Y(n4936) );
  BUFX2 U548 ( .A(n2883), .Y(n4937) );
  BUFX2 U549 ( .A(n2870), .Y(n4938) );
  BUFX2 U550 ( .A(n2863), .Y(n4939) );
  BUFX2 U551 ( .A(n2856), .Y(n4940) );
  BUFX2 U552 ( .A(n2849), .Y(n4941) );
  BUFX2 U553 ( .A(n2836), .Y(n4942) );
  BUFX2 U554 ( .A(n2829), .Y(n4943) );
  BUFX2 U555 ( .A(n2822), .Y(n4944) );
  BUFX2 U556 ( .A(n2815), .Y(n4945) );
  BUFX2 U557 ( .A(n2802), .Y(n4946) );
  BUFX2 U558 ( .A(n2795), .Y(n4947) );
  BUFX2 U559 ( .A(n2788), .Y(n4948) );
  BUFX2 U560 ( .A(n2781), .Y(n4949) );
  BUFX2 U561 ( .A(n2768), .Y(n4950) );
  BUFX2 U562 ( .A(n2761), .Y(n4951) );
  BUFX2 U563 ( .A(n2754), .Y(n4952) );
  BUFX2 U564 ( .A(n2747), .Y(n4953) );
  BUFX2 U565 ( .A(n2734), .Y(n4954) );
  BUFX2 U566 ( .A(n2727), .Y(n4955) );
  BUFX2 U567 ( .A(n2720), .Y(n4956) );
  BUFX2 U568 ( .A(n2713), .Y(n4957) );
  BUFX2 U569 ( .A(n2700), .Y(n4958) );
  BUFX2 U570 ( .A(n2693), .Y(n4959) );
  BUFX2 U571 ( .A(n2686), .Y(n4960) );
  BUFX2 U572 ( .A(n2679), .Y(n4961) );
  BUFX2 U573 ( .A(n2666), .Y(n4962) );
  BUFX2 U574 ( .A(n2659), .Y(n4963) );
  BUFX2 U575 ( .A(n2652), .Y(n4964) );
  BUFX2 U576 ( .A(n2645), .Y(n4965) );
  BUFX2 U577 ( .A(n2632), .Y(n4966) );
  BUFX2 U578 ( .A(n2625), .Y(n4967) );
  BUFX2 U579 ( .A(n2618), .Y(n4968) );
  BUFX2 U580 ( .A(n2611), .Y(n4969) );
  BUFX2 U581 ( .A(n1532), .Y(n4970) );
  BUFX2 U582 ( .A(n1525), .Y(n4971) );
  BUFX2 U583 ( .A(n1518), .Y(n4972) );
  BUFX2 U584 ( .A(n1511), .Y(n4973) );
  BUFX2 U585 ( .A(n1498), .Y(n4974) );
  BUFX2 U586 ( .A(n1491), .Y(n4975) );
  BUFX2 U587 ( .A(n1484), .Y(n4976) );
  BUFX2 U588 ( .A(n1477), .Y(n4977) );
  BUFX2 U589 ( .A(n1464), .Y(n4978) );
  BUFX2 U590 ( .A(n1457), .Y(n4979) );
  BUFX2 U591 ( .A(n1450), .Y(n4980) );
  BUFX2 U592 ( .A(n1443), .Y(n4981) );
  BUFX2 U593 ( .A(n1430), .Y(n4982) );
  BUFX2 U594 ( .A(n1423), .Y(n4983) );
  BUFX2 U595 ( .A(n1416), .Y(n4984) );
  BUFX2 U596 ( .A(n1409), .Y(n4985) );
  BUFX2 U597 ( .A(n1396), .Y(n4986) );
  BUFX2 U598 ( .A(n1389), .Y(n4987) );
  BUFX2 U599 ( .A(n1382), .Y(n4988) );
  BUFX2 U600 ( .A(n1375), .Y(n4989) );
  BUFX2 U601 ( .A(n1362), .Y(n4990) );
  BUFX2 U602 ( .A(n1355), .Y(n4991) );
  BUFX2 U603 ( .A(n1348), .Y(n4992) );
  BUFX2 U604 ( .A(n1341), .Y(n4993) );
  BUFX2 U605 ( .A(n1328), .Y(n4994) );
  BUFX2 U606 ( .A(n1321), .Y(n4995) );
  BUFX2 U607 ( .A(n1314), .Y(n4996) );
  BUFX2 U608 ( .A(n1307), .Y(n4997) );
  BUFX2 U609 ( .A(n1294), .Y(n4998) );
  BUFX2 U610 ( .A(n1287), .Y(n4999) );
  BUFX2 U611 ( .A(n1280), .Y(n5000) );
  BUFX2 U612 ( .A(n1273), .Y(n5001) );
  BUFX2 U613 ( .A(n1260), .Y(n5002) );
  BUFX2 U614 ( .A(n1253), .Y(n5003) );
  BUFX2 U615 ( .A(n1246), .Y(n5004) );
  BUFX2 U616 ( .A(n1239), .Y(n5005) );
  BUFX2 U617 ( .A(n1226), .Y(n5006) );
  BUFX2 U618 ( .A(n1219), .Y(n5007) );
  BUFX2 U619 ( .A(n1212), .Y(n5008) );
  BUFX2 U620 ( .A(n1205), .Y(n5009) );
  BUFX2 U621 ( .A(n1192), .Y(n5010) );
  BUFX2 U622 ( .A(n1185), .Y(n5011) );
  BUFX2 U623 ( .A(n1178), .Y(n5012) );
  BUFX2 U624 ( .A(n1171), .Y(n5013) );
  BUFX2 U625 ( .A(n1158), .Y(n5014) );
  BUFX2 U626 ( .A(n1151), .Y(n5015) );
  BUFX2 U627 ( .A(n1144), .Y(n5016) );
  BUFX2 U628 ( .A(n1137), .Y(n5017) );
  BUFX2 U629 ( .A(n1123), .Y(n5018) );
  BUFX2 U630 ( .A(n1115), .Y(n5019) );
  BUFX2 U631 ( .A(n1107), .Y(n5020) );
  BUFX2 U632 ( .A(n1093), .Y(n5021) );
  BUFX2 U633 ( .A(n3284), .Y(n5022) );
  BUFX2 U634 ( .A(n3277), .Y(n5023) );
  BUFX2 U635 ( .A(n3269), .Y(n5024) );
  BUFX2 U636 ( .A(n3261), .Y(n5025) );
  BUFX2 U637 ( .A(n3247), .Y(n5026) );
  BUFX2 U638 ( .A(n3240), .Y(n5027) );
  BUFX2 U639 ( .A(n3233), .Y(n5028) );
  BUFX2 U640 ( .A(n3226), .Y(n5029) );
  BUFX2 U641 ( .A(n3213), .Y(n5030) );
  BUFX2 U642 ( .A(n3206), .Y(n5031) );
  BUFX2 U643 ( .A(n3199), .Y(n5032) );
  BUFX2 U644 ( .A(n3192), .Y(n5033) );
  BUFX2 U645 ( .A(n3179), .Y(n5034) );
  BUFX2 U646 ( .A(n3172), .Y(n5035) );
  BUFX2 U647 ( .A(n3165), .Y(n5036) );
  BUFX2 U648 ( .A(n3158), .Y(n5037) );
  BUFX2 U649 ( .A(n3145), .Y(n5038) );
  BUFX2 U650 ( .A(n3138), .Y(n5039) );
  BUFX2 U651 ( .A(n3131), .Y(n5040) );
  BUFX2 U652 ( .A(n3124), .Y(n5041) );
  BUFX2 U653 ( .A(n3111), .Y(n5042) );
  BUFX2 U654 ( .A(n3104), .Y(n5043) );
  BUFX2 U655 ( .A(n3097), .Y(n5044) );
  BUFX2 U656 ( .A(n3090), .Y(n5045) );
  BUFX2 U657 ( .A(n3077), .Y(n5046) );
  BUFX2 U658 ( .A(n3070), .Y(n5047) );
  BUFX2 U659 ( .A(n3063), .Y(n5048) );
  BUFX2 U660 ( .A(n3056), .Y(n5049) );
  BUFX2 U661 ( .A(n3043), .Y(n5050) );
  BUFX2 U662 ( .A(n3036), .Y(n5051) );
  BUFX2 U663 ( .A(n3029), .Y(n5052) );
  BUFX2 U664 ( .A(n3022), .Y(n5053) );
  BUFX2 U665 ( .A(n3009), .Y(n5054) );
  BUFX2 U666 ( .A(n3002), .Y(n5055) );
  BUFX2 U667 ( .A(n2995), .Y(n5056) );
  BUFX2 U668 ( .A(n2988), .Y(n5057) );
  BUFX2 U669 ( .A(n2975), .Y(n5058) );
  BUFX2 U670 ( .A(n2968), .Y(n5059) );
  BUFX2 U671 ( .A(n2961), .Y(n5060) );
  BUFX2 U672 ( .A(n2954), .Y(n5061) );
  BUFX2 U673 ( .A(n2941), .Y(n5062) );
  BUFX2 U674 ( .A(n2934), .Y(n5063) );
  BUFX2 U675 ( .A(n2927), .Y(n5064) );
  BUFX2 U676 ( .A(n2920), .Y(n5065) );
  BUFX2 U677 ( .A(n2907), .Y(n5066) );
  BUFX2 U678 ( .A(n2900), .Y(n5067) );
  BUFX2 U679 ( .A(n2893), .Y(n5068) );
  BUFX2 U680 ( .A(n2886), .Y(n5069) );
  BUFX2 U681 ( .A(n2873), .Y(n5070) );
  BUFX2 U682 ( .A(n2866), .Y(n5071) );
  BUFX2 U683 ( .A(n2859), .Y(n5072) );
  BUFX2 U684 ( .A(n2852), .Y(n5073) );
  BUFX2 U685 ( .A(n2839), .Y(n5074) );
  BUFX2 U686 ( .A(n2832), .Y(n5075) );
  BUFX2 U687 ( .A(n2825), .Y(n5076) );
  BUFX2 U688 ( .A(n2818), .Y(n5077) );
  BUFX2 U689 ( .A(n2805), .Y(n5078) );
  BUFX2 U690 ( .A(n2798), .Y(n5079) );
  BUFX2 U691 ( .A(n2791), .Y(n5080) );
  BUFX2 U692 ( .A(n2784), .Y(n5081) );
  BUFX2 U693 ( .A(n2771), .Y(n5082) );
  BUFX2 U694 ( .A(n2764), .Y(n5083) );
  BUFX2 U695 ( .A(n2757), .Y(n5084) );
  BUFX2 U696 ( .A(n2750), .Y(n5085) );
  BUFX2 U697 ( .A(n2737), .Y(n5086) );
  BUFX2 U698 ( .A(n2730), .Y(n5087) );
  BUFX2 U699 ( .A(n2723), .Y(n5088) );
  BUFX2 U700 ( .A(n2716), .Y(n5089) );
  BUFX2 U701 ( .A(n2703), .Y(n5090) );
  BUFX2 U702 ( .A(n2696), .Y(n5091) );
  BUFX2 U703 ( .A(n2689), .Y(n5092) );
  BUFX2 U704 ( .A(n2682), .Y(n5093) );
  BUFX2 U705 ( .A(n2669), .Y(n5094) );
  BUFX2 U706 ( .A(n2662), .Y(n5095) );
  BUFX2 U707 ( .A(n2655), .Y(n5096) );
  BUFX2 U708 ( .A(n2648), .Y(n5097) );
  BUFX2 U709 ( .A(n2635), .Y(n5098) );
  BUFX2 U710 ( .A(n2628), .Y(n5099) );
  BUFX2 U711 ( .A(n2621), .Y(n5100) );
  BUFX2 U712 ( .A(n2614), .Y(n5101) );
  BUFX2 U713 ( .A(n1535), .Y(n5102) );
  BUFX2 U714 ( .A(n1528), .Y(n5103) );
  BUFX2 U715 ( .A(n1521), .Y(n5104) );
  BUFX2 U716 ( .A(n1514), .Y(n5105) );
  BUFX2 U717 ( .A(n1501), .Y(n5106) );
  BUFX2 U718 ( .A(n1494), .Y(n5107) );
  BUFX2 U719 ( .A(n1487), .Y(n5108) );
  BUFX2 U720 ( .A(n1480), .Y(n5109) );
  BUFX2 U721 ( .A(n1467), .Y(n5110) );
  BUFX2 U722 ( .A(n1460), .Y(n5111) );
  BUFX2 U723 ( .A(n1453), .Y(n5112) );
  BUFX2 U724 ( .A(n1446), .Y(n5113) );
  BUFX2 U725 ( .A(n1433), .Y(n5114) );
  BUFX2 U726 ( .A(n1426), .Y(n5115) );
  BUFX2 U727 ( .A(n1419), .Y(n5116) );
  BUFX2 U728 ( .A(n1412), .Y(n5117) );
  BUFX2 U729 ( .A(n1399), .Y(n5118) );
  BUFX2 U730 ( .A(n1392), .Y(n5119) );
  BUFX2 U731 ( .A(n1385), .Y(n5120) );
  BUFX2 U732 ( .A(n1378), .Y(n5121) );
  BUFX2 U733 ( .A(n1365), .Y(n5122) );
  BUFX2 U734 ( .A(n1358), .Y(n5123) );
  BUFX2 U735 ( .A(n1351), .Y(n5124) );
  BUFX2 U736 ( .A(n1344), .Y(n5125) );
  BUFX2 U737 ( .A(n1331), .Y(n5126) );
  BUFX2 U738 ( .A(n1324), .Y(n5127) );
  BUFX2 U739 ( .A(n1317), .Y(n5128) );
  BUFX2 U740 ( .A(n1310), .Y(n5129) );
  BUFX2 U741 ( .A(n1297), .Y(n5130) );
  BUFX2 U742 ( .A(n1290), .Y(n5131) );
  BUFX2 U743 ( .A(n1283), .Y(n5132) );
  BUFX2 U744 ( .A(n1276), .Y(n5133) );
  BUFX2 U745 ( .A(n1263), .Y(n5134) );
  BUFX2 U746 ( .A(n1256), .Y(n5135) );
  BUFX2 U747 ( .A(n1249), .Y(n5136) );
  BUFX2 U748 ( .A(n1242), .Y(n5137) );
  BUFX2 U749 ( .A(n1229), .Y(n5138) );
  BUFX2 U750 ( .A(n1222), .Y(n5139) );
  BUFX2 U751 ( .A(n1215), .Y(n5140) );
  BUFX2 U752 ( .A(n1208), .Y(n5141) );
  BUFX2 U753 ( .A(n1195), .Y(n5142) );
  BUFX2 U754 ( .A(n1188), .Y(n5143) );
  BUFX2 U755 ( .A(n1181), .Y(n5144) );
  BUFX2 U756 ( .A(n1174), .Y(n5145) );
  BUFX2 U757 ( .A(n1161), .Y(n5146) );
  BUFX2 U758 ( .A(n1154), .Y(n5147) );
  BUFX2 U759 ( .A(n1147), .Y(n5148) );
  BUFX2 U760 ( .A(n1140), .Y(n5149) );
  BUFX2 U761 ( .A(n1127), .Y(n5150) );
  BUFX2 U762 ( .A(n1119), .Y(n5151) );
  BUFX2 U763 ( .A(n1111), .Y(n5152) );
  BUFX2 U764 ( .A(n1098), .Y(n5153) );
  AND2X1 U765 ( .A(n1124), .B(n6810), .Y(n3296) );
  INVX1 U766 ( .A(n3296), .Y(n5154) );
  AND2X1 U767 ( .A(data_out[0]), .B(n3299), .Y(n3250) );
  INVX1 U768 ( .A(n3250), .Y(n5155) );
  AND2X1 U769 ( .A(data_out[1]), .B(n3299), .Y(n3216) );
  INVX1 U770 ( .A(n3216), .Y(n5156) );
  AND2X1 U771 ( .A(data_out[2]), .B(n3299), .Y(n3182) );
  INVX1 U772 ( .A(n3182), .Y(n5157) );
  AND2X1 U773 ( .A(data_out[3]), .B(n3299), .Y(n3148) );
  INVX1 U774 ( .A(n3148), .Y(n5158) );
  AND2X1 U775 ( .A(data_out[4]), .B(n3299), .Y(n3114) );
  INVX1 U776 ( .A(n3114), .Y(n5159) );
  AND2X1 U777 ( .A(data_out[5]), .B(n3299), .Y(n3080) );
  INVX1 U778 ( .A(n3080), .Y(n5160) );
  AND2X1 U779 ( .A(data_out[6]), .B(n3299), .Y(n3046) );
  INVX1 U780 ( .A(n3046), .Y(n5161) );
  AND2X1 U781 ( .A(data_out[7]), .B(n3299), .Y(n3012) );
  INVX1 U782 ( .A(n3012), .Y(n5162) );
  AND2X1 U783 ( .A(data_out[8]), .B(n3299), .Y(n2978) );
  INVX1 U784 ( .A(n2978), .Y(n5163) );
  AND2X1 U785 ( .A(data_out[9]), .B(n3299), .Y(n2944) );
  INVX1 U786 ( .A(n2944), .Y(n5164) );
  AND2X1 U787 ( .A(data_out[10]), .B(n3299), .Y(n2910) );
  INVX1 U788 ( .A(n2910), .Y(n5165) );
  AND2X1 U789 ( .A(data_out[11]), .B(n3299), .Y(n2876) );
  INVX1 U790 ( .A(n2876), .Y(n5166) );
  AND2X1 U791 ( .A(data_out[24]), .B(n3299), .Y(n2842) );
  INVX1 U792 ( .A(n2842), .Y(n5167) );
  AND2X1 U793 ( .A(data_out[26]), .B(n3299), .Y(n2808) );
  INVX1 U794 ( .A(n2808), .Y(n5168) );
  AND2X1 U795 ( .A(data_out[28]), .B(n3299), .Y(n2774) );
  INVX1 U796 ( .A(n2774), .Y(n5169) );
  AND2X1 U797 ( .A(data_out[30]), .B(n3299), .Y(n2740) );
  INVX1 U798 ( .A(n2740), .Y(n5170) );
  AND2X1 U799 ( .A(data_out[32]), .B(n3299), .Y(n2706) );
  INVX1 U800 ( .A(n2706), .Y(n5171) );
  AND2X1 U801 ( .A(data_out[12]), .B(n3299), .Y(n2672) );
  INVX1 U802 ( .A(n2672), .Y(n5172) );
  AND2X1 U803 ( .A(data_out[13]), .B(n3299), .Y(n2638) );
  INVX1 U804 ( .A(n2638), .Y(n5173) );
  AND2X1 U805 ( .A(data_out[14]), .B(n3299), .Y(n2604) );
  INVX1 U806 ( .A(n2604), .Y(n5174) );
  AND2X1 U807 ( .A(data_out[15]), .B(n3299), .Y(n1504) );
  INVX1 U808 ( .A(n1504), .Y(n5175) );
  AND2X1 U809 ( .A(data_out[16]), .B(n3299), .Y(n1470) );
  INVX1 U810 ( .A(n1470), .Y(n5176) );
  AND2X1 U811 ( .A(data_out[17]), .B(n3299), .Y(n1436) );
  INVX1 U812 ( .A(n1436), .Y(n5177) );
  AND2X1 U813 ( .A(data_out[18]), .B(n3299), .Y(n1402) );
  INVX1 U814 ( .A(n1402), .Y(n5178) );
  AND2X1 U815 ( .A(data_out[19]), .B(n3299), .Y(n1368) );
  INVX1 U816 ( .A(n1368), .Y(n5179) );
  AND2X1 U817 ( .A(data_out[20]), .B(n3299), .Y(n1334) );
  INVX1 U818 ( .A(n1334), .Y(n5180) );
  AND2X1 U819 ( .A(data_out[21]), .B(n3299), .Y(n1300) );
  INVX1 U820 ( .A(n1300), .Y(n5181) );
  AND2X1 U821 ( .A(data_out[22]), .B(n3299), .Y(n1266) );
  INVX1 U822 ( .A(n1266), .Y(n5182) );
  AND2X1 U823 ( .A(data_out[23]), .B(n3299), .Y(n1232) );
  INVX1 U824 ( .A(n1232), .Y(n5183) );
  AND2X1 U825 ( .A(data_out[25]), .B(n3299), .Y(n1198) );
  INVX1 U826 ( .A(n1198), .Y(n5184) );
  AND2X1 U827 ( .A(data_out[27]), .B(n3299), .Y(n1164) );
  INVX1 U828 ( .A(n1164), .Y(n5185) );
  AND2X1 U829 ( .A(data_out[29]), .B(n3299), .Y(n1130) );
  INVX1 U830 ( .A(n1130), .Y(n5186) );
  AND2X1 U831 ( .A(data_out[31]), .B(n3299), .Y(n1086) );
  INVX1 U832 ( .A(n1086), .Y(n5187) );
  BUFX2 U833 ( .A(n3304), .Y(n5188) );
  AND2X1 U834 ( .A(n6822), .B(n7520), .Y(n3285) );
  INVX1 U835 ( .A(n3285), .Y(n5189) );
  AND2X1 U836 ( .A(n6810), .B(n7421), .Y(n3282) );
  INVX1 U837 ( .A(n3282), .Y(n5190) );
  AND2X1 U838 ( .A(n6822), .B(n7784), .Y(n3278) );
  INVX1 U839 ( .A(n3278), .Y(n5191) );
  AND2X1 U840 ( .A(n6811), .B(n7685), .Y(n3274) );
  INVX1 U841 ( .A(n3274), .Y(n5192) );
  AND2X1 U842 ( .A(n6822), .B(n6992), .Y(n3270) );
  INVX1 U843 ( .A(n3270), .Y(n5193) );
  AND2X1 U844 ( .A(n6810), .B(n6893), .Y(n3266) );
  INVX1 U845 ( .A(n3266), .Y(n5194) );
  AND2X1 U846 ( .A(n6822), .B(n7256), .Y(n3262) );
  INVX1 U847 ( .A(n3262), .Y(n5195) );
  AND2X1 U848 ( .A(n6810), .B(n7157), .Y(n3258) );
  INVX1 U849 ( .A(n3258), .Y(n5196) );
  AND2X1 U850 ( .A(n6822), .B(n7519), .Y(n3248) );
  INVX1 U851 ( .A(n3248), .Y(n5197) );
  AND2X1 U852 ( .A(n6811), .B(n7420), .Y(n3245) );
  INVX1 U853 ( .A(n3245), .Y(n5198) );
  AND2X1 U854 ( .A(n6822), .B(n7783), .Y(n3241) );
  INVX1 U855 ( .A(n3241), .Y(n5199) );
  AND2X1 U856 ( .A(n6811), .B(n7684), .Y(n3238) );
  INVX1 U857 ( .A(n3238), .Y(n5200) );
  AND2X1 U858 ( .A(n6822), .B(n6991), .Y(n3234) );
  INVX1 U859 ( .A(n3234), .Y(n5201) );
  AND2X1 U860 ( .A(n6811), .B(n6892), .Y(n3231) );
  INVX1 U861 ( .A(n3231), .Y(n5202) );
  AND2X1 U862 ( .A(n6822), .B(n7255), .Y(n3227) );
  INVX1 U863 ( .A(n3227), .Y(n5203) );
  AND2X1 U864 ( .A(n6811), .B(n7156), .Y(n3224) );
  INVX1 U865 ( .A(n3224), .Y(n5204) );
  AND2X1 U866 ( .A(n6822), .B(n7518), .Y(n3214) );
  INVX1 U867 ( .A(n3214), .Y(n5205) );
  AND2X1 U868 ( .A(n6811), .B(n7419), .Y(n3211) );
  INVX1 U869 ( .A(n3211), .Y(n5206) );
  AND2X1 U870 ( .A(n6822), .B(n7782), .Y(n3207) );
  INVX1 U871 ( .A(n3207), .Y(n5207) );
  AND2X1 U872 ( .A(n6811), .B(n7683), .Y(n3204) );
  INVX1 U873 ( .A(n3204), .Y(n5208) );
  AND2X1 U874 ( .A(n6822), .B(n6990), .Y(n3200) );
  INVX1 U875 ( .A(n3200), .Y(n5209) );
  AND2X1 U876 ( .A(n6810), .B(n6891), .Y(n3197) );
  INVX1 U877 ( .A(n3197), .Y(n5210) );
  AND2X1 U878 ( .A(n6822), .B(n7254), .Y(n3193) );
  INVX1 U879 ( .A(n3193), .Y(n5211) );
  AND2X1 U880 ( .A(n6811), .B(n7155), .Y(n3190) );
  INVX1 U881 ( .A(n3190), .Y(n5212) );
  AND2X1 U882 ( .A(n6821), .B(n7517), .Y(n3180) );
  INVX1 U883 ( .A(n3180), .Y(n5213) );
  AND2X1 U884 ( .A(n6811), .B(n7418), .Y(n3177) );
  INVX1 U885 ( .A(n3177), .Y(n5214) );
  AND2X1 U886 ( .A(n6821), .B(n7781), .Y(n3173) );
  INVX1 U887 ( .A(n3173), .Y(n5215) );
  AND2X1 U888 ( .A(n6811), .B(n7682), .Y(n3170) );
  INVX1 U889 ( .A(n3170), .Y(n5216) );
  AND2X1 U890 ( .A(n6821), .B(n6989), .Y(n3166) );
  INVX1 U891 ( .A(n3166), .Y(n5217) );
  AND2X1 U892 ( .A(n6811), .B(n6890), .Y(n3163) );
  INVX1 U893 ( .A(n3163), .Y(n5218) );
  AND2X1 U894 ( .A(n6821), .B(n7253), .Y(n3159) );
  INVX1 U895 ( .A(n3159), .Y(n5219) );
  AND2X1 U896 ( .A(n6811), .B(n7154), .Y(n3156) );
  INVX1 U897 ( .A(n3156), .Y(n5220) );
  AND2X1 U898 ( .A(n6821), .B(n7516), .Y(n3146) );
  INVX1 U899 ( .A(n3146), .Y(n5221) );
  AND2X1 U900 ( .A(n6811), .B(n7417), .Y(n3143) );
  INVX1 U901 ( .A(n3143), .Y(n5222) );
  AND2X1 U902 ( .A(n6821), .B(n7780), .Y(n3139) );
  INVX1 U903 ( .A(n3139), .Y(n5223) );
  AND2X1 U904 ( .A(n6811), .B(n7681), .Y(n3136) );
  INVX1 U905 ( .A(n3136), .Y(n5224) );
  AND2X1 U906 ( .A(n6821), .B(n6988), .Y(n3132) );
  INVX1 U907 ( .A(n3132), .Y(n5225) );
  AND2X1 U908 ( .A(n6811), .B(n6889), .Y(n3129) );
  INVX1 U909 ( .A(n3129), .Y(n5226) );
  AND2X1 U910 ( .A(n6821), .B(n7252), .Y(n3125) );
  INVX1 U911 ( .A(n3125), .Y(n5227) );
  AND2X1 U912 ( .A(n6811), .B(n7153), .Y(n3122) );
  INVX1 U913 ( .A(n3122), .Y(n5228) );
  AND2X1 U914 ( .A(n6821), .B(n7515), .Y(n3112) );
  INVX1 U915 ( .A(n3112), .Y(n5229) );
  AND2X1 U916 ( .A(n6811), .B(n7416), .Y(n3109) );
  INVX1 U917 ( .A(n3109), .Y(n5230) );
  AND2X1 U918 ( .A(n6821), .B(n7779), .Y(n3105) );
  INVX1 U919 ( .A(n3105), .Y(n5231) );
  AND2X1 U920 ( .A(n6811), .B(n7680), .Y(n3102) );
  INVX1 U921 ( .A(n3102), .Y(n5232) );
  AND2X1 U922 ( .A(n6821), .B(n6987), .Y(n3098) );
  INVX1 U923 ( .A(n3098), .Y(n5233) );
  AND2X1 U924 ( .A(n6811), .B(n6888), .Y(n3095) );
  INVX1 U925 ( .A(n3095), .Y(n5234) );
  AND2X1 U926 ( .A(n6821), .B(n7251), .Y(n3091) );
  INVX1 U927 ( .A(n3091), .Y(n5235) );
  AND2X1 U928 ( .A(n6811), .B(n7152), .Y(n3088) );
  INVX1 U929 ( .A(n3088), .Y(n5236) );
  AND2X1 U930 ( .A(n6820), .B(n7514), .Y(n3078) );
  INVX1 U931 ( .A(n3078), .Y(n5237) );
  AND2X1 U932 ( .A(n6811), .B(n7415), .Y(n3075) );
  INVX1 U933 ( .A(n3075), .Y(n5238) );
  AND2X1 U934 ( .A(n6820), .B(n7778), .Y(n3071) );
  INVX1 U935 ( .A(n3071), .Y(n5239) );
  AND2X1 U936 ( .A(n6811), .B(n7679), .Y(n3068) );
  INVX1 U937 ( .A(n3068), .Y(n5240) );
  AND2X1 U938 ( .A(n6820), .B(n6986), .Y(n3064) );
  INVX1 U939 ( .A(n3064), .Y(n5241) );
  AND2X1 U940 ( .A(n6811), .B(n6887), .Y(n3061) );
  INVX1 U941 ( .A(n3061), .Y(n5242) );
  AND2X1 U942 ( .A(n6820), .B(n7250), .Y(n3057) );
  INVX1 U943 ( .A(n3057), .Y(n5243) );
  AND2X1 U944 ( .A(n6811), .B(n7151), .Y(n3054) );
  INVX1 U945 ( .A(n3054), .Y(n5244) );
  AND2X1 U946 ( .A(n6820), .B(n7513), .Y(n3044) );
  INVX1 U947 ( .A(n3044), .Y(n5245) );
  AND2X1 U948 ( .A(n6811), .B(n7414), .Y(n3041) );
  INVX1 U949 ( .A(n3041), .Y(n5246) );
  AND2X1 U950 ( .A(n6820), .B(n7777), .Y(n3037) );
  INVX1 U951 ( .A(n3037), .Y(n5247) );
  AND2X1 U952 ( .A(n6811), .B(n7678), .Y(n3034) );
  INVX1 U953 ( .A(n3034), .Y(n5248) );
  AND2X1 U954 ( .A(n6820), .B(n6985), .Y(n3030) );
  INVX1 U955 ( .A(n3030), .Y(n5249) );
  AND2X1 U956 ( .A(n6811), .B(n6886), .Y(n3027) );
  INVX1 U957 ( .A(n3027), .Y(n5250) );
  AND2X1 U958 ( .A(n6820), .B(n7249), .Y(n3023) );
  INVX1 U959 ( .A(n3023), .Y(n5251) );
  AND2X1 U960 ( .A(n6811), .B(n7150), .Y(n3020) );
  INVX1 U961 ( .A(n3020), .Y(n5252) );
  AND2X1 U962 ( .A(n6820), .B(n7512), .Y(n3010) );
  INVX1 U963 ( .A(n3010), .Y(n5253) );
  AND2X1 U964 ( .A(n6811), .B(n7413), .Y(n3007) );
  INVX1 U965 ( .A(n3007), .Y(n5254) );
  AND2X1 U966 ( .A(n6820), .B(n7776), .Y(n3003) );
  INVX1 U967 ( .A(n3003), .Y(n5255) );
  AND2X1 U968 ( .A(n6810), .B(n7677), .Y(n3000) );
  INVX1 U969 ( .A(n3000), .Y(n5256) );
  AND2X1 U970 ( .A(n6820), .B(n6984), .Y(n2996) );
  INVX1 U971 ( .A(n2996), .Y(n5257) );
  AND2X1 U972 ( .A(n6810), .B(n6885), .Y(n2993) );
  INVX1 U973 ( .A(n2993), .Y(n5258) );
  AND2X1 U974 ( .A(n6820), .B(n7248), .Y(n2989) );
  INVX1 U975 ( .A(n2989), .Y(n5259) );
  AND2X1 U976 ( .A(n6810), .B(n7149), .Y(n2986) );
  INVX1 U977 ( .A(n2986), .Y(n5260) );
  AND2X1 U978 ( .A(n6820), .B(n7511), .Y(n2976) );
  INVX1 U979 ( .A(n2976), .Y(n5261) );
  AND2X1 U980 ( .A(n6810), .B(n7412), .Y(n2973) );
  INVX1 U981 ( .A(n2973), .Y(n5262) );
  AND2X1 U982 ( .A(n6822), .B(n7775), .Y(n2969) );
  INVX1 U983 ( .A(n2969), .Y(n5263) );
  AND2X1 U984 ( .A(n6811), .B(n7676), .Y(n2966) );
  INVX1 U985 ( .A(n2966), .Y(n5264) );
  AND2X1 U986 ( .A(n6820), .B(n6983), .Y(n2962) );
  INVX1 U987 ( .A(n2962), .Y(n5265) );
  AND2X1 U988 ( .A(n6811), .B(n6884), .Y(n2959) );
  INVX1 U989 ( .A(n2959), .Y(n5266) );
  AND2X1 U990 ( .A(n6822), .B(n7247), .Y(n2955) );
  INVX1 U991 ( .A(n2955), .Y(n5267) );
  AND2X1 U992 ( .A(n6811), .B(n7148), .Y(n2952) );
  INVX1 U993 ( .A(n2952), .Y(n5268) );
  AND2X1 U994 ( .A(n6821), .B(n7510), .Y(n2942) );
  INVX1 U995 ( .A(n2942), .Y(n5269) );
  AND2X1 U996 ( .A(n6811), .B(n7411), .Y(n2939) );
  INVX1 U997 ( .A(n2939), .Y(n5270) );
  AND2X1 U998 ( .A(n6820), .B(n7774), .Y(n2935) );
  INVX1 U999 ( .A(n2935), .Y(n5271) );
  AND2X1 U1000 ( .A(n6810), .B(n7675), .Y(n2932) );
  INVX1 U1001 ( .A(n2932), .Y(n5272) );
  AND2X1 U1002 ( .A(n6821), .B(n6982), .Y(n2928) );
  INVX1 U1003 ( .A(n2928), .Y(n5273) );
  AND2X1 U1004 ( .A(n6810), .B(n6883), .Y(n2925) );
  INVX1 U1005 ( .A(n2925), .Y(n5274) );
  AND2X1 U1006 ( .A(n6820), .B(n7246), .Y(n2921) );
  INVX1 U1007 ( .A(n2921), .Y(n5275) );
  AND2X1 U1008 ( .A(n6810), .B(n7147), .Y(n2918) );
  INVX1 U1009 ( .A(n2918), .Y(n5276) );
  AND2X1 U1010 ( .A(n6822), .B(n7509), .Y(n2908) );
  INVX1 U1011 ( .A(n2908), .Y(n5277) );
  AND2X1 U1012 ( .A(n6810), .B(n7410), .Y(n2905) );
  INVX1 U1013 ( .A(n2905), .Y(n5278) );
  AND2X1 U1014 ( .A(n6821), .B(n7773), .Y(n2901) );
  INVX1 U1015 ( .A(n2901), .Y(n5279) );
  AND2X1 U1016 ( .A(n6811), .B(n7674), .Y(n2898) );
  INVX1 U1017 ( .A(n2898), .Y(n5280) );
  AND2X1 U1018 ( .A(n6822), .B(n6981), .Y(n2894) );
  INVX1 U1019 ( .A(n2894), .Y(n5281) );
  AND2X1 U1020 ( .A(n6811), .B(n6882), .Y(n2891) );
  INVX1 U1021 ( .A(n2891), .Y(n5282) );
  AND2X1 U1022 ( .A(n6821), .B(n7245), .Y(n2887) );
  INVX1 U1023 ( .A(n2887), .Y(n5283) );
  AND2X1 U1024 ( .A(n6811), .B(n7146), .Y(n2884) );
  INVX1 U1025 ( .A(n2884), .Y(n5284) );
  AND2X1 U1026 ( .A(n6821), .B(n7496), .Y(n2874) );
  INVX1 U1027 ( .A(n2874), .Y(n5285) );
  AND2X1 U1028 ( .A(n6810), .B(n7397), .Y(n2871) );
  INVX1 U1029 ( .A(n2871), .Y(n5286) );
  AND2X1 U1030 ( .A(n6820), .B(n7760), .Y(n2867) );
  INVX1 U1031 ( .A(n2867), .Y(n5287) );
  AND2X1 U1032 ( .A(n6810), .B(n7661), .Y(n2864) );
  INVX1 U1033 ( .A(n2864), .Y(n5288) );
  AND2X1 U1034 ( .A(n6822), .B(n6968), .Y(n2860) );
  INVX1 U1035 ( .A(n2860), .Y(n5289) );
  AND2X1 U1036 ( .A(n6810), .B(n6869), .Y(n2857) );
  INVX1 U1037 ( .A(n2857), .Y(n5290) );
  AND2X1 U1038 ( .A(n6820), .B(n7232), .Y(n2853) );
  INVX1 U1039 ( .A(n2853), .Y(n5291) );
  AND2X1 U1040 ( .A(n6810), .B(n7133), .Y(n2850) );
  INVX1 U1041 ( .A(n2850), .Y(n5292) );
  AND2X1 U1042 ( .A(n6822), .B(n7494), .Y(n2840) );
  INVX1 U1043 ( .A(n2840), .Y(n5293) );
  AND2X1 U1044 ( .A(n6810), .B(n7395), .Y(n2837) );
  INVX1 U1045 ( .A(n2837), .Y(n5294) );
  AND2X1 U1046 ( .A(n6820), .B(n7758), .Y(n2833) );
  INVX1 U1047 ( .A(n2833), .Y(n5295) );
  AND2X1 U1048 ( .A(n6810), .B(n7659), .Y(n2830) );
  INVX1 U1049 ( .A(n2830), .Y(n5296) );
  AND2X1 U1050 ( .A(n6822), .B(n6966), .Y(n2826) );
  INVX1 U1051 ( .A(n2826), .Y(n5297) );
  AND2X1 U1052 ( .A(n6810), .B(n6867), .Y(n2823) );
  INVX1 U1053 ( .A(n2823), .Y(n5298) );
  AND2X1 U1054 ( .A(n6822), .B(n7230), .Y(n2819) );
  INVX1 U1055 ( .A(n2819), .Y(n5299) );
  AND2X1 U1056 ( .A(n6810), .B(n7131), .Y(n2816) );
  INVX1 U1057 ( .A(n2816), .Y(n5300) );
  AND2X1 U1058 ( .A(n6822), .B(n7492), .Y(n2806) );
  INVX1 U1059 ( .A(n2806), .Y(n5301) );
  AND2X1 U1060 ( .A(n6810), .B(n7393), .Y(n2803) );
  INVX1 U1061 ( .A(n2803), .Y(n5302) );
  AND2X1 U1062 ( .A(n6821), .B(n7756), .Y(n2799) );
  INVX1 U1063 ( .A(n2799), .Y(n5303) );
  AND2X1 U1064 ( .A(n6810), .B(n7657), .Y(n2796) );
  INVX1 U1065 ( .A(n2796), .Y(n5304) );
  AND2X1 U1066 ( .A(n6820), .B(n6964), .Y(n2792) );
  INVX1 U1067 ( .A(n2792), .Y(n5305) );
  AND2X1 U1068 ( .A(n6810), .B(n6865), .Y(n2789) );
  INVX1 U1069 ( .A(n2789), .Y(n5306) );
  AND2X1 U1070 ( .A(n6820), .B(n7228), .Y(n2785) );
  INVX1 U1071 ( .A(n2785), .Y(n5307) );
  AND2X1 U1072 ( .A(n6810), .B(n7129), .Y(n2782) );
  INVX1 U1073 ( .A(n2782), .Y(n5308) );
  AND2X1 U1074 ( .A(n6820), .B(n7490), .Y(n2772) );
  INVX1 U1075 ( .A(n2772), .Y(n5309) );
  AND2X1 U1076 ( .A(n6810), .B(n7391), .Y(n2769) );
  INVX1 U1077 ( .A(n2769), .Y(n5310) );
  AND2X1 U1078 ( .A(n6821), .B(n7754), .Y(n2765) );
  INVX1 U1079 ( .A(n2765), .Y(n5311) );
  AND2X1 U1080 ( .A(n6810), .B(n7655), .Y(n2762) );
  INVX1 U1081 ( .A(n2762), .Y(n5312) );
  AND2X1 U1082 ( .A(n6822), .B(n6962), .Y(n2758) );
  INVX1 U1083 ( .A(n2758), .Y(n5313) );
  AND2X1 U1084 ( .A(n6810), .B(n6863), .Y(n2755) );
  INVX1 U1085 ( .A(n2755), .Y(n5314) );
  AND2X1 U1086 ( .A(n6822), .B(n7226), .Y(n2751) );
  INVX1 U1087 ( .A(n2751), .Y(n5315) );
  AND2X1 U1088 ( .A(n6810), .B(n7127), .Y(n2748) );
  INVX1 U1089 ( .A(n2748), .Y(n5316) );
  AND2X1 U1090 ( .A(n6821), .B(n7488), .Y(n2738) );
  INVX1 U1091 ( .A(n2738), .Y(n5317) );
  AND2X1 U1092 ( .A(n6810), .B(n7389), .Y(n2735) );
  INVX1 U1093 ( .A(n2735), .Y(n5318) );
  AND2X1 U1094 ( .A(n6822), .B(n7752), .Y(n2731) );
  INVX1 U1095 ( .A(n2731), .Y(n5319) );
  AND2X1 U1096 ( .A(n6810), .B(n7653), .Y(n2728) );
  INVX1 U1097 ( .A(n2728), .Y(n5320) );
  AND2X1 U1098 ( .A(n6820), .B(n6960), .Y(n2724) );
  INVX1 U1099 ( .A(n2724), .Y(n5321) );
  AND2X1 U1100 ( .A(n6811), .B(n6861), .Y(n2721) );
  INVX1 U1101 ( .A(n2721), .Y(n5322) );
  AND2X1 U1102 ( .A(n6821), .B(n7224), .Y(n2717) );
  INVX1 U1103 ( .A(n2717), .Y(n5323) );
  AND2X1 U1104 ( .A(n6810), .B(n7125), .Y(n2714) );
  INVX1 U1105 ( .A(n2714), .Y(n5324) );
  AND2X1 U1106 ( .A(n6822), .B(n7508), .Y(n2704) );
  INVX1 U1107 ( .A(n2704), .Y(n5325) );
  AND2X1 U1108 ( .A(n6810), .B(n7409), .Y(n2701) );
  INVX1 U1109 ( .A(n2701), .Y(n5326) );
  AND2X1 U1110 ( .A(n6821), .B(n7772), .Y(n2697) );
  INVX1 U1111 ( .A(n2697), .Y(n5327) );
  AND2X1 U1112 ( .A(n6810), .B(n7673), .Y(n2694) );
  INVX1 U1113 ( .A(n2694), .Y(n5328) );
  AND2X1 U1114 ( .A(n6821), .B(n6980), .Y(n2690) );
  INVX1 U1115 ( .A(n2690), .Y(n5329) );
  AND2X1 U1116 ( .A(n6811), .B(n6881), .Y(n2687) );
  INVX1 U1117 ( .A(n2687), .Y(n5330) );
  AND2X1 U1118 ( .A(n6821), .B(n7244), .Y(n2683) );
  INVX1 U1119 ( .A(n2683), .Y(n5331) );
  AND2X1 U1120 ( .A(n6811), .B(n7145), .Y(n2680) );
  INVX1 U1121 ( .A(n2680), .Y(n5332) );
  AND2X1 U1122 ( .A(n1103), .B(n7507), .Y(n2670) );
  INVX1 U1123 ( .A(n2670), .Y(n5333) );
  AND2X1 U1124 ( .A(n6810), .B(n7408), .Y(n2667) );
  INVX1 U1125 ( .A(n2667), .Y(n5334) );
  AND2X1 U1126 ( .A(n1103), .B(n7771), .Y(n2663) );
  INVX1 U1127 ( .A(n2663), .Y(n5335) );
  AND2X1 U1128 ( .A(n6811), .B(n7672), .Y(n2660) );
  INVX1 U1129 ( .A(n2660), .Y(n5336) );
  AND2X1 U1130 ( .A(n1103), .B(n6979), .Y(n2656) );
  INVX1 U1131 ( .A(n2656), .Y(n5337) );
  AND2X1 U1132 ( .A(n6811), .B(n6880), .Y(n2653) );
  INVX1 U1133 ( .A(n2653), .Y(n5338) );
  AND2X1 U1134 ( .A(n1103), .B(n7243), .Y(n2649) );
  INVX1 U1135 ( .A(n2649), .Y(n5339) );
  AND2X1 U1136 ( .A(n6811), .B(n7144), .Y(n2646) );
  INVX1 U1137 ( .A(n2646), .Y(n5340) );
  AND2X1 U1138 ( .A(n1103), .B(n7506), .Y(n2636) );
  INVX1 U1139 ( .A(n2636), .Y(n5341) );
  AND2X1 U1140 ( .A(n6811), .B(n7407), .Y(n2633) );
  INVX1 U1141 ( .A(n2633), .Y(n5342) );
  AND2X1 U1142 ( .A(n1103), .B(n7770), .Y(n2629) );
  INVX1 U1143 ( .A(n2629), .Y(n5343) );
  AND2X1 U1144 ( .A(n6811), .B(n7671), .Y(n2626) );
  INVX1 U1145 ( .A(n2626), .Y(n5344) );
  AND2X1 U1146 ( .A(n1103), .B(n6978), .Y(n2622) );
  INVX1 U1147 ( .A(n2622), .Y(n5345) );
  AND2X1 U1148 ( .A(n6810), .B(n6879), .Y(n2619) );
  INVX1 U1149 ( .A(n2619), .Y(n5346) );
  AND2X1 U1150 ( .A(n1103), .B(n7242), .Y(n2615) );
  INVX1 U1151 ( .A(n2615), .Y(n5347) );
  AND2X1 U1152 ( .A(n6810), .B(n7143), .Y(n2612) );
  INVX1 U1153 ( .A(n2612), .Y(n5348) );
  AND2X1 U1154 ( .A(n6820), .B(n7505), .Y(n1536) );
  INVX1 U1155 ( .A(n1536), .Y(n5349) );
  AND2X1 U1156 ( .A(n6811), .B(n7406), .Y(n1533) );
  INVX1 U1157 ( .A(n1533), .Y(n5350) );
  AND2X1 U1158 ( .A(n1103), .B(n7769), .Y(n1529) );
  INVX1 U1159 ( .A(n1529), .Y(n5351) );
  AND2X1 U1160 ( .A(n6811), .B(n7670), .Y(n1526) );
  INVX1 U1163 ( .A(n1526), .Y(n5352) );
  AND2X1 U1166 ( .A(n1103), .B(n6977), .Y(n1522) );
  INVX1 U1169 ( .A(n1522), .Y(n5353) );
  AND2X1 U1171 ( .A(n6810), .B(n6878), .Y(n1519) );
  INVX1 U1174 ( .A(n1519), .Y(n5354) );
  AND2X1 U1177 ( .A(n1103), .B(n7241), .Y(n1515) );
  INVX1 U1179 ( .A(n1515), .Y(n5355) );
  AND2X1 U1182 ( .A(n6811), .B(n7142), .Y(n1512) );
  INVX1 U1185 ( .A(n1512), .Y(n5356) );
  AND2X1 U1189 ( .A(n1103), .B(n7504), .Y(n1502) );
  INVX1 U1192 ( .A(n1502), .Y(n5357) );
  AND2X1 U1194 ( .A(n6810), .B(n7405), .Y(n1499) );
  INVX1 U1197 ( .A(n1499), .Y(n5358) );
  AND2X1 U1200 ( .A(n1103), .B(n7768), .Y(n1495) );
  INVX1 U1203 ( .A(n1495), .Y(n5359) );
  AND2X1 U1205 ( .A(n6810), .B(n7669), .Y(n1492) );
  INVX1 U1208 ( .A(n1492), .Y(n5360) );
  AND2X1 U1211 ( .A(n1103), .B(n6976), .Y(n1488) );
  INVX1 U1213 ( .A(n1488), .Y(n5361) );
  AND2X1 U1216 ( .A(n6811), .B(n6877), .Y(n1485) );
  INVX1 U1219 ( .A(n1485), .Y(n5362) );
  AND2X1 U1223 ( .A(n1103), .B(n7240), .Y(n1481) );
  INVX1 U1226 ( .A(n1481), .Y(n5363) );
  AND2X1 U1228 ( .A(n6811), .B(n7141), .Y(n1478) );
  INVX1 U1231 ( .A(n1478), .Y(n5364) );
  AND2X1 U1234 ( .A(n1103), .B(n7503), .Y(n1468) );
  INVX1 U1237 ( .A(n1468), .Y(n5365) );
  AND2X1 U1239 ( .A(n6810), .B(n7404), .Y(n1465) );
  INVX1 U1242 ( .A(n1465), .Y(n5366) );
  AND2X1 U1245 ( .A(n1103), .B(n7767), .Y(n1461) );
  INVX1 U1247 ( .A(n1461), .Y(n5367) );
  AND2X1 U1250 ( .A(n6810), .B(n7668), .Y(n1458) );
  INVX1 U1253 ( .A(n1458), .Y(n5368) );
  AND2X1 U1257 ( .A(n1103), .B(n6975), .Y(n1454) );
  INVX1 U1260 ( .A(n1454), .Y(n5369) );
  AND2X1 U1262 ( .A(n6811), .B(n6876), .Y(n1451) );
  INVX1 U1265 ( .A(n1451), .Y(n5370) );
  AND2X1 U1268 ( .A(n1103), .B(n7239), .Y(n1447) );
  INVX1 U1271 ( .A(n1447), .Y(n5371) );
  AND2X1 U1273 ( .A(n6810), .B(n7140), .Y(n1444) );
  INVX1 U1276 ( .A(n1444), .Y(n5372) );
  AND2X1 U1279 ( .A(n1103), .B(n7502), .Y(n1434) );
  INVX1 U1281 ( .A(n1434), .Y(n5373) );
  AND2X1 U1284 ( .A(n6811), .B(n7403), .Y(n1431) );
  INVX1 U1287 ( .A(n1431), .Y(n5374) );
  AND2X1 U1291 ( .A(n1103), .B(n7766), .Y(n1427) );
  INVX1 U1294 ( .A(n1427), .Y(n5375) );
  AND2X1 U1296 ( .A(n6811), .B(n7667), .Y(n1424) );
  INVX1 U1299 ( .A(n1424), .Y(n5376) );
  AND2X1 U1302 ( .A(n1103), .B(n6974), .Y(n1420) );
  INVX1 U1305 ( .A(n1420), .Y(n5377) );
  AND2X1 U1307 ( .A(n6810), .B(n6875), .Y(n1417) );
  INVX1 U1310 ( .A(n1417), .Y(n5378) );
  AND2X1 U1313 ( .A(n1103), .B(n7238), .Y(n1413) );
  INVX1 U1315 ( .A(n1413), .Y(n5379) );
  AND2X1 U1318 ( .A(n6810), .B(n7139), .Y(n1410) );
  INVX1 U1321 ( .A(n1410), .Y(n5380) );
  AND2X1 U1325 ( .A(n1103), .B(n7501), .Y(n1400) );
  INVX1 U1328 ( .A(n1400), .Y(n5381) );
  AND2X1 U1330 ( .A(n6810), .B(n7402), .Y(n1397) );
  INVX1 U1333 ( .A(n1397), .Y(n5382) );
  AND2X1 U1336 ( .A(n1103), .B(n7765), .Y(n1393) );
  INVX1 U1339 ( .A(n1393), .Y(n5383) );
  AND2X1 U1341 ( .A(n6810), .B(n7666), .Y(n1390) );
  INVX1 U1344 ( .A(n1390), .Y(n5384) );
  AND2X1 U1347 ( .A(n1103), .B(n6973), .Y(n1386) );
  INVX1 U1349 ( .A(n1386), .Y(n5385) );
  AND2X1 U1352 ( .A(n6810), .B(n6874), .Y(n1383) );
  INVX1 U1355 ( .A(n1383), .Y(n5386) );
  AND2X1 U1359 ( .A(n1103), .B(n7237), .Y(n1379) );
  INVX1 U1362 ( .A(n1379), .Y(n5387) );
  AND2X1 U1364 ( .A(n6811), .B(n7138), .Y(n1376) );
  INVX1 U1367 ( .A(n1376), .Y(n5388) );
  AND2X1 U1370 ( .A(n1103), .B(n7500), .Y(n1366) );
  INVX1 U1373 ( .A(n1366), .Y(n5389) );
  AND2X1 U1375 ( .A(n6811), .B(n7401), .Y(n1363) );
  INVX1 U1378 ( .A(n1363), .Y(n5390) );
  AND2X1 U1381 ( .A(n1103), .B(n7764), .Y(n1359) );
  INVX1 U1383 ( .A(n1359), .Y(n5391) );
  AND2X1 U1386 ( .A(n6810), .B(n7665), .Y(n1356) );
  INVX1 U1389 ( .A(n1356), .Y(n5392) );
  AND2X1 U1393 ( .A(n1103), .B(n6972), .Y(n1352) );
  INVX1 U1396 ( .A(n1352), .Y(n5393) );
  AND2X1 U1398 ( .A(n6810), .B(n6873), .Y(n1349) );
  INVX1 U1401 ( .A(n1349), .Y(n5394) );
  AND2X1 U1404 ( .A(n1103), .B(n7236), .Y(n1345) );
  INVX1 U1407 ( .A(n1345), .Y(n5395) );
  AND2X1 U1409 ( .A(n6811), .B(n7137), .Y(n1342) );
  INVX1 U1412 ( .A(n1342), .Y(n5396) );
  AND2X1 U1415 ( .A(n1103), .B(n7499), .Y(n1332) );
  INVX1 U1417 ( .A(n1332), .Y(n5397) );
  AND2X1 U1420 ( .A(n6810), .B(n7400), .Y(n1329) );
  INVX1 U1423 ( .A(n1329), .Y(n5398) );
  AND2X1 U1427 ( .A(n1103), .B(n7763), .Y(n1325) );
  INVX1 U1430 ( .A(n1325), .Y(n5399) );
  AND2X1 U1432 ( .A(n6811), .B(n7664), .Y(n1322) );
  INVX1 U1435 ( .A(n1322), .Y(n5400) );
  AND2X1 U1438 ( .A(n1103), .B(n6971), .Y(n1318) );
  INVX1 U1441 ( .A(n1318), .Y(n5401) );
  AND2X1 U1443 ( .A(n6810), .B(n6872), .Y(n1315) );
  INVX1 U1446 ( .A(n1315), .Y(n5402) );
  AND2X1 U1449 ( .A(n1103), .B(n7235), .Y(n1311) );
  INVX1 U1451 ( .A(n1311), .Y(n5403) );
  AND2X1 U1454 ( .A(n6811), .B(n7136), .Y(n1308) );
  INVX1 U1457 ( .A(n1308), .Y(n5404) );
  AND2X1 U1461 ( .A(n1103), .B(n7498), .Y(n1298) );
  INVX1 U1464 ( .A(n1298), .Y(n5405) );
  AND2X1 U1466 ( .A(n6811), .B(n7399), .Y(n1295) );
  INVX1 U1469 ( .A(n1295), .Y(n5406) );
  AND2X1 U1472 ( .A(n1103), .B(n7762), .Y(n1291) );
  INVX1 U1475 ( .A(n1291), .Y(n5407) );
  AND2X1 U1477 ( .A(n6811), .B(n7663), .Y(n1288) );
  INVX1 U1480 ( .A(n1288), .Y(n5408) );
  AND2X1 U1483 ( .A(n1103), .B(n6970), .Y(n1284) );
  INVX1 U1485 ( .A(n1284), .Y(n5409) );
  AND2X1 U1488 ( .A(n6811), .B(n6871), .Y(n1281) );
  INVX1 U1491 ( .A(n1281), .Y(n5410) );
  AND2X1 U1495 ( .A(n1103), .B(n7234), .Y(n1277) );
  INVX1 U1498 ( .A(n1277), .Y(n5411) );
  AND2X1 U1500 ( .A(n6810), .B(n7135), .Y(n1274) );
  INVX1 U1503 ( .A(n1274), .Y(n5412) );
  AND2X1 U1506 ( .A(n1103), .B(n7497), .Y(n1264) );
  INVX1 U1509 ( .A(n1264), .Y(n5413) );
  AND2X1 U1511 ( .A(n6810), .B(n7398), .Y(n1261) );
  INVX1 U1514 ( .A(n1261), .Y(n5414) );
  AND2X1 U1517 ( .A(n1103), .B(n7761), .Y(n1257) );
  INVX1 U1519 ( .A(n1257), .Y(n5415) );
  AND2X1 U1522 ( .A(n6811), .B(n7662), .Y(n1254) );
  INVX1 U1525 ( .A(n1254), .Y(n5416) );
  AND2X1 U1529 ( .A(n1103), .B(n6969), .Y(n1250) );
  INVX1 U1532 ( .A(n1250), .Y(n5417) );
  AND2X1 U1534 ( .A(n6810), .B(n6870), .Y(n1247) );
  INVX1 U1537 ( .A(n1247), .Y(n5418) );
  AND2X1 U1540 ( .A(n1103), .B(n7233), .Y(n1243) );
  INVX1 U1543 ( .A(n1243), .Y(n5419) );
  AND2X1 U1545 ( .A(n6810), .B(n7134), .Y(n1240) );
  INVX1 U1548 ( .A(n1240), .Y(n5420) );
  AND2X1 U1551 ( .A(n1103), .B(n7495), .Y(n1230) );
  INVX1 U1553 ( .A(n1230), .Y(n5421) );
  AND2X1 U1556 ( .A(n6811), .B(n7396), .Y(n1227) );
  INVX1 U1559 ( .A(n1227), .Y(n5422) );
  AND2X1 U1563 ( .A(n1103), .B(n7759), .Y(n1223) );
  INVX1 U1566 ( .A(n1223), .Y(n5423) );
  AND2X1 U1568 ( .A(n6810), .B(n7660), .Y(n1220) );
  INVX1 U1571 ( .A(n1220), .Y(n5424) );
  AND2X1 U1574 ( .A(n1103), .B(n6967), .Y(n1216) );
  INVX1 U1577 ( .A(n1216), .Y(n5425) );
  AND2X1 U1579 ( .A(n6810), .B(n6868), .Y(n1213) );
  INVX1 U1582 ( .A(n1213), .Y(n5426) );
  AND2X1 U1585 ( .A(n1103), .B(n7231), .Y(n1209) );
  INVX1 U1587 ( .A(n1209), .Y(n5427) );
  AND2X1 U1590 ( .A(n6810), .B(n7132), .Y(n1206) );
  INVX1 U1593 ( .A(n1206), .Y(n5428) );
  AND2X1 U1597 ( .A(n1103), .B(n7493), .Y(n1196) );
  INVX1 U1600 ( .A(n1196), .Y(n5429) );
  AND2X1 U1602 ( .A(n6810), .B(n7394), .Y(n1193) );
  INVX1 U1605 ( .A(n1193), .Y(n5430) );
  AND2X1 U1608 ( .A(n1103), .B(n7757), .Y(n1189) );
  INVX1 U1611 ( .A(n1189), .Y(n5431) );
  AND2X1 U1613 ( .A(n6810), .B(n7658), .Y(n1186) );
  INVX1 U1616 ( .A(n1186), .Y(n5432) );
  AND2X1 U1619 ( .A(n1103), .B(n6965), .Y(n1182) );
  INVX1 U1621 ( .A(n1182), .Y(n5433) );
  AND2X1 U1624 ( .A(n6810), .B(n6866), .Y(n1179) );
  INVX1 U1627 ( .A(n1179), .Y(n5434) );
  AND2X1 U1631 ( .A(n1103), .B(n7229), .Y(n1175) );
  INVX1 U1634 ( .A(n1175), .Y(n5435) );
  AND2X1 U1636 ( .A(n6811), .B(n7130), .Y(n1172) );
  INVX1 U1639 ( .A(n1172), .Y(n5436) );
  AND2X1 U1642 ( .A(n1103), .B(n7491), .Y(n1162) );
  INVX1 U1645 ( .A(n1162), .Y(n5437) );
  AND2X1 U1647 ( .A(n6810), .B(n7392), .Y(n1159) );
  INVX1 U1650 ( .A(n1159), .Y(n5438) );
  AND2X1 U1653 ( .A(n1103), .B(n7755), .Y(n1155) );
  INVX1 U1655 ( .A(n1155), .Y(n5439) );
  AND2X1 U1658 ( .A(n6811), .B(n7656), .Y(n1152) );
  INVX1 U1661 ( .A(n1152), .Y(n5440) );
  AND2X1 U1665 ( .A(n1103), .B(n6963), .Y(n1148) );
  INVX1 U1668 ( .A(n1148), .Y(n5441) );
  AND2X1 U1670 ( .A(n6811), .B(n6864), .Y(n1145) );
  INVX1 U1673 ( .A(n1145), .Y(n5442) );
  AND2X1 U1676 ( .A(n1103), .B(n7227), .Y(n1141) );
  INVX1 U1679 ( .A(n1141), .Y(n5443) );
  AND2X1 U1681 ( .A(n6810), .B(n7128), .Y(n1138) );
  INVX1 U1684 ( .A(n1138), .Y(n5444) );
  AND2X1 U1687 ( .A(n1103), .B(n7489), .Y(n1128) );
  INVX1 U1689 ( .A(n1128), .Y(n5445) );
  AND2X1 U1692 ( .A(n6811), .B(n7390), .Y(n1125) );
  INVX1 U1695 ( .A(n1125), .Y(n5446) );
  AND2X1 U1699 ( .A(n1103), .B(n7753), .Y(n1120) );
  INVX1 U1702 ( .A(n1120), .Y(n5447) );
  AND2X1 U1704 ( .A(n6810), .B(n7654), .Y(n1117) );
  INVX1 U1707 ( .A(n1117), .Y(n5448) );
  AND2X1 U1710 ( .A(n1103), .B(n6961), .Y(n1112) );
  INVX1 U1713 ( .A(n1112), .Y(n5449) );
  AND2X1 U1715 ( .A(n6811), .B(n6862), .Y(n1109) );
  INVX1 U1718 ( .A(n1109), .Y(n5450) );
  AND2X1 U1721 ( .A(n1103), .B(n7225), .Y(n1099) );
  INVX1 U1723 ( .A(n1099), .Y(n5451) );
  AND2X1 U1726 ( .A(n6810), .B(n7126), .Y(n1094) );
  INVX1 U1729 ( .A(n1094), .Y(n5452) );
  BUFX2 U1733 ( .A(n3297), .Y(n5453) );
  BUFX2 U1736 ( .A(n3286), .Y(n5454) );
  BUFX2 U1738 ( .A(n3283), .Y(n5455) );
  BUFX2 U1741 ( .A(n3279), .Y(n5456) );
  BUFX2 U1744 ( .A(n3275), .Y(n5457) );
  BUFX2 U1747 ( .A(n3271), .Y(n5458) );
  BUFX2 U1749 ( .A(n3267), .Y(n5459) );
  BUFX2 U1752 ( .A(n3263), .Y(n5460) );
  BUFX2 U1755 ( .A(n3259), .Y(n5461) );
  BUFX2 U1757 ( .A(n3249), .Y(n5462) );
  BUFX2 U1760 ( .A(n3246), .Y(n5463) );
  BUFX2 U1763 ( .A(n3242), .Y(n5464) );
  BUFX2 U1767 ( .A(n3239), .Y(n5465) );
  BUFX2 U1770 ( .A(n3235), .Y(n5466) );
  BUFX2 U1772 ( .A(n3232), .Y(n5467) );
  BUFX2 U1775 ( .A(n3228), .Y(n5468) );
  BUFX2 U1778 ( .A(n3225), .Y(n5469) );
  BUFX2 U1781 ( .A(n3215), .Y(n5470) );
  BUFX2 U1783 ( .A(n3212), .Y(n5471) );
  BUFX2 U1786 ( .A(n3208), .Y(n5472) );
  BUFX2 U1789 ( .A(n3205), .Y(n5473) );
  BUFX2 U1791 ( .A(n3201), .Y(n5474) );
  BUFX2 U1794 ( .A(n3198), .Y(n5475) );
  BUFX2 U1797 ( .A(n3194), .Y(n5476) );
  BUFX2 U1801 ( .A(n3191), .Y(n5477) );
  BUFX2 U1804 ( .A(n3181), .Y(n5478) );
  BUFX2 U1806 ( .A(n3178), .Y(n5479) );
  BUFX2 U1809 ( .A(n3174), .Y(n5480) );
  BUFX2 U1812 ( .A(n3171), .Y(n5481) );
  BUFX2 U1815 ( .A(n3167), .Y(n5482) );
  BUFX2 U1817 ( .A(n3164), .Y(n5483) );
  BUFX2 U1820 ( .A(n3160), .Y(n5484) );
  BUFX2 U1823 ( .A(n3157), .Y(n5485) );
  BUFX2 U1825 ( .A(n3147), .Y(n5486) );
  BUFX2 U1828 ( .A(n3144), .Y(n5487) );
  BUFX2 U1831 ( .A(n3140), .Y(n5488) );
  BUFX2 U1835 ( .A(n3137), .Y(n5489) );
  BUFX2 U1838 ( .A(n3133), .Y(n5490) );
  BUFX2 U1840 ( .A(n3130), .Y(n5491) );
  BUFX2 U1843 ( .A(n3126), .Y(n5492) );
  BUFX2 U1846 ( .A(n3123), .Y(n5493) );
  BUFX2 U1849 ( .A(n3113), .Y(n5494) );
  BUFX2 U1851 ( .A(n3110), .Y(n5495) );
  BUFX2 U1854 ( .A(n3106), .Y(n5496) );
  BUFX2 U1857 ( .A(n3103), .Y(n5497) );
  BUFX2 U1859 ( .A(n3099), .Y(n5498) );
  BUFX2 U1862 ( .A(n3096), .Y(n5499) );
  BUFX2 U1865 ( .A(n3092), .Y(n5500) );
  BUFX2 U1869 ( .A(n3089), .Y(n5501) );
  BUFX2 U1872 ( .A(n3079), .Y(n5502) );
  BUFX2 U1874 ( .A(n3076), .Y(n5503) );
  BUFX2 U1877 ( .A(n3072), .Y(n5504) );
  BUFX2 U1880 ( .A(n3069), .Y(n5505) );
  BUFX2 U1883 ( .A(n3065), .Y(n5506) );
  BUFX2 U1885 ( .A(n3062), .Y(n5507) );
  BUFX2 U1888 ( .A(n3058), .Y(n5508) );
  BUFX2 U1891 ( .A(n3055), .Y(n5509) );
  BUFX2 U1893 ( .A(n3045), .Y(n5510) );
  BUFX2 U1896 ( .A(n3042), .Y(n5511) );
  BUFX2 U1899 ( .A(n3038), .Y(n5512) );
  BUFX2 U1903 ( .A(n3035), .Y(n5513) );
  BUFX2 U1906 ( .A(n3031), .Y(n5514) );
  BUFX2 U1908 ( .A(n3028), .Y(n5515) );
  BUFX2 U1911 ( .A(n3024), .Y(n5516) );
  BUFX2 U1914 ( .A(n3021), .Y(n5517) );
  BUFX2 U1917 ( .A(n3011), .Y(n5518) );
  BUFX2 U1919 ( .A(n3008), .Y(n5519) );
  BUFX2 U1922 ( .A(n3004), .Y(n5520) );
  BUFX2 U1925 ( .A(n3001), .Y(n5521) );
  BUFX2 U1927 ( .A(n2997), .Y(n5522) );
  BUFX2 U1930 ( .A(n2994), .Y(n5523) );
  BUFX2 U1933 ( .A(n2990), .Y(n5524) );
  BUFX2 U1937 ( .A(n2987), .Y(n5525) );
  BUFX2 U1940 ( .A(n2977), .Y(n5526) );
  BUFX2 U1942 ( .A(n2974), .Y(n5527) );
  BUFX2 U1945 ( .A(n2970), .Y(n5528) );
  BUFX2 U1948 ( .A(n2967), .Y(n5529) );
  BUFX2 U1951 ( .A(n2963), .Y(n5530) );
  BUFX2 U1953 ( .A(n2960), .Y(n5531) );
  BUFX2 U1956 ( .A(n2956), .Y(n5532) );
  BUFX2 U1959 ( .A(n2953), .Y(n5533) );
  BUFX2 U1961 ( .A(n2943), .Y(n5534) );
  BUFX2 U1964 ( .A(n2940), .Y(n5535) );
  BUFX2 U1967 ( .A(n2936), .Y(n5536) );
  BUFX2 U1971 ( .A(n2933), .Y(n5537) );
  BUFX2 U1974 ( .A(n2929), .Y(n5538) );
  BUFX2 U1976 ( .A(n2926), .Y(n5539) );
  BUFX2 U1979 ( .A(n2922), .Y(n5540) );
  BUFX2 U1982 ( .A(n2919), .Y(n5541) );
  BUFX2 U1985 ( .A(n2909), .Y(n5542) );
  BUFX2 U1987 ( .A(n2906), .Y(n5543) );
  BUFX2 U1990 ( .A(n2902), .Y(n5544) );
  BUFX2 U1993 ( .A(n2899), .Y(n5545) );
  BUFX2 U1995 ( .A(n2895), .Y(n5546) );
  BUFX2 U1998 ( .A(n2892), .Y(n5547) );
  BUFX2 U2001 ( .A(n2888), .Y(n5548) );
  BUFX2 U2005 ( .A(n2885), .Y(n5549) );
  BUFX2 U2008 ( .A(n2875), .Y(n5550) );
  BUFX2 U2010 ( .A(n2872), .Y(n5551) );
  BUFX2 U2013 ( .A(n2868), .Y(n5552) );
  BUFX2 U2016 ( .A(n2865), .Y(n5553) );
  BUFX2 U2019 ( .A(n2861), .Y(n5554) );
  BUFX2 U2021 ( .A(n2858), .Y(n5555) );
  BUFX2 U2024 ( .A(n2854), .Y(n5556) );
  BUFX2 U2027 ( .A(n2851), .Y(n5557) );
  BUFX2 U2029 ( .A(n2841), .Y(n5558) );
  BUFX2 U2032 ( .A(n2838), .Y(n5559) );
  BUFX2 U2035 ( .A(n2834), .Y(n5560) );
  BUFX2 U2039 ( .A(n2831), .Y(n5561) );
  BUFX2 U2042 ( .A(n2827), .Y(n5562) );
  BUFX2 U2044 ( .A(n2824), .Y(n5563) );
  BUFX2 U2047 ( .A(n2820), .Y(n5564) );
  BUFX2 U2050 ( .A(n2817), .Y(n5565) );
  BUFX2 U2053 ( .A(n2807), .Y(n5566) );
  BUFX2 U2055 ( .A(n2804), .Y(n5567) );
  BUFX2 U2058 ( .A(n2800), .Y(n5568) );
  BUFX2 U2061 ( .A(n2797), .Y(n5569) );
  BUFX2 U2063 ( .A(n2793), .Y(n5570) );
  BUFX2 U2066 ( .A(n2790), .Y(n5571) );
  BUFX2 U2069 ( .A(n2786), .Y(n5572) );
  BUFX2 U2073 ( .A(n2783), .Y(n5573) );
  BUFX2 U2076 ( .A(n2773), .Y(n5574) );
  BUFX2 U2078 ( .A(n2770), .Y(n5575) );
  BUFX2 U2081 ( .A(n2766), .Y(n5576) );
  BUFX2 U2084 ( .A(n2763), .Y(n5577) );
  BUFX2 U2087 ( .A(n2759), .Y(n5578) );
  BUFX2 U2089 ( .A(n2756), .Y(n5579) );
  BUFX2 U2092 ( .A(n2752), .Y(n5580) );
  BUFX2 U2095 ( .A(n2749), .Y(n5581) );
  BUFX2 U2097 ( .A(n2739), .Y(n5582) );
  BUFX2 U2100 ( .A(n2736), .Y(n5583) );
  BUFX2 U2103 ( .A(n2732), .Y(n5584) );
  BUFX2 U2107 ( .A(n2729), .Y(n5585) );
  BUFX2 U2110 ( .A(n2725), .Y(n5586) );
  BUFX2 U2112 ( .A(n2722), .Y(n5587) );
  BUFX2 U2115 ( .A(n2718), .Y(n5588) );
  BUFX2 U2118 ( .A(n2715), .Y(n5589) );
  BUFX2 U2121 ( .A(n2705), .Y(n5590) );
  BUFX2 U2123 ( .A(n2702), .Y(n5591) );
  BUFX2 U2126 ( .A(n2698), .Y(n5592) );
  BUFX2 U2129 ( .A(n2695), .Y(n5593) );
  BUFX2 U2131 ( .A(n2691), .Y(n5594) );
  BUFX2 U2134 ( .A(n2688), .Y(n5595) );
  BUFX2 U2137 ( .A(n2684), .Y(n5596) );
  BUFX2 U2141 ( .A(n2681), .Y(n5597) );
  BUFX2 U2144 ( .A(n2671), .Y(n5598) );
  BUFX2 U2146 ( .A(n2668), .Y(n5599) );
  BUFX2 U2149 ( .A(n2664), .Y(n5600) );
  BUFX2 U2152 ( .A(n2661), .Y(n5601) );
  BUFX2 U2155 ( .A(n2657), .Y(n5602) );
  BUFX2 U2157 ( .A(n2654), .Y(n5603) );
  BUFX2 U2160 ( .A(n2650), .Y(n5604) );
  BUFX2 U2163 ( .A(n2647), .Y(n5605) );
  BUFX2 U2165 ( .A(n2637), .Y(n5606) );
  BUFX2 U2168 ( .A(n2634), .Y(n5607) );
  BUFX2 U2171 ( .A(n2630), .Y(n5608) );
  BUFX2 U2175 ( .A(n2627), .Y(n5609) );
  BUFX2 U2178 ( .A(n2623), .Y(n5610) );
  BUFX2 U2180 ( .A(n2620), .Y(n5611) );
  BUFX2 U2183 ( .A(n2616), .Y(n5612) );
  BUFX2 U2186 ( .A(n2613), .Y(n5613) );
  BUFX2 U2189 ( .A(n1537), .Y(n5614) );
  BUFX2 U2191 ( .A(n1534), .Y(n5615) );
  BUFX2 U2194 ( .A(n1530), .Y(n5616) );
  BUFX2 U2197 ( .A(n1527), .Y(n5617) );
  BUFX2 U2199 ( .A(n1523), .Y(n5618) );
  BUFX2 U2202 ( .A(n1520), .Y(n5619) );
  BUFX2 U2205 ( .A(n1516), .Y(n5620) );
  BUFX2 U2209 ( .A(n1513), .Y(n5621) );
  BUFX2 U2212 ( .A(n1503), .Y(n5622) );
  BUFX2 U2214 ( .A(n1500), .Y(n5623) );
  BUFX2 U2217 ( .A(n1496), .Y(n5624) );
  BUFX2 U2220 ( .A(n1493), .Y(n5625) );
  BUFX2 U2223 ( .A(n1489), .Y(n5626) );
  BUFX2 U2225 ( .A(n1486), .Y(n5627) );
  BUFX2 U2228 ( .A(n1482), .Y(n5628) );
  BUFX2 U2231 ( .A(n1479), .Y(n5629) );
  BUFX2 U2233 ( .A(n1469), .Y(n5630) );
  BUFX2 U2236 ( .A(n1466), .Y(n5631) );
  BUFX2 U2239 ( .A(n1462), .Y(n5632) );
  BUFX2 U2243 ( .A(n1459), .Y(n5633) );
  BUFX2 U2246 ( .A(n1455), .Y(n5634) );
  BUFX2 U2248 ( .A(n1452), .Y(n5635) );
  BUFX2 U2251 ( .A(n1448), .Y(n5636) );
  BUFX2 U2254 ( .A(n1445), .Y(n5637) );
  BUFX2 U2257 ( .A(n1435), .Y(n5638) );
  BUFX2 U2259 ( .A(n1432), .Y(n5639) );
  BUFX2 U2262 ( .A(n1428), .Y(n5640) );
  BUFX2 U2265 ( .A(n1425), .Y(n5641) );
  BUFX2 U2267 ( .A(n1421), .Y(n5642) );
  BUFX2 U2270 ( .A(n1418), .Y(n5643) );
  BUFX2 U2274 ( .A(n1414), .Y(n5644) );
  BUFX2 U2279 ( .A(n1411), .Y(n5645) );
  BUFX2 U2282 ( .A(n1401), .Y(n5646) );
  BUFX2 U2284 ( .A(n1398), .Y(n5647) );
  BUFX2 U2291 ( .A(n1394), .Y(n5648) );
  BUFX2 U2292 ( .A(n1391), .Y(n5649) );
  BUFX2 U2295 ( .A(n1387), .Y(n5650) );
  BUFX2 U2305 ( .A(n1384), .Y(n5651) );
  BUFX2 U2306 ( .A(n1380), .Y(n5652) );
  BUFX2 U2307 ( .A(n1377), .Y(n5653) );
  BUFX2 U2312 ( .A(n1367), .Y(n5654) );
  BUFX2 U2322 ( .A(n1364), .Y(n5655) );
  BUFX2 U2323 ( .A(n1360), .Y(n5656) );
  BUFX2 U2325 ( .A(n1357), .Y(n5657) );
  BUFX2 U2327 ( .A(n1353), .Y(n5658) );
  BUFX2 U2329 ( .A(n1350), .Y(n5659) );
  BUFX2 U2331 ( .A(n1346), .Y(n5660) );
  BUFX2 U2333 ( .A(n1343), .Y(n5661) );
  BUFX2 U2335 ( .A(n1333), .Y(n5662) );
  BUFX2 U2337 ( .A(n1330), .Y(n5663) );
  BUFX2 U2339 ( .A(n1326), .Y(n5664) );
  BUFX2 U2341 ( .A(n1323), .Y(n5665) );
  BUFX2 U2343 ( .A(n1319), .Y(n5666) );
  BUFX2 U2345 ( .A(n1316), .Y(n5667) );
  BUFX2 U2347 ( .A(n1312), .Y(n5668) );
  BUFX2 U2349 ( .A(n1309), .Y(n5669) );
  BUFX2 U2351 ( .A(n1299), .Y(n5670) );
  BUFX2 U2353 ( .A(n1296), .Y(n5671) );
  BUFX2 U2355 ( .A(n1292), .Y(n5672) );
  BUFX2 U2357 ( .A(n1289), .Y(n5673) );
  BUFX2 U2359 ( .A(n1285), .Y(n5674) );
  BUFX2 U2361 ( .A(n1282), .Y(n5675) );
  BUFX2 U2363 ( .A(n1278), .Y(n5676) );
  BUFX2 U2365 ( .A(n1275), .Y(n5677) );
  BUFX2 U2367 ( .A(n1265), .Y(n5678) );
  BUFX2 U2369 ( .A(n1262), .Y(n5679) );
  BUFX2 U2371 ( .A(n1258), .Y(n5680) );
  BUFX2 U2373 ( .A(n1255), .Y(n5681) );
  BUFX2 U2375 ( .A(n1251), .Y(n5682) );
  BUFX2 U2377 ( .A(n1248), .Y(n5683) );
  BUFX2 U2379 ( .A(n1244), .Y(n5684) );
  BUFX2 U2381 ( .A(n1241), .Y(n5685) );
  BUFX2 U2383 ( .A(n1231), .Y(n5686) );
  BUFX2 U2385 ( .A(n1228), .Y(n5687) );
  BUFX2 U2387 ( .A(n1224), .Y(n5688) );
  BUFX2 U2389 ( .A(n1221), .Y(n5689) );
  BUFX2 U2392 ( .A(n1217), .Y(n5690) );
  BUFX2 U2394 ( .A(n1214), .Y(n5691) );
  BUFX2 U2396 ( .A(n1210), .Y(n5692) );
  BUFX2 U2398 ( .A(n1207), .Y(n5693) );
  BUFX2 U2400 ( .A(n1197), .Y(n5694) );
  BUFX2 U2402 ( .A(n1194), .Y(n5695) );
  BUFX2 U2404 ( .A(n1190), .Y(n5696) );
  BUFX2 U2406 ( .A(n1187), .Y(n5697) );
  BUFX2 U2408 ( .A(n1183), .Y(n5698) );
  BUFX2 U2410 ( .A(n1180), .Y(n5699) );
  BUFX2 U2412 ( .A(n1176), .Y(n5700) );
  BUFX2 U2414 ( .A(n1173), .Y(n5701) );
  BUFX2 U2416 ( .A(n1163), .Y(n5702) );
  BUFX2 U2418 ( .A(n1160), .Y(n5703) );
  BUFX2 U2420 ( .A(n1156), .Y(n5704) );
  BUFX2 U2422 ( .A(n1153), .Y(n5705) );
  BUFX2 U2424 ( .A(n1149), .Y(n5706) );
  BUFX2 U2426 ( .A(n1146), .Y(n5707) );
  BUFX2 U2428 ( .A(n1142), .Y(n5708) );
  BUFX2 U2430 ( .A(n1139), .Y(n5709) );
  BUFX2 U2432 ( .A(n1129), .Y(n5710) );
  BUFX2 U2434 ( .A(n1126), .Y(n5711) );
  BUFX2 U2436 ( .A(n1121), .Y(n5712) );
  BUFX2 U2438 ( .A(n1118), .Y(n5713) );
  BUFX2 U2440 ( .A(n1113), .Y(n5714) );
  BUFX2 U2442 ( .A(n1110), .Y(n5715) );
  BUFX2 U2444 ( .A(n1100), .Y(n5716) );
  BUFX2 U2446 ( .A(n1095), .Y(n5717) );
  INVX1 U2448 ( .A(n3253), .Y(n5718) );
  INVX1 U2450 ( .A(n3219), .Y(n5719) );
  INVX1 U2452 ( .A(n3185), .Y(n5720) );
  INVX1 U2454 ( .A(n3151), .Y(n5721) );
  INVX1 U2456 ( .A(n3117), .Y(n5722) );
  INVX1 U2459 ( .A(n3083), .Y(n5723) );
  INVX1 U2461 ( .A(n3049), .Y(n5724) );
  INVX1 U2463 ( .A(n3015), .Y(n5725) );
  INVX1 U2465 ( .A(n2981), .Y(n5726) );
  INVX1 U2467 ( .A(n2947), .Y(n5727) );
  INVX1 U2469 ( .A(n2913), .Y(n5728) );
  INVX1 U2471 ( .A(n2879), .Y(n5729) );
  INVX1 U2473 ( .A(n2845), .Y(n5730) );
  INVX1 U2475 ( .A(n2811), .Y(n5731) );
  INVX1 U2477 ( .A(n2777), .Y(n5732) );
  INVX1 U2479 ( .A(n2743), .Y(n5733) );
  INVX1 U2481 ( .A(n2709), .Y(n5734) );
  INVX1 U2483 ( .A(n2675), .Y(n5735) );
  INVX1 U2485 ( .A(n2641), .Y(n5736) );
  INVX1 U2487 ( .A(n2607), .Y(n5737) );
  INVX1 U2489 ( .A(n1507), .Y(n5738) );
  INVX1 U2491 ( .A(n1473), .Y(n5739) );
  INVX1 U2493 ( .A(n1439), .Y(n5740) );
  INVX1 U2495 ( .A(n1405), .Y(n5741) );
  INVX1 U2497 ( .A(n1371), .Y(n5742) );
  INVX1 U2499 ( .A(n1337), .Y(n5743) );
  INVX1 U2501 ( .A(n1303), .Y(n5744) );
  INVX1 U2503 ( .A(n1269), .Y(n5745) );
  INVX1 U2505 ( .A(n1235), .Y(n5746) );
  INVX1 U2507 ( .A(n1201), .Y(n5747) );
  INVX1 U2509 ( .A(n1167), .Y(n5748) );
  INVX1 U2511 ( .A(n1133), .Y(n5749) );
  INVX1 U2513 ( .A(n1089), .Y(n5750) );
  INVX1 U2515 ( .A(n3254), .Y(n5751) );
  INVX1 U2517 ( .A(n3220), .Y(n5752) );
  INVX1 U2519 ( .A(n3186), .Y(n5753) );
  INVX1 U2521 ( .A(n3152), .Y(n5754) );
  INVX1 U2523 ( .A(n3118), .Y(n5755) );
  INVX1 U2526 ( .A(n3084), .Y(n5756) );
  INVX1 U2528 ( .A(n3050), .Y(n5757) );
  INVX1 U2530 ( .A(n3016), .Y(n5758) );
  INVX1 U2532 ( .A(n2982), .Y(n5759) );
  INVX1 U2534 ( .A(n2948), .Y(n5760) );
  INVX1 U2536 ( .A(n2914), .Y(n5761) );
  INVX1 U2538 ( .A(n2880), .Y(n5762) );
  INVX1 U2540 ( .A(n2846), .Y(n5763) );
  INVX1 U2542 ( .A(n2812), .Y(n5764) );
  INVX1 U2544 ( .A(n2778), .Y(n5765) );
  INVX1 U2546 ( .A(n2744), .Y(n5766) );
  INVX1 U2548 ( .A(n2710), .Y(n5767) );
  INVX1 U2550 ( .A(n2676), .Y(n5768) );
  INVX1 U2552 ( .A(n2642), .Y(n5769) );
  INVX1 U2554 ( .A(n2608), .Y(n5770) );
  INVX1 U2556 ( .A(n1508), .Y(n5771) );
  INVX1 U2558 ( .A(n1474), .Y(n5772) );
  INVX1 U2560 ( .A(n1440), .Y(n5773) );
  INVX1 U2562 ( .A(n1406), .Y(n5774) );
  INVX1 U2564 ( .A(n1372), .Y(n5775) );
  INVX1 U2566 ( .A(n1338), .Y(n5776) );
  INVX1 U2568 ( .A(n1304), .Y(n5777) );
  INVX1 U2570 ( .A(n1270), .Y(n5778) );
  INVX1 U2572 ( .A(n1236), .Y(n5779) );
  INVX1 U2574 ( .A(n1202), .Y(n5780) );
  INVX1 U2576 ( .A(n1168), .Y(n5781) );
  INVX1 U2578 ( .A(n1134), .Y(n5782) );
  INVX1 U2580 ( .A(n1090), .Y(n5783) );
  INVX1 U2582 ( .A(n3255), .Y(n5784) );
  INVX1 U2584 ( .A(n3221), .Y(n5785) );
  INVX1 U2586 ( .A(n3187), .Y(n5786) );
  INVX1 U2588 ( .A(n3153), .Y(n5787) );
  INVX1 U2590 ( .A(n3119), .Y(n5788) );
  INVX1 U2593 ( .A(n3085), .Y(n5789) );
  INVX1 U2595 ( .A(n3051), .Y(n5790) );
  INVX1 U2597 ( .A(n3017), .Y(n5791) );
  INVX1 U2599 ( .A(n2983), .Y(n5792) );
  INVX1 U2601 ( .A(n2949), .Y(n5793) );
  INVX1 U2603 ( .A(n2915), .Y(n5794) );
  INVX1 U2605 ( .A(n2881), .Y(n5795) );
  INVX1 U2607 ( .A(n2847), .Y(n5796) );
  INVX1 U2609 ( .A(n2813), .Y(n5797) );
  INVX1 U2611 ( .A(n2779), .Y(n5798) );
  INVX1 U2613 ( .A(n2745), .Y(n5799) );
  INVX1 U2615 ( .A(n2711), .Y(n5800) );
  INVX1 U2617 ( .A(n2677), .Y(n5801) );
  INVX1 U2619 ( .A(n2643), .Y(n5802) );
  INVX1 U2621 ( .A(n2609), .Y(n5803) );
  INVX1 U2623 ( .A(n1509), .Y(n5804) );
  INVX1 U2625 ( .A(n1475), .Y(n5805) );
  INVX1 U2627 ( .A(n1441), .Y(n5806) );
  INVX1 U2629 ( .A(n1407), .Y(n5807) );
  INVX1 U2631 ( .A(n1373), .Y(n5808) );
  INVX1 U2633 ( .A(n1339), .Y(n5809) );
  INVX1 U2635 ( .A(n1305), .Y(n5810) );
  INVX1 U2637 ( .A(n1271), .Y(n5811) );
  INVX1 U2639 ( .A(n1237), .Y(n5812) );
  INVX1 U2641 ( .A(n1203), .Y(n5813) );
  INVX1 U2643 ( .A(n1169), .Y(n5814) );
  INVX1 U2645 ( .A(n1135), .Y(n5815) );
  INVX1 U2647 ( .A(n1091), .Y(n5816) );
  BUFX2 U2649 ( .A(n3301), .Y(n5817) );
  AND2X1 U2651 ( .A(n3357), .B(n3323), .Y(n3356) );
  INVX1 U2653 ( .A(n3356), .Y(n5818) );
  AND2X1 U2655 ( .A(n3381), .B(n3323), .Y(n3380) );
  INVX1 U2657 ( .A(n3380), .Y(n5819) );
  AND2X1 U2660 ( .A(n3355), .B(n3391), .Y(n3407) );
  INVX1 U2662 ( .A(n3407), .Y(n5820) );
  AND2X1 U2664 ( .A(n3379), .B(n3391), .Y(n3419) );
  INVX1 U2666 ( .A(n3419), .Y(n5821) );
  AND2X1 U2668 ( .A(n3353), .B(n3426), .Y(n3441) );
  INVX1 U2670 ( .A(n3441), .Y(n5822) );
  AND2X1 U2672 ( .A(n3377), .B(n3426), .Y(n3453) );
  INVX1 U2674 ( .A(n3453), .Y(n5823) );
  AND2X1 U2676 ( .A(n3349), .B(n3461), .Y(n3474) );
  INVX1 U2678 ( .A(n3474), .Y(n5824) );
  AND2X1 U2680 ( .A(n3375), .B(n3461), .Y(n3487) );
  INVX1 U2682 ( .A(n3487), .Y(n5825) );
  AND2X1 U2684 ( .A(n3345), .B(n3496), .Y(n3507) );
  INVX1 U2686 ( .A(n3507), .Y(n5826) );
  AND2X1 U2688 ( .A(n3373), .B(n3496), .Y(n3521) );
  INVX1 U2690 ( .A(n3521), .Y(n5827) );
  AND2X1 U2692 ( .A(n3351), .B(n3530), .Y(n3544) );
  INVX1 U2694 ( .A(n3544), .Y(n5828) );
  AND2X1 U2696 ( .A(n3371), .B(n3530), .Y(n3554) );
  INVX1 U2698 ( .A(n3554), .Y(n5829) );
  AND2X1 U2700 ( .A(n3329), .B(n3565), .Y(n3568) );
  INVX1 U2702 ( .A(n3568), .Y(n5830) );
  AND2X1 U2704 ( .A(n3369), .B(n3565), .Y(n3588) );
  INVX1 U2706 ( .A(n3588), .Y(n5831) );
  AND2X1 U2708 ( .A(n3327), .B(n3600), .Y(n3602) );
  INVX1 U2710 ( .A(n3602), .Y(n5832) );
  AND2X1 U2712 ( .A(n3367), .B(n3600), .Y(n3622) );
  INVX1 U2714 ( .A(n3622), .Y(n5833) );
  AND2X1 U2716 ( .A(n3347), .B(n3635), .Y(n3647) );
  INVX1 U2718 ( .A(n3647), .Y(n5834) );
  AND2X1 U2720 ( .A(n3325), .B(n3670), .Y(n3671) );
  INVX1 U2722 ( .A(n3671), .Y(n5835) );
  AND2X1 U2724 ( .A(n3341), .B(n3670), .Y(n3679) );
  INVX1 U2727 ( .A(n3679), .Y(n5836) );
  AND2X1 U2729 ( .A(n3339), .B(n3704), .Y(n3712) );
  INVX1 U2731 ( .A(n3712), .Y(n5837) );
  AND2X1 U2733 ( .A(n3337), .B(n3738), .Y(n3745) );
  INVX1 U2735 ( .A(n3745), .Y(n5838) );
  AND2X1 U2737 ( .A(n3357), .B(n3772), .Y(n3789) );
  INVX1 U2739 ( .A(n3789), .Y(n5839) );
  AND2X1 U2741 ( .A(n3381), .B(n3772), .Y(n3801) );
  INVX1 U2743 ( .A(n3801), .Y(n5840) );
  AND2X1 U2745 ( .A(n3355), .B(n3806), .Y(n3822) );
  INVX1 U2747 ( .A(n3822), .Y(n5841) );
  AND2X1 U2749 ( .A(n3379), .B(n3806), .Y(n3834) );
  INVX1 U2751 ( .A(n3834), .Y(n5842) );
  AND2X1 U2753 ( .A(n3353), .B(n3840), .Y(n3855) );
  INVX1 U2755 ( .A(n3855), .Y(n5843) );
  AND2X1 U2757 ( .A(n3377), .B(n3840), .Y(n3867) );
  INVX1 U2759 ( .A(n3867), .Y(n5844) );
  AND2X1 U2761 ( .A(n3349), .B(n3874), .Y(n3887) );
  INVX1 U2763 ( .A(n3887), .Y(n5845) );
  AND2X1 U2765 ( .A(n3375), .B(n3874), .Y(n3900) );
  INVX1 U2767 ( .A(n3900), .Y(n5846) );
  AND2X1 U2769 ( .A(n3345), .B(n3908), .Y(n3919) );
  INVX1 U2771 ( .A(n3919), .Y(n5847) );
  AND2X1 U2773 ( .A(n3373), .B(n3908), .Y(n3933) );
  INVX1 U2775 ( .A(n3933), .Y(n5848) );
  AND2X1 U2777 ( .A(n3351), .B(n3943), .Y(n3957) );
  INVX1 U2779 ( .A(n3957), .Y(n5849) );
  AND2X1 U2781 ( .A(n3371), .B(n3943), .Y(n3967) );
  INVX1 U2783 ( .A(n3967), .Y(n5850) );
  AND2X1 U2785 ( .A(n3329), .B(n3977), .Y(n3980) );
  INVX1 U2787 ( .A(n3980), .Y(n5851) );
  AND2X1 U2789 ( .A(n3369), .B(n3977), .Y(n4000) );
  INVX1 U2791 ( .A(n4000), .Y(n5852) );
  AND2X1 U2794 ( .A(n3327), .B(n4011), .Y(n4013) );
  INVX1 U2796 ( .A(n4013), .Y(n5853) );
  AND2X1 U2798 ( .A(n3367), .B(n4011), .Y(n4033) );
  INVX1 U2800 ( .A(n4033), .Y(n5854) );
  AND2X1 U2802 ( .A(n3347), .B(n4045), .Y(n4057) );
  INVX1 U2804 ( .A(n4057), .Y(n5855) );
  AND2X1 U2806 ( .A(n3325), .B(n4079), .Y(n4080) );
  INVX1 U2808 ( .A(n4080), .Y(n5856) );
  AND2X1 U2810 ( .A(n3341), .B(n4079), .Y(n4088) );
  INVX1 U2812 ( .A(n4088), .Y(n5857) );
  AND2X1 U2814 ( .A(n3339), .B(n4113), .Y(n4121) );
  INVX1 U2816 ( .A(n4121), .Y(n5858) );
  AND2X1 U2818 ( .A(n3337), .B(n4147), .Y(n4154) );
  INVX1 U2820 ( .A(n4154), .Y(n5859) );
  AND2X1 U2822 ( .A(n3345), .B(n4181), .Y(n4192) );
  INVX1 U2824 ( .A(n4192), .Y(n5860) );
  AND2X1 U2826 ( .A(n3373), .B(n4181), .Y(n4206) );
  INVX1 U2828 ( .A(n4206), .Y(n5861) );
  AND2X1 U2830 ( .A(n3351), .B(n4216), .Y(n4230) );
  INVX1 U2832 ( .A(n4230), .Y(n5862) );
  AND2X1 U2834 ( .A(n3371), .B(n4216), .Y(n4240) );
  INVX1 U2836 ( .A(n4240), .Y(n5863) );
  AND2X1 U2838 ( .A(n3329), .B(n4250), .Y(n4253) );
  INVX1 U2840 ( .A(n4253), .Y(n5864) );
  AND2X1 U2842 ( .A(n3369), .B(n4250), .Y(n4273) );
  INVX1 U2844 ( .A(n4273), .Y(n5865) );
  AND2X1 U2846 ( .A(n3327), .B(n4284), .Y(n4286) );
  INVX1 U2848 ( .A(n4286), .Y(n5866) );
  AND2X1 U2850 ( .A(n3367), .B(n4284), .Y(n4306) );
  INVX1 U2852 ( .A(n4306), .Y(n5867) );
  AND2X1 U2854 ( .A(n3347), .B(n4318), .Y(n4330) );
  INVX1 U2856 ( .A(n4330), .Y(n5868) );
  AND2X1 U2858 ( .A(n3325), .B(n4352), .Y(n4353) );
  INVX1 U2862 ( .A(n4353), .Y(n5869) );
  AND2X1 U2864 ( .A(n3341), .B(n4352), .Y(n4361) );
  INVX1 U2866 ( .A(n4361), .Y(n5870) );
  AND2X1 U2868 ( .A(n3339), .B(n4386), .Y(n4394) );
  INVX1 U2870 ( .A(n4394), .Y(n5871) );
  AND2X1 U2872 ( .A(n3337), .B(n4420), .Y(n4427) );
  INVX1 U2874 ( .A(n4427), .Y(n5872) );
  AND2X1 U2876 ( .A(n3355), .B(n3323), .Y(n3354) );
  INVX1 U2878 ( .A(n3354), .Y(n5873) );
  AND2X1 U2880 ( .A(n3379), .B(n3323), .Y(n3378) );
  INVX1 U2882 ( .A(n3378), .Y(n5874) );
  AND2X1 U2884 ( .A(n3357), .B(n3391), .Y(n3408) );
  INVX1 U2886 ( .A(n3408), .Y(n5875) );
  AND2X1 U2888 ( .A(n3381), .B(n3391), .Y(n3420) );
  INVX1 U2890 ( .A(n3420), .Y(n5876) );
  AND2X1 U2892 ( .A(n3349), .B(n3426), .Y(n3439) );
  INVX1 U2894 ( .A(n3439), .Y(n5877) );
  AND2X1 U2896 ( .A(n3375), .B(n3426), .Y(n3452) );
  INVX1 U2898 ( .A(n3452), .Y(n5878) );
  AND2X1 U2900 ( .A(n3353), .B(n3461), .Y(n3476) );
  INVX1 U2902 ( .A(n3476), .Y(n5879) );
  AND2X1 U2904 ( .A(n3377), .B(n3461), .Y(n3488) );
  INVX1 U2906 ( .A(n3488), .Y(n5880) );
  AND2X1 U2908 ( .A(n3351), .B(n3496), .Y(n3510) );
  INVX1 U2910 ( .A(n3510), .Y(n5881) );
  AND2X1 U2912 ( .A(n3371), .B(n3496), .Y(n3520) );
  INVX1 U2914 ( .A(n3520), .Y(n5882) );
  AND2X1 U2916 ( .A(n3345), .B(n3530), .Y(n3541) );
  INVX1 U2918 ( .A(n3541), .Y(n5883) );
  AND2X1 U2920 ( .A(n3373), .B(n3530), .Y(n3555) );
  INVX1 U2922 ( .A(n3555), .Y(n5884) );
  AND2X1 U2924 ( .A(n3327), .B(n3565), .Y(n3567) );
  INVX1 U2926 ( .A(n3567), .Y(n5885) );
  AND2X1 U2929 ( .A(n3367), .B(n3565), .Y(n3587) );
  INVX1 U2931 ( .A(n3587), .Y(n5886) );
  AND2X1 U2933 ( .A(n3329), .B(n3600), .Y(n3603) );
  INVX1 U2935 ( .A(n3603), .Y(n5887) );
  AND2X1 U2937 ( .A(n3369), .B(n3600), .Y(n3623) );
  INVX1 U2939 ( .A(n3623), .Y(n5888) );
  AND2X1 U2941 ( .A(n3325), .B(n3635), .Y(n3636) );
  INVX1 U2943 ( .A(n3636), .Y(n5889) );
  AND2X1 U2945 ( .A(n3341), .B(n3635), .Y(n3644) );
  INVX1 U2947 ( .A(n3644), .Y(n5890) );
  AND2X1 U2949 ( .A(n3347), .B(n3670), .Y(n3682) );
  INVX1 U2951 ( .A(n3682), .Y(n5891) );
  AND2X1 U2953 ( .A(n3337), .B(n3704), .Y(n3711) );
  INVX1 U2955 ( .A(n3711), .Y(n5892) );
  AND2X1 U2957 ( .A(n3339), .B(n3738), .Y(n3746) );
  INVX1 U2959 ( .A(n3746), .Y(n5893) );
  AND2X1 U2961 ( .A(n3355), .B(n3772), .Y(n3788) );
  INVX1 U2963 ( .A(n3788), .Y(n5894) );
  AND2X1 U2965 ( .A(n3379), .B(n3772), .Y(n3800) );
  INVX1 U2967 ( .A(n3800), .Y(n5895) );
  AND2X1 U2969 ( .A(n3357), .B(n3806), .Y(n3823) );
  INVX1 U2971 ( .A(n3823), .Y(n5896) );
  AND2X1 U2973 ( .A(n3381), .B(n3806), .Y(n3835) );
  INVX1 U2975 ( .A(n3835), .Y(n5897) );
  AND2X1 U2977 ( .A(n3349), .B(n3840), .Y(n3853) );
  INVX1 U2979 ( .A(n3853), .Y(n5898) );
  AND2X1 U2981 ( .A(n3375), .B(n3840), .Y(n3866) );
  INVX1 U2983 ( .A(n3866), .Y(n5899) );
  AND2X1 U2985 ( .A(n3353), .B(n3874), .Y(n3889) );
  INVX1 U2987 ( .A(n3889), .Y(n5900) );
  AND2X1 U2989 ( .A(n3377), .B(n3874), .Y(n3901) );
  INVX1 U2991 ( .A(n3901), .Y(n5901) );
  AND2X1 U2993 ( .A(n3351), .B(n3908), .Y(n3922) );
  INVX1 U2996 ( .A(n3922), .Y(n5902) );
  AND2X1 U2998 ( .A(n3371), .B(n3908), .Y(n3932) );
  INVX1 U3000 ( .A(n3932), .Y(n5903) );
  AND2X1 U3002 ( .A(n3345), .B(n3943), .Y(n3954) );
  INVX1 U3004 ( .A(n3954), .Y(n5904) );
  AND2X1 U3006 ( .A(n3373), .B(n3943), .Y(n3968) );
  INVX1 U3008 ( .A(n3968), .Y(n5905) );
  AND2X1 U3010 ( .A(n3327), .B(n3977), .Y(n3979) );
  INVX1 U3012 ( .A(n3979), .Y(n5906) );
  AND2X1 U3014 ( .A(n3367), .B(n3977), .Y(n3999) );
  INVX1 U3016 ( .A(n3999), .Y(n5907) );
  AND2X1 U3018 ( .A(n3329), .B(n4011), .Y(n4014) );
  INVX1 U3020 ( .A(n4014), .Y(n5908) );
  AND2X1 U3022 ( .A(n3369), .B(n4011), .Y(n4034) );
  INVX1 U3024 ( .A(n4034), .Y(n5909) );
  AND2X1 U3026 ( .A(n3325), .B(n4045), .Y(n4046) );
  INVX1 U3028 ( .A(n4046), .Y(n5910) );
  AND2X1 U3030 ( .A(n3341), .B(n4045), .Y(n4054) );
  INVX1 U3032 ( .A(n4054), .Y(n5911) );
  AND2X1 U3034 ( .A(n3347), .B(n4079), .Y(n4091) );
  INVX1 U3036 ( .A(n4091), .Y(n5912) );
  AND2X1 U3038 ( .A(n3337), .B(n4113), .Y(n4120) );
  INVX1 U3040 ( .A(n4120), .Y(n5913) );
  AND2X1 U3042 ( .A(n3339), .B(n4147), .Y(n4155) );
  INVX1 U3044 ( .A(n4155), .Y(n5914) );
  AND2X1 U3046 ( .A(n3351), .B(n4181), .Y(n4195) );
  INVX1 U3048 ( .A(n4195), .Y(n5915) );
  AND2X1 U3050 ( .A(n3371), .B(n4181), .Y(n4205) );
  INVX1 U3052 ( .A(n4205), .Y(n5916) );
  AND2X1 U3054 ( .A(n3345), .B(n4216), .Y(n4227) );
  INVX1 U3056 ( .A(n4227), .Y(n5917) );
  AND2X1 U3058 ( .A(n3373), .B(n4216), .Y(n4241) );
  INVX1 U3060 ( .A(n4241), .Y(n5918) );
  AND2X1 U3063 ( .A(n3327), .B(n4250), .Y(n4252) );
  INVX1 U3065 ( .A(n4252), .Y(n5919) );
  AND2X1 U3067 ( .A(n3367), .B(n4250), .Y(n4272) );
  INVX1 U3069 ( .A(n4272), .Y(n5920) );
  AND2X1 U3071 ( .A(n3329), .B(n4284), .Y(n4287) );
  INVX1 U3073 ( .A(n4287), .Y(n5921) );
  AND2X1 U3075 ( .A(n3369), .B(n4284), .Y(n4307) );
  INVX1 U3077 ( .A(n4307), .Y(n5922) );
  AND2X1 U3079 ( .A(n3325), .B(n4318), .Y(n4319) );
  INVX1 U3081 ( .A(n4319), .Y(n5923) );
  AND2X1 U3083 ( .A(n3341), .B(n4318), .Y(n4327) );
  INVX1 U3085 ( .A(n4327), .Y(n5924) );
  AND2X1 U3087 ( .A(n3347), .B(n4352), .Y(n4364) );
  INVX1 U3089 ( .A(n4364), .Y(n5925) );
  AND2X1 U3091 ( .A(n3337), .B(n4386), .Y(n4393) );
  INVX1 U3093 ( .A(n4393), .Y(n5926) );
  AND2X1 U3095 ( .A(n3339), .B(n4420), .Y(n4428) );
  INVX1 U3097 ( .A(n4428), .Y(n5927) );
  AND2X1 U3099 ( .A(n3353), .B(n3323), .Y(n3352) );
  INVX1 U3101 ( .A(n3352), .Y(n5928) );
  AND2X1 U3103 ( .A(n3377), .B(n3323), .Y(n3376) );
  INVX1 U3105 ( .A(n3376), .Y(n5929) );
  AND2X1 U3107 ( .A(n3349), .B(n3391), .Y(n3404) );
  INVX1 U3109 ( .A(n3404), .Y(n5930) );
  AND2X1 U3111 ( .A(n3375), .B(n3391), .Y(n3417) );
  INVX1 U3113 ( .A(n3417), .Y(n5931) );
  AND2X1 U3115 ( .A(n3357), .B(n3426), .Y(n3443) );
  INVX1 U3117 ( .A(n3443), .Y(n5932) );
  AND2X1 U3119 ( .A(n3381), .B(n3426), .Y(n3455) );
  INVX1 U3121 ( .A(n3455), .Y(n5933) );
  AND2X1 U3123 ( .A(n3355), .B(n3461), .Y(n3477) );
  INVX1 U3125 ( .A(n3477), .Y(n5934) );
  AND2X1 U3127 ( .A(n3379), .B(n3461), .Y(n3489) );
  INVX1 U3130 ( .A(n3489), .Y(n5935) );
  AND2X1 U3132 ( .A(n3329), .B(n3496), .Y(n3499) );
  INVX1 U3134 ( .A(n3499), .Y(n5936) );
  AND2X1 U3136 ( .A(n3369), .B(n3496), .Y(n3519) );
  INVX1 U3138 ( .A(n3519), .Y(n5937) );
  AND2X1 U3140 ( .A(n3327), .B(n3530), .Y(n3532) );
  INVX1 U3142 ( .A(n3532), .Y(n5938) );
  AND2X1 U3144 ( .A(n3367), .B(n3530), .Y(n3552) );
  INVX1 U3146 ( .A(n3552), .Y(n5939) );
  AND2X1 U3148 ( .A(n3345), .B(n3565), .Y(n3576) );
  INVX1 U3150 ( .A(n3576), .Y(n5940) );
  AND2X1 U3152 ( .A(n3373), .B(n3565), .Y(n3590) );
  INVX1 U3154 ( .A(n3590), .Y(n5941) );
  AND2X1 U3156 ( .A(n3351), .B(n3600), .Y(n3614) );
  INVX1 U3158 ( .A(n3614), .Y(n5942) );
  AND2X1 U3160 ( .A(n3371), .B(n3600), .Y(n3624) );
  INVX1 U3162 ( .A(n3624), .Y(n5943) );
  AND2X1 U3164 ( .A(n3339), .B(n3635), .Y(n3643) );
  INVX1 U3166 ( .A(n3643), .Y(n5944) );
  AND2X1 U3168 ( .A(n3337), .B(n3670), .Y(n3677) );
  INVX1 U3170 ( .A(n3677), .Y(n5945) );
  AND2X1 U3172 ( .A(n3347), .B(n3704), .Y(n3716) );
  INVX1 U3174 ( .A(n3716), .Y(n5946) );
  AND2X1 U3176 ( .A(n3325), .B(n3738), .Y(n3739) );
  INVX1 U3178 ( .A(n3739), .Y(n5947) );
  AND2X1 U3180 ( .A(n3341), .B(n3738), .Y(n3747) );
  INVX1 U3182 ( .A(n3747), .Y(n5948) );
  AND2X1 U3184 ( .A(n3353), .B(n3772), .Y(n3787) );
  INVX1 U3186 ( .A(n3787), .Y(n5949) );
  AND2X1 U3188 ( .A(n3377), .B(n3772), .Y(n3799) );
  INVX1 U3190 ( .A(n3799), .Y(n5950) );
  AND2X1 U3192 ( .A(n3349), .B(n3806), .Y(n3819) );
  INVX1 U3194 ( .A(n3819), .Y(n5951) );
  AND2X1 U3197 ( .A(n3375), .B(n3806), .Y(n3832) );
  INVX1 U3199 ( .A(n3832), .Y(n5952) );
  AND2X1 U3201 ( .A(n3357), .B(n3840), .Y(n3857) );
  INVX1 U3203 ( .A(n3857), .Y(n5953) );
  AND2X1 U3205 ( .A(n3381), .B(n3840), .Y(n3869) );
  INVX1 U3207 ( .A(n3869), .Y(n5954) );
  AND2X1 U3209 ( .A(n3355), .B(n3874), .Y(n3890) );
  INVX1 U3211 ( .A(n3890), .Y(n5955) );
  AND2X1 U3213 ( .A(n3379), .B(n3874), .Y(n3902) );
  INVX1 U3215 ( .A(n3902), .Y(n5956) );
  AND2X1 U3217 ( .A(n3329), .B(n3908), .Y(n3911) );
  INVX1 U3219 ( .A(n3911), .Y(n5957) );
  AND2X1 U3221 ( .A(n3369), .B(n3908), .Y(n3931) );
  INVX1 U3223 ( .A(n3931), .Y(n5958) );
  AND2X1 U3225 ( .A(n3327), .B(n3943), .Y(n3945) );
  INVX1 U3227 ( .A(n3945), .Y(n5959) );
  AND2X1 U3229 ( .A(n3367), .B(n3943), .Y(n3965) );
  INVX1 U3231 ( .A(n3965), .Y(n5960) );
  AND2X1 U3233 ( .A(n3345), .B(n3977), .Y(n3988) );
  INVX1 U3235 ( .A(n3988), .Y(n5961) );
  AND2X1 U3237 ( .A(n3373), .B(n3977), .Y(n4002) );
  INVX1 U3239 ( .A(n4002), .Y(n5962) );
  AND2X1 U3241 ( .A(n3351), .B(n4011), .Y(n4025) );
  INVX1 U3243 ( .A(n4025), .Y(n5963) );
  AND2X1 U3245 ( .A(n3371), .B(n4011), .Y(n4035) );
  INVX1 U3247 ( .A(n4035), .Y(n5964) );
  AND2X1 U3249 ( .A(n3339), .B(n4045), .Y(n4053) );
  INVX1 U3251 ( .A(n4053), .Y(n5965) );
  AND2X1 U3253 ( .A(n3337), .B(n4079), .Y(n4086) );
  INVX1 U3255 ( .A(n4086), .Y(n5966) );
  AND2X1 U3257 ( .A(n3347), .B(n4113), .Y(n4125) );
  INVX1 U3259 ( .A(n4125), .Y(n5967) );
  AND2X1 U3261 ( .A(n3325), .B(n4147), .Y(n4148) );
  INVX1 U3264 ( .A(n4148), .Y(n5968) );
  AND2X1 U3266 ( .A(n3341), .B(n4147), .Y(n4156) );
  INVX1 U3268 ( .A(n4156), .Y(n5969) );
  AND2X1 U3270 ( .A(n3329), .B(n4181), .Y(n4184) );
  INVX1 U3272 ( .A(n4184), .Y(n5970) );
  AND2X1 U3274 ( .A(n3369), .B(n4181), .Y(n4204) );
  INVX1 U3276 ( .A(n4204), .Y(n5971) );
  AND2X1 U3278 ( .A(n3327), .B(n4216), .Y(n4218) );
  INVX1 U3280 ( .A(n4218), .Y(n5972) );
  AND2X1 U3282 ( .A(n3367), .B(n4216), .Y(n4238) );
  INVX1 U3284 ( .A(n4238), .Y(n5973) );
  AND2X1 U3286 ( .A(n3345), .B(n4250), .Y(n4261) );
  INVX1 U3288 ( .A(n4261), .Y(n5974) );
  AND2X1 U3290 ( .A(n3373), .B(n4250), .Y(n4275) );
  INVX1 U3292 ( .A(n4275), .Y(n5975) );
  AND2X1 U3294 ( .A(n3351), .B(n4284), .Y(n4298) );
  INVX1 U3296 ( .A(n4298), .Y(n5976) );
  AND2X1 U3298 ( .A(n3371), .B(n4284), .Y(n4308) );
  INVX1 U3300 ( .A(n4308), .Y(n5977) );
  AND2X1 U3302 ( .A(n3339), .B(n4318), .Y(n4326) );
  INVX1 U3304 ( .A(n4326), .Y(n5978) );
  AND2X1 U3306 ( .A(n3337), .B(n4352), .Y(n4359) );
  INVX1 U3308 ( .A(n4359), .Y(n5979) );
  AND2X1 U3310 ( .A(n3347), .B(n4386), .Y(n4398) );
  INVX1 U3312 ( .A(n4398), .Y(n5980) );
  AND2X1 U3314 ( .A(n3325), .B(n4420), .Y(n4421) );
  INVX1 U3316 ( .A(n4421), .Y(n5981) );
  AND2X1 U3318 ( .A(n3341), .B(n4420), .Y(n4429) );
  INVX1 U3320 ( .A(n4429), .Y(n5982) );
  AND2X1 U3322 ( .A(n3349), .B(n3323), .Y(n3348) );
  INVX1 U3324 ( .A(n3348), .Y(n5983) );
  AND2X1 U3326 ( .A(n3375), .B(n3323), .Y(n3374) );
  INVX1 U3328 ( .A(n3374), .Y(n5984) );
  AND2X1 U3331 ( .A(n3353), .B(n3391), .Y(n3406) );
  INVX1 U3333 ( .A(n3406), .Y(n5985) );
  AND2X1 U3335 ( .A(n3377), .B(n3391), .Y(n3418) );
  INVX1 U3337 ( .A(n3418), .Y(n5986) );
  AND2X1 U3339 ( .A(n3355), .B(n3426), .Y(n3442) );
  INVX1 U3341 ( .A(n3442), .Y(n5987) );
  AND2X1 U3343 ( .A(n3379), .B(n3426), .Y(n3454) );
  INVX1 U3345 ( .A(n3454), .Y(n5988) );
  AND2X1 U3347 ( .A(n3357), .B(n3461), .Y(n3478) );
  INVX1 U3349 ( .A(n3478), .Y(n5989) );
  AND2X1 U3351 ( .A(n3381), .B(n3461), .Y(n3490) );
  INVX1 U3353 ( .A(n3490), .Y(n5990) );
  AND2X1 U3355 ( .A(n3327), .B(n3496), .Y(n3498) );
  INVX1 U3357 ( .A(n3498), .Y(n5991) );
  AND2X1 U3359 ( .A(n3367), .B(n3496), .Y(n3518) );
  INVX1 U3361 ( .A(n3518), .Y(n5992) );
  AND2X1 U3363 ( .A(n3329), .B(n3530), .Y(n3533) );
  INVX1 U3365 ( .A(n3533), .Y(n5993) );
  AND2X1 U3367 ( .A(n3369), .B(n3530), .Y(n3553) );
  INVX1 U3369 ( .A(n3553), .Y(n5994) );
  AND2X1 U3371 ( .A(n3351), .B(n3565), .Y(n3579) );
  INVX1 U3373 ( .A(n3579), .Y(n5995) );
  AND2X1 U3375 ( .A(n3371), .B(n3565), .Y(n3589) );
  INVX1 U3377 ( .A(n3589), .Y(n5996) );
  AND2X1 U3379 ( .A(n3345), .B(n3600), .Y(n3611) );
  INVX1 U3381 ( .A(n3611), .Y(n5997) );
  AND2X1 U3383 ( .A(n3373), .B(n3600), .Y(n3625) );
  INVX1 U3385 ( .A(n3625), .Y(n5998) );
  AND2X1 U3387 ( .A(n3337), .B(n3635), .Y(n3642) );
  INVX1 U3389 ( .A(n3642), .Y(n5999) );
  AND2X1 U3391 ( .A(n3339), .B(n3670), .Y(n3678) );
  INVX1 U3393 ( .A(n3678), .Y(n6000) );
  AND2X1 U3395 ( .A(n3325), .B(n3704), .Y(n3705) );
  INVX1 U3399 ( .A(n3705), .Y(n6001) );
  AND2X1 U3401 ( .A(n3341), .B(n3704), .Y(n3713) );
  INVX1 U3403 ( .A(n3713), .Y(n6002) );
  AND2X1 U3405 ( .A(n3347), .B(n3738), .Y(n3750) );
  INVX1 U3407 ( .A(n3750), .Y(n6003) );
  AND2X1 U3409 ( .A(n3349), .B(n3772), .Y(n3785) );
  INVX1 U3411 ( .A(n3785), .Y(n6004) );
  AND2X1 U3413 ( .A(n3375), .B(n3772), .Y(n3798) );
  INVX1 U3415 ( .A(n3798), .Y(n6005) );
  AND2X1 U3417 ( .A(n3353), .B(n3806), .Y(n3821) );
  INVX1 U3419 ( .A(n3821), .Y(n6006) );
  AND2X1 U3421 ( .A(n3377), .B(n3806), .Y(n3833) );
  INVX1 U3423 ( .A(n3833), .Y(n6007) );
  AND2X1 U3425 ( .A(n3355), .B(n3840), .Y(n3856) );
  INVX1 U3427 ( .A(n3856), .Y(n6008) );
  AND2X1 U3429 ( .A(n3379), .B(n3840), .Y(n3868) );
  INVX1 U3431 ( .A(n3868), .Y(n6009) );
  AND2X1 U3433 ( .A(n3357), .B(n3874), .Y(n3891) );
  INVX1 U3435 ( .A(n3891), .Y(n6010) );
  AND2X1 U3437 ( .A(n3381), .B(n3874), .Y(n3903) );
  INVX1 U3439 ( .A(n3903), .Y(n6011) );
  AND2X1 U3441 ( .A(n3327), .B(n3908), .Y(n3910) );
  INVX1 U3443 ( .A(n3910), .Y(n6012) );
  AND2X1 U3445 ( .A(n3367), .B(n3908), .Y(n3930) );
  INVX1 U3447 ( .A(n3930), .Y(n6013) );
  AND2X1 U3449 ( .A(n3329), .B(n3943), .Y(n3946) );
  INVX1 U3451 ( .A(n3946), .Y(n6014) );
  AND2X1 U3453 ( .A(n3369), .B(n3943), .Y(n3966) );
  INVX1 U3455 ( .A(n3966), .Y(n6015) );
  AND2X1 U3457 ( .A(n3351), .B(n3977), .Y(n3991) );
  INVX1 U3459 ( .A(n3991), .Y(n6016) );
  AND2X1 U3461 ( .A(n3371), .B(n3977), .Y(n4001) );
  INVX1 U3463 ( .A(n4001), .Y(n6017) );
  AND2X1 U3466 ( .A(n3345), .B(n4011), .Y(n4022) );
  INVX1 U3468 ( .A(n4022), .Y(n6018) );
  AND2X1 U3470 ( .A(n3373), .B(n4011), .Y(n4036) );
  INVX1 U3472 ( .A(n4036), .Y(n6019) );
  AND2X1 U3474 ( .A(n3337), .B(n4045), .Y(n4052) );
  INVX1 U3476 ( .A(n4052), .Y(n6020) );
  AND2X1 U3478 ( .A(n3339), .B(n4079), .Y(n4087) );
  INVX1 U3480 ( .A(n4087), .Y(n6021) );
  AND2X1 U3482 ( .A(n3325), .B(n4113), .Y(n4114) );
  INVX1 U3484 ( .A(n4114), .Y(n6022) );
  AND2X1 U3486 ( .A(n3341), .B(n4113), .Y(n4122) );
  INVX1 U3488 ( .A(n4122), .Y(n6023) );
  AND2X1 U3490 ( .A(n3347), .B(n4147), .Y(n4159) );
  INVX1 U3492 ( .A(n4159), .Y(n6024) );
  AND2X1 U3494 ( .A(n3327), .B(n4181), .Y(n4183) );
  INVX1 U3496 ( .A(n4183), .Y(n6025) );
  AND2X1 U3498 ( .A(n3367), .B(n4181), .Y(n4203) );
  INVX1 U3500 ( .A(n4203), .Y(n6026) );
  AND2X1 U3502 ( .A(n3329), .B(n4216), .Y(n4219) );
  INVX1 U3504 ( .A(n4219), .Y(n6027) );
  AND2X1 U3506 ( .A(n3369), .B(n4216), .Y(n4239) );
  INVX1 U3508 ( .A(n4239), .Y(n6028) );
  AND2X1 U3510 ( .A(n3351), .B(n4250), .Y(n4264) );
  INVX1 U3512 ( .A(n4264), .Y(n6029) );
  AND2X1 U3514 ( .A(n3371), .B(n4250), .Y(n4274) );
  INVX1 U3516 ( .A(n4274), .Y(n6030) );
  AND2X1 U3518 ( .A(n3345), .B(n4284), .Y(n4295) );
  INVX1 U3520 ( .A(n4295), .Y(n6031) );
  AND2X1 U3522 ( .A(n3373), .B(n4284), .Y(n4309) );
  INVX1 U3524 ( .A(n4309), .Y(n6032) );
  AND2X1 U3526 ( .A(n3337), .B(n4318), .Y(n4325) );
  INVX1 U3528 ( .A(n4325), .Y(n6033) );
  AND2X1 U3530 ( .A(n3339), .B(n4352), .Y(n4360) );
  INVX1 U3533 ( .A(n4360), .Y(n6034) );
  AND2X1 U3535 ( .A(n3325), .B(n4386), .Y(n4387) );
  INVX1 U3537 ( .A(n4387), .Y(n6035) );
  AND2X1 U3539 ( .A(n3341), .B(n4386), .Y(n4395) );
  INVX1 U3541 ( .A(n4395), .Y(n6036) );
  AND2X1 U3543 ( .A(n3347), .B(n4420), .Y(n4432) );
  INVX1 U3545 ( .A(n4432), .Y(n6037) );
  AND2X1 U3547 ( .A(n3343), .B(n3323), .Y(n3342) );
  INVX1 U3549 ( .A(n3342), .Y(n6038) );
  AND2X1 U3551 ( .A(n3365), .B(n3323), .Y(n3364) );
  INVX1 U3553 ( .A(n3364), .Y(n6039) );
  AND2X1 U3555 ( .A(n3389), .B(n3323), .Y(n3388) );
  INVX1 U3557 ( .A(n3388), .Y(n6040) );
  AND2X1 U3559 ( .A(n3363), .B(n3391), .Y(n3411) );
  INVX1 U3561 ( .A(n3411), .Y(n6041) );
  AND2X1 U3563 ( .A(n3387), .B(n3391), .Y(n3423) );
  INVX1 U3565 ( .A(n3423), .Y(n6042) );
  AND2X1 U3567 ( .A(n3361), .B(n3426), .Y(n3445) );
  INVX1 U3569 ( .A(n3445), .Y(n6043) );
  AND2X1 U3571 ( .A(n3385), .B(n3426), .Y(n3457) );
  INVX1 U3573 ( .A(n3457), .Y(n6044) );
  AND2X1 U3575 ( .A(n3359), .B(n3461), .Y(n3479) );
  INVX1 U3577 ( .A(n3479), .Y(n6045) );
  AND2X1 U3579 ( .A(n3383), .B(n3461), .Y(n3491) );
  INVX1 U3581 ( .A(n3491), .Y(n6046) );
  AND2X1 U3583 ( .A(n3347), .B(n3496), .Y(n3508) );
  INVX1 U3585 ( .A(n3508), .Y(n6047) );
  AND2X1 U3587 ( .A(n3325), .B(n3530), .Y(n3531) );
  INVX1 U3589 ( .A(n3531), .Y(n6048) );
  AND2X1 U3591 ( .A(n3341), .B(n3530), .Y(n3539) );
  INVX1 U3593 ( .A(n3539), .Y(n6049) );
  AND2X1 U3595 ( .A(n3339), .B(n3565), .Y(n3573) );
  INVX1 U3597 ( .A(n3573), .Y(n6050) );
  AND2X1 U3600 ( .A(n3337), .B(n3600), .Y(n3607) );
  INVX1 U3602 ( .A(n3607), .Y(n6051) );
  AND2X1 U3604 ( .A(n3345), .B(n3635), .Y(n3646) );
  INVX1 U3606 ( .A(n3646), .Y(n6052) );
  AND2X1 U3608 ( .A(n3373), .B(n3635), .Y(n3660) );
  INVX1 U3610 ( .A(n3660), .Y(n6053) );
  AND2X1 U3612 ( .A(n3351), .B(n3670), .Y(n3684) );
  INVX1 U3614 ( .A(n3684), .Y(n6054) );
  AND2X1 U3616 ( .A(n3371), .B(n3670), .Y(n3694) );
  INVX1 U3618 ( .A(n3694), .Y(n6055) );
  AND2X1 U3620 ( .A(n3329), .B(n3704), .Y(n3707) );
  INVX1 U3622 ( .A(n3707), .Y(n6056) );
  AND2X1 U3624 ( .A(n3369), .B(n3704), .Y(n3727) );
  INVX1 U3626 ( .A(n3727), .Y(n6057) );
  AND2X1 U3628 ( .A(n3327), .B(n3738), .Y(n3740) );
  INVX1 U3630 ( .A(n3740), .Y(n6058) );
  AND2X1 U3632 ( .A(n3367), .B(n3738), .Y(n3760) );
  INVX1 U3634 ( .A(n3760), .Y(n6059) );
  AND2X1 U3636 ( .A(n3343), .B(n3772), .Y(n3782) );
  INVX1 U3638 ( .A(n3782), .Y(n6060) );
  AND2X1 U3640 ( .A(n3365), .B(n3772), .Y(n3793) );
  INVX1 U3642 ( .A(n3793), .Y(n6061) );
  AND2X1 U3644 ( .A(n3389), .B(n3772), .Y(n3805) );
  INVX1 U3646 ( .A(n3805), .Y(n6062) );
  AND2X1 U3648 ( .A(n3363), .B(n3806), .Y(n3826) );
  INVX1 U3650 ( .A(n3826), .Y(n6063) );
  AND2X1 U3652 ( .A(n3387), .B(n3806), .Y(n3838) );
  INVX1 U3654 ( .A(n3838), .Y(n6064) );
  AND2X1 U3656 ( .A(n3361), .B(n3840), .Y(n3859) );
  INVX1 U3658 ( .A(n3859), .Y(n6065) );
  AND2X1 U3660 ( .A(n3385), .B(n3840), .Y(n3871) );
  INVX1 U3662 ( .A(n3871), .Y(n6066) );
  AND2X1 U3664 ( .A(n3359), .B(n3874), .Y(n3892) );
  INVX1 U3667 ( .A(n3892), .Y(n6067) );
  AND2X1 U3669 ( .A(n3383), .B(n3874), .Y(n3904) );
  INVX1 U3671 ( .A(n3904), .Y(n6068) );
  AND2X1 U3673 ( .A(n3347), .B(n3908), .Y(n3920) );
  INVX1 U3675 ( .A(n3920), .Y(n6069) );
  AND2X1 U3677 ( .A(n3325), .B(n3943), .Y(n3944) );
  INVX1 U3679 ( .A(n3944), .Y(n6070) );
  AND2X1 U3681 ( .A(n3341), .B(n3943), .Y(n3952) );
  INVX1 U3683 ( .A(n3952), .Y(n6071) );
  AND2X1 U3685 ( .A(n3339), .B(n3977), .Y(n3985) );
  INVX1 U3687 ( .A(n3985), .Y(n6072) );
  AND2X1 U3689 ( .A(n3337), .B(n4011), .Y(n4018) );
  INVX1 U3691 ( .A(n4018), .Y(n6073) );
  AND2X1 U3693 ( .A(n3345), .B(n4045), .Y(n4056) );
  INVX1 U3695 ( .A(n4056), .Y(n6074) );
  AND2X1 U3697 ( .A(n3373), .B(n4045), .Y(n4070) );
  INVX1 U3699 ( .A(n4070), .Y(n6075) );
  AND2X1 U3701 ( .A(n3351), .B(n4079), .Y(n4093) );
  INVX1 U3703 ( .A(n4093), .Y(n6076) );
  AND2X1 U3705 ( .A(n3371), .B(n4079), .Y(n4103) );
  INVX1 U3707 ( .A(n4103), .Y(n6077) );
  AND2X1 U3709 ( .A(n3329), .B(n4113), .Y(n4116) );
  INVX1 U3711 ( .A(n4116), .Y(n6078) );
  AND2X1 U3713 ( .A(n3369), .B(n4113), .Y(n4136) );
  INVX1 U3715 ( .A(n4136), .Y(n6079) );
  AND2X1 U3717 ( .A(n3327), .B(n4147), .Y(n4149) );
  INVX1 U3719 ( .A(n4149), .Y(n6080) );
  AND2X1 U3721 ( .A(n3367), .B(n4147), .Y(n4169) );
  INVX1 U3723 ( .A(n4169), .Y(n6081) );
  AND2X1 U3725 ( .A(n3347), .B(n4181), .Y(n4193) );
  INVX1 U3727 ( .A(n4193), .Y(n6082) );
  AND2X1 U3729 ( .A(n3325), .B(n4216), .Y(n4217) );
  INVX1 U3731 ( .A(n4217), .Y(n6083) );
  AND2X1 U3734 ( .A(n3341), .B(n4216), .Y(n4225) );
  INVX1 U3736 ( .A(n4225), .Y(n6084) );
  AND2X1 U3738 ( .A(n3339), .B(n4250), .Y(n4258) );
  INVX1 U3740 ( .A(n4258), .Y(n6085) );
  AND2X1 U3742 ( .A(n3337), .B(n4284), .Y(n4291) );
  INVX1 U3744 ( .A(n4291), .Y(n6086) );
  AND2X1 U3746 ( .A(n3345), .B(n4318), .Y(n4329) );
  INVX1 U3748 ( .A(n4329), .Y(n6087) );
  AND2X1 U3750 ( .A(n3373), .B(n4318), .Y(n4343) );
  INVX1 U3752 ( .A(n4343), .Y(n6088) );
  AND2X1 U3754 ( .A(n3351), .B(n4352), .Y(n4366) );
  INVX1 U3756 ( .A(n4366), .Y(n6089) );
  AND2X1 U3758 ( .A(n3371), .B(n4352), .Y(n4376) );
  INVX1 U3760 ( .A(n4376), .Y(n6090) );
  AND2X1 U3762 ( .A(n3329), .B(n4386), .Y(n4389) );
  INVX1 U3764 ( .A(n4389), .Y(n6091) );
  AND2X1 U3766 ( .A(n3369), .B(n4386), .Y(n4409) );
  INVX1 U3768 ( .A(n4409), .Y(n6092) );
  AND2X1 U3770 ( .A(n3327), .B(n4420), .Y(n4422) );
  INVX1 U3772 ( .A(n4422), .Y(n6093) );
  AND2X1 U3774 ( .A(n3367), .B(n4420), .Y(n4442) );
  INVX1 U3776 ( .A(n4442), .Y(n6094) );
  AND2X1 U3778 ( .A(n3363), .B(n3323), .Y(n3362) );
  INVX1 U3780 ( .A(n3362), .Y(n6095) );
  AND2X1 U3782 ( .A(n3387), .B(n3323), .Y(n3386) );
  INVX1 U3784 ( .A(n3386), .Y(n6096) );
  AND2X1 U3786 ( .A(n3343), .B(n3391), .Y(n3401) );
  INVX1 U3788 ( .A(n3401), .Y(n6097) );
  AND2X1 U3790 ( .A(n3365), .B(n3391), .Y(n3412) );
  INVX1 U3792 ( .A(n3412), .Y(n6098) );
  AND2X1 U3794 ( .A(n3389), .B(n3391), .Y(n3424) );
  INVX1 U3796 ( .A(n3424), .Y(n6099) );
  AND2X1 U3798 ( .A(n3359), .B(n3426), .Y(n3444) );
  INVX1 U3801 ( .A(n3444), .Y(n6100) );
  AND2X1 U3803 ( .A(n3383), .B(n3426), .Y(n3456) );
  INVX1 U3805 ( .A(n3456), .Y(n6101) );
  AND2X1 U3807 ( .A(n3361), .B(n3461), .Y(n3480) );
  INVX1 U3809 ( .A(n3480), .Y(n6102) );
  AND2X1 U3811 ( .A(n3385), .B(n3461), .Y(n3492) );
  INVX1 U3813 ( .A(n3492), .Y(n6103) );
  AND2X1 U3815 ( .A(n3325), .B(n3496), .Y(n3497) );
  INVX1 U3817 ( .A(n3497), .Y(n6104) );
  AND2X1 U3819 ( .A(n3341), .B(n3496), .Y(n3505) );
  INVX1 U3821 ( .A(n3505), .Y(n6105) );
  AND2X1 U3823 ( .A(n3347), .B(n3530), .Y(n3542) );
  INVX1 U3825 ( .A(n3542), .Y(n6106) );
  AND2X1 U3827 ( .A(n3337), .B(n3565), .Y(n3572) );
  INVX1 U3829 ( .A(n3572), .Y(n6107) );
  AND2X1 U3831 ( .A(n3339), .B(n3600), .Y(n3608) );
  INVX1 U3833 ( .A(n3608), .Y(n6108) );
  AND2X1 U3835 ( .A(n3351), .B(n3635), .Y(n3649) );
  INVX1 U3837 ( .A(n3649), .Y(n6109) );
  AND2X1 U3839 ( .A(n3371), .B(n3635), .Y(n3659) );
  INVX1 U3841 ( .A(n3659), .Y(n6110) );
  AND2X1 U3843 ( .A(n3345), .B(n3670), .Y(n3681) );
  INVX1 U3845 ( .A(n3681), .Y(n6111) );
  AND2X1 U3847 ( .A(n3373), .B(n3670), .Y(n3695) );
  INVX1 U3849 ( .A(n3695), .Y(n6112) );
  AND2X1 U3851 ( .A(n3327), .B(n3704), .Y(n3706) );
  INVX1 U3853 ( .A(n3706), .Y(n6113) );
  AND2X1 U3855 ( .A(n3367), .B(n3704), .Y(n3726) );
  INVX1 U3857 ( .A(n3726), .Y(n6114) );
  AND2X1 U3859 ( .A(n3329), .B(n3738), .Y(n3741) );
  INVX1 U3861 ( .A(n3741), .Y(n6115) );
  AND2X1 U3863 ( .A(n3369), .B(n3738), .Y(n3761) );
  INVX1 U3865 ( .A(n3761), .Y(n6116) );
  AND2X1 U3868 ( .A(n3363), .B(n3772), .Y(n3792) );
  INVX1 U3870 ( .A(n3792), .Y(n6117) );
  AND2X1 U3872 ( .A(n3387), .B(n3772), .Y(n3804) );
  INVX1 U3874 ( .A(n3804), .Y(n6118) );
  AND2X1 U3876 ( .A(n3343), .B(n3806), .Y(n3816) );
  INVX1 U3878 ( .A(n3816), .Y(n6119) );
  AND2X1 U3880 ( .A(n3365), .B(n3806), .Y(n3827) );
  INVX1 U3882 ( .A(n3827), .Y(n6120) );
  AND2X1 U3884 ( .A(n3389), .B(n3806), .Y(n3839) );
  INVX1 U3886 ( .A(n3839), .Y(n6121) );
  AND2X1 U3888 ( .A(n3359), .B(n3840), .Y(n3858) );
  INVX1 U3890 ( .A(n3858), .Y(n6122) );
  AND2X1 U3892 ( .A(n3383), .B(n3840), .Y(n3870) );
  INVX1 U3894 ( .A(n3870), .Y(n6123) );
  AND2X1 U3896 ( .A(n3361), .B(n3874), .Y(n3893) );
  INVX1 U3898 ( .A(n3893), .Y(n6124) );
  AND2X1 U3900 ( .A(n3385), .B(n3874), .Y(n3905) );
  INVX1 U3902 ( .A(n3905), .Y(n6125) );
  AND2X1 U3904 ( .A(n3325), .B(n3908), .Y(n3909) );
  INVX1 U3906 ( .A(n3909), .Y(n6126) );
  AND2X1 U3908 ( .A(n3341), .B(n3908), .Y(n3917) );
  INVX1 U3910 ( .A(n3917), .Y(n6127) );
  AND2X1 U3912 ( .A(n3347), .B(n3943), .Y(n3955) );
  INVX1 U3914 ( .A(n3955), .Y(n6128) );
  AND2X1 U3916 ( .A(n3337), .B(n3977), .Y(n3984) );
  INVX1 U3918 ( .A(n3984), .Y(n6129) );
  AND2X1 U3920 ( .A(n3339), .B(n4011), .Y(n4019) );
  INVX1 U3922 ( .A(n4019), .Y(n6130) );
  AND2X1 U3924 ( .A(n3351), .B(n4045), .Y(n4059) );
  INVX1 U3926 ( .A(n4059), .Y(n6131) );
  AND2X1 U3928 ( .A(n3371), .B(n4045), .Y(n4069) );
  INVX1 U3930 ( .A(n4069), .Y(n6132) );
  AND2X1 U3932 ( .A(n3345), .B(n4079), .Y(n4090) );
  INVX1 U3936 ( .A(n4090), .Y(n6133) );
  AND2X1 U3938 ( .A(n3373), .B(n4079), .Y(n4104) );
  INVX1 U3940 ( .A(n4104), .Y(n6134) );
  AND2X1 U3942 ( .A(n3327), .B(n4113), .Y(n4115) );
  INVX1 U3944 ( .A(n4115), .Y(n6135) );
  AND2X1 U3946 ( .A(n3367), .B(n4113), .Y(n4135) );
  INVX1 U3948 ( .A(n4135), .Y(n6136) );
  AND2X1 U3950 ( .A(n3329), .B(n4147), .Y(n4150) );
  INVX1 U3952 ( .A(n4150), .Y(n6137) );
  AND2X1 U3954 ( .A(n3369), .B(n4147), .Y(n4170) );
  INVX1 U3956 ( .A(n4170), .Y(n6138) );
  AND2X1 U3958 ( .A(n3325), .B(n4181), .Y(n4182) );
  INVX1 U3960 ( .A(n4182), .Y(n6139) );
  AND2X1 U3962 ( .A(n3341), .B(n4181), .Y(n4190) );
  INVX1 U3964 ( .A(n4190), .Y(n6140) );
  AND2X1 U3966 ( .A(n3347), .B(n4216), .Y(n4228) );
  INVX1 U3968 ( .A(n4228), .Y(n6141) );
  AND2X1 U3970 ( .A(n3337), .B(n4250), .Y(n4257) );
  INVX1 U3972 ( .A(n4257), .Y(n6142) );
  AND2X1 U3974 ( .A(n3339), .B(n4284), .Y(n4292) );
  INVX1 U3976 ( .A(n4292), .Y(n6143) );
  AND2X1 U3978 ( .A(n3351), .B(n4318), .Y(n4332) );
  INVX1 U3980 ( .A(n4332), .Y(n6144) );
  AND2X1 U3982 ( .A(n3371), .B(n4318), .Y(n4342) );
  INVX1 U3984 ( .A(n4342), .Y(n6145) );
  AND2X1 U3986 ( .A(n3345), .B(n4352), .Y(n4363) );
  INVX1 U3988 ( .A(n4363), .Y(n6146) );
  AND2X1 U3990 ( .A(n3373), .B(n4352), .Y(n4377) );
  INVX1 U3992 ( .A(n4377), .Y(n6147) );
  AND2X1 U3994 ( .A(n3327), .B(n4386), .Y(n4388) );
  INVX1 U3996 ( .A(n4388), .Y(n6148) );
  AND2X1 U3998 ( .A(n3367), .B(n4386), .Y(n4408) );
  INVX1 U4000 ( .A(n4408), .Y(n6149) );
  AND2X1 U4004 ( .A(n3329), .B(n4420), .Y(n4423) );
  INVX1 U4006 ( .A(n4423), .Y(n6150) );
  AND2X1 U4008 ( .A(n3369), .B(n4420), .Y(n4443) );
  INVX1 U4010 ( .A(n4443), .Y(n6151) );
  AND2X1 U4012 ( .A(n3361), .B(n3323), .Y(n3360) );
  INVX1 U4014 ( .A(n3360), .Y(n6152) );
  AND2X1 U4016 ( .A(n3385), .B(n3323), .Y(n3384) );
  INVX1 U4018 ( .A(n3384), .Y(n6153) );
  AND2X1 U4020 ( .A(n3359), .B(n3391), .Y(n3409) );
  INVX1 U4022 ( .A(n3409), .Y(n6154) );
  AND2X1 U4024 ( .A(n3383), .B(n3391), .Y(n3421) );
  INVX1 U4026 ( .A(n3421), .Y(n6155) );
  AND2X1 U4028 ( .A(n3343), .B(n3426), .Y(n3436) );
  INVX1 U4030 ( .A(n3436), .Y(n6156) );
  AND2X1 U4032 ( .A(n3365), .B(n3426), .Y(n3447) );
  INVX1 U4034 ( .A(n3447), .Y(n6157) );
  AND2X1 U4036 ( .A(n3389), .B(n3426), .Y(n3459) );
  INVX1 U4038 ( .A(n3459), .Y(n6158) );
  AND2X1 U4040 ( .A(n3363), .B(n3461), .Y(n3481) );
  INVX1 U4042 ( .A(n3481), .Y(n6159) );
  AND2X1 U4044 ( .A(n3387), .B(n3461), .Y(n3493) );
  INVX1 U4046 ( .A(n3493), .Y(n6160) );
  AND2X1 U4048 ( .A(n3339), .B(n3496), .Y(n3504) );
  INVX1 U4050 ( .A(n3504), .Y(n6161) );
  AND2X1 U4052 ( .A(n3337), .B(n3530), .Y(n3537) );
  INVX1 U4054 ( .A(n3537), .Y(n6162) );
  AND2X1 U4056 ( .A(n3347), .B(n3565), .Y(n3577) );
  INVX1 U4058 ( .A(n3577), .Y(n6163) );
  AND2X1 U4060 ( .A(n3325), .B(n3600), .Y(n3601) );
  INVX1 U4062 ( .A(n3601), .Y(n6164) );
  AND2X1 U4064 ( .A(n3341), .B(n3600), .Y(n3609) );
  INVX1 U4066 ( .A(n3609), .Y(n6165) );
  AND2X1 U4068 ( .A(n3329), .B(n3635), .Y(n3638) );
  INVX1 U4072 ( .A(n3638), .Y(n6166) );
  AND2X1 U4074 ( .A(n3369), .B(n3635), .Y(n3658) );
  INVX1 U4076 ( .A(n3658), .Y(n6167) );
  AND2X1 U4078 ( .A(n3327), .B(n3670), .Y(n3672) );
  INVX1 U4080 ( .A(n3672), .Y(n6168) );
  AND2X1 U4082 ( .A(n3367), .B(n3670), .Y(n3692) );
  INVX1 U4084 ( .A(n3692), .Y(n6169) );
  AND2X1 U4086 ( .A(n3345), .B(n3704), .Y(n3715) );
  INVX1 U4088 ( .A(n3715), .Y(n6170) );
  AND2X1 U4090 ( .A(n3373), .B(n3704), .Y(n3729) );
  INVX1 U4092 ( .A(n3729), .Y(n6171) );
  AND2X1 U4094 ( .A(n3351), .B(n3738), .Y(n3752) );
  INVX1 U4096 ( .A(n3752), .Y(n6172) );
  AND2X1 U4098 ( .A(n3371), .B(n3738), .Y(n3762) );
  INVX1 U4100 ( .A(n3762), .Y(n6173) );
  AND2X1 U4102 ( .A(n3361), .B(n3772), .Y(n3791) );
  INVX1 U4104 ( .A(n3791), .Y(n6174) );
  AND2X1 U4106 ( .A(n3385), .B(n3772), .Y(n3803) );
  INVX1 U4108 ( .A(n3803), .Y(n6175) );
  AND2X1 U4110 ( .A(n3359), .B(n3806), .Y(n3824) );
  INVX1 U4112 ( .A(n3824), .Y(n6176) );
  AND2X1 U4114 ( .A(n3383), .B(n3806), .Y(n3836) );
  INVX1 U4116 ( .A(n3836), .Y(n6177) );
  AND2X1 U4118 ( .A(n3343), .B(n3840), .Y(n3850) );
  INVX1 U4120 ( .A(n3850), .Y(n6178) );
  AND2X1 U4122 ( .A(n3365), .B(n3840), .Y(n3861) );
  INVX1 U4124 ( .A(n3861), .Y(n6179) );
  AND2X1 U4126 ( .A(n3389), .B(n3840), .Y(n3873) );
  INVX1 U4128 ( .A(n3873), .Y(n6180) );
  AND2X1 U4130 ( .A(n3363), .B(n3874), .Y(n3894) );
  INVX1 U4132 ( .A(n3894), .Y(n6181) );
  AND2X1 U4134 ( .A(n3387), .B(n3874), .Y(n3906) );
  INVX1 U4136 ( .A(n3906), .Y(n6182) );
  AND2X1 U4140 ( .A(n3339), .B(n3908), .Y(n3916) );
  INVX1 U4142 ( .A(n3916), .Y(n6183) );
  AND2X1 U4144 ( .A(n3337), .B(n3943), .Y(n3950) );
  INVX1 U4146 ( .A(n3950), .Y(n6184) );
  AND2X1 U4148 ( .A(n3347), .B(n3977), .Y(n3989) );
  INVX1 U4150 ( .A(n3989), .Y(n6185) );
  AND2X1 U4152 ( .A(n3325), .B(n4011), .Y(n4012) );
  INVX1 U4154 ( .A(n4012), .Y(n6186) );
  AND2X1 U4156 ( .A(n3341), .B(n4011), .Y(n4020) );
  INVX1 U4158 ( .A(n4020), .Y(n6187) );
  AND2X1 U4160 ( .A(n3329), .B(n4045), .Y(n4048) );
  INVX1 U4162 ( .A(n4048), .Y(n6188) );
  AND2X1 U4164 ( .A(n3369), .B(n4045), .Y(n4068) );
  INVX1 U4166 ( .A(n4068), .Y(n6189) );
  AND2X1 U4168 ( .A(n3327), .B(n4079), .Y(n4081) );
  INVX1 U4170 ( .A(n4081), .Y(n6190) );
  AND2X1 U4172 ( .A(n3367), .B(n4079), .Y(n4101) );
  INVX1 U4174 ( .A(n4101), .Y(n6191) );
  AND2X1 U4176 ( .A(n3345), .B(n4113), .Y(n4124) );
  INVX1 U4178 ( .A(n4124), .Y(n6192) );
  AND2X1 U4180 ( .A(n3373), .B(n4113), .Y(n4138) );
  INVX1 U4182 ( .A(n4138), .Y(n6193) );
  AND2X1 U4184 ( .A(n3351), .B(n4147), .Y(n4161) );
  INVX1 U4186 ( .A(n4161), .Y(n6194) );
  AND2X1 U4188 ( .A(n3371), .B(n4147), .Y(n4171) );
  INVX1 U4190 ( .A(n4171), .Y(n6195) );
  AND2X1 U4192 ( .A(n3339), .B(n4181), .Y(n4189) );
  INVX1 U4194 ( .A(n4189), .Y(n6196) );
  AND2X1 U4196 ( .A(n3337), .B(n4216), .Y(n4223) );
  INVX1 U4198 ( .A(n4223), .Y(n6197) );
  AND2X1 U4200 ( .A(n3347), .B(n4250), .Y(n4262) );
  INVX1 U4202 ( .A(n4262), .Y(n6198) );
  AND2X1 U4204 ( .A(n3325), .B(n4284), .Y(n4285) );
  INVX1 U4208 ( .A(n4285), .Y(n6199) );
  AND2X1 U4210 ( .A(n3341), .B(n4284), .Y(n4293) );
  INVX1 U4212 ( .A(n4293), .Y(n6200) );
  AND2X1 U4214 ( .A(n3329), .B(n4318), .Y(n4321) );
  INVX1 U4216 ( .A(n4321), .Y(n6201) );
  AND2X1 U4218 ( .A(n3369), .B(n4318), .Y(n4341) );
  INVX1 U4220 ( .A(n4341), .Y(n6202) );
  AND2X1 U4222 ( .A(n3327), .B(n4352), .Y(n4354) );
  INVX1 U4224 ( .A(n4354), .Y(n6203) );
  AND2X1 U4226 ( .A(n3367), .B(n4352), .Y(n4374) );
  INVX1 U4228 ( .A(n4374), .Y(n6204) );
  AND2X1 U4230 ( .A(n3345), .B(n4386), .Y(n4397) );
  INVX1 U4232 ( .A(n4397), .Y(n6205) );
  AND2X1 U4234 ( .A(n3373), .B(n4386), .Y(n4411) );
  INVX1 U4236 ( .A(n4411), .Y(n6206) );
  AND2X1 U4238 ( .A(n3351), .B(n4420), .Y(n4434) );
  INVX1 U4240 ( .A(n4434), .Y(n6207) );
  AND2X1 U4242 ( .A(n3371), .B(n4420), .Y(n4444) );
  INVX1 U4244 ( .A(n4444), .Y(n6208) );
  AND2X1 U4246 ( .A(n3359), .B(n3323), .Y(n3358) );
  INVX1 U4248 ( .A(n3358), .Y(n6209) );
  AND2X1 U4250 ( .A(n3383), .B(n3323), .Y(n3382) );
  INVX1 U4252 ( .A(n3382), .Y(n6210) );
  AND2X1 U4254 ( .A(n3361), .B(n3391), .Y(n3410) );
  INVX1 U4256 ( .A(n3410), .Y(n6211) );
  AND2X1 U4258 ( .A(n3385), .B(n3391), .Y(n3422) );
  INVX1 U4260 ( .A(n3422), .Y(n6212) );
  AND2X1 U4262 ( .A(n3363), .B(n3426), .Y(n3446) );
  INVX1 U4264 ( .A(n3446), .Y(n6213) );
  AND2X1 U4266 ( .A(n3387), .B(n3426), .Y(n3458) );
  INVX1 U4268 ( .A(n3458), .Y(n6214) );
  AND2X1 U4270 ( .A(n3343), .B(n3461), .Y(n3471) );
  INVX1 U4272 ( .A(n3471), .Y(n6215) );
  AND2X1 U4276 ( .A(n3365), .B(n3461), .Y(n3482) );
  INVX1 U4278 ( .A(n3482), .Y(n6216) );
  AND2X1 U4280 ( .A(n3389), .B(n3461), .Y(n3494) );
  INVX1 U4282 ( .A(n3494), .Y(n6217) );
  AND2X1 U4284 ( .A(n3337), .B(n3496), .Y(n3503) );
  INVX1 U4286 ( .A(n3503), .Y(n6218) );
  AND2X1 U4288 ( .A(n3339), .B(n3530), .Y(n3538) );
  INVX1 U4290 ( .A(n3538), .Y(n6219) );
  AND2X1 U4292 ( .A(n3325), .B(n3565), .Y(n3566) );
  INVX1 U4294 ( .A(n3566), .Y(n6220) );
  AND2X1 U4296 ( .A(n3341), .B(n3565), .Y(n3574) );
  INVX1 U4298 ( .A(n3574), .Y(n6221) );
  AND2X1 U4300 ( .A(n3347), .B(n3600), .Y(n3612) );
  INVX1 U4302 ( .A(n3612), .Y(n6222) );
  AND2X1 U4304 ( .A(n3327), .B(n3635), .Y(n3637) );
  INVX1 U4306 ( .A(n3637), .Y(n6223) );
  AND2X1 U4308 ( .A(n3367), .B(n3635), .Y(n3657) );
  INVX1 U4310 ( .A(n3657), .Y(n6224) );
  AND2X1 U4312 ( .A(n3329), .B(n3670), .Y(n3673) );
  INVX1 U4314 ( .A(n3673), .Y(n6225) );
  AND2X1 U4316 ( .A(n3369), .B(n3670), .Y(n3693) );
  INVX1 U4318 ( .A(n3693), .Y(n6226) );
  AND2X1 U4320 ( .A(n3351), .B(n3704), .Y(n3718) );
  INVX1 U4322 ( .A(n3718), .Y(n6227) );
  AND2X1 U4324 ( .A(n3371), .B(n3704), .Y(n3728) );
  INVX1 U4326 ( .A(n3728), .Y(n6228) );
  AND2X1 U4328 ( .A(n3345), .B(n3738), .Y(n3749) );
  INVX1 U4330 ( .A(n3749), .Y(n6229) );
  AND2X1 U4332 ( .A(n3373), .B(n3738), .Y(n3763) );
  INVX1 U4334 ( .A(n3763), .Y(n6230) );
  AND2X1 U4336 ( .A(n3359), .B(n3772), .Y(n3790) );
  INVX1 U4338 ( .A(n3790), .Y(n6231) );
  AND2X1 U4340 ( .A(n3383), .B(n3772), .Y(n3802) );
  INVX1 U4344 ( .A(n3802), .Y(n6232) );
  AND2X1 U4346 ( .A(n3361), .B(n3806), .Y(n3825) );
  INVX1 U4348 ( .A(n3825), .Y(n6233) );
  AND2X1 U4350 ( .A(n3385), .B(n3806), .Y(n3837) );
  INVX1 U4352 ( .A(n3837), .Y(n6234) );
  AND2X1 U4354 ( .A(n3363), .B(n3840), .Y(n3860) );
  INVX1 U4356 ( .A(n3860), .Y(n6235) );
  AND2X1 U4358 ( .A(n3387), .B(n3840), .Y(n3872) );
  INVX1 U4360 ( .A(n3872), .Y(n6236) );
  AND2X1 U4362 ( .A(n3343), .B(n3874), .Y(n3884) );
  INVX1 U4364 ( .A(n3884), .Y(n6237) );
  AND2X1 U4366 ( .A(n3365), .B(n3874), .Y(n3895) );
  INVX1 U4368 ( .A(n3895), .Y(n6238) );
  AND2X1 U4370 ( .A(n3389), .B(n3874), .Y(n3907) );
  INVX1 U4372 ( .A(n3907), .Y(n6239) );
  AND2X1 U4374 ( .A(n3337), .B(n3908), .Y(n3915) );
  INVX1 U4376 ( .A(n3915), .Y(n6240) );
  AND2X1 U4378 ( .A(n3339), .B(n3943), .Y(n3951) );
  INVX1 U4380 ( .A(n3951), .Y(n6241) );
  AND2X1 U4382 ( .A(n3325), .B(n3977), .Y(n3978) );
  INVX1 U4384 ( .A(n3978), .Y(n6242) );
  AND2X1 U4386 ( .A(n3341), .B(n3977), .Y(n3986) );
  INVX1 U4388 ( .A(n3986), .Y(n6243) );
  AND2X1 U4390 ( .A(n3347), .B(n4011), .Y(n4023) );
  INVX1 U4392 ( .A(n4023), .Y(n6244) );
  AND2X1 U4394 ( .A(n3327), .B(n4045), .Y(n4047) );
  INVX1 U4396 ( .A(n4047), .Y(n6245) );
  AND2X1 U4398 ( .A(n3367), .B(n4045), .Y(n4067) );
  INVX1 U4400 ( .A(n4067), .Y(n6246) );
  AND2X1 U4402 ( .A(n3329), .B(n4079), .Y(n4082) );
  INVX1 U4404 ( .A(n4082), .Y(n6247) );
  AND2X1 U4406 ( .A(n3369), .B(n4079), .Y(n4102) );
  INVX1 U4408 ( .A(n4102), .Y(n6248) );
  AND2X1 U4412 ( .A(n3351), .B(n4113), .Y(n4127) );
  INVX1 U4414 ( .A(n4127), .Y(n6249) );
  AND2X1 U4416 ( .A(n3371), .B(n4113), .Y(n4137) );
  INVX1 U4418 ( .A(n4137), .Y(n6250) );
  AND2X1 U4420 ( .A(n3345), .B(n4147), .Y(n4158) );
  INVX1 U4422 ( .A(n4158), .Y(n6251) );
  AND2X1 U4424 ( .A(n3373), .B(n4147), .Y(n4172) );
  INVX1 U4426 ( .A(n4172), .Y(n6252) );
  AND2X1 U4428 ( .A(n3337), .B(n4181), .Y(n4188) );
  INVX1 U4430 ( .A(n4188), .Y(n6253) );
  AND2X1 U4432 ( .A(n3339), .B(n4216), .Y(n4224) );
  INVX1 U4434 ( .A(n4224), .Y(n6254) );
  AND2X1 U4436 ( .A(n3325), .B(n4250), .Y(n4251) );
  INVX1 U4438 ( .A(n4251), .Y(n6255) );
  AND2X1 U4440 ( .A(n3341), .B(n4250), .Y(n4259) );
  INVX1 U4442 ( .A(n4259), .Y(n6256) );
  AND2X1 U4444 ( .A(n3347), .B(n4284), .Y(n4296) );
  INVX1 U4446 ( .A(n4296), .Y(n6257) );
  AND2X1 U4448 ( .A(n3327), .B(n4318), .Y(n4320) );
  INVX1 U4450 ( .A(n4320), .Y(n6258) );
  AND2X1 U4452 ( .A(n3367), .B(n4318), .Y(n4340) );
  INVX1 U4454 ( .A(n4340), .Y(n6259) );
  AND2X1 U4456 ( .A(n3329), .B(n4352), .Y(n4355) );
  INVX1 U4458 ( .A(n4355), .Y(n6260) );
  AND2X1 U4460 ( .A(n3369), .B(n4352), .Y(n4375) );
  INVX1 U4462 ( .A(n4375), .Y(n6261) );
  AND2X1 U4464 ( .A(n3351), .B(n4386), .Y(n4400) );
  INVX1 U4466 ( .A(n4400), .Y(n6262) );
  AND2X1 U4468 ( .A(n3371), .B(n4386), .Y(n4410) );
  INVX1 U4470 ( .A(n4410), .Y(n6263) );
  AND2X1 U4472 ( .A(n3345), .B(n4420), .Y(n4431) );
  INVX1 U4474 ( .A(n4431), .Y(n6264) );
  AND2X1 U4476 ( .A(n3373), .B(n4420), .Y(n4445) );
  INVX1 U4495 ( .A(n4445), .Y(n6265) );
  BUFX2 U4496 ( .A(n3316), .Y(n6266) );
  AND2X1 U4497 ( .A(n3347), .B(n3323), .Y(n3346) );
  INVX1 U4498 ( .A(n3346), .Y(n6267) );
  AND2X1 U4499 ( .A(n3325), .B(n3391), .Y(n3392) );
  INVX1 U4500 ( .A(n3392), .Y(n6268) );
  AND2X1 U4501 ( .A(n3341), .B(n3391), .Y(n3400) );
  INVX1 U4502 ( .A(n3400), .Y(n6269) );
  AND2X1 U4503 ( .A(n3339), .B(n3426), .Y(n3434) );
  INVX1 U4504 ( .A(n3434), .Y(n6270) );
  AND2X1 U4505 ( .A(n3337), .B(n3461), .Y(n3468) );
  INVX1 U4506 ( .A(n3468), .Y(n6271) );
  AND2X1 U4507 ( .A(n3343), .B(n3496), .Y(n3506) );
  INVX1 U4508 ( .A(n3506), .Y(n6272) );
  AND2X1 U4509 ( .A(n3365), .B(n3496), .Y(n3517) );
  INVX1 U4510 ( .A(n3517), .Y(n6273) );
  AND2X1 U4511 ( .A(n3389), .B(n3496), .Y(n3529) );
  INVX1 U4512 ( .A(n3529), .Y(n6274) );
  AND2X1 U4513 ( .A(n3363), .B(n3530), .Y(n3550) );
  INVX1 U4514 ( .A(n3550), .Y(n6275) );
  AND2X1 U4515 ( .A(n3387), .B(n3530), .Y(n3562) );
  INVX1 U4516 ( .A(n3562), .Y(n6276) );
  AND2X1 U4517 ( .A(n3361), .B(n3565), .Y(n3584) );
  INVX1 U4518 ( .A(n3584), .Y(n6277) );
  AND2X1 U4519 ( .A(n3385), .B(n3565), .Y(n3596) );
  INVX1 U4520 ( .A(n3596), .Y(n6278) );
  AND2X1 U4521 ( .A(n3359), .B(n3600), .Y(n3618) );
  INVX1 U4522 ( .A(n3618), .Y(n6279) );
  AND2X1 U4523 ( .A(n3383), .B(n3600), .Y(n3630) );
  INVX1 U4524 ( .A(n3630), .Y(n6280) );
  AND2X1 U4525 ( .A(n3357), .B(n3635), .Y(n3652) );
  INVX1 U4526 ( .A(n3652), .Y(n6281) );
  AND2X1 U4527 ( .A(n3381), .B(n3635), .Y(n3664) );
  INVX1 U4528 ( .A(n3664), .Y(n6282) );
  AND2X1 U4529 ( .A(n3355), .B(n3670), .Y(n3686) );
  INVX1 U4530 ( .A(n3686), .Y(n6283) );
  AND2X1 U4531 ( .A(n3379), .B(n3670), .Y(n3698) );
  INVX1 U4532 ( .A(n3698), .Y(n6284) );
  AND2X1 U4533 ( .A(n3353), .B(n3704), .Y(n3719) );
  INVX1 U4534 ( .A(n3719), .Y(n6285) );
  AND2X1 U4535 ( .A(n3377), .B(n3704), .Y(n3731) );
  INVX1 U4536 ( .A(n3731), .Y(n6286) );
  AND2X1 U4537 ( .A(n3349), .B(n3738), .Y(n3751) );
  INVX1 U4538 ( .A(n3751), .Y(n6287) );
  AND2X1 U4539 ( .A(n3375), .B(n3738), .Y(n3764) );
  INVX1 U4540 ( .A(n3764), .Y(n6288) );
  AND2X1 U4541 ( .A(n3347), .B(n3772), .Y(n3784) );
  INVX1 U4542 ( .A(n3784), .Y(n6289) );
  AND2X1 U4543 ( .A(n3325), .B(n3806), .Y(n3807) );
  INVX1 U4544 ( .A(n3807), .Y(n6290) );
  AND2X1 U4545 ( .A(n3341), .B(n3806), .Y(n3815) );
  INVX1 U4546 ( .A(n3815), .Y(n6291) );
  AND2X1 U4547 ( .A(n3339), .B(n3840), .Y(n3848) );
  INVX1 U4548 ( .A(n3848), .Y(n6292) );
  AND2X1 U4549 ( .A(n3337), .B(n3874), .Y(n3881) );
  INVX1 U4550 ( .A(n3881), .Y(n6293) );
  AND2X1 U4551 ( .A(n3343), .B(n3908), .Y(n3918) );
  INVX1 U4552 ( .A(n3918), .Y(n6294) );
  AND2X1 U4553 ( .A(n3365), .B(n3908), .Y(n3929) );
  INVX1 U4554 ( .A(n3929), .Y(n6295) );
  AND2X1 U4555 ( .A(n3389), .B(n3908), .Y(n3941) );
  INVX1 U4556 ( .A(n3941), .Y(n6296) );
  AND2X1 U4557 ( .A(n3363), .B(n3943), .Y(n3963) );
  INVX1 U4558 ( .A(n3963), .Y(n6297) );
  AND2X1 U4559 ( .A(n3387), .B(n3943), .Y(n3975) );
  INVX1 U4560 ( .A(n3975), .Y(n6298) );
  AND2X1 U4561 ( .A(n3361), .B(n3977), .Y(n3996) );
  INVX1 U4562 ( .A(n3996), .Y(n6299) );
  AND2X1 U4563 ( .A(n3385), .B(n3977), .Y(n4008) );
  INVX1 U4564 ( .A(n4008), .Y(n6300) );
  AND2X1 U4565 ( .A(n3359), .B(n4011), .Y(n4029) );
  INVX1 U4566 ( .A(n4029), .Y(n6301) );
  AND2X1 U4567 ( .A(n3383), .B(n4011), .Y(n4041) );
  INVX1 U4568 ( .A(n4041), .Y(n6302) );
  AND2X1 U4569 ( .A(n3357), .B(n4045), .Y(n4062) );
  INVX1 U4570 ( .A(n4062), .Y(n6303) );
  AND2X1 U4571 ( .A(n3381), .B(n4045), .Y(n4074) );
  INVX1 U4572 ( .A(n4074), .Y(n6304) );
  AND2X1 U4573 ( .A(n3355), .B(n4079), .Y(n4095) );
  INVX1 U4574 ( .A(n4095), .Y(n6305) );
  AND2X1 U4575 ( .A(n3379), .B(n4079), .Y(n4107) );
  INVX1 U4576 ( .A(n4107), .Y(n6306) );
  AND2X1 U4577 ( .A(n3353), .B(n4113), .Y(n4128) );
  INVX1 U4578 ( .A(n4128), .Y(n6307) );
  AND2X1 U4579 ( .A(n3377), .B(n4113), .Y(n4140) );
  INVX1 U4580 ( .A(n4140), .Y(n6308) );
  AND2X1 U4581 ( .A(n3349), .B(n4147), .Y(n4160) );
  INVX1 U4582 ( .A(n4160), .Y(n6309) );
  AND2X1 U4583 ( .A(n3375), .B(n4147), .Y(n4173) );
  INVX1 U4584 ( .A(n4173), .Y(n6310) );
  AND2X1 U4585 ( .A(n3343), .B(n4181), .Y(n4191) );
  INVX1 U4586 ( .A(n4191), .Y(n6311) );
  AND2X1 U4587 ( .A(n3365), .B(n4181), .Y(n4202) );
  INVX1 U4588 ( .A(n4202), .Y(n6312) );
  AND2X1 U4589 ( .A(n3389), .B(n4181), .Y(n4214) );
  INVX1 U4590 ( .A(n4214), .Y(n6313) );
  AND2X1 U4591 ( .A(n3363), .B(n4216), .Y(n4236) );
  INVX1 U4592 ( .A(n4236), .Y(n6314) );
  AND2X1 U4593 ( .A(n3387), .B(n4216), .Y(n4248) );
  INVX1 U4594 ( .A(n4248), .Y(n6315) );
  AND2X1 U4595 ( .A(n3361), .B(n4250), .Y(n4269) );
  INVX1 U4596 ( .A(n4269), .Y(n6316) );
  AND2X1 U4597 ( .A(n3385), .B(n4250), .Y(n4281) );
  INVX1 U4598 ( .A(n4281), .Y(n6317) );
  AND2X1 U4599 ( .A(n3359), .B(n4284), .Y(n4302) );
  INVX1 U4600 ( .A(n4302), .Y(n6318) );
  AND2X1 U4601 ( .A(n3383), .B(n4284), .Y(n4314) );
  INVX1 U4602 ( .A(n4314), .Y(n6319) );
  AND2X1 U4603 ( .A(n3357), .B(n4318), .Y(n4335) );
  INVX1 U4604 ( .A(n4335), .Y(n6320) );
  AND2X1 U4605 ( .A(n3381), .B(n4318), .Y(n4347) );
  INVX1 U4606 ( .A(n4347), .Y(n6321) );
  AND2X1 U4607 ( .A(n3355), .B(n4352), .Y(n4368) );
  INVX1 U4608 ( .A(n4368), .Y(n6322) );
  AND2X1 U4609 ( .A(n3379), .B(n4352), .Y(n4380) );
  INVX1 U4610 ( .A(n4380), .Y(n6323) );
  AND2X1 U4611 ( .A(n3353), .B(n4386), .Y(n4401) );
  INVX1 U4612 ( .A(n4401), .Y(n6324) );
  AND2X1 U4613 ( .A(n3377), .B(n4386), .Y(n4413) );
  INVX1 U4614 ( .A(n4413), .Y(n6325) );
  AND2X1 U4615 ( .A(n3349), .B(n4420), .Y(n4433) );
  INVX1 U4616 ( .A(n4433), .Y(n6326) );
  AND2X1 U4617 ( .A(n3375), .B(n4420), .Y(n4446) );
  INVX1 U4618 ( .A(n4446), .Y(n6327) );
  BUFX2 U4619 ( .A(n3318), .Y(n6328) );
  AND2X1 U4620 ( .A(n3325), .B(n3323), .Y(n3324) );
  INVX1 U4621 ( .A(n3324), .Y(n6329) );
  AND2X1 U4622 ( .A(n3341), .B(n3323), .Y(n3340) );
  INVX1 U4623 ( .A(n3340), .Y(n6330) );
  AND2X1 U4624 ( .A(n3347), .B(n3391), .Y(n3403) );
  INVX1 U4625 ( .A(n3403), .Y(n6331) );
  AND2X1 U4626 ( .A(n3337), .B(n3426), .Y(n3433) );
  INVX1 U4627 ( .A(n3433), .Y(n6332) );
  AND2X1 U4628 ( .A(n3339), .B(n3461), .Y(n3469) );
  INVX1 U4629 ( .A(n3469), .Y(n6333) );
  AND2X1 U4630 ( .A(n3363), .B(n3496), .Y(n3516) );
  INVX1 U4631 ( .A(n3516), .Y(n6334) );
  AND2X1 U4632 ( .A(n3387), .B(n3496), .Y(n3528) );
  INVX1 U4633 ( .A(n3528), .Y(n6335) );
  AND2X1 U4634 ( .A(n3343), .B(n3530), .Y(n3540) );
  INVX1 U4635 ( .A(n3540), .Y(n6336) );
  AND2X1 U4636 ( .A(n3365), .B(n3530), .Y(n3551) );
  INVX1 U4637 ( .A(n3551), .Y(n6337) );
  AND2X1 U4638 ( .A(n3389), .B(n3530), .Y(n3563) );
  INVX1 U4639 ( .A(n3563), .Y(n6338) );
  AND2X1 U4640 ( .A(n3359), .B(n3565), .Y(n3583) );
  INVX1 U4641 ( .A(n3583), .Y(n6339) );
  AND2X1 U4642 ( .A(n3383), .B(n3565), .Y(n3595) );
  INVX1 U4643 ( .A(n3595), .Y(n6340) );
  AND2X1 U4644 ( .A(n3361), .B(n3600), .Y(n3619) );
  INVX1 U4645 ( .A(n3619), .Y(n6341) );
  AND2X1 U4646 ( .A(n3385), .B(n3600), .Y(n3631) );
  INVX1 U4647 ( .A(n3631), .Y(n6342) );
  AND2X1 U4648 ( .A(n3355), .B(n3635), .Y(n3651) );
  INVX1 U4649 ( .A(n3651), .Y(n6343) );
  AND2X1 U4650 ( .A(n3379), .B(n3635), .Y(n3663) );
  INVX1 U4651 ( .A(n3663), .Y(n6344) );
  AND2X1 U4652 ( .A(n3357), .B(n3670), .Y(n3687) );
  INVX1 U4653 ( .A(n3687), .Y(n6345) );
  AND2X1 U4654 ( .A(n3381), .B(n3670), .Y(n3699) );
  INVX1 U4655 ( .A(n3699), .Y(n6346) );
  AND2X1 U4656 ( .A(n3349), .B(n3704), .Y(n3717) );
  INVX1 U4657 ( .A(n3717), .Y(n6347) );
  AND2X1 U4658 ( .A(n3375), .B(n3704), .Y(n3730) );
  INVX1 U4659 ( .A(n3730), .Y(n6348) );
  AND2X1 U4660 ( .A(n3353), .B(n3738), .Y(n3753) );
  INVX1 U4661 ( .A(n3753), .Y(n6349) );
  AND2X1 U4662 ( .A(n3377), .B(n3738), .Y(n3765) );
  INVX1 U4663 ( .A(n3765), .Y(n6350) );
  AND2X1 U4664 ( .A(n3325), .B(n3772), .Y(n3773) );
  INVX1 U4665 ( .A(n3773), .Y(n6351) );
  AND2X1 U4666 ( .A(n3341), .B(n3772), .Y(n3781) );
  INVX1 U4667 ( .A(n3781), .Y(n6352) );
  AND2X1 U4668 ( .A(n3347), .B(n3806), .Y(n3818) );
  INVX1 U4669 ( .A(n3818), .Y(n6353) );
  AND2X1 U4670 ( .A(n3337), .B(n3840), .Y(n3847) );
  INVX1 U4671 ( .A(n3847), .Y(n6354) );
  AND2X1 U4672 ( .A(n3339), .B(n3874), .Y(n3882) );
  INVX1 U4673 ( .A(n3882), .Y(n6355) );
  AND2X1 U4674 ( .A(n3363), .B(n3908), .Y(n3928) );
  INVX1 U4675 ( .A(n3928), .Y(n6356) );
  AND2X1 U4676 ( .A(n3387), .B(n3908), .Y(n3940) );
  INVX1 U4677 ( .A(n3940), .Y(n6357) );
  AND2X1 U4678 ( .A(n3343), .B(n3943), .Y(n3953) );
  INVX1 U4679 ( .A(n3953), .Y(n6358) );
  AND2X1 U4680 ( .A(n3365), .B(n3943), .Y(n3964) );
  INVX1 U4681 ( .A(n3964), .Y(n6359) );
  AND2X1 U4682 ( .A(n3389), .B(n3943), .Y(n3976) );
  INVX1 U4683 ( .A(n3976), .Y(n6360) );
  AND2X1 U4684 ( .A(n3359), .B(n3977), .Y(n3995) );
  INVX1 U4685 ( .A(n3995), .Y(n6361) );
  AND2X1 U4686 ( .A(n3383), .B(n3977), .Y(n4007) );
  INVX1 U4687 ( .A(n4007), .Y(n6362) );
  AND2X1 U4688 ( .A(n3361), .B(n4011), .Y(n4030) );
  INVX1 U4689 ( .A(n4030), .Y(n6363) );
  AND2X1 U4690 ( .A(n3385), .B(n4011), .Y(n4042) );
  INVX1 U4691 ( .A(n4042), .Y(n6364) );
  AND2X1 U4692 ( .A(n3355), .B(n4045), .Y(n4061) );
  INVX1 U4693 ( .A(n4061), .Y(n6365) );
  AND2X1 U4694 ( .A(n3379), .B(n4045), .Y(n4073) );
  INVX1 U4695 ( .A(n4073), .Y(n6366) );
  AND2X1 U4696 ( .A(n3357), .B(n4079), .Y(n4096) );
  INVX1 U4697 ( .A(n4096), .Y(n6367) );
  AND2X1 U4698 ( .A(n3381), .B(n4079), .Y(n4108) );
  INVX1 U4699 ( .A(n4108), .Y(n6368) );
  AND2X1 U4700 ( .A(n3349), .B(n4113), .Y(n4126) );
  INVX1 U4701 ( .A(n4126), .Y(n6369) );
  AND2X1 U4702 ( .A(n3375), .B(n4113), .Y(n4139) );
  INVX1 U4703 ( .A(n4139), .Y(n6370) );
  AND2X1 U4704 ( .A(n3353), .B(n4147), .Y(n4162) );
  INVX1 U4705 ( .A(n4162), .Y(n6371) );
  AND2X1 U4706 ( .A(n3377), .B(n4147), .Y(n4174) );
  INVX1 U4707 ( .A(n4174), .Y(n6372) );
  AND2X1 U4708 ( .A(n3363), .B(n4181), .Y(n4201) );
  INVX1 U4709 ( .A(n4201), .Y(n6373) );
  AND2X1 U4710 ( .A(n3387), .B(n4181), .Y(n4213) );
  INVX1 U4711 ( .A(n4213), .Y(n6374) );
  AND2X1 U4712 ( .A(n3343), .B(n4216), .Y(n4226) );
  INVX1 U4713 ( .A(n4226), .Y(n6375) );
  AND2X1 U4714 ( .A(n3365), .B(n4216), .Y(n4237) );
  INVX1 U4715 ( .A(n4237), .Y(n6376) );
  AND2X1 U4716 ( .A(n3389), .B(n4216), .Y(n4249) );
  INVX1 U4717 ( .A(n4249), .Y(n6377) );
  AND2X1 U4718 ( .A(n3359), .B(n4250), .Y(n4268) );
  INVX1 U4719 ( .A(n4268), .Y(n6378) );
  AND2X1 U4720 ( .A(n3383), .B(n4250), .Y(n4280) );
  INVX1 U4721 ( .A(n4280), .Y(n6379) );
  AND2X1 U4722 ( .A(n3361), .B(n4284), .Y(n4303) );
  INVX1 U4723 ( .A(n4303), .Y(n6380) );
  AND2X1 U4724 ( .A(n3385), .B(n4284), .Y(n4315) );
  INVX1 U4725 ( .A(n4315), .Y(n6381) );
  AND2X1 U4726 ( .A(n3355), .B(n4318), .Y(n4334) );
  INVX1 U4727 ( .A(n4334), .Y(n6382) );
  AND2X1 U4728 ( .A(n3379), .B(n4318), .Y(n4346) );
  INVX1 U4729 ( .A(n4346), .Y(n6383) );
  AND2X1 U4730 ( .A(n3357), .B(n4352), .Y(n4369) );
  INVX1 U4731 ( .A(n4369), .Y(n6384) );
  AND2X1 U4732 ( .A(n3381), .B(n4352), .Y(n4381) );
  INVX1 U4733 ( .A(n4381), .Y(n6385) );
  AND2X1 U4734 ( .A(n3349), .B(n4386), .Y(n4399) );
  INVX1 U4735 ( .A(n4399), .Y(n6386) );
  AND2X1 U4736 ( .A(n3375), .B(n4386), .Y(n4412) );
  INVX1 U4737 ( .A(n4412), .Y(n6387) );
  AND2X1 U4738 ( .A(n3353), .B(n4420), .Y(n4435) );
  INVX1 U4739 ( .A(n4435), .Y(n6388) );
  AND2X1 U4740 ( .A(n3377), .B(n4420), .Y(n4447) );
  INVX1 U4741 ( .A(n4447), .Y(n6389) );
  BUFX2 U4742 ( .A(n4456), .Y(n6390) );
  BUFX2 U4743 ( .A(n4459), .Y(n6391) );
  AND2X1 U4744 ( .A(n3339), .B(n3323), .Y(n3338) );
  INVX1 U4745 ( .A(n3338), .Y(n6392) );
  AND2X1 U4746 ( .A(n3337), .B(n3391), .Y(n3398) );
  INVX1 U4747 ( .A(n3398), .Y(n6393) );
  AND2X1 U4748 ( .A(n3347), .B(n3426), .Y(n3438) );
  INVX1 U4749 ( .A(n3438), .Y(n6394) );
  AND2X1 U4750 ( .A(n3325), .B(n3461), .Y(n3462) );
  INVX1 U4751 ( .A(n3462), .Y(n6395) );
  AND2X1 U4752 ( .A(n3341), .B(n3461), .Y(n3470) );
  INVX1 U4753 ( .A(n3470), .Y(n6396) );
  AND2X1 U4754 ( .A(n3361), .B(n3496), .Y(n3515) );
  INVX1 U4755 ( .A(n3515), .Y(n6397) );
  AND2X1 U4756 ( .A(n3385), .B(n3496), .Y(n3527) );
  INVX1 U4757 ( .A(n3527), .Y(n6398) );
  AND2X1 U4758 ( .A(n3359), .B(n3530), .Y(n3548) );
  INVX1 U4759 ( .A(n3548), .Y(n6399) );
  AND2X1 U4760 ( .A(n3383), .B(n3530), .Y(n3560) );
  INVX1 U4761 ( .A(n3560), .Y(n6400) );
  AND2X1 U4762 ( .A(n3343), .B(n3565), .Y(n3575) );
  INVX1 U4763 ( .A(n3575), .Y(n6401) );
  AND2X1 U4764 ( .A(n3365), .B(n3565), .Y(n3586) );
  INVX1 U4765 ( .A(n3586), .Y(n6402) );
  AND2X1 U4766 ( .A(n3389), .B(n3565), .Y(n3598) );
  INVX1 U4767 ( .A(n3598), .Y(n6403) );
  AND2X1 U4768 ( .A(n3363), .B(n3600), .Y(n3620) );
  INVX1 U4769 ( .A(n3620), .Y(n6404) );
  AND2X1 U4770 ( .A(n3387), .B(n3600), .Y(n3632) );
  INVX1 U4771 ( .A(n3632), .Y(n6405) );
  AND2X1 U4772 ( .A(n3353), .B(n3635), .Y(n3650) );
  INVX1 U4773 ( .A(n3650), .Y(n6406) );
  AND2X1 U4774 ( .A(n3377), .B(n3635), .Y(n3662) );
  INVX1 U4775 ( .A(n3662), .Y(n6407) );
  AND2X1 U4776 ( .A(n3349), .B(n3670), .Y(n3683) );
  INVX1 U4777 ( .A(n3683), .Y(n6408) );
  AND2X1 U4778 ( .A(n3375), .B(n3670), .Y(n3696) );
  INVX1 U4779 ( .A(n3696), .Y(n6409) );
  AND2X1 U4780 ( .A(n3357), .B(n3704), .Y(n3721) );
  INVX1 U4781 ( .A(n3721), .Y(n6410) );
  AND2X1 U4782 ( .A(n3381), .B(n3704), .Y(n3733) );
  INVX1 U4783 ( .A(n3733), .Y(n6411) );
  AND2X1 U4784 ( .A(n3355), .B(n3738), .Y(n3754) );
  INVX1 U4785 ( .A(n3754), .Y(n6412) );
  AND2X1 U4786 ( .A(n3379), .B(n3738), .Y(n3766) );
  INVX1 U4787 ( .A(n3766), .Y(n6413) );
  AND2X1 U4788 ( .A(n3339), .B(n3772), .Y(n3780) );
  INVX1 U4789 ( .A(n3780), .Y(n6414) );
  AND2X1 U4790 ( .A(n3337), .B(n3806), .Y(n3813) );
  INVX1 U4791 ( .A(n3813), .Y(n6415) );
  AND2X1 U4792 ( .A(n3347), .B(n3840), .Y(n3852) );
  INVX1 U4793 ( .A(n3852), .Y(n6416) );
  AND2X1 U4794 ( .A(n3325), .B(n3874), .Y(n3875) );
  INVX1 U4795 ( .A(n3875), .Y(n6417) );
  AND2X1 U4796 ( .A(n3341), .B(n3874), .Y(n3883) );
  INVX1 U4797 ( .A(n3883), .Y(n6418) );
  AND2X1 U4798 ( .A(n3361), .B(n3908), .Y(n3927) );
  INVX1 U4799 ( .A(n3927), .Y(n6419) );
  AND2X1 U4800 ( .A(n3385), .B(n3908), .Y(n3939) );
  INVX1 U4801 ( .A(n3939), .Y(n6420) );
  AND2X1 U4802 ( .A(n3359), .B(n3943), .Y(n3961) );
  INVX1 U4803 ( .A(n3961), .Y(n6421) );
  AND2X1 U4804 ( .A(n3383), .B(n3943), .Y(n3973) );
  INVX1 U4805 ( .A(n3973), .Y(n6422) );
  AND2X1 U4806 ( .A(n3343), .B(n3977), .Y(n3987) );
  INVX1 U4807 ( .A(n3987), .Y(n6423) );
  AND2X1 U4808 ( .A(n3365), .B(n3977), .Y(n3998) );
  INVX1 U4809 ( .A(n3998), .Y(n6424) );
  AND2X1 U4810 ( .A(n3389), .B(n3977), .Y(n4010) );
  INVX1 U4811 ( .A(n4010), .Y(n6425) );
  AND2X1 U4812 ( .A(n3363), .B(n4011), .Y(n4031) );
  INVX1 U4813 ( .A(n4031), .Y(n6426) );
  AND2X1 U4814 ( .A(n3387), .B(n4011), .Y(n4043) );
  INVX1 U4815 ( .A(n4043), .Y(n6427) );
  AND2X1 U4816 ( .A(n3353), .B(n4045), .Y(n4060) );
  INVX1 U4817 ( .A(n4060), .Y(n6428) );
  AND2X1 U4818 ( .A(n3377), .B(n4045), .Y(n4072) );
  INVX1 U4819 ( .A(n4072), .Y(n6429) );
  AND2X1 U4820 ( .A(n3349), .B(n4079), .Y(n4092) );
  INVX1 U4821 ( .A(n4092), .Y(n6430) );
  AND2X1 U4822 ( .A(n3375), .B(n4079), .Y(n4105) );
  INVX1 U4823 ( .A(n4105), .Y(n6431) );
  AND2X1 U4824 ( .A(n3357), .B(n4113), .Y(n4130) );
  INVX1 U4825 ( .A(n4130), .Y(n6432) );
  AND2X1 U4826 ( .A(n3381), .B(n4113), .Y(n4142) );
  INVX1 U4827 ( .A(n4142), .Y(n6433) );
  AND2X1 U4828 ( .A(n3355), .B(n4147), .Y(n4163) );
  INVX1 U4829 ( .A(n4163), .Y(n6434) );
  AND2X1 U4830 ( .A(n3379), .B(n4147), .Y(n4175) );
  INVX1 U4831 ( .A(n4175), .Y(n6435) );
  AND2X1 U4832 ( .A(n3361), .B(n4181), .Y(n4200) );
  INVX1 U4833 ( .A(n4200), .Y(n6436) );
  AND2X1 U4834 ( .A(n3385), .B(n4181), .Y(n4212) );
  INVX1 U4835 ( .A(n4212), .Y(n6437) );
  AND2X1 U4836 ( .A(n3359), .B(n4216), .Y(n4234) );
  INVX1 U4837 ( .A(n4234), .Y(n6438) );
  AND2X1 U4838 ( .A(n3383), .B(n4216), .Y(n4246) );
  INVX1 U4839 ( .A(n4246), .Y(n6439) );
  AND2X1 U4840 ( .A(n3343), .B(n4250), .Y(n4260) );
  INVX1 U4841 ( .A(n4260), .Y(n6440) );
  AND2X1 U4842 ( .A(n3365), .B(n4250), .Y(n4271) );
  INVX1 U4843 ( .A(n4271), .Y(n6441) );
  AND2X1 U4844 ( .A(n3389), .B(n4250), .Y(n4283) );
  INVX1 U4845 ( .A(n4283), .Y(n6442) );
  AND2X1 U4846 ( .A(n3363), .B(n4284), .Y(n4304) );
  INVX1 U4847 ( .A(n4304), .Y(n6443) );
  AND2X1 U4848 ( .A(n3387), .B(n4284), .Y(n4316) );
  INVX1 U4849 ( .A(n4316), .Y(n6444) );
  AND2X1 U4850 ( .A(n3353), .B(n4318), .Y(n4333) );
  INVX1 U4851 ( .A(n4333), .Y(n6445) );
  AND2X1 U4852 ( .A(n3377), .B(n4318), .Y(n4345) );
  INVX1 U4853 ( .A(n4345), .Y(n6446) );
  AND2X1 U4854 ( .A(n3349), .B(n4352), .Y(n4365) );
  INVX1 U4855 ( .A(n4365), .Y(n6447) );
  AND2X1 U4856 ( .A(n3375), .B(n4352), .Y(n4378) );
  INVX1 U4857 ( .A(n4378), .Y(n6448) );
  AND2X1 U4858 ( .A(n3357), .B(n4386), .Y(n4403) );
  INVX1 U4859 ( .A(n4403), .Y(n6449) );
  AND2X1 U4860 ( .A(n3381), .B(n4386), .Y(n4415) );
  INVX1 U4861 ( .A(n4415), .Y(n6450) );
  AND2X1 U4862 ( .A(n3355), .B(n4420), .Y(n4436) );
  INVX1 U4863 ( .A(n4436), .Y(n6451) );
  AND2X1 U4864 ( .A(n3379), .B(n4420), .Y(n4448) );
  INVX1 U4865 ( .A(n4448), .Y(n6452) );
  BUFX2 U4866 ( .A(n3321), .Y(n6453) );
  BUFX2 U4867 ( .A(n3460), .Y(n6454) );
  BUFX2 U4868 ( .A(n3564), .Y(n6455) );
  AND2X1 U4869 ( .A(n3276), .B(n6853), .Y(n3300) );
  INVX1 U4870 ( .A(n3300), .Y(n6456) );
  AND2X1 U4871 ( .A(n3337), .B(n3323), .Y(n3336) );
  INVX1 U4872 ( .A(n3336), .Y(n6457) );
  AND2X1 U4873 ( .A(n3339), .B(n3391), .Y(n3399) );
  INVX1 U4874 ( .A(n3399), .Y(n6458) );
  AND2X1 U4875 ( .A(n3325), .B(n3426), .Y(n3427) );
  INVX1 U4876 ( .A(n3427), .Y(n6459) );
  AND2X1 U4877 ( .A(n3341), .B(n3426), .Y(n3435) );
  INVX1 U4878 ( .A(n3435), .Y(n6460) );
  AND2X1 U4879 ( .A(n3347), .B(n3461), .Y(n3473) );
  INVX1 U4880 ( .A(n3473), .Y(n6461) );
  AND2X1 U4881 ( .A(n3359), .B(n3496), .Y(n3514) );
  INVX1 U4882 ( .A(n3514), .Y(n6462) );
  AND2X1 U4883 ( .A(n3383), .B(n3496), .Y(n3526) );
  INVX1 U4884 ( .A(n3526), .Y(n6463) );
  AND2X1 U4885 ( .A(n3361), .B(n3530), .Y(n3549) );
  INVX1 U4886 ( .A(n3549), .Y(n6464) );
  AND2X1 U4887 ( .A(n3385), .B(n3530), .Y(n3561) );
  INVX1 U4888 ( .A(n3561), .Y(n6465) );
  AND2X1 U4889 ( .A(n3363), .B(n3565), .Y(n3585) );
  INVX1 U4890 ( .A(n3585), .Y(n6466) );
  AND2X1 U4891 ( .A(n3387), .B(n3565), .Y(n3597) );
  INVX1 U4892 ( .A(n3597), .Y(n6467) );
  AND2X1 U4893 ( .A(n3343), .B(n3600), .Y(n3610) );
  INVX1 U4894 ( .A(n3610), .Y(n6468) );
  AND2X1 U4895 ( .A(n3365), .B(n3600), .Y(n3621) );
  INVX1 U4896 ( .A(n3621), .Y(n6469) );
  AND2X1 U4897 ( .A(n3389), .B(n3600), .Y(n3633) );
  INVX1 U4898 ( .A(n3633), .Y(n6470) );
  AND2X1 U4899 ( .A(n3349), .B(n3635), .Y(n3648) );
  INVX1 U4900 ( .A(n3648), .Y(n6471) );
  AND2X1 U4901 ( .A(n3375), .B(n3635), .Y(n3661) );
  INVX1 U4902 ( .A(n3661), .Y(n6472) );
  AND2X1 U4903 ( .A(n3353), .B(n3670), .Y(n3685) );
  INVX1 U4904 ( .A(n3685), .Y(n6473) );
  AND2X1 U4905 ( .A(n3377), .B(n3670), .Y(n3697) );
  INVX1 U4906 ( .A(n3697), .Y(n6474) );
  AND2X1 U4907 ( .A(n3355), .B(n3704), .Y(n3720) );
  INVX1 U4908 ( .A(n3720), .Y(n6475) );
  AND2X1 U4909 ( .A(n3379), .B(n3704), .Y(n3732) );
  INVX1 U4910 ( .A(n3732), .Y(n6476) );
  AND2X1 U4911 ( .A(n3357), .B(n3738), .Y(n3755) );
  INVX1 U4912 ( .A(n3755), .Y(n6477) );
  AND2X1 U4913 ( .A(n3381), .B(n3738), .Y(n3767) );
  INVX1 U4914 ( .A(n3767), .Y(n6478) );
  AND2X1 U4915 ( .A(n3337), .B(n3772), .Y(n3779) );
  INVX1 U4916 ( .A(n3779), .Y(n6479) );
  AND2X1 U4917 ( .A(n3339), .B(n3806), .Y(n3814) );
  INVX1 U4918 ( .A(n3814), .Y(n6480) );
  AND2X1 U4919 ( .A(n3325), .B(n3840), .Y(n3841) );
  INVX1 U4920 ( .A(n3841), .Y(n6481) );
  AND2X1 U4921 ( .A(n3341), .B(n3840), .Y(n3849) );
  INVX1 U4922 ( .A(n3849), .Y(n6482) );
  AND2X1 U4923 ( .A(n3347), .B(n3874), .Y(n3886) );
  INVX1 U4924 ( .A(n3886), .Y(n6483) );
  AND2X1 U4925 ( .A(n3359), .B(n3908), .Y(n3926) );
  INVX1 U4926 ( .A(n3926), .Y(n6484) );
  AND2X1 U4927 ( .A(n3383), .B(n3908), .Y(n3938) );
  INVX1 U4928 ( .A(n3938), .Y(n6485) );
  AND2X1 U4929 ( .A(n3361), .B(n3943), .Y(n3962) );
  INVX1 U4930 ( .A(n3962), .Y(n6486) );
  AND2X1 U4931 ( .A(n3385), .B(n3943), .Y(n3974) );
  INVX1 U4932 ( .A(n3974), .Y(n6487) );
  AND2X1 U4933 ( .A(n3363), .B(n3977), .Y(n3997) );
  INVX1 U4934 ( .A(n3997), .Y(n6488) );
  AND2X1 U4935 ( .A(n3387), .B(n3977), .Y(n4009) );
  INVX1 U4936 ( .A(n4009), .Y(n6489) );
  AND2X1 U4937 ( .A(n3343), .B(n4011), .Y(n4021) );
  INVX1 U4938 ( .A(n4021), .Y(n6490) );
  AND2X1 U4939 ( .A(n3365), .B(n4011), .Y(n4032) );
  INVX1 U4940 ( .A(n4032), .Y(n6491) );
  AND2X1 U4941 ( .A(n3389), .B(n4011), .Y(n4044) );
  INVX1 U4942 ( .A(n4044), .Y(n6492) );
  AND2X1 U4943 ( .A(n3349), .B(n4045), .Y(n4058) );
  INVX1 U4944 ( .A(n4058), .Y(n6493) );
  AND2X1 U4945 ( .A(n3375), .B(n4045), .Y(n4071) );
  INVX1 U4946 ( .A(n4071), .Y(n6494) );
  AND2X1 U4947 ( .A(n3353), .B(n4079), .Y(n4094) );
  INVX1 U4948 ( .A(n4094), .Y(n6495) );
  AND2X1 U4949 ( .A(n3377), .B(n4079), .Y(n4106) );
  INVX1 U4950 ( .A(n4106), .Y(n6496) );
  AND2X1 U4951 ( .A(n3355), .B(n4113), .Y(n4129) );
  INVX1 U4952 ( .A(n4129), .Y(n6497) );
  AND2X1 U4953 ( .A(n3379), .B(n4113), .Y(n4141) );
  INVX1 U4954 ( .A(n4141), .Y(n6498) );
  AND2X1 U4955 ( .A(n3357), .B(n4147), .Y(n4164) );
  INVX1 U4956 ( .A(n4164), .Y(n6499) );
  AND2X1 U4957 ( .A(n3381), .B(n4147), .Y(n4176) );
  INVX1 U4958 ( .A(n4176), .Y(n6500) );
  AND2X1 U4959 ( .A(n3359), .B(n4181), .Y(n4199) );
  INVX1 U4960 ( .A(n4199), .Y(n6501) );
  AND2X1 U4961 ( .A(n3383), .B(n4181), .Y(n4211) );
  INVX1 U4962 ( .A(n4211), .Y(n6502) );
  AND2X1 U4963 ( .A(n3361), .B(n4216), .Y(n4235) );
  INVX1 U4964 ( .A(n4235), .Y(n6503) );
  AND2X1 U4965 ( .A(n3385), .B(n4216), .Y(n4247) );
  INVX1 U4966 ( .A(n4247), .Y(n6504) );
  AND2X1 U4967 ( .A(n3363), .B(n4250), .Y(n4270) );
  INVX1 U4968 ( .A(n4270), .Y(n6505) );
  AND2X1 U4969 ( .A(n3387), .B(n4250), .Y(n4282) );
  INVX1 U4970 ( .A(n4282), .Y(n6506) );
  AND2X1 U4971 ( .A(n3343), .B(n4284), .Y(n4294) );
  INVX1 U4972 ( .A(n4294), .Y(n6507) );
  AND2X1 U4973 ( .A(n3365), .B(n4284), .Y(n4305) );
  INVX1 U4974 ( .A(n4305), .Y(n6508) );
  AND2X1 U4975 ( .A(n3389), .B(n4284), .Y(n4317) );
  INVX1 U4976 ( .A(n4317), .Y(n6509) );
  AND2X1 U4977 ( .A(n3349), .B(n4318), .Y(n4331) );
  INVX1 U4978 ( .A(n4331), .Y(n6510) );
  AND2X1 U4979 ( .A(n3375), .B(n4318), .Y(n4344) );
  INVX1 U4980 ( .A(n4344), .Y(n6511) );
  AND2X1 U4981 ( .A(n3353), .B(n4352), .Y(n4367) );
  INVX1 U4982 ( .A(n4367), .Y(n6512) );
  AND2X1 U4983 ( .A(n3377), .B(n4352), .Y(n4379) );
  INVX1 U4984 ( .A(n4379), .Y(n6513) );
  AND2X1 U4985 ( .A(n3355), .B(n4386), .Y(n4402) );
  INVX1 U4986 ( .A(n4402), .Y(n6514) );
  AND2X1 U4987 ( .A(n3379), .B(n4386), .Y(n4414) );
  INVX1 U4988 ( .A(n4414), .Y(n6515) );
  AND2X1 U4989 ( .A(n3357), .B(n4420), .Y(n4437) );
  INVX1 U4990 ( .A(n4437), .Y(n6516) );
  AND2X1 U4991 ( .A(n3381), .B(n4420), .Y(n4449) );
  INVX1 U4992 ( .A(n4449), .Y(n6517) );
  BUFX2 U4993 ( .A(n3313), .Y(n6518) );
  BUFX2 U4994 ( .A(n3312), .Y(n6519) );
  OR2X1 U4995 ( .A(n6860), .B(wr_ptr[4]), .Y(n3314) );
  INVX1 U4996 ( .A(n3314), .Y(n6520) );
  BUFX2 U4997 ( .A(n3425), .Y(n6521) );
  BUFX2 U4998 ( .A(n3599), .Y(n6522) );
  AND2X1 U4999 ( .A(n3345), .B(n3323), .Y(n3344) );
  INVX1 U5000 ( .A(n3344), .Y(n6523) );
  AND2X1 U5001 ( .A(n3373), .B(n3323), .Y(n3372) );
  INVX1 U5002 ( .A(n3372), .Y(n6524) );
  AND2X1 U5003 ( .A(n3351), .B(n3391), .Y(n3405) );
  INVX1 U5004 ( .A(n3405), .Y(n6525) );
  AND2X1 U5005 ( .A(n3371), .B(n3391), .Y(n3415) );
  INVX1 U5006 ( .A(n3415), .Y(n6526) );
  AND2X1 U5007 ( .A(n3329), .B(n3426), .Y(n3429) );
  INVX1 U5008 ( .A(n3429), .Y(n6527) );
  AND2X1 U5009 ( .A(n3369), .B(n3426), .Y(n3449) );
  INVX1 U5010 ( .A(n3449), .Y(n6528) );
  AND2X1 U5011 ( .A(n3327), .B(n3461), .Y(n3463) );
  INVX1 U5012 ( .A(n3463), .Y(n6529) );
  AND2X1 U5013 ( .A(n3367), .B(n3461), .Y(n3483) );
  INVX1 U5014 ( .A(n3483), .Y(n6530) );
  AND2X1 U5015 ( .A(n3357), .B(n3496), .Y(n3513) );
  INVX1 U5016 ( .A(n3513), .Y(n6531) );
  AND2X1 U5017 ( .A(n3381), .B(n3496), .Y(n3525) );
  INVX1 U5018 ( .A(n3525), .Y(n6532) );
  AND2X1 U5019 ( .A(n3355), .B(n3530), .Y(n3546) );
  INVX1 U5020 ( .A(n3546), .Y(n6533) );
  AND2X1 U5021 ( .A(n3379), .B(n3530), .Y(n3558) );
  INVX1 U5022 ( .A(n3558), .Y(n6534) );
  AND2X1 U5023 ( .A(n3353), .B(n3565), .Y(n3580) );
  INVX1 U5024 ( .A(n3580), .Y(n6535) );
  AND2X1 U5025 ( .A(n3377), .B(n3565), .Y(n3592) );
  INVX1 U5026 ( .A(n3592), .Y(n6536) );
  AND2X1 U5027 ( .A(n3349), .B(n3600), .Y(n3613) );
  INVX1 U5028 ( .A(n3613), .Y(n6537) );
  AND2X1 U5029 ( .A(n3375), .B(n3600), .Y(n3626) );
  INVX1 U5030 ( .A(n3626), .Y(n6538) );
  AND2X1 U5031 ( .A(n3343), .B(n3635), .Y(n3645) );
  INVX1 U5032 ( .A(n3645), .Y(n6539) );
  AND2X1 U5033 ( .A(n3365), .B(n3635), .Y(n3656) );
  INVX1 U5034 ( .A(n3656), .Y(n6540) );
  AND2X1 U5035 ( .A(n3389), .B(n3635), .Y(n3668) );
  INVX1 U5036 ( .A(n3668), .Y(n6541) );
  AND2X1 U5037 ( .A(n3363), .B(n3670), .Y(n3690) );
  INVX1 U5038 ( .A(n3690), .Y(n6542) );
  AND2X1 U5039 ( .A(n3387), .B(n3670), .Y(n3702) );
  INVX1 U5040 ( .A(n3702), .Y(n6543) );
  AND2X1 U5041 ( .A(n3361), .B(n3704), .Y(n3723) );
  INVX1 U5042 ( .A(n3723), .Y(n6544) );
  AND2X1 U5043 ( .A(n3385), .B(n3704), .Y(n3735) );
  INVX1 U5044 ( .A(n3735), .Y(n6545) );
  AND2X1 U5045 ( .A(n3359), .B(n3738), .Y(n3756) );
  INVX1 U5046 ( .A(n3756), .Y(n6546) );
  AND2X1 U5047 ( .A(n3383), .B(n3738), .Y(n3768) );
  INVX1 U5048 ( .A(n3768), .Y(n6547) );
  AND2X1 U5049 ( .A(n3345), .B(n3772), .Y(n3783) );
  INVX1 U5050 ( .A(n3783), .Y(n6548) );
  AND2X1 U5051 ( .A(n3373), .B(n3772), .Y(n3797) );
  INVX1 U5052 ( .A(n3797), .Y(n6549) );
  AND2X1 U5053 ( .A(n3351), .B(n3806), .Y(n3820) );
  INVX1 U5054 ( .A(n3820), .Y(n6550) );
  AND2X1 U5055 ( .A(n3371), .B(n3806), .Y(n3830) );
  INVX1 U5056 ( .A(n3830), .Y(n6551) );
  AND2X1 U5057 ( .A(n3329), .B(n3840), .Y(n3843) );
  INVX1 U5058 ( .A(n3843), .Y(n6552) );
  AND2X1 U5059 ( .A(n3369), .B(n3840), .Y(n3863) );
  INVX1 U5060 ( .A(n3863), .Y(n6553) );
  AND2X1 U5061 ( .A(n3327), .B(n3874), .Y(n3876) );
  INVX1 U5062 ( .A(n3876), .Y(n6554) );
  AND2X1 U5063 ( .A(n3367), .B(n3874), .Y(n3896) );
  INVX1 U5064 ( .A(n3896), .Y(n6555) );
  AND2X1 U5065 ( .A(n3357), .B(n3908), .Y(n3925) );
  INVX1 U5066 ( .A(n3925), .Y(n6556) );
  AND2X1 U5067 ( .A(n3381), .B(n3908), .Y(n3937) );
  INVX1 U5068 ( .A(n3937), .Y(n6557) );
  AND2X1 U5069 ( .A(n3355), .B(n3943), .Y(n3959) );
  INVX1 U5070 ( .A(n3959), .Y(n6558) );
  AND2X1 U5071 ( .A(n3379), .B(n3943), .Y(n3971) );
  INVX1 U5072 ( .A(n3971), .Y(n6559) );
  AND2X1 U5073 ( .A(n3353), .B(n3977), .Y(n3992) );
  INVX1 U5074 ( .A(n3992), .Y(n6560) );
  AND2X1 U5075 ( .A(n3377), .B(n3977), .Y(n4004) );
  INVX1 U5076 ( .A(n4004), .Y(n6561) );
  AND2X1 U5077 ( .A(n3349), .B(n4011), .Y(n4024) );
  INVX1 U5078 ( .A(n4024), .Y(n6562) );
  AND2X1 U5079 ( .A(n3375), .B(n4011), .Y(n4037) );
  INVX1 U5080 ( .A(n4037), .Y(n6563) );
  AND2X1 U5081 ( .A(n3343), .B(n4045), .Y(n4055) );
  INVX1 U5082 ( .A(n4055), .Y(n6564) );
  AND2X1 U5083 ( .A(n3365), .B(n4045), .Y(n4066) );
  INVX1 U5084 ( .A(n4066), .Y(n6565) );
  AND2X1 U5085 ( .A(n3389), .B(n4045), .Y(n4078) );
  INVX1 U5086 ( .A(n4078), .Y(n6566) );
  AND2X1 U5087 ( .A(n3363), .B(n4079), .Y(n4099) );
  INVX1 U5088 ( .A(n4099), .Y(n6567) );
  AND2X1 U5089 ( .A(n3387), .B(n4079), .Y(n4111) );
  INVX1 U5090 ( .A(n4111), .Y(n6568) );
  AND2X1 U5091 ( .A(n3361), .B(n4113), .Y(n4132) );
  INVX1 U5092 ( .A(n4132), .Y(n6569) );
  AND2X1 U5093 ( .A(n3385), .B(n4113), .Y(n4144) );
  INVX1 U5094 ( .A(n4144), .Y(n6570) );
  AND2X1 U5095 ( .A(n3359), .B(n4147), .Y(n4165) );
  INVX1 U5096 ( .A(n4165), .Y(n6571) );
  AND2X1 U5097 ( .A(n3383), .B(n4147), .Y(n4177) );
  INVX1 U5098 ( .A(n4177), .Y(n6572) );
  AND2X1 U5099 ( .A(n3357), .B(n4181), .Y(n4198) );
  INVX1 U5100 ( .A(n4198), .Y(n6573) );
  AND2X1 U5101 ( .A(n3381), .B(n4181), .Y(n4210) );
  INVX1 U5102 ( .A(n4210), .Y(n6574) );
  AND2X1 U5103 ( .A(n3355), .B(n4216), .Y(n4232) );
  INVX1 U5104 ( .A(n4232), .Y(n6575) );
  AND2X1 U5105 ( .A(n3379), .B(n4216), .Y(n4244) );
  INVX1 U5106 ( .A(n4244), .Y(n6576) );
  AND2X1 U5107 ( .A(n3353), .B(n4250), .Y(n4265) );
  INVX1 U5108 ( .A(n4265), .Y(n6577) );
  AND2X1 U5109 ( .A(n3377), .B(n4250), .Y(n4277) );
  INVX1 U5110 ( .A(n4277), .Y(n6578) );
  AND2X1 U5111 ( .A(n3349), .B(n4284), .Y(n4297) );
  INVX1 U5112 ( .A(n4297), .Y(n6579) );
  AND2X1 U5113 ( .A(n3375), .B(n4284), .Y(n4310) );
  INVX1 U5114 ( .A(n4310), .Y(n6580) );
  AND2X1 U5115 ( .A(n3343), .B(n4318), .Y(n4328) );
  INVX1 U5116 ( .A(n4328), .Y(n6581) );
  AND2X1 U5117 ( .A(n3365), .B(n4318), .Y(n4339) );
  INVX1 U5118 ( .A(n4339), .Y(n6582) );
  AND2X1 U5119 ( .A(n3389), .B(n4318), .Y(n4351) );
  INVX1 U5120 ( .A(n4351), .Y(n6583) );
  AND2X1 U5121 ( .A(n3363), .B(n4352), .Y(n4372) );
  INVX1 U5122 ( .A(n4372), .Y(n6584) );
  AND2X1 U5123 ( .A(n3387), .B(n4352), .Y(n4384) );
  INVX1 U5124 ( .A(n4384), .Y(n6585) );
  AND2X1 U5125 ( .A(n3361), .B(n4386), .Y(n4405) );
  INVX1 U5126 ( .A(n4405), .Y(n6586) );
  AND2X1 U5127 ( .A(n3385), .B(n4386), .Y(n4417) );
  INVX1 U5128 ( .A(n4417), .Y(n6587) );
  AND2X1 U5129 ( .A(n3359), .B(n4420), .Y(n4438) );
  INVX1 U5130 ( .A(n4438), .Y(n6588) );
  AND2X1 U5131 ( .A(n3383), .B(n4420), .Y(n4450) );
  INVX1 U5132 ( .A(n4450), .Y(n6589) );
  INVX1 U5133 ( .A(n3299), .Y(n6590) );
  INVX1 U5134 ( .A(n3306), .Y(n6591) );
  BUFX2 U5135 ( .A(n4624), .Y(empty_bar) );
  BUFX2 U5136 ( .A(n3634), .Y(n6593) );
  BUFX2 U5137 ( .A(n3322), .Y(n6594) );
  AND2X1 U5138 ( .A(n3351), .B(n3323), .Y(n3350) );
  INVX1 U5139 ( .A(n3350), .Y(n6595) );
  AND2X1 U5140 ( .A(n3371), .B(n3323), .Y(n3370) );
  INVX1 U5141 ( .A(n3370), .Y(n6596) );
  AND2X1 U5142 ( .A(n3345), .B(n3391), .Y(n3402) );
  INVX1 U5143 ( .A(n3402), .Y(n6597) );
  AND2X1 U5144 ( .A(n3373), .B(n3391), .Y(n3416) );
  INVX1 U5145 ( .A(n3416), .Y(n6598) );
  AND2X1 U5146 ( .A(n3327), .B(n3426), .Y(n3428) );
  INVX1 U5147 ( .A(n3428), .Y(n6599) );
  AND2X1 U5148 ( .A(n3367), .B(n3426), .Y(n3448) );
  INVX1 U5149 ( .A(n3448), .Y(n6600) );
  AND2X1 U5150 ( .A(n3329), .B(n3461), .Y(n3464) );
  INVX1 U5151 ( .A(n3464), .Y(n6601) );
  AND2X1 U5152 ( .A(n3369), .B(n3461), .Y(n3484) );
  INVX1 U5153 ( .A(n3484), .Y(n6602) );
  AND2X1 U5154 ( .A(n3355), .B(n3496), .Y(n3512) );
  INVX1 U5155 ( .A(n3512), .Y(n6603) );
  AND2X1 U5156 ( .A(n3379), .B(n3496), .Y(n3524) );
  INVX1 U5157 ( .A(n3524), .Y(n6604) );
  AND2X1 U5158 ( .A(n3357), .B(n3530), .Y(n3547) );
  INVX1 U5159 ( .A(n3547), .Y(n6605) );
  AND2X1 U5160 ( .A(n3381), .B(n3530), .Y(n3559) );
  INVX1 U5161 ( .A(n3559), .Y(n6606) );
  AND2X1 U5162 ( .A(n3349), .B(n3565), .Y(n3578) );
  INVX1 U5163 ( .A(n3578), .Y(n6607) );
  AND2X1 U5164 ( .A(n3375), .B(n3565), .Y(n3591) );
  INVX1 U5165 ( .A(n3591), .Y(n6608) );
  AND2X1 U5166 ( .A(n3353), .B(n3600), .Y(n3615) );
  INVX1 U5167 ( .A(n3615), .Y(n6609) );
  AND2X1 U5168 ( .A(n3377), .B(n3600), .Y(n3627) );
  INVX1 U5169 ( .A(n3627), .Y(n6610) );
  AND2X1 U5170 ( .A(n3363), .B(n3635), .Y(n3655) );
  INVX1 U5171 ( .A(n3655), .Y(n6611) );
  AND2X1 U5172 ( .A(n3387), .B(n3635), .Y(n3667) );
  INVX1 U5173 ( .A(n3667), .Y(n6612) );
  AND2X1 U5174 ( .A(n3343), .B(n3670), .Y(n3680) );
  INVX1 U5175 ( .A(n3680), .Y(n6613) );
  AND2X1 U5176 ( .A(n3365), .B(n3670), .Y(n3691) );
  INVX1 U5177 ( .A(n3691), .Y(n6614) );
  AND2X1 U5178 ( .A(n3389), .B(n3670), .Y(n3703) );
  INVX1 U5179 ( .A(n3703), .Y(n6615) );
  AND2X1 U5180 ( .A(n3359), .B(n3704), .Y(n3722) );
  INVX1 U5181 ( .A(n3722), .Y(n6616) );
  AND2X1 U5182 ( .A(n3383), .B(n3704), .Y(n3734) );
  INVX1 U5183 ( .A(n3734), .Y(n6617) );
  AND2X1 U5184 ( .A(n3361), .B(n3738), .Y(n3757) );
  INVX1 U5185 ( .A(n3757), .Y(n6618) );
  AND2X1 U5186 ( .A(n3385), .B(n3738), .Y(n3769) );
  INVX1 U5187 ( .A(n3769), .Y(n6619) );
  AND2X1 U5188 ( .A(n3351), .B(n3772), .Y(n3786) );
  INVX1 U5189 ( .A(n3786), .Y(n6620) );
  AND2X1 U5190 ( .A(n3371), .B(n3772), .Y(n3796) );
  INVX1 U5191 ( .A(n3796), .Y(n6621) );
  AND2X1 U5192 ( .A(n3345), .B(n3806), .Y(n3817) );
  INVX1 U5193 ( .A(n3817), .Y(n6622) );
  AND2X1 U5194 ( .A(n3373), .B(n3806), .Y(n3831) );
  INVX1 U5195 ( .A(n3831), .Y(n6623) );
  AND2X1 U5196 ( .A(n3327), .B(n3840), .Y(n3842) );
  INVX1 U5197 ( .A(n3842), .Y(n6624) );
  AND2X1 U5198 ( .A(n3367), .B(n3840), .Y(n3862) );
  INVX1 U5199 ( .A(n3862), .Y(n6625) );
  AND2X1 U5200 ( .A(n3329), .B(n3874), .Y(n3877) );
  INVX1 U5201 ( .A(n3877), .Y(n6626) );
  AND2X1 U5202 ( .A(n3369), .B(n3874), .Y(n3897) );
  INVX1 U5203 ( .A(n3897), .Y(n6627) );
  AND2X1 U5204 ( .A(n3355), .B(n3908), .Y(n3924) );
  INVX1 U5205 ( .A(n3924), .Y(n6628) );
  AND2X1 U5206 ( .A(n3379), .B(n3908), .Y(n3936) );
  INVX1 U5207 ( .A(n3936), .Y(n6629) );
  AND2X1 U5208 ( .A(n3357), .B(n3943), .Y(n3960) );
  INVX1 U5209 ( .A(n3960), .Y(n6630) );
  AND2X1 U5210 ( .A(n3381), .B(n3943), .Y(n3972) );
  INVX1 U5211 ( .A(n3972), .Y(n6631) );
  AND2X1 U5212 ( .A(n3349), .B(n3977), .Y(n3990) );
  INVX1 U5213 ( .A(n3990), .Y(n6632) );
  AND2X1 U5214 ( .A(n3375), .B(n3977), .Y(n4003) );
  INVX1 U5215 ( .A(n4003), .Y(n6633) );
  AND2X1 U5216 ( .A(n3353), .B(n4011), .Y(n4026) );
  INVX1 U5217 ( .A(n4026), .Y(n6634) );
  AND2X1 U5218 ( .A(n3377), .B(n4011), .Y(n4038) );
  INVX1 U5219 ( .A(n4038), .Y(n6635) );
  AND2X1 U5220 ( .A(n3363), .B(n4045), .Y(n4065) );
  INVX1 U5221 ( .A(n4065), .Y(n6636) );
  AND2X1 U5222 ( .A(n3387), .B(n4045), .Y(n4077) );
  INVX1 U5223 ( .A(n4077), .Y(n6637) );
  AND2X1 U5224 ( .A(n3343), .B(n4079), .Y(n4089) );
  INVX1 U5225 ( .A(n4089), .Y(n6638) );
  AND2X1 U5226 ( .A(n3365), .B(n4079), .Y(n4100) );
  INVX1 U5227 ( .A(n4100), .Y(n6639) );
  AND2X1 U5228 ( .A(n3389), .B(n4079), .Y(n4112) );
  INVX1 U5229 ( .A(n4112), .Y(n6640) );
  AND2X1 U5230 ( .A(n3359), .B(n4113), .Y(n4131) );
  INVX1 U5231 ( .A(n4131), .Y(n6641) );
  AND2X1 U5232 ( .A(n3383), .B(n4113), .Y(n4143) );
  INVX1 U5233 ( .A(n4143), .Y(n6642) );
  AND2X1 U5234 ( .A(n3361), .B(n4147), .Y(n4166) );
  INVX1 U5235 ( .A(n4166), .Y(n6643) );
  AND2X1 U5236 ( .A(n3385), .B(n4147), .Y(n4178) );
  INVX1 U5237 ( .A(n4178), .Y(n6644) );
  AND2X1 U5238 ( .A(n3355), .B(n4181), .Y(n4197) );
  INVX1 U5239 ( .A(n4197), .Y(n6645) );
  AND2X1 U5240 ( .A(n3379), .B(n4181), .Y(n4209) );
  INVX1 U5241 ( .A(n4209), .Y(n6646) );
  AND2X1 U5242 ( .A(n3357), .B(n4216), .Y(n4233) );
  INVX1 U5243 ( .A(n4233), .Y(n6647) );
  AND2X1 U5244 ( .A(n3381), .B(n4216), .Y(n4245) );
  INVX1 U5245 ( .A(n4245), .Y(n6648) );
  AND2X1 U5246 ( .A(n3349), .B(n4250), .Y(n4263) );
  INVX1 U5247 ( .A(n4263), .Y(n6649) );
  AND2X1 U5248 ( .A(n3375), .B(n4250), .Y(n4276) );
  INVX1 U5249 ( .A(n4276), .Y(n6650) );
  AND2X1 U5250 ( .A(n3353), .B(n4284), .Y(n4299) );
  INVX1 U5251 ( .A(n4299), .Y(n6651) );
  AND2X1 U5252 ( .A(n3377), .B(n4284), .Y(n4311) );
  INVX1 U5253 ( .A(n4311), .Y(n6652) );
  AND2X1 U5254 ( .A(n3363), .B(n4318), .Y(n4338) );
  INVX1 U5255 ( .A(n4338), .Y(n6653) );
  AND2X1 U5256 ( .A(n3387), .B(n4318), .Y(n4350) );
  INVX1 U5257 ( .A(n4350), .Y(n6654) );
  AND2X1 U5258 ( .A(n3343), .B(n4352), .Y(n4362) );
  INVX1 U5259 ( .A(n4362), .Y(n6655) );
  AND2X1 U5260 ( .A(n3365), .B(n4352), .Y(n4373) );
  INVX1 U5261 ( .A(n4373), .Y(n6656) );
  AND2X1 U5262 ( .A(n3389), .B(n4352), .Y(n4385) );
  INVX1 U5263 ( .A(n4385), .Y(n6657) );
  AND2X1 U5264 ( .A(n3359), .B(n4386), .Y(n4404) );
  INVX1 U5265 ( .A(n4404), .Y(n6658) );
  AND2X1 U5266 ( .A(n3383), .B(n4386), .Y(n4416) );
  INVX1 U5267 ( .A(n4416), .Y(n6659) );
  AND2X1 U5268 ( .A(n3361), .B(n4420), .Y(n4439) );
  INVX1 U5269 ( .A(n4439), .Y(n6660) );
  AND2X1 U5270 ( .A(n3385), .B(n4420), .Y(n4451) );
  INVX1 U5271 ( .A(n4451), .Y(n6661) );
  INVX1 U5272 ( .A(n3276), .Y(n6662) );
  BUFX2 U5273 ( .A(n3291), .Y(n6663) );
  BUFX2 U5274 ( .A(n4455), .Y(n6664) );
  BUFX2 U5275 ( .A(n3495), .Y(n6665) );
  BUFX2 U5276 ( .A(n3320), .Y(n6666) );
  AND2X1 U5277 ( .A(n3329), .B(n3323), .Y(n3328) );
  INVX1 U5278 ( .A(n3328), .Y(n6667) );
  AND2X1 U5279 ( .A(n3369), .B(n3323), .Y(n3368) );
  INVX1 U5280 ( .A(n3368), .Y(n6668) );
  AND2X1 U5281 ( .A(n3327), .B(n3391), .Y(n3393) );
  INVX1 U5282 ( .A(n3393), .Y(n6669) );
  AND2X1 U5283 ( .A(n3367), .B(n3391), .Y(n3413) );
  INVX1 U5284 ( .A(n3413), .Y(n6670) );
  AND2X1 U5285 ( .A(n3345), .B(n3426), .Y(n3437) );
  INVX1 U5286 ( .A(n3437), .Y(n6671) );
  AND2X1 U5287 ( .A(n3373), .B(n3426), .Y(n3451) );
  INVX1 U5288 ( .A(n3451), .Y(n6672) );
  AND2X1 U5289 ( .A(n3351), .B(n3461), .Y(n3475) );
  INVX1 U5290 ( .A(n3475), .Y(n6673) );
  AND2X1 U5291 ( .A(n3371), .B(n3461), .Y(n3485) );
  INVX1 U5292 ( .A(n3485), .Y(n6674) );
  AND2X1 U5293 ( .A(n3353), .B(n3496), .Y(n3511) );
  INVX1 U5294 ( .A(n3511), .Y(n6675) );
  AND2X1 U5295 ( .A(n3377), .B(n3496), .Y(n3523) );
  INVX1 U5296 ( .A(n3523), .Y(n6676) );
  AND2X1 U5297 ( .A(n3349), .B(n3530), .Y(n3543) );
  INVX1 U5298 ( .A(n3543), .Y(n6677) );
  AND2X1 U5299 ( .A(n3375), .B(n3530), .Y(n3556) );
  INVX1 U5300 ( .A(n3556), .Y(n6678) );
  AND2X1 U5301 ( .A(n3357), .B(n3565), .Y(n3582) );
  INVX1 U5302 ( .A(n3582), .Y(n6679) );
  AND2X1 U5303 ( .A(n3381), .B(n3565), .Y(n3594) );
  INVX1 U5304 ( .A(n3594), .Y(n6680) );
  AND2X1 U5305 ( .A(n3355), .B(n3600), .Y(n3616) );
  INVX1 U5306 ( .A(n3616), .Y(n6681) );
  AND2X1 U5307 ( .A(n3379), .B(n3600), .Y(n3628) );
  INVX1 U5308 ( .A(n3628), .Y(n6682) );
  AND2X1 U5309 ( .A(n3361), .B(n3635), .Y(n3654) );
  INVX1 U5310 ( .A(n3654), .Y(n6683) );
  AND2X1 U5311 ( .A(n3385), .B(n3635), .Y(n3666) );
  INVX1 U5312 ( .A(n3666), .Y(n6684) );
  AND2X1 U5313 ( .A(n3359), .B(n3670), .Y(n3688) );
  INVX1 U5314 ( .A(n3688), .Y(n6685) );
  AND2X1 U5315 ( .A(n3383), .B(n3670), .Y(n3700) );
  INVX1 U5316 ( .A(n3700), .Y(n6686) );
  AND2X1 U5317 ( .A(n3343), .B(n3704), .Y(n3714) );
  INVX1 U5318 ( .A(n3714), .Y(n6687) );
  AND2X1 U5319 ( .A(n3365), .B(n3704), .Y(n3725) );
  INVX1 U5320 ( .A(n3725), .Y(n6688) );
  AND2X1 U5321 ( .A(n3389), .B(n3704), .Y(n3737) );
  INVX1 U5322 ( .A(n3737), .Y(n6689) );
  AND2X1 U5323 ( .A(n3363), .B(n3738), .Y(n3758) );
  INVX1 U5324 ( .A(n3758), .Y(n6690) );
  AND2X1 U5325 ( .A(n3387), .B(n3738), .Y(n3770) );
  INVX1 U5326 ( .A(n3770), .Y(n6691) );
  AND2X1 U5327 ( .A(n3329), .B(n3772), .Y(n3775) );
  INVX1 U5328 ( .A(n3775), .Y(n6692) );
  AND2X1 U5329 ( .A(n3369), .B(n3772), .Y(n3795) );
  INVX1 U5330 ( .A(n3795), .Y(n6693) );
  AND2X1 U5331 ( .A(n3327), .B(n3806), .Y(n3808) );
  INVX1 U5332 ( .A(n3808), .Y(n6694) );
  AND2X1 U5333 ( .A(n3367), .B(n3806), .Y(n3828) );
  INVX1 U5334 ( .A(n3828), .Y(n6695) );
  AND2X1 U5335 ( .A(n3345), .B(n3840), .Y(n3851) );
  INVX1 U5336 ( .A(n3851), .Y(n6696) );
  AND2X1 U5337 ( .A(n3373), .B(n3840), .Y(n3865) );
  INVX1 U5338 ( .A(n3865), .Y(n6697) );
  AND2X1 U5339 ( .A(n3351), .B(n3874), .Y(n3888) );
  INVX1 U5340 ( .A(n3888), .Y(n6698) );
  AND2X1 U5341 ( .A(n3371), .B(n3874), .Y(n3898) );
  INVX1 U5342 ( .A(n3898), .Y(n6699) );
  AND2X1 U5343 ( .A(n3353), .B(n3908), .Y(n3923) );
  INVX1 U5344 ( .A(n3923), .Y(n6700) );
  AND2X1 U5345 ( .A(n3377), .B(n3908), .Y(n3935) );
  INVX1 U5346 ( .A(n3935), .Y(n6701) );
  AND2X1 U5347 ( .A(n3349), .B(n3943), .Y(n3956) );
  INVX1 U5348 ( .A(n3956), .Y(n6702) );
  AND2X1 U5349 ( .A(n3375), .B(n3943), .Y(n3969) );
  INVX1 U5350 ( .A(n3969), .Y(n6703) );
  AND2X1 U5351 ( .A(n3357), .B(n3977), .Y(n3994) );
  INVX1 U5352 ( .A(n3994), .Y(n6704) );
  AND2X1 U5353 ( .A(n3381), .B(n3977), .Y(n4006) );
  INVX1 U5354 ( .A(n4006), .Y(n6705) );
  AND2X1 U5355 ( .A(n3355), .B(n4011), .Y(n4027) );
  INVX1 U5356 ( .A(n4027), .Y(n6706) );
  AND2X1 U5357 ( .A(n3379), .B(n4011), .Y(n4039) );
  INVX1 U5358 ( .A(n4039), .Y(n6707) );
  AND2X1 U5359 ( .A(n3361), .B(n4045), .Y(n4064) );
  INVX1 U5360 ( .A(n4064), .Y(n6708) );
  AND2X1 U5361 ( .A(n3385), .B(n4045), .Y(n4076) );
  INVX1 U5362 ( .A(n4076), .Y(n6709) );
  AND2X1 U5363 ( .A(n3359), .B(n4079), .Y(n4097) );
  INVX1 U5364 ( .A(n4097), .Y(n6710) );
  AND2X1 U5365 ( .A(n3383), .B(n4079), .Y(n4109) );
  INVX1 U5366 ( .A(n4109), .Y(n6711) );
  AND2X1 U5367 ( .A(n3343), .B(n4113), .Y(n4123) );
  INVX1 U5368 ( .A(n4123), .Y(n6712) );
  AND2X1 U5369 ( .A(n3365), .B(n4113), .Y(n4134) );
  INVX1 U5370 ( .A(n4134), .Y(n6713) );
  AND2X1 U5371 ( .A(n3389), .B(n4113), .Y(n4146) );
  INVX1 U5372 ( .A(n4146), .Y(n6714) );
  AND2X1 U5373 ( .A(n3363), .B(n4147), .Y(n4167) );
  INVX1 U5374 ( .A(n4167), .Y(n6715) );
  AND2X1 U5375 ( .A(n3387), .B(n4147), .Y(n4179) );
  INVX1 U5376 ( .A(n4179), .Y(n6716) );
  AND2X1 U5377 ( .A(n3353), .B(n4181), .Y(n4196) );
  INVX1 U5378 ( .A(n4196), .Y(n6717) );
  AND2X1 U5379 ( .A(n3377), .B(n4181), .Y(n4208) );
  INVX1 U5380 ( .A(n4208), .Y(n6718) );
  AND2X1 U5381 ( .A(n3349), .B(n4216), .Y(n4229) );
  INVX1 U5382 ( .A(n4229), .Y(n6719) );
  AND2X1 U5383 ( .A(n3375), .B(n4216), .Y(n4242) );
  INVX1 U5384 ( .A(n4242), .Y(n6720) );
  AND2X1 U5385 ( .A(n3357), .B(n4250), .Y(n4267) );
  INVX1 U5386 ( .A(n4267), .Y(n6721) );
  AND2X1 U5387 ( .A(n3381), .B(n4250), .Y(n4279) );
  INVX1 U5388 ( .A(n4279), .Y(n6722) );
  AND2X1 U5389 ( .A(n3355), .B(n4284), .Y(n4300) );
  INVX1 U5390 ( .A(n4300), .Y(n6723) );
  AND2X1 U5391 ( .A(n3379), .B(n4284), .Y(n4312) );
  INVX1 U5392 ( .A(n4312), .Y(n6724) );
  AND2X1 U5393 ( .A(n3361), .B(n4318), .Y(n4337) );
  INVX1 U5394 ( .A(n4337), .Y(n6725) );
  AND2X1 U5395 ( .A(n3385), .B(n4318), .Y(n4349) );
  INVX1 U5396 ( .A(n4349), .Y(n6726) );
  AND2X1 U5397 ( .A(n3359), .B(n4352), .Y(n4370) );
  INVX1 U5398 ( .A(n4370), .Y(n6727) );
  AND2X1 U5399 ( .A(n3383), .B(n4352), .Y(n4382) );
  INVX1 U5400 ( .A(n4382), .Y(n6728) );
  AND2X1 U5401 ( .A(n3343), .B(n4386), .Y(n4396) );
  INVX1 U5402 ( .A(n4396), .Y(n6729) );
  AND2X1 U5403 ( .A(n3365), .B(n4386), .Y(n4407) );
  INVX1 U5404 ( .A(n4407), .Y(n6730) );
  AND2X1 U5405 ( .A(n3389), .B(n4386), .Y(n4419) );
  INVX1 U5406 ( .A(n4419), .Y(n6731) );
  AND2X1 U5407 ( .A(n3363), .B(n4420), .Y(n4440) );
  INVX1 U5408 ( .A(n4440), .Y(n6732) );
  AND2X1 U5409 ( .A(n3387), .B(n4420), .Y(n4452) );
  INVX1 U5410 ( .A(n4452), .Y(n6733) );
  BUFX2 U5411 ( .A(n3298), .Y(n6734) );
  AND2X1 U5412 ( .A(n6842), .B(n7917), .Y(n3295) );
  INVX1 U5413 ( .A(n3295), .Y(n6735) );
  BUFX2 U5414 ( .A(n3669), .Y(n6736) );
  BUFX2 U5415 ( .A(n3942), .Y(n6737) );
  AND2X1 U5416 ( .A(n3327), .B(n3323), .Y(n3326) );
  INVX1 U5417 ( .A(n3326), .Y(n6738) );
  AND2X1 U5418 ( .A(n3367), .B(n3323), .Y(n3366) );
  INVX1 U5419 ( .A(n3366), .Y(n6739) );
  AND2X1 U5420 ( .A(n3329), .B(n3391), .Y(n3394) );
  INVX1 U5421 ( .A(n3394), .Y(n6740) );
  AND2X1 U5422 ( .A(n3369), .B(n3391), .Y(n3414) );
  INVX1 U5423 ( .A(n3414), .Y(n6741) );
  AND2X1 U5424 ( .A(n3351), .B(n3426), .Y(n3440) );
  INVX1 U5425 ( .A(n3440), .Y(n6742) );
  AND2X1 U5426 ( .A(n3371), .B(n3426), .Y(n3450) );
  INVX1 U5427 ( .A(n3450), .Y(n6743) );
  AND2X1 U5428 ( .A(n3345), .B(n3461), .Y(n3472) );
  INVX1 U5429 ( .A(n3472), .Y(n6744) );
  AND2X1 U5430 ( .A(n3373), .B(n3461), .Y(n3486) );
  INVX1 U5431 ( .A(n3486), .Y(n6745) );
  AND2X1 U5432 ( .A(n3349), .B(n3496), .Y(n3509) );
  INVX1 U5433 ( .A(n3509), .Y(n6746) );
  AND2X1 U5434 ( .A(n3375), .B(n3496), .Y(n3522) );
  INVX1 U5435 ( .A(n3522), .Y(n6747) );
  AND2X1 U5436 ( .A(n3353), .B(n3530), .Y(n3545) );
  INVX1 U5437 ( .A(n3545), .Y(n6748) );
  AND2X1 U5438 ( .A(n3377), .B(n3530), .Y(n3557) );
  INVX1 U5439 ( .A(n3557), .Y(n6749) );
  AND2X1 U5440 ( .A(n3355), .B(n3565), .Y(n3581) );
  INVX1 U5441 ( .A(n3581), .Y(n6750) );
  AND2X1 U5442 ( .A(n3379), .B(n3565), .Y(n3593) );
  INVX1 U5443 ( .A(n3593), .Y(n6751) );
  AND2X1 U5444 ( .A(n3357), .B(n3600), .Y(n3617) );
  INVX1 U5445 ( .A(n3617), .Y(n6752) );
  AND2X1 U5446 ( .A(n3381), .B(n3600), .Y(n3629) );
  INVX1 U5447 ( .A(n3629), .Y(n6753) );
  AND2X1 U5448 ( .A(n3359), .B(n3635), .Y(n3653) );
  INVX1 U5449 ( .A(n3653), .Y(n6754) );
  AND2X1 U5450 ( .A(n3383), .B(n3635), .Y(n3665) );
  INVX1 U5451 ( .A(n3665), .Y(n6755) );
  AND2X1 U5452 ( .A(n3361), .B(n3670), .Y(n3689) );
  INVX1 U5453 ( .A(n3689), .Y(n6756) );
  AND2X1 U5454 ( .A(n3385), .B(n3670), .Y(n3701) );
  INVX1 U5455 ( .A(n3701), .Y(n6757) );
  AND2X1 U5456 ( .A(n3363), .B(n3704), .Y(n3724) );
  INVX1 U5457 ( .A(n3724), .Y(n6758) );
  AND2X1 U5458 ( .A(n3387), .B(n3704), .Y(n3736) );
  INVX1 U5459 ( .A(n3736), .Y(n6759) );
  AND2X1 U5460 ( .A(n3343), .B(n3738), .Y(n3748) );
  INVX1 U5461 ( .A(n3748), .Y(n6760) );
  AND2X1 U5462 ( .A(n3365), .B(n3738), .Y(n3759) );
  INVX1 U5463 ( .A(n3759), .Y(n6761) );
  AND2X1 U5464 ( .A(n3389), .B(n3738), .Y(n3771) );
  INVX1 U5465 ( .A(n3771), .Y(n6762) );
  AND2X1 U5466 ( .A(n3327), .B(n3772), .Y(n3774) );
  INVX1 U5467 ( .A(n3774), .Y(n6763) );
  AND2X1 U5468 ( .A(n3367), .B(n3772), .Y(n3794) );
  INVX1 U5469 ( .A(n3794), .Y(n6764) );
  AND2X1 U5470 ( .A(n3329), .B(n3806), .Y(n3809) );
  INVX1 U5471 ( .A(n3809), .Y(n6765) );
  AND2X1 U5472 ( .A(n3369), .B(n3806), .Y(n3829) );
  INVX1 U5473 ( .A(n3829), .Y(n6766) );
  AND2X1 U5474 ( .A(n3351), .B(n3840), .Y(n3854) );
  INVX1 U5475 ( .A(n3854), .Y(n6767) );
  AND2X1 U5476 ( .A(n3371), .B(n3840), .Y(n3864) );
  INVX1 U5477 ( .A(n3864), .Y(n6768) );
  AND2X1 U5478 ( .A(n3345), .B(n3874), .Y(n3885) );
  INVX1 U5479 ( .A(n3885), .Y(n6769) );
  AND2X1 U5480 ( .A(n3373), .B(n3874), .Y(n3899) );
  INVX1 U5481 ( .A(n3899), .Y(n6770) );
  AND2X1 U5482 ( .A(n3349), .B(n3908), .Y(n3921) );
  INVX1 U5483 ( .A(n3921), .Y(n6771) );
  AND2X1 U5484 ( .A(n3375), .B(n3908), .Y(n3934) );
  INVX1 U5485 ( .A(n3934), .Y(n6772) );
  AND2X1 U5486 ( .A(n3353), .B(n3943), .Y(n3958) );
  INVX1 U5487 ( .A(n3958), .Y(n6773) );
  AND2X1 U5488 ( .A(n3377), .B(n3943), .Y(n3970) );
  INVX1 U5489 ( .A(n3970), .Y(n6774) );
  AND2X1 U5490 ( .A(n3355), .B(n3977), .Y(n3993) );
  INVX1 U5491 ( .A(n3993), .Y(n6775) );
  AND2X1 U5492 ( .A(n3379), .B(n3977), .Y(n4005) );
  INVX1 U5493 ( .A(n4005), .Y(n6776) );
  AND2X1 U5494 ( .A(n3357), .B(n4011), .Y(n4028) );
  INVX1 U5495 ( .A(n4028), .Y(n6777) );
  AND2X1 U5496 ( .A(n3381), .B(n4011), .Y(n4040) );
  INVX1 U5497 ( .A(n4040), .Y(n6778) );
  AND2X1 U5498 ( .A(n3359), .B(n4045), .Y(n4063) );
  INVX1 U5499 ( .A(n4063), .Y(n6779) );
  AND2X1 U5500 ( .A(n3383), .B(n4045), .Y(n4075) );
  INVX1 U5501 ( .A(n4075), .Y(n6780) );
  AND2X1 U5502 ( .A(n3361), .B(n4079), .Y(n4098) );
  INVX1 U5503 ( .A(n4098), .Y(n6781) );
  AND2X1 U5504 ( .A(n3385), .B(n4079), .Y(n4110) );
  INVX1 U5505 ( .A(n4110), .Y(n6782) );
  AND2X1 U5506 ( .A(n3363), .B(n4113), .Y(n4133) );
  INVX1 U5507 ( .A(n4133), .Y(n6783) );
  AND2X1 U5508 ( .A(n3387), .B(n4113), .Y(n4145) );
  INVX1 U5509 ( .A(n4145), .Y(n6784) );
  AND2X1 U5510 ( .A(n3343), .B(n4147), .Y(n4157) );
  INVX1 U5511 ( .A(n4157), .Y(n6785) );
  AND2X1 U5512 ( .A(n3365), .B(n4147), .Y(n4168) );
  INVX1 U5513 ( .A(n4168), .Y(n6786) );
  AND2X1 U5514 ( .A(n3389), .B(n4147), .Y(n4180) );
  INVX1 U5515 ( .A(n4180), .Y(n6787) );
  AND2X1 U5516 ( .A(n3349), .B(n4181), .Y(n4194) );
  INVX1 U5517 ( .A(n4194), .Y(n6788) );
  AND2X1 U5518 ( .A(n3375), .B(n4181), .Y(n4207) );
  INVX1 U5519 ( .A(n4207), .Y(n6789) );
  AND2X1 U5520 ( .A(n3353), .B(n4216), .Y(n4231) );
  INVX1 U5521 ( .A(n4231), .Y(n6790) );
  AND2X1 U5522 ( .A(n3377), .B(n4216), .Y(n4243) );
  INVX1 U5523 ( .A(n4243), .Y(n6791) );
  AND2X1 U5524 ( .A(n3355), .B(n4250), .Y(n4266) );
  INVX1 U5525 ( .A(n4266), .Y(n6792) );
  AND2X1 U5526 ( .A(n3379), .B(n4250), .Y(n4278) );
  INVX1 U5527 ( .A(n4278), .Y(n6793) );
  AND2X1 U5528 ( .A(n3357), .B(n4284), .Y(n4301) );
  INVX1 U5529 ( .A(n4301), .Y(n6794) );
  AND2X1 U5530 ( .A(n3381), .B(n4284), .Y(n4313) );
  INVX1 U5531 ( .A(n4313), .Y(n6795) );
  AND2X1 U5532 ( .A(n3359), .B(n4318), .Y(n4336) );
  INVX1 U5533 ( .A(n4336), .Y(n6796) );
  AND2X1 U5534 ( .A(n3383), .B(n4318), .Y(n4348) );
  INVX1 U5535 ( .A(n4348), .Y(n6797) );
  AND2X1 U5536 ( .A(n3361), .B(n4352), .Y(n4371) );
  INVX1 U5537 ( .A(n4371), .Y(n6798) );
  AND2X1 U5538 ( .A(n3385), .B(n4352), .Y(n4383) );
  INVX1 U5539 ( .A(n4383), .Y(n6799) );
  AND2X1 U5540 ( .A(n3363), .B(n4386), .Y(n4406) );
  INVX1 U5541 ( .A(n4406), .Y(n6800) );
  AND2X1 U5542 ( .A(n3387), .B(n4386), .Y(n4418) );
  INVX1 U5543 ( .A(n4418), .Y(n6801) );
  AND2X1 U5544 ( .A(n3343), .B(n4420), .Y(n4430) );
  INVX1 U5545 ( .A(n4430), .Y(n6802) );
  AND2X1 U5546 ( .A(n3365), .B(n4420), .Y(n4441) );
  INVX1 U5547 ( .A(n4441), .Y(n6803) );
  AND2X1 U5548 ( .A(n3389), .B(n4420), .Y(n4453) );
  INVX1 U5549 ( .A(n4453), .Y(n6804) );
  AND2X1 U5550 ( .A(n3268), .B(n6856), .Y(n3260) );
  INVX1 U5551 ( .A(n3260), .Y(n6805) );
  AND2X1 U5552 ( .A(n12), .B(n6849), .Y(n4458) );
  INVX1 U5553 ( .A(n4458), .Y(n6806) );
  INVX1 U5554 ( .A(n3293), .Y(n6807) );
  BUFX2 U5555 ( .A(n3390), .Y(n6808) );
  BUFX2 U5556 ( .A(n4215), .Y(n6809) );
  INVX1 U5557 ( .A(n6819), .Y(n6816) );
  INVX1 U5558 ( .A(n6819), .Y(n6817) );
  INVX1 U5559 ( .A(n6844), .Y(n6842) );
  INVX1 U5560 ( .A(n6832), .Y(n6835) );
  INVX1 U5561 ( .A(n6832), .Y(n6836) );
  INVX1 U5562 ( .A(n6734), .Y(n6811) );
  INVX1 U5563 ( .A(n6734), .Y(n6810) );
  INVX1 U5564 ( .A(n6819), .Y(n6818) );
  INVX1 U5565 ( .A(n6815), .Y(n6814) );
  INVX1 U5566 ( .A(n6815), .Y(n6813) );
  INVX1 U5567 ( .A(n6815), .Y(n6812) );
  INVX1 U5568 ( .A(n1104), .Y(n6819) );
  INVX1 U5569 ( .A(n1105), .Y(n6815) );
  INVX1 U5570 ( .A(n1103), .Y(n6823) );
  INVX1 U5571 ( .A(n6844), .Y(n6843) );
  INVX1 U5572 ( .A(n6823), .Y(n6822) );
  INVX1 U5573 ( .A(n6823), .Y(n6821) );
  INVX1 U5574 ( .A(n6823), .Y(n6820) );
  INVX1 U5575 ( .A(reset), .Y(n6844) );
  INVX1 U5576 ( .A(n6841), .Y(n6840) );
  INVX1 U5577 ( .A(n6841), .Y(n6838) );
  INVX1 U5578 ( .A(n6831), .Y(n6829) );
  INVX1 U5579 ( .A(n6841), .Y(n6839) );
  INVX1 U5580 ( .A(n6831), .Y(n6828) );
  INVX1 U5581 ( .A(n6831), .Y(n6830) );
  INVX1 U5582 ( .A(n6827), .Y(n6826) );
  INVX1 U5583 ( .A(n6827), .Y(n6825) );
  INVX1 U5584 ( .A(n6827), .Y(n6824) );
  INVX1 U5585 ( .A(n6841), .Y(n6837) );
  INVX1 U5586 ( .A(n6832), .Y(n6833) );
  INVX1 U5587 ( .A(n6832), .Y(n6834) );
  INVX1 U5588 ( .A(n1096), .Y(n6841) );
  INVX1 U5589 ( .A(n1101), .Y(n6831) );
  INVX1 U5590 ( .A(n1102), .Y(n6827) );
  INVX1 U5591 ( .A(n3315), .Y(n6851) );
  INVX1 U5592 ( .A(n6594), .Y(n6852) );
  AND2X1 U5593 ( .A(n3288), .B(n6853), .Y(n1104) );
  AND2X1 U5594 ( .A(n3289), .B(n6853), .Y(n1105) );
  AND2X1 U5595 ( .A(n3287), .B(n6853), .Y(n1103) );
  AND2X1 U5596 ( .A(n6854), .B(n6855), .Y(n3288) );
  INVX1 U5597 ( .A(n6390), .Y(n6848) );
  INVX1 U5598 ( .A(n3290), .Y(fillcount[5]) );
  AND2X1 U5599 ( .A(n3276), .B(n16), .Y(n3268) );
  AND2X1 U5600 ( .A(n3268), .B(n15), .Y(n1108) );
  AND2X1 U5601 ( .A(n3289), .B(n12), .Y(n1096) );
  AND2X1 U5602 ( .A(n3288), .B(n12), .Y(n1101) );
  AND2X1 U5603 ( .A(n3287), .B(n12), .Y(n1102) );
  INVX1 U5604 ( .A(put), .Y(n7917) );
  INVX1 U5605 ( .A(wr_ptr[0]), .Y(n6849) );
  INVX1 U5606 ( .A(wr_ptr[3]), .Y(n6860) );
  INVX1 U5607 ( .A(n3317), .Y(n6850) );
  INVX1 U5608 ( .A(wr_ptr[2]), .Y(n6859) );
  INVX1 U5609 ( .A(n13), .Y(n6854) );
  INVX1 U5610 ( .A(n1097), .Y(n6832) );
  INVX1 U5611 ( .A(wr_ptr[4]), .Y(n6857) );
  INVX1 U5612 ( .A(n12), .Y(n6853) );
  INVX1 U5613 ( .A(n15), .Y(n6856) );
  INVX1 U5614 ( .A(n14), .Y(n6855) );
  INVX1 U5615 ( .A(wr_ptr[1]), .Y(n6858) );
  AND2X1 U5616 ( .A(n14), .B(n6854), .Y(n3287) );
  AND2X1 U5617 ( .A(n13), .B(n6855), .Y(n3289) );
  INVX1 U5618 ( .A(mem[726]), .Y(n7190) );
  INVX1 U5619 ( .A(mem[693]), .Y(n7223) );
  INVX1 U5620 ( .A(mem[594]), .Y(n7322) );
  INVX1 U5621 ( .A(mem[990]), .Y(n6926) );
  INVX1 U5622 ( .A(mem[957]), .Y(n6959) );
  INVX1 U5623 ( .A(mem[858]), .Y(n7058) );
  INVX1 U5624 ( .A(mem[198]), .Y(n7718) );
  INVX1 U5625 ( .A(mem[165]), .Y(n7751) );
  INVX1 U5626 ( .A(mem[66]), .Y(n7850) );
  INVX1 U5627 ( .A(mem[727]), .Y(n7189) );
  INVX1 U5628 ( .A(mem[694]), .Y(n7222) );
  INVX1 U5629 ( .A(mem[595]), .Y(n7321) );
  INVX1 U5630 ( .A(mem[991]), .Y(n6925) );
  INVX1 U5631 ( .A(mem[958]), .Y(n6958) );
  INVX1 U5632 ( .A(mem[859]), .Y(n7057) );
  INVX1 U5633 ( .A(mem[199]), .Y(n7717) );
  INVX1 U5634 ( .A(mem[166]), .Y(n7750) );
  INVX1 U5635 ( .A(mem[67]), .Y(n7849) );
  INVX1 U5636 ( .A(mem[728]), .Y(n7188) );
  INVX1 U5637 ( .A(mem[695]), .Y(n7221) );
  INVX1 U5638 ( .A(mem[596]), .Y(n7320) );
  INVX1 U5639 ( .A(mem[992]), .Y(n6924) );
  INVX1 U5640 ( .A(mem[959]), .Y(n6957) );
  INVX1 U5641 ( .A(mem[860]), .Y(n7056) );
  INVX1 U5642 ( .A(mem[200]), .Y(n7716) );
  INVX1 U5643 ( .A(mem[167]), .Y(n7749) );
  INVX1 U5644 ( .A(mem[68]), .Y(n7848) );
  INVX1 U5645 ( .A(mem[729]), .Y(n7187) );
  INVX1 U5646 ( .A(mem[696]), .Y(n7220) );
  INVX1 U5647 ( .A(mem[597]), .Y(n7319) );
  INVX1 U5648 ( .A(mem[993]), .Y(n6923) );
  INVX1 U5649 ( .A(mem[960]), .Y(n6956) );
  INVX1 U5650 ( .A(mem[861]), .Y(n7055) );
  INVX1 U5651 ( .A(mem[201]), .Y(n7715) );
  INVX1 U5652 ( .A(mem[168]), .Y(n7748) );
  INVX1 U5653 ( .A(mem[69]), .Y(n7847) );
  INVX1 U5654 ( .A(mem[730]), .Y(n7186) );
  INVX1 U5655 ( .A(mem[697]), .Y(n7219) );
  INVX1 U5656 ( .A(mem[598]), .Y(n7318) );
  INVX1 U5657 ( .A(mem[994]), .Y(n6922) );
  INVX1 U5658 ( .A(mem[961]), .Y(n6955) );
  INVX1 U5659 ( .A(mem[862]), .Y(n7054) );
  INVX1 U5660 ( .A(mem[202]), .Y(n7714) );
  INVX1 U5661 ( .A(mem[169]), .Y(n7747) );
  INVX1 U5662 ( .A(mem[70]), .Y(n7846) );
  INVX1 U5663 ( .A(mem[731]), .Y(n7185) );
  INVX1 U5664 ( .A(mem[698]), .Y(n7218) );
  INVX1 U5665 ( .A(mem[599]), .Y(n7317) );
  INVX1 U5666 ( .A(mem[995]), .Y(n6921) );
  INVX1 U5667 ( .A(mem[962]), .Y(n6954) );
  INVX1 U5668 ( .A(mem[863]), .Y(n7053) );
  INVX1 U5669 ( .A(mem[203]), .Y(n7713) );
  INVX1 U5670 ( .A(mem[170]), .Y(n7746) );
  INVX1 U5671 ( .A(mem[71]), .Y(n7845) );
  INVX1 U5672 ( .A(mem[732]), .Y(n7184) );
  INVX1 U5673 ( .A(mem[699]), .Y(n7217) );
  INVX1 U5674 ( .A(mem[600]), .Y(n7316) );
  INVX1 U5675 ( .A(mem[996]), .Y(n6920) );
  INVX1 U5676 ( .A(mem[963]), .Y(n6953) );
  INVX1 U5677 ( .A(mem[864]), .Y(n7052) );
  INVX1 U5678 ( .A(mem[204]), .Y(n7712) );
  INVX1 U5679 ( .A(mem[171]), .Y(n7745) );
  INVX1 U5680 ( .A(mem[72]), .Y(n7844) );
  INVX1 U5681 ( .A(mem[733]), .Y(n7183) );
  INVX1 U5682 ( .A(mem[700]), .Y(n7216) );
  INVX1 U5683 ( .A(mem[601]), .Y(n7315) );
  INVX1 U5684 ( .A(mem[997]), .Y(n6919) );
  INVX1 U5685 ( .A(mem[964]), .Y(n6952) );
  INVX1 U5686 ( .A(mem[865]), .Y(n7051) );
  INVX1 U5687 ( .A(mem[205]), .Y(n7711) );
  INVX1 U5688 ( .A(mem[172]), .Y(n7744) );
  INVX1 U5689 ( .A(mem[73]), .Y(n7843) );
  INVX1 U5690 ( .A(mem[734]), .Y(n7182) );
  INVX1 U5691 ( .A(mem[701]), .Y(n7215) );
  INVX1 U5692 ( .A(mem[602]), .Y(n7314) );
  INVX1 U5693 ( .A(mem[998]), .Y(n6918) );
  INVX1 U5694 ( .A(mem[965]), .Y(n6951) );
  INVX1 U5695 ( .A(mem[866]), .Y(n7050) );
  INVX1 U5696 ( .A(mem[206]), .Y(n7710) );
  INVX1 U5697 ( .A(mem[173]), .Y(n7743) );
  INVX1 U5698 ( .A(mem[74]), .Y(n7842) );
  INVX1 U5699 ( .A(mem[735]), .Y(n7181) );
  INVX1 U5700 ( .A(mem[702]), .Y(n7214) );
  INVX1 U5701 ( .A(mem[603]), .Y(n7313) );
  INVX1 U5702 ( .A(mem[999]), .Y(n6917) );
  INVX1 U5703 ( .A(mem[966]), .Y(n6950) );
  INVX1 U5704 ( .A(mem[867]), .Y(n7049) );
  INVX1 U5705 ( .A(mem[207]), .Y(n7709) );
  INVX1 U5706 ( .A(mem[174]), .Y(n7742) );
  INVX1 U5707 ( .A(mem[75]), .Y(n7841) );
  INVX1 U5708 ( .A(mem[736]), .Y(n7180) );
  INVX1 U5709 ( .A(mem[703]), .Y(n7213) );
  INVX1 U5710 ( .A(mem[604]), .Y(n7312) );
  INVX1 U5711 ( .A(mem[1000]), .Y(n6916) );
  INVX1 U5712 ( .A(mem[967]), .Y(n6949) );
  INVX1 U5713 ( .A(mem[868]), .Y(n7048) );
  INVX1 U5714 ( .A(mem[208]), .Y(n7708) );
  INVX1 U5715 ( .A(mem[175]), .Y(n7741) );
  INVX1 U5716 ( .A(mem[76]), .Y(n7840) );
  INVX1 U5717 ( .A(mem[737]), .Y(n7179) );
  INVX1 U5718 ( .A(mem[704]), .Y(n7212) );
  INVX1 U5719 ( .A(mem[605]), .Y(n7311) );
  INVX1 U5720 ( .A(mem[1001]), .Y(n6915) );
  INVX1 U5721 ( .A(mem[968]), .Y(n6948) );
  INVX1 U5722 ( .A(mem[869]), .Y(n7047) );
  INVX1 U5723 ( .A(mem[209]), .Y(n7707) );
  INVX1 U5724 ( .A(mem[176]), .Y(n7740) );
  INVX1 U5725 ( .A(mem[77]), .Y(n7839) );
  INVX1 U5726 ( .A(mem[738]), .Y(n7178) );
  INVX1 U5727 ( .A(mem[705]), .Y(n7211) );
  INVX1 U5728 ( .A(mem[606]), .Y(n7310) );
  INVX1 U5729 ( .A(mem[1002]), .Y(n6914) );
  INVX1 U5730 ( .A(mem[969]), .Y(n6947) );
  INVX1 U5731 ( .A(mem[870]), .Y(n7046) );
  INVX1 U5732 ( .A(mem[210]), .Y(n7706) );
  INVX1 U5733 ( .A(mem[177]), .Y(n7739) );
  INVX1 U5734 ( .A(mem[78]), .Y(n7838) );
  INVX1 U5735 ( .A(mem[739]), .Y(n7177) );
  INVX1 U5736 ( .A(mem[706]), .Y(n7210) );
  INVX1 U5737 ( .A(mem[607]), .Y(n7309) );
  INVX1 U5738 ( .A(mem[1003]), .Y(n6913) );
  INVX1 U5739 ( .A(mem[970]), .Y(n6946) );
  INVX1 U5740 ( .A(mem[871]), .Y(n7045) );
  INVX1 U5741 ( .A(mem[211]), .Y(n7705) );
  INVX1 U5742 ( .A(mem[178]), .Y(n7738) );
  INVX1 U5743 ( .A(mem[79]), .Y(n7837) );
  INVX1 U5744 ( .A(mem[740]), .Y(n7176) );
  INVX1 U5745 ( .A(mem[707]), .Y(n7209) );
  INVX1 U5746 ( .A(mem[608]), .Y(n7308) );
  INVX1 U5747 ( .A(mem[1004]), .Y(n6912) );
  INVX1 U5748 ( .A(mem[971]), .Y(n6945) );
  INVX1 U5749 ( .A(mem[872]), .Y(n7044) );
  INVX1 U5750 ( .A(mem[212]), .Y(n7704) );
  INVX1 U5751 ( .A(mem[179]), .Y(n7737) );
  INVX1 U5752 ( .A(mem[80]), .Y(n7836) );
  INVX1 U5753 ( .A(mem[741]), .Y(n7175) );
  INVX1 U5754 ( .A(mem[708]), .Y(n7208) );
  INVX1 U5755 ( .A(mem[609]), .Y(n7307) );
  INVX1 U5756 ( .A(mem[1005]), .Y(n6911) );
  INVX1 U5757 ( .A(mem[972]), .Y(n6944) );
  INVX1 U5758 ( .A(mem[873]), .Y(n7043) );
  INVX1 U5759 ( .A(mem[213]), .Y(n7703) );
  INVX1 U5760 ( .A(mem[180]), .Y(n7736) );
  INVX1 U5761 ( .A(mem[81]), .Y(n7835) );
  INVX1 U5762 ( .A(mem[742]), .Y(n7174) );
  INVX1 U5763 ( .A(mem[709]), .Y(n7207) );
  INVX1 U5764 ( .A(mem[610]), .Y(n7306) );
  INVX1 U5765 ( .A(mem[1006]), .Y(n6910) );
  INVX1 U5766 ( .A(mem[973]), .Y(n6943) );
  INVX1 U5767 ( .A(mem[874]), .Y(n7042) );
  INVX1 U5768 ( .A(mem[214]), .Y(n7702) );
  INVX1 U5769 ( .A(mem[181]), .Y(n7735) );
  INVX1 U5770 ( .A(mem[82]), .Y(n7834) );
  INVX1 U5771 ( .A(mem[743]), .Y(n7173) );
  INVX1 U5772 ( .A(mem[710]), .Y(n7206) );
  INVX1 U5773 ( .A(mem[611]), .Y(n7305) );
  INVX1 U5774 ( .A(mem[1007]), .Y(n6909) );
  INVX1 U5775 ( .A(mem[974]), .Y(n6942) );
  INVX1 U5776 ( .A(mem[875]), .Y(n7041) );
  INVX1 U5777 ( .A(mem[215]), .Y(n7701) );
  INVX1 U5778 ( .A(mem[182]), .Y(n7734) );
  INVX1 U5779 ( .A(mem[83]), .Y(n7833) );
  INVX1 U5780 ( .A(mem[744]), .Y(n7172) );
  INVX1 U5781 ( .A(mem[711]), .Y(n7205) );
  INVX1 U5782 ( .A(mem[612]), .Y(n7304) );
  INVX1 U5783 ( .A(mem[1008]), .Y(n6908) );
  INVX1 U5784 ( .A(mem[975]), .Y(n6941) );
  INVX1 U5785 ( .A(mem[876]), .Y(n7040) );
  INVX1 U5786 ( .A(mem[216]), .Y(n7700) );
  INVX1 U5787 ( .A(mem[183]), .Y(n7733) );
  INVX1 U5788 ( .A(mem[84]), .Y(n7832) );
  INVX1 U5789 ( .A(mem[745]), .Y(n7171) );
  INVX1 U5790 ( .A(mem[712]), .Y(n7204) );
  INVX1 U5791 ( .A(mem[613]), .Y(n7303) );
  INVX1 U5792 ( .A(mem[1009]), .Y(n6907) );
  INVX1 U5793 ( .A(mem[976]), .Y(n6940) );
  INVX1 U5794 ( .A(mem[877]), .Y(n7039) );
  INVX1 U5795 ( .A(mem[217]), .Y(n7699) );
  INVX1 U5796 ( .A(mem[184]), .Y(n7732) );
  INVX1 U5797 ( .A(mem[85]), .Y(n7831) );
  INVX1 U5798 ( .A(mem[746]), .Y(n7170) );
  INVX1 U5799 ( .A(mem[713]), .Y(n7203) );
  INVX1 U5800 ( .A(mem[614]), .Y(n7302) );
  INVX1 U5801 ( .A(mem[1010]), .Y(n6906) );
  INVX1 U5802 ( .A(mem[977]), .Y(n6939) );
  INVX1 U5803 ( .A(mem[878]), .Y(n7038) );
  INVX1 U5804 ( .A(mem[218]), .Y(n7698) );
  INVX1 U5805 ( .A(mem[185]), .Y(n7731) );
  INVX1 U5806 ( .A(mem[86]), .Y(n7830) );
  INVX1 U5807 ( .A(mem[747]), .Y(n7169) );
  INVX1 U5808 ( .A(mem[714]), .Y(n7202) );
  INVX1 U5809 ( .A(mem[615]), .Y(n7301) );
  INVX1 U5810 ( .A(mem[1011]), .Y(n6905) );
  INVX1 U5811 ( .A(mem[978]), .Y(n6938) );
  INVX1 U5812 ( .A(mem[879]), .Y(n7037) );
  INVX1 U5813 ( .A(mem[219]), .Y(n7697) );
  INVX1 U5814 ( .A(mem[186]), .Y(n7730) );
  INVX1 U5815 ( .A(mem[87]), .Y(n7829) );
  INVX1 U5816 ( .A(mem[748]), .Y(n7168) );
  INVX1 U5817 ( .A(mem[715]), .Y(n7201) );
  INVX1 U5818 ( .A(mem[616]), .Y(n7300) );
  INVX1 U5819 ( .A(mem[1012]), .Y(n6904) );
  INVX1 U5820 ( .A(mem[979]), .Y(n6937) );
  INVX1 U5821 ( .A(mem[880]), .Y(n7036) );
  INVX1 U5822 ( .A(mem[220]), .Y(n7696) );
  INVX1 U5823 ( .A(mem[187]), .Y(n7729) );
  INVX1 U5824 ( .A(mem[88]), .Y(n7828) );
  INVX1 U5825 ( .A(mem[749]), .Y(n7167) );
  INVX1 U5826 ( .A(mem[716]), .Y(n7200) );
  INVX1 U5827 ( .A(mem[617]), .Y(n7299) );
  INVX1 U5828 ( .A(mem[1013]), .Y(n6903) );
  INVX1 U5829 ( .A(mem[980]), .Y(n6936) );
  INVX1 U5830 ( .A(mem[881]), .Y(n7035) );
  INVX1 U5831 ( .A(mem[221]), .Y(n7695) );
  INVX1 U5832 ( .A(mem[188]), .Y(n7728) );
  INVX1 U5833 ( .A(mem[89]), .Y(n7827) );
  INVX1 U5834 ( .A(mem[750]), .Y(n7166) );
  INVX1 U5835 ( .A(mem[717]), .Y(n7199) );
  INVX1 U5836 ( .A(mem[618]), .Y(n7298) );
  INVX1 U5837 ( .A(mem[1014]), .Y(n6902) );
  INVX1 U5838 ( .A(mem[981]), .Y(n6935) );
  INVX1 U5839 ( .A(mem[882]), .Y(n7034) );
  INVX1 U5840 ( .A(mem[222]), .Y(n7694) );
  INVX1 U5841 ( .A(mem[189]), .Y(n7727) );
  INVX1 U5842 ( .A(mem[90]), .Y(n7826) );
  INVX1 U5843 ( .A(mem[751]), .Y(n7165) );
  INVX1 U5844 ( .A(mem[718]), .Y(n7198) );
  INVX1 U5845 ( .A(mem[619]), .Y(n7297) );
  INVX1 U5846 ( .A(mem[1015]), .Y(n6901) );
  INVX1 U5847 ( .A(mem[982]), .Y(n6934) );
  INVX1 U5848 ( .A(mem[883]), .Y(n7033) );
  INVX1 U5849 ( .A(mem[223]), .Y(n7693) );
  INVX1 U5850 ( .A(mem[190]), .Y(n7726) );
  INVX1 U5851 ( .A(mem[91]), .Y(n7825) );
  INVX1 U5852 ( .A(mem[752]), .Y(n7164) );
  INVX1 U5853 ( .A(mem[719]), .Y(n7197) );
  INVX1 U5854 ( .A(mem[620]), .Y(n7296) );
  INVX1 U5855 ( .A(mem[1016]), .Y(n6900) );
  INVX1 U5856 ( .A(mem[983]), .Y(n6933) );
  INVX1 U5857 ( .A(mem[884]), .Y(n7032) );
  INVX1 U5858 ( .A(mem[224]), .Y(n7692) );
  INVX1 U5859 ( .A(mem[191]), .Y(n7725) );
  INVX1 U5860 ( .A(mem[92]), .Y(n7824) );
  INVX1 U5861 ( .A(mem[753]), .Y(n7163) );
  INVX1 U5862 ( .A(mem[720]), .Y(n7196) );
  INVX1 U5863 ( .A(mem[621]), .Y(n7295) );
  INVX1 U5864 ( .A(mem[1017]), .Y(n6899) );
  INVX1 U5865 ( .A(mem[984]), .Y(n6932) );
  INVX1 U5866 ( .A(mem[885]), .Y(n7031) );
  INVX1 U5867 ( .A(mem[225]), .Y(n7691) );
  INVX1 U5868 ( .A(mem[192]), .Y(n7724) );
  INVX1 U5869 ( .A(mem[93]), .Y(n7823) );
  INVX1 U5870 ( .A(mem[754]), .Y(n7162) );
  INVX1 U5871 ( .A(mem[721]), .Y(n7195) );
  INVX1 U5872 ( .A(mem[622]), .Y(n7294) );
  INVX1 U5873 ( .A(mem[1018]), .Y(n6898) );
  INVX1 U5874 ( .A(mem[985]), .Y(n6931) );
  INVX1 U5875 ( .A(mem[886]), .Y(n7030) );
  INVX1 U5876 ( .A(mem[226]), .Y(n7690) );
  INVX1 U5877 ( .A(mem[193]), .Y(n7723) );
  INVX1 U5878 ( .A(mem[94]), .Y(n7822) );
  INVX1 U5879 ( .A(mem[755]), .Y(n7161) );
  INVX1 U5880 ( .A(mem[722]), .Y(n7194) );
  INVX1 U5881 ( .A(mem[623]), .Y(n7293) );
  INVX1 U5882 ( .A(mem[1019]), .Y(n6897) );
  INVX1 U5883 ( .A(mem[986]), .Y(n6930) );
  INVX1 U5884 ( .A(mem[887]), .Y(n7029) );
  INVX1 U5885 ( .A(mem[227]), .Y(n7689) );
  INVX1 U5886 ( .A(mem[194]), .Y(n7722) );
  INVX1 U5887 ( .A(mem[95]), .Y(n7821) );
  INVX1 U5888 ( .A(mem[756]), .Y(n7160) );
  INVX1 U5889 ( .A(mem[723]), .Y(n7193) );
  INVX1 U5890 ( .A(mem[624]), .Y(n7292) );
  INVX1 U5891 ( .A(mem[1020]), .Y(n6896) );
  INVX1 U5892 ( .A(mem[987]), .Y(n6929) );
  INVX1 U5893 ( .A(mem[888]), .Y(n7028) );
  INVX1 U5894 ( .A(mem[228]), .Y(n7688) );
  INVX1 U5895 ( .A(mem[195]), .Y(n7721) );
  INVX1 U5896 ( .A(mem[96]), .Y(n7820) );
  INVX1 U5897 ( .A(mem[757]), .Y(n7159) );
  INVX1 U5898 ( .A(mem[724]), .Y(n7192) );
  INVX1 U5899 ( .A(mem[625]), .Y(n7291) );
  INVX1 U5900 ( .A(mem[1021]), .Y(n6895) );
  INVX1 U5901 ( .A(mem[988]), .Y(n6928) );
  INVX1 U5902 ( .A(mem[889]), .Y(n7027) );
  INVX1 U5903 ( .A(mem[229]), .Y(n7687) );
  INVX1 U5904 ( .A(mem[196]), .Y(n7720) );
  INVX1 U5905 ( .A(mem[97]), .Y(n7819) );
  INVX1 U5906 ( .A(mem[758]), .Y(n7158) );
  INVX1 U5907 ( .A(mem[725]), .Y(n7191) );
  INVX1 U5908 ( .A(mem[626]), .Y(n7290) );
  INVX1 U5909 ( .A(mem[1022]), .Y(n6894) );
  INVX1 U5910 ( .A(mem[989]), .Y(n6927) );
  INVX1 U5911 ( .A(mem[890]), .Y(n7026) );
  INVX1 U5912 ( .A(mem[230]), .Y(n7686) );
  INVX1 U5913 ( .A(mem[197]), .Y(n7719) );
  INVX1 U5914 ( .A(mem[98]), .Y(n7818) );
  INVX1 U5915 ( .A(mem[462]), .Y(n7454) );
  INVX1 U5916 ( .A(mem[429]), .Y(n7487) );
  INVX1 U5917 ( .A(mem[330]), .Y(n7586) );
  INVX1 U5918 ( .A(mem[463]), .Y(n7453) );
  INVX1 U5919 ( .A(mem[430]), .Y(n7486) );
  INVX1 U5920 ( .A(mem[331]), .Y(n7585) );
  INVX1 U5921 ( .A(mem[464]), .Y(n7452) );
  INVX1 U5922 ( .A(mem[431]), .Y(n7485) );
  INVX1 U5923 ( .A(mem[332]), .Y(n7584) );
  INVX1 U5924 ( .A(mem[465]), .Y(n7451) );
  INVX1 U5925 ( .A(mem[432]), .Y(n7484) );
  INVX1 U5926 ( .A(mem[333]), .Y(n7583) );
  INVX1 U5927 ( .A(mem[466]), .Y(n7450) );
  INVX1 U5928 ( .A(mem[433]), .Y(n7483) );
  INVX1 U5929 ( .A(mem[334]), .Y(n7582) );
  INVX1 U5930 ( .A(mem[467]), .Y(n7449) );
  INVX1 U5931 ( .A(mem[434]), .Y(n7482) );
  INVX1 U5932 ( .A(mem[335]), .Y(n7581) );
  INVX1 U5933 ( .A(mem[468]), .Y(n7448) );
  INVX1 U5934 ( .A(mem[435]), .Y(n7481) );
  INVX1 U5935 ( .A(mem[336]), .Y(n7580) );
  INVX1 U5936 ( .A(mem[469]), .Y(n7447) );
  INVX1 U5937 ( .A(mem[436]), .Y(n7480) );
  INVX1 U5938 ( .A(mem[337]), .Y(n7579) );
  INVX1 U5939 ( .A(mem[470]), .Y(n7446) );
  INVX1 U5940 ( .A(mem[437]), .Y(n7479) );
  INVX1 U5941 ( .A(mem[338]), .Y(n7578) );
  INVX1 U5942 ( .A(mem[471]), .Y(n7445) );
  INVX1 U5943 ( .A(mem[438]), .Y(n7478) );
  INVX1 U5944 ( .A(mem[339]), .Y(n7577) );
  INVX1 U5945 ( .A(mem[472]), .Y(n7444) );
  INVX1 U5946 ( .A(mem[439]), .Y(n7477) );
  INVX1 U5947 ( .A(mem[340]), .Y(n7576) );
  INVX1 U5948 ( .A(mem[473]), .Y(n7443) );
  INVX1 U5949 ( .A(mem[440]), .Y(n7476) );
  INVX1 U5950 ( .A(mem[341]), .Y(n7575) );
  INVX1 U5951 ( .A(mem[474]), .Y(n7442) );
  INVX1 U5952 ( .A(mem[441]), .Y(n7475) );
  INVX1 U5953 ( .A(mem[342]), .Y(n7574) );
  INVX1 U5954 ( .A(mem[475]), .Y(n7441) );
  INVX1 U5955 ( .A(mem[442]), .Y(n7474) );
  INVX1 U5956 ( .A(mem[343]), .Y(n7573) );
  INVX1 U5957 ( .A(mem[476]), .Y(n7440) );
  INVX1 U5958 ( .A(mem[443]), .Y(n7473) );
  INVX1 U5959 ( .A(mem[344]), .Y(n7572) );
  INVX1 U5960 ( .A(mem[477]), .Y(n7439) );
  INVX1 U5961 ( .A(mem[444]), .Y(n7472) );
  INVX1 U5962 ( .A(mem[345]), .Y(n7571) );
  INVX1 U5963 ( .A(mem[478]), .Y(n7438) );
  INVX1 U5964 ( .A(mem[445]), .Y(n7471) );
  INVX1 U5965 ( .A(mem[346]), .Y(n7570) );
  INVX1 U5966 ( .A(mem[479]), .Y(n7437) );
  INVX1 U5967 ( .A(mem[446]), .Y(n7470) );
  INVX1 U5968 ( .A(mem[347]), .Y(n7569) );
  INVX1 U5969 ( .A(mem[480]), .Y(n7436) );
  INVX1 U5970 ( .A(mem[447]), .Y(n7469) );
  INVX1 U5971 ( .A(mem[348]), .Y(n7568) );
  INVX1 U5972 ( .A(mem[481]), .Y(n7435) );
  INVX1 U5973 ( .A(mem[448]), .Y(n7468) );
  INVX1 U5974 ( .A(mem[349]), .Y(n7567) );
  INVX1 U5975 ( .A(mem[482]), .Y(n7434) );
  INVX1 U5976 ( .A(mem[449]), .Y(n7467) );
  INVX1 U5977 ( .A(mem[350]), .Y(n7566) );
  INVX1 U5978 ( .A(mem[483]), .Y(n7433) );
  INVX1 U5979 ( .A(mem[450]), .Y(n7466) );
  INVX1 U5980 ( .A(mem[351]), .Y(n7565) );
  INVX1 U5981 ( .A(mem[484]), .Y(n7432) );
  INVX1 U5982 ( .A(mem[451]), .Y(n7465) );
  INVX1 U5983 ( .A(mem[352]), .Y(n7564) );
  INVX1 U5984 ( .A(mem[485]), .Y(n7431) );
  INVX1 U5985 ( .A(mem[452]), .Y(n7464) );
  INVX1 U5986 ( .A(mem[353]), .Y(n7563) );
  INVX1 U5987 ( .A(mem[486]), .Y(n7430) );
  INVX1 U5988 ( .A(mem[453]), .Y(n7463) );
  INVX1 U5989 ( .A(mem[354]), .Y(n7562) );
  INVX1 U5990 ( .A(mem[487]), .Y(n7429) );
  INVX1 U5991 ( .A(mem[454]), .Y(n7462) );
  INVX1 U5992 ( .A(mem[355]), .Y(n7561) );
  INVX1 U5993 ( .A(mem[488]), .Y(n7428) );
  INVX1 U5994 ( .A(mem[455]), .Y(n7461) );
  INVX1 U5995 ( .A(mem[356]), .Y(n7560) );
  INVX1 U5996 ( .A(mem[489]), .Y(n7427) );
  INVX1 U5997 ( .A(mem[456]), .Y(n7460) );
  INVX1 U5998 ( .A(mem[357]), .Y(n7559) );
  INVX1 U5999 ( .A(mem[490]), .Y(n7426) );
  INVX1 U6000 ( .A(mem[457]), .Y(n7459) );
  INVX1 U6001 ( .A(mem[358]), .Y(n7558) );
  INVX1 U6002 ( .A(mem[491]), .Y(n7425) );
  INVX1 U6003 ( .A(mem[458]), .Y(n7458) );
  INVX1 U6004 ( .A(mem[359]), .Y(n7557) );
  INVX1 U6005 ( .A(mem[492]), .Y(n7424) );
  INVX1 U6006 ( .A(mem[459]), .Y(n7457) );
  INVX1 U6007 ( .A(mem[360]), .Y(n7556) );
  INVX1 U6008 ( .A(mem[493]), .Y(n7423) );
  INVX1 U6009 ( .A(mem[460]), .Y(n7456) );
  INVX1 U6010 ( .A(mem[361]), .Y(n7555) );
  INVX1 U6011 ( .A(mem[494]), .Y(n7422) );
  INVX1 U6012 ( .A(mem[461]), .Y(n7455) );
  INVX1 U6013 ( .A(mem[362]), .Y(n7554) );
  INVX1 U6014 ( .A(mem[627]), .Y(n7289) );
  INVX1 U6015 ( .A(mem[561]), .Y(n7355) );
  INVX1 U6016 ( .A(mem[528]), .Y(n7388) );
  INVX1 U6017 ( .A(mem[891]), .Y(n7025) );
  INVX1 U6018 ( .A(mem[825]), .Y(n7091) );
  INVX1 U6019 ( .A(mem[792]), .Y(n7124) );
  INVX1 U6020 ( .A(mem[99]), .Y(n7817) );
  INVX1 U6021 ( .A(mem[33]), .Y(n7883) );
  INVX1 U6022 ( .A(mem[0]), .Y(n7916) );
  INVX1 U6023 ( .A(mem[628]), .Y(n7288) );
  INVX1 U6024 ( .A(mem[562]), .Y(n7354) );
  INVX1 U6025 ( .A(mem[529]), .Y(n7387) );
  INVX1 U6026 ( .A(mem[892]), .Y(n7024) );
  INVX1 U6027 ( .A(mem[826]), .Y(n7090) );
  INVX1 U6028 ( .A(mem[793]), .Y(n7123) );
  INVX1 U6029 ( .A(mem[100]), .Y(n7816) );
  INVX1 U6030 ( .A(mem[34]), .Y(n7882) );
  INVX1 U6031 ( .A(mem[1]), .Y(n7915) );
  INVX1 U6032 ( .A(mem[629]), .Y(n7287) );
  INVX1 U6033 ( .A(mem[563]), .Y(n7353) );
  INVX1 U6034 ( .A(mem[530]), .Y(n7386) );
  INVX1 U6035 ( .A(mem[893]), .Y(n7023) );
  INVX1 U6036 ( .A(mem[827]), .Y(n7089) );
  INVX1 U6037 ( .A(mem[794]), .Y(n7122) );
  INVX1 U6038 ( .A(mem[101]), .Y(n7815) );
  INVX1 U6039 ( .A(mem[35]), .Y(n7881) );
  INVX1 U6040 ( .A(mem[2]), .Y(n7914) );
  INVX1 U6041 ( .A(mem[630]), .Y(n7286) );
  INVX1 U6042 ( .A(mem[564]), .Y(n7352) );
  INVX1 U6043 ( .A(mem[531]), .Y(n7385) );
  INVX1 U6044 ( .A(mem[894]), .Y(n7022) );
  INVX1 U6045 ( .A(mem[828]), .Y(n7088) );
  INVX1 U6046 ( .A(mem[795]), .Y(n7121) );
  INVX1 U6047 ( .A(mem[102]), .Y(n7814) );
  INVX1 U6048 ( .A(mem[36]), .Y(n7880) );
  INVX1 U6049 ( .A(mem[3]), .Y(n7913) );
  INVX1 U6050 ( .A(mem[631]), .Y(n7285) );
  INVX1 U6051 ( .A(mem[565]), .Y(n7351) );
  INVX1 U6052 ( .A(mem[532]), .Y(n7384) );
  INVX1 U6053 ( .A(mem[895]), .Y(n7021) );
  INVX1 U6054 ( .A(mem[829]), .Y(n7087) );
  INVX1 U6055 ( .A(mem[796]), .Y(n7120) );
  INVX1 U6056 ( .A(mem[103]), .Y(n7813) );
  INVX1 U6057 ( .A(mem[37]), .Y(n7879) );
  INVX1 U6058 ( .A(mem[4]), .Y(n7912) );
  INVX1 U6059 ( .A(mem[632]), .Y(n7284) );
  INVX1 U6060 ( .A(mem[566]), .Y(n7350) );
  INVX1 U6061 ( .A(mem[533]), .Y(n7383) );
  INVX1 U6062 ( .A(mem[896]), .Y(n7020) );
  INVX1 U6063 ( .A(mem[830]), .Y(n7086) );
  INVX1 U6064 ( .A(mem[797]), .Y(n7119) );
  INVX1 U6065 ( .A(mem[104]), .Y(n7812) );
  INVX1 U6066 ( .A(mem[38]), .Y(n7878) );
  INVX1 U6067 ( .A(mem[5]), .Y(n7911) );
  INVX1 U6068 ( .A(mem[633]), .Y(n7283) );
  INVX1 U6069 ( .A(mem[567]), .Y(n7349) );
  INVX1 U6070 ( .A(mem[534]), .Y(n7382) );
  INVX1 U6071 ( .A(mem[897]), .Y(n7019) );
  INVX1 U6072 ( .A(mem[831]), .Y(n7085) );
  INVX1 U6073 ( .A(mem[798]), .Y(n7118) );
  INVX1 U6074 ( .A(mem[105]), .Y(n7811) );
  INVX1 U6075 ( .A(mem[39]), .Y(n7877) );
  INVX1 U6076 ( .A(mem[6]), .Y(n7910) );
  INVX1 U6077 ( .A(mem[634]), .Y(n7282) );
  INVX1 U6078 ( .A(mem[568]), .Y(n7348) );
  INVX1 U6079 ( .A(mem[535]), .Y(n7381) );
  INVX1 U6080 ( .A(mem[898]), .Y(n7018) );
  INVX1 U6081 ( .A(mem[832]), .Y(n7084) );
  INVX1 U6082 ( .A(mem[799]), .Y(n7117) );
  INVX1 U6083 ( .A(mem[106]), .Y(n7810) );
  INVX1 U6084 ( .A(mem[40]), .Y(n7876) );
  INVX1 U6085 ( .A(mem[7]), .Y(n7909) );
  INVX1 U6086 ( .A(mem[635]), .Y(n7281) );
  INVX1 U6087 ( .A(mem[569]), .Y(n7347) );
  INVX1 U6088 ( .A(mem[536]), .Y(n7380) );
  INVX1 U6089 ( .A(mem[899]), .Y(n7017) );
  INVX1 U6090 ( .A(mem[833]), .Y(n7083) );
  INVX1 U6091 ( .A(mem[800]), .Y(n7116) );
  INVX1 U6092 ( .A(mem[107]), .Y(n7809) );
  INVX1 U6093 ( .A(mem[41]), .Y(n7875) );
  INVX1 U6094 ( .A(mem[8]), .Y(n7908) );
  INVX1 U6095 ( .A(mem[636]), .Y(n7280) );
  INVX1 U6096 ( .A(mem[570]), .Y(n7346) );
  INVX1 U6097 ( .A(mem[537]), .Y(n7379) );
  INVX1 U6098 ( .A(mem[900]), .Y(n7016) );
  INVX1 U6099 ( .A(mem[834]), .Y(n7082) );
  INVX1 U6100 ( .A(mem[801]), .Y(n7115) );
  INVX1 U6101 ( .A(mem[108]), .Y(n7808) );
  INVX1 U6102 ( .A(mem[42]), .Y(n7874) );
  INVX1 U6103 ( .A(mem[9]), .Y(n7907) );
  INVX1 U6104 ( .A(mem[637]), .Y(n7279) );
  INVX1 U6105 ( .A(mem[571]), .Y(n7345) );
  INVX1 U6106 ( .A(mem[538]), .Y(n7378) );
  INVX1 U6107 ( .A(mem[901]), .Y(n7015) );
  INVX1 U6108 ( .A(mem[835]), .Y(n7081) );
  INVX1 U6109 ( .A(mem[802]), .Y(n7114) );
  INVX1 U6110 ( .A(mem[109]), .Y(n7807) );
  INVX1 U6111 ( .A(mem[43]), .Y(n7873) );
  INVX1 U6112 ( .A(mem[10]), .Y(n7906) );
  INVX1 U6113 ( .A(mem[638]), .Y(n7278) );
  INVX1 U6114 ( .A(mem[572]), .Y(n7344) );
  INVX1 U6115 ( .A(mem[539]), .Y(n7377) );
  INVX1 U6116 ( .A(mem[902]), .Y(n7014) );
  INVX1 U6117 ( .A(mem[836]), .Y(n7080) );
  INVX1 U6118 ( .A(mem[803]), .Y(n7113) );
  INVX1 U6119 ( .A(mem[110]), .Y(n7806) );
  INVX1 U6120 ( .A(mem[44]), .Y(n7872) );
  INVX1 U6121 ( .A(mem[11]), .Y(n7905) );
  INVX1 U6122 ( .A(mem[639]), .Y(n7277) );
  INVX1 U6123 ( .A(mem[573]), .Y(n7343) );
  INVX1 U6124 ( .A(mem[540]), .Y(n7376) );
  INVX1 U6125 ( .A(mem[903]), .Y(n7013) );
  INVX1 U6126 ( .A(mem[837]), .Y(n7079) );
  INVX1 U6127 ( .A(mem[804]), .Y(n7112) );
  INVX1 U6128 ( .A(mem[111]), .Y(n7805) );
  INVX1 U6129 ( .A(mem[45]), .Y(n7871) );
  INVX1 U6130 ( .A(mem[12]), .Y(n7904) );
  INVX1 U6131 ( .A(mem[640]), .Y(n7276) );
  INVX1 U6132 ( .A(mem[574]), .Y(n7342) );
  INVX1 U6133 ( .A(mem[541]), .Y(n7375) );
  INVX1 U6134 ( .A(mem[904]), .Y(n7012) );
  INVX1 U6135 ( .A(mem[838]), .Y(n7078) );
  INVX1 U6136 ( .A(mem[805]), .Y(n7111) );
  INVX1 U6137 ( .A(mem[112]), .Y(n7804) );
  INVX1 U6138 ( .A(mem[46]), .Y(n7870) );
  INVX1 U6139 ( .A(mem[13]), .Y(n7903) );
  INVX1 U6140 ( .A(mem[641]), .Y(n7275) );
  INVX1 U6141 ( .A(mem[575]), .Y(n7341) );
  INVX1 U6142 ( .A(mem[542]), .Y(n7374) );
  INVX1 U6143 ( .A(mem[905]), .Y(n7011) );
  INVX1 U6144 ( .A(mem[839]), .Y(n7077) );
  INVX1 U6145 ( .A(mem[806]), .Y(n7110) );
  INVX1 U6146 ( .A(mem[113]), .Y(n7803) );
  INVX1 U6147 ( .A(mem[47]), .Y(n7869) );
  INVX1 U6148 ( .A(mem[14]), .Y(n7902) );
  INVX1 U6149 ( .A(mem[642]), .Y(n7274) );
  INVX1 U6150 ( .A(mem[576]), .Y(n7340) );
  INVX1 U6151 ( .A(mem[543]), .Y(n7373) );
  INVX1 U6152 ( .A(mem[906]), .Y(n7010) );
  INVX1 U6153 ( .A(mem[840]), .Y(n7076) );
  INVX1 U6154 ( .A(mem[807]), .Y(n7109) );
  INVX1 U6155 ( .A(mem[114]), .Y(n7802) );
  INVX1 U6156 ( .A(mem[48]), .Y(n7868) );
  INVX1 U6157 ( .A(mem[15]), .Y(n7901) );
  INVX1 U6158 ( .A(mem[643]), .Y(n7273) );
  INVX1 U6159 ( .A(mem[577]), .Y(n7339) );
  INVX1 U6160 ( .A(mem[544]), .Y(n7372) );
  INVX1 U6161 ( .A(mem[907]), .Y(n7009) );
  INVX1 U6162 ( .A(mem[841]), .Y(n7075) );
  INVX1 U6163 ( .A(mem[808]), .Y(n7108) );
  INVX1 U6164 ( .A(mem[115]), .Y(n7801) );
  INVX1 U6165 ( .A(mem[49]), .Y(n7867) );
  INVX1 U6166 ( .A(mem[16]), .Y(n7900) );
  INVX1 U6167 ( .A(mem[644]), .Y(n7272) );
  INVX1 U6168 ( .A(mem[578]), .Y(n7338) );
  INVX1 U6169 ( .A(mem[545]), .Y(n7371) );
  INVX1 U6170 ( .A(mem[908]), .Y(n7008) );
  INVX1 U6171 ( .A(mem[842]), .Y(n7074) );
  INVX1 U6172 ( .A(mem[809]), .Y(n7107) );
  INVX1 U6173 ( .A(mem[116]), .Y(n7800) );
  INVX1 U6174 ( .A(mem[50]), .Y(n7866) );
  INVX1 U6175 ( .A(mem[17]), .Y(n7899) );
  INVX1 U6176 ( .A(mem[645]), .Y(n7271) );
  INVX1 U6177 ( .A(mem[579]), .Y(n7337) );
  INVX1 U6178 ( .A(mem[546]), .Y(n7370) );
  INVX1 U6179 ( .A(mem[909]), .Y(n7007) );
  INVX1 U6180 ( .A(mem[843]), .Y(n7073) );
  INVX1 U6181 ( .A(mem[810]), .Y(n7106) );
  INVX1 U6182 ( .A(mem[117]), .Y(n7799) );
  INVX1 U6183 ( .A(mem[51]), .Y(n7865) );
  INVX1 U6184 ( .A(mem[18]), .Y(n7898) );
  INVX1 U6185 ( .A(mem[646]), .Y(n7270) );
  INVX1 U6186 ( .A(mem[580]), .Y(n7336) );
  INVX1 U6187 ( .A(mem[547]), .Y(n7369) );
  INVX1 U6188 ( .A(mem[910]), .Y(n7006) );
  INVX1 U6189 ( .A(mem[844]), .Y(n7072) );
  INVX1 U6190 ( .A(mem[811]), .Y(n7105) );
  INVX1 U6191 ( .A(mem[118]), .Y(n7798) );
  INVX1 U6192 ( .A(mem[52]), .Y(n7864) );
  INVX1 U6193 ( .A(mem[19]), .Y(n7897) );
  INVX1 U6194 ( .A(mem[647]), .Y(n7269) );
  INVX1 U6195 ( .A(mem[581]), .Y(n7335) );
  INVX1 U6196 ( .A(mem[548]), .Y(n7368) );
  INVX1 U6197 ( .A(mem[911]), .Y(n7005) );
  INVX1 U6198 ( .A(mem[845]), .Y(n7071) );
  INVX1 U6199 ( .A(mem[812]), .Y(n7104) );
  INVX1 U6200 ( .A(mem[119]), .Y(n7797) );
  INVX1 U6201 ( .A(mem[53]), .Y(n7863) );
  INVX1 U6202 ( .A(mem[20]), .Y(n7896) );
  INVX1 U6203 ( .A(mem[648]), .Y(n7268) );
  INVX1 U6204 ( .A(mem[582]), .Y(n7334) );
  INVX1 U6205 ( .A(mem[549]), .Y(n7367) );
  INVX1 U6206 ( .A(mem[912]), .Y(n7004) );
  INVX1 U6207 ( .A(mem[846]), .Y(n7070) );
  INVX1 U6208 ( .A(mem[813]), .Y(n7103) );
  INVX1 U6209 ( .A(mem[120]), .Y(n7796) );
  INVX1 U6210 ( .A(mem[54]), .Y(n7862) );
  INVX1 U6211 ( .A(mem[21]), .Y(n7895) );
  INVX1 U6212 ( .A(mem[649]), .Y(n7267) );
  INVX1 U6213 ( .A(mem[583]), .Y(n7333) );
  INVX1 U6214 ( .A(mem[550]), .Y(n7366) );
  INVX1 U6215 ( .A(mem[913]), .Y(n7003) );
  INVX1 U6216 ( .A(mem[847]), .Y(n7069) );
  INVX1 U6217 ( .A(mem[814]), .Y(n7102) );
  INVX1 U6218 ( .A(mem[121]), .Y(n7795) );
  INVX1 U6219 ( .A(mem[55]), .Y(n7861) );
  INVX1 U6220 ( .A(mem[22]), .Y(n7894) );
  INVX1 U6221 ( .A(mem[650]), .Y(n7266) );
  INVX1 U6222 ( .A(mem[584]), .Y(n7332) );
  INVX1 U6223 ( .A(mem[551]), .Y(n7365) );
  INVX1 U6224 ( .A(mem[914]), .Y(n7002) );
  INVX1 U6225 ( .A(mem[848]), .Y(n7068) );
  INVX1 U6226 ( .A(mem[815]), .Y(n7101) );
  INVX1 U6227 ( .A(mem[122]), .Y(n7794) );
  INVX1 U6228 ( .A(mem[56]), .Y(n7860) );
  INVX1 U6229 ( .A(mem[23]), .Y(n7893) );
  INVX1 U6230 ( .A(mem[651]), .Y(n7265) );
  INVX1 U6231 ( .A(mem[585]), .Y(n7331) );
  INVX1 U6232 ( .A(mem[552]), .Y(n7364) );
  INVX1 U6233 ( .A(mem[915]), .Y(n7001) );
  INVX1 U6234 ( .A(mem[849]), .Y(n7067) );
  INVX1 U6235 ( .A(mem[816]), .Y(n7100) );
  INVX1 U6236 ( .A(mem[123]), .Y(n7793) );
  INVX1 U6237 ( .A(mem[57]), .Y(n7859) );
  INVX1 U6238 ( .A(mem[24]), .Y(n7892) );
  INVX1 U6239 ( .A(mem[652]), .Y(n7264) );
  INVX1 U6240 ( .A(mem[586]), .Y(n7330) );
  INVX1 U6241 ( .A(mem[553]), .Y(n7363) );
  INVX1 U6242 ( .A(mem[916]), .Y(n7000) );
  INVX1 U6243 ( .A(mem[850]), .Y(n7066) );
  INVX1 U6244 ( .A(mem[817]), .Y(n7099) );
  INVX1 U6245 ( .A(mem[124]), .Y(n7792) );
  INVX1 U6246 ( .A(mem[58]), .Y(n7858) );
  INVX1 U6247 ( .A(mem[25]), .Y(n7891) );
  INVX1 U6248 ( .A(mem[653]), .Y(n7263) );
  INVX1 U6249 ( .A(mem[587]), .Y(n7329) );
  INVX1 U6250 ( .A(mem[554]), .Y(n7362) );
  INVX1 U6251 ( .A(mem[917]), .Y(n6999) );
  INVX1 U6252 ( .A(mem[851]), .Y(n7065) );
  INVX1 U6253 ( .A(mem[818]), .Y(n7098) );
  INVX1 U6254 ( .A(mem[125]), .Y(n7791) );
  INVX1 U6255 ( .A(mem[59]), .Y(n7857) );
  INVX1 U6256 ( .A(mem[26]), .Y(n7890) );
  INVX1 U6257 ( .A(mem[654]), .Y(n7262) );
  INVX1 U6258 ( .A(mem[588]), .Y(n7328) );
  INVX1 U6259 ( .A(mem[555]), .Y(n7361) );
  INVX1 U6260 ( .A(mem[918]), .Y(n6998) );
  INVX1 U6261 ( .A(mem[852]), .Y(n7064) );
  INVX1 U6262 ( .A(mem[819]), .Y(n7097) );
  INVX1 U6263 ( .A(mem[126]), .Y(n7790) );
  INVX1 U6264 ( .A(mem[60]), .Y(n7856) );
  INVX1 U6265 ( .A(mem[27]), .Y(n7889) );
  INVX1 U6266 ( .A(mem[655]), .Y(n7261) );
  INVX1 U6267 ( .A(mem[589]), .Y(n7327) );
  INVX1 U6268 ( .A(mem[556]), .Y(n7360) );
  INVX1 U6269 ( .A(mem[919]), .Y(n6997) );
  INVX1 U6270 ( .A(mem[853]), .Y(n7063) );
  INVX1 U6271 ( .A(mem[820]), .Y(n7096) );
  INVX1 U6272 ( .A(mem[127]), .Y(n7789) );
  INVX1 U6273 ( .A(mem[61]), .Y(n7855) );
  INVX1 U6274 ( .A(mem[28]), .Y(n7888) );
  INVX1 U6275 ( .A(mem[656]), .Y(n7260) );
  INVX1 U6276 ( .A(mem[590]), .Y(n7326) );
  INVX1 U6277 ( .A(mem[557]), .Y(n7359) );
  INVX1 U6278 ( .A(mem[920]), .Y(n6996) );
  INVX1 U6279 ( .A(mem[854]), .Y(n7062) );
  INVX1 U6280 ( .A(mem[821]), .Y(n7095) );
  INVX1 U6281 ( .A(mem[128]), .Y(n7788) );
  INVX1 U6282 ( .A(mem[62]), .Y(n7854) );
  INVX1 U6283 ( .A(mem[29]), .Y(n7887) );
  INVX1 U6284 ( .A(mem[657]), .Y(n7259) );
  INVX1 U6285 ( .A(mem[591]), .Y(n7325) );
  INVX1 U6286 ( .A(mem[558]), .Y(n7358) );
  INVX1 U6287 ( .A(mem[921]), .Y(n6995) );
  INVX1 U6288 ( .A(mem[855]), .Y(n7061) );
  INVX1 U6289 ( .A(mem[822]), .Y(n7094) );
  INVX1 U6290 ( .A(mem[129]), .Y(n7787) );
  INVX1 U6291 ( .A(mem[63]), .Y(n7853) );
  INVX1 U6292 ( .A(mem[30]), .Y(n7886) );
  INVX1 U6293 ( .A(mem[658]), .Y(n7258) );
  INVX1 U6294 ( .A(mem[592]), .Y(n7324) );
  INVX1 U6295 ( .A(mem[559]), .Y(n7357) );
  INVX1 U6296 ( .A(mem[922]), .Y(n6994) );
  INVX1 U6297 ( .A(mem[856]), .Y(n7060) );
  INVX1 U6298 ( .A(mem[823]), .Y(n7093) );
  INVX1 U6299 ( .A(mem[130]), .Y(n7786) );
  INVX1 U6300 ( .A(mem[64]), .Y(n7852) );
  INVX1 U6301 ( .A(mem[31]), .Y(n7885) );
  INVX1 U6302 ( .A(mem[659]), .Y(n7257) );
  INVX1 U6303 ( .A(mem[593]), .Y(n7323) );
  INVX1 U6304 ( .A(mem[560]), .Y(n7356) );
  INVX1 U6305 ( .A(mem[923]), .Y(n6993) );
  INVX1 U6306 ( .A(mem[857]), .Y(n7059) );
  INVX1 U6307 ( .A(mem[824]), .Y(n7092) );
  INVX1 U6308 ( .A(mem[131]), .Y(n7785) );
  INVX1 U6309 ( .A(mem[65]), .Y(n7851) );
  INVX1 U6310 ( .A(mem[32]), .Y(n7884) );
  INVX1 U6311 ( .A(mem[363]), .Y(n7553) );
  INVX1 U6312 ( .A(mem[297]), .Y(n7619) );
  INVX1 U6313 ( .A(mem[264]), .Y(n7652) );
  INVX1 U6314 ( .A(mem[364]), .Y(n7552) );
  INVX1 U6315 ( .A(mem[298]), .Y(n7618) );
  INVX1 U6316 ( .A(mem[265]), .Y(n7651) );
  INVX1 U6317 ( .A(mem[365]), .Y(n7551) );
  INVX1 U6318 ( .A(mem[299]), .Y(n7617) );
  INVX1 U6319 ( .A(mem[266]), .Y(n7650) );
  INVX1 U6320 ( .A(mem[366]), .Y(n7550) );
  INVX1 U6321 ( .A(mem[300]), .Y(n7616) );
  INVX1 U6322 ( .A(mem[267]), .Y(n7649) );
  INVX1 U6323 ( .A(mem[367]), .Y(n7549) );
  INVX1 U6324 ( .A(mem[301]), .Y(n7615) );
  INVX1 U6325 ( .A(mem[268]), .Y(n7648) );
  INVX1 U6326 ( .A(mem[368]), .Y(n7548) );
  INVX1 U6327 ( .A(mem[302]), .Y(n7614) );
  INVX1 U6328 ( .A(mem[269]), .Y(n7647) );
  INVX1 U6329 ( .A(mem[369]), .Y(n7547) );
  INVX1 U6330 ( .A(mem[303]), .Y(n7613) );
  INVX1 U6331 ( .A(mem[270]), .Y(n7646) );
  INVX1 U6332 ( .A(mem[370]), .Y(n7546) );
  INVX1 U6333 ( .A(mem[304]), .Y(n7612) );
  INVX1 U6334 ( .A(mem[271]), .Y(n7645) );
  INVX1 U6335 ( .A(mem[371]), .Y(n7545) );
  INVX1 U6336 ( .A(mem[305]), .Y(n7611) );
  INVX1 U6337 ( .A(mem[272]), .Y(n7644) );
  INVX1 U6338 ( .A(mem[372]), .Y(n7544) );
  INVX1 U6339 ( .A(mem[306]), .Y(n7610) );
  INVX1 U6340 ( .A(mem[273]), .Y(n7643) );
  INVX1 U6341 ( .A(mem[373]), .Y(n7543) );
  INVX1 U6342 ( .A(mem[307]), .Y(n7609) );
  INVX1 U6343 ( .A(mem[274]), .Y(n7642) );
  INVX1 U6344 ( .A(mem[374]), .Y(n7542) );
  INVX1 U6345 ( .A(mem[308]), .Y(n7608) );
  INVX1 U6346 ( .A(mem[275]), .Y(n7641) );
  INVX1 U6347 ( .A(mem[375]), .Y(n7541) );
  INVX1 U6348 ( .A(mem[309]), .Y(n7607) );
  INVX1 U6349 ( .A(mem[276]), .Y(n7640) );
  INVX1 U6350 ( .A(mem[376]), .Y(n7540) );
  INVX1 U6351 ( .A(mem[310]), .Y(n7606) );
  INVX1 U6352 ( .A(mem[277]), .Y(n7639) );
  INVX1 U6353 ( .A(mem[377]), .Y(n7539) );
  INVX1 U6354 ( .A(mem[311]), .Y(n7605) );
  INVX1 U6355 ( .A(mem[278]), .Y(n7638) );
  INVX1 U6356 ( .A(mem[378]), .Y(n7538) );
  INVX1 U6357 ( .A(mem[312]), .Y(n7604) );
  INVX1 U6358 ( .A(mem[279]), .Y(n7637) );
  INVX1 U6359 ( .A(mem[379]), .Y(n7537) );
  INVX1 U6360 ( .A(mem[313]), .Y(n7603) );
  INVX1 U6361 ( .A(mem[280]), .Y(n7636) );
  INVX1 U6362 ( .A(mem[380]), .Y(n7536) );
  INVX1 U6363 ( .A(mem[314]), .Y(n7602) );
  INVX1 U6364 ( .A(mem[281]), .Y(n7635) );
  INVX1 U6365 ( .A(mem[381]), .Y(n7535) );
  INVX1 U6366 ( .A(mem[315]), .Y(n7601) );
  INVX1 U6367 ( .A(mem[282]), .Y(n7634) );
  INVX1 U6368 ( .A(mem[382]), .Y(n7534) );
  INVX1 U6369 ( .A(mem[316]), .Y(n7600) );
  INVX1 U6370 ( .A(mem[283]), .Y(n7633) );
  INVX1 U6371 ( .A(mem[383]), .Y(n7533) );
  INVX1 U6372 ( .A(mem[317]), .Y(n7599) );
  INVX1 U6373 ( .A(mem[284]), .Y(n7632) );
  INVX1 U6374 ( .A(mem[384]), .Y(n7532) );
  INVX1 U6375 ( .A(mem[318]), .Y(n7598) );
  INVX1 U6376 ( .A(mem[285]), .Y(n7631) );
  INVX1 U6377 ( .A(mem[385]), .Y(n7531) );
  INVX1 U6378 ( .A(mem[319]), .Y(n7597) );
  INVX1 U6379 ( .A(mem[286]), .Y(n7630) );
  INVX1 U6380 ( .A(mem[386]), .Y(n7530) );
  INVX1 U6381 ( .A(mem[320]), .Y(n7596) );
  INVX1 U6382 ( .A(mem[287]), .Y(n7629) );
  INVX1 U6383 ( .A(mem[387]), .Y(n7529) );
  INVX1 U6384 ( .A(mem[321]), .Y(n7595) );
  INVX1 U6385 ( .A(mem[288]), .Y(n7628) );
  INVX1 U6386 ( .A(mem[388]), .Y(n7528) );
  INVX1 U6387 ( .A(mem[322]), .Y(n7594) );
  INVX1 U6388 ( .A(mem[289]), .Y(n7627) );
  INVX1 U6389 ( .A(mem[389]), .Y(n7527) );
  INVX1 U6390 ( .A(mem[323]), .Y(n7593) );
  INVX1 U6391 ( .A(mem[290]), .Y(n7626) );
  INVX1 U6392 ( .A(mem[390]), .Y(n7526) );
  INVX1 U6393 ( .A(mem[324]), .Y(n7592) );
  INVX1 U6394 ( .A(mem[291]), .Y(n7625) );
  INVX1 U6395 ( .A(mem[391]), .Y(n7525) );
  INVX1 U6396 ( .A(mem[325]), .Y(n7591) );
  INVX1 U6397 ( .A(mem[292]), .Y(n7624) );
  INVX1 U6398 ( .A(mem[392]), .Y(n7524) );
  INVX1 U6399 ( .A(mem[326]), .Y(n7590) );
  INVX1 U6400 ( .A(mem[293]), .Y(n7623) );
  INVX1 U6401 ( .A(mem[393]), .Y(n7523) );
  INVX1 U6402 ( .A(mem[327]), .Y(n7589) );
  INVX1 U6403 ( .A(mem[294]), .Y(n7622) );
  INVX1 U6404 ( .A(mem[394]), .Y(n7522) );
  INVX1 U6405 ( .A(mem[328]), .Y(n7588) );
  INVX1 U6406 ( .A(mem[295]), .Y(n7621) );
  INVX1 U6407 ( .A(mem[395]), .Y(n7521) );
  INVX1 U6408 ( .A(mem[329]), .Y(n7587) );
  INVX1 U6409 ( .A(mem[296]), .Y(n7620) );
  INVX1 U6410 ( .A(mem[759]), .Y(n7157) );
  INVX1 U6411 ( .A(mem[660]), .Y(n7256) );
  INVX1 U6412 ( .A(mem[1023]), .Y(n6893) );
  INVX1 U6413 ( .A(mem[924]), .Y(n6992) );
  INVX1 U6414 ( .A(mem[231]), .Y(n7685) );
  INVX1 U6415 ( .A(mem[132]), .Y(n7784) );
  INVX1 U6416 ( .A(mem[760]), .Y(n7156) );
  INVX1 U6417 ( .A(mem[661]), .Y(n7255) );
  INVX1 U6418 ( .A(mem[1024]), .Y(n6892) );
  INVX1 U6419 ( .A(mem[925]), .Y(n6991) );
  INVX1 U6420 ( .A(mem[232]), .Y(n7684) );
  INVX1 U6421 ( .A(mem[133]), .Y(n7783) );
  INVX1 U6422 ( .A(mem[761]), .Y(n7155) );
  INVX1 U6423 ( .A(mem[662]), .Y(n7254) );
  INVX1 U6424 ( .A(mem[1025]), .Y(n6891) );
  INVX1 U6425 ( .A(mem[926]), .Y(n6990) );
  INVX1 U6426 ( .A(mem[233]), .Y(n7683) );
  INVX1 U6427 ( .A(mem[134]), .Y(n7782) );
  INVX1 U6428 ( .A(mem[762]), .Y(n7154) );
  INVX1 U6429 ( .A(mem[663]), .Y(n7253) );
  INVX1 U6430 ( .A(mem[1026]), .Y(n6890) );
  INVX1 U6431 ( .A(mem[927]), .Y(n6989) );
  INVX1 U6432 ( .A(mem[234]), .Y(n7682) );
  INVX1 U6433 ( .A(mem[135]), .Y(n7781) );
  INVX1 U6434 ( .A(mem[763]), .Y(n7153) );
  INVX1 U6435 ( .A(mem[664]), .Y(n7252) );
  INVX1 U6436 ( .A(mem[1027]), .Y(n6889) );
  INVX1 U6437 ( .A(mem[928]), .Y(n6988) );
  INVX1 U6438 ( .A(mem[235]), .Y(n7681) );
  INVX1 U6439 ( .A(mem[136]), .Y(n7780) );
  INVX1 U6440 ( .A(mem[764]), .Y(n7152) );
  INVX1 U6441 ( .A(mem[665]), .Y(n7251) );
  INVX1 U6442 ( .A(mem[1028]), .Y(n6888) );
  INVX1 U6443 ( .A(mem[929]), .Y(n6987) );
  INVX1 U6444 ( .A(mem[236]), .Y(n7680) );
  INVX1 U6445 ( .A(mem[137]), .Y(n7779) );
  INVX1 U6446 ( .A(mem[765]), .Y(n7151) );
  INVX1 U6447 ( .A(mem[666]), .Y(n7250) );
  INVX1 U6448 ( .A(mem[1029]), .Y(n6887) );
  INVX1 U6449 ( .A(mem[930]), .Y(n6986) );
  INVX1 U6450 ( .A(mem[237]), .Y(n7679) );
  INVX1 U6451 ( .A(mem[138]), .Y(n7778) );
  INVX1 U6452 ( .A(mem[766]), .Y(n7150) );
  INVX1 U6453 ( .A(mem[667]), .Y(n7249) );
  INVX1 U6454 ( .A(mem[1030]), .Y(n6886) );
  INVX1 U6455 ( .A(mem[931]), .Y(n6985) );
  INVX1 U6456 ( .A(mem[238]), .Y(n7678) );
  INVX1 U6457 ( .A(mem[139]), .Y(n7777) );
  INVX1 U6458 ( .A(mem[767]), .Y(n7149) );
  INVX1 U6459 ( .A(mem[668]), .Y(n7248) );
  INVX1 U6460 ( .A(mem[1031]), .Y(n6885) );
  INVX1 U6461 ( .A(mem[932]), .Y(n6984) );
  INVX1 U6462 ( .A(mem[239]), .Y(n7677) );
  INVX1 U6463 ( .A(mem[140]), .Y(n7776) );
  INVX1 U6464 ( .A(mem[768]), .Y(n7148) );
  INVX1 U6465 ( .A(mem[669]), .Y(n7247) );
  INVX1 U6466 ( .A(mem[1032]), .Y(n6884) );
  INVX1 U6467 ( .A(mem[933]), .Y(n6983) );
  INVX1 U6468 ( .A(mem[240]), .Y(n7676) );
  INVX1 U6469 ( .A(mem[141]), .Y(n7775) );
  INVX1 U6470 ( .A(mem[769]), .Y(n7147) );
  INVX1 U6471 ( .A(mem[670]), .Y(n7246) );
  INVX1 U6472 ( .A(mem[1033]), .Y(n6883) );
  INVX1 U6473 ( .A(mem[934]), .Y(n6982) );
  INVX1 U6474 ( .A(mem[241]), .Y(n7675) );
  INVX1 U6475 ( .A(mem[142]), .Y(n7774) );
  INVX1 U6476 ( .A(mem[770]), .Y(n7146) );
  INVX1 U6477 ( .A(mem[671]), .Y(n7245) );
  INVX1 U6478 ( .A(mem[1034]), .Y(n6882) );
  INVX1 U6479 ( .A(mem[935]), .Y(n6981) );
  INVX1 U6480 ( .A(mem[242]), .Y(n7674) );
  INVX1 U6481 ( .A(mem[143]), .Y(n7773) );
  INVX1 U6482 ( .A(mem[771]), .Y(n7145) );
  INVX1 U6483 ( .A(mem[672]), .Y(n7244) );
  INVX1 U6484 ( .A(mem[1035]), .Y(n6881) );
  INVX1 U6485 ( .A(mem[936]), .Y(n6980) );
  INVX1 U6486 ( .A(mem[243]), .Y(n7673) );
  INVX1 U6487 ( .A(mem[144]), .Y(n7772) );
  INVX1 U6488 ( .A(mem[772]), .Y(n7144) );
  INVX1 U6489 ( .A(mem[673]), .Y(n7243) );
  INVX1 U6490 ( .A(mem[1036]), .Y(n6880) );
  INVX1 U6491 ( .A(mem[937]), .Y(n6979) );
  INVX1 U6492 ( .A(mem[244]), .Y(n7672) );
  INVX1 U6493 ( .A(mem[145]), .Y(n7771) );
  INVX1 U6494 ( .A(mem[773]), .Y(n7143) );
  INVX1 U6495 ( .A(mem[674]), .Y(n7242) );
  INVX1 U6496 ( .A(mem[1037]), .Y(n6879) );
  INVX1 U6497 ( .A(mem[938]), .Y(n6978) );
  INVX1 U6498 ( .A(mem[245]), .Y(n7671) );
  INVX1 U6499 ( .A(mem[146]), .Y(n7770) );
  INVX1 U6500 ( .A(mem[774]), .Y(n7142) );
  INVX1 U6501 ( .A(mem[675]), .Y(n7241) );
  INVX1 U6502 ( .A(mem[1038]), .Y(n6878) );
  INVX1 U6503 ( .A(mem[939]), .Y(n6977) );
  INVX1 U6504 ( .A(mem[246]), .Y(n7670) );
  INVX1 U6505 ( .A(mem[147]), .Y(n7769) );
  INVX1 U6506 ( .A(mem[775]), .Y(n7141) );
  INVX1 U6507 ( .A(mem[676]), .Y(n7240) );
  INVX1 U6508 ( .A(mem[1039]), .Y(n6877) );
  INVX1 U6509 ( .A(mem[940]), .Y(n6976) );
  INVX1 U6510 ( .A(mem[247]), .Y(n7669) );
  INVX1 U6511 ( .A(mem[148]), .Y(n7768) );
  INVX1 U6512 ( .A(mem[776]), .Y(n7140) );
  INVX1 U6513 ( .A(mem[677]), .Y(n7239) );
  INVX1 U6514 ( .A(mem[1040]), .Y(n6876) );
  INVX1 U6515 ( .A(mem[941]), .Y(n6975) );
  INVX1 U6516 ( .A(mem[248]), .Y(n7668) );
  INVX1 U6517 ( .A(mem[149]), .Y(n7767) );
  INVX1 U6518 ( .A(mem[777]), .Y(n7139) );
  INVX1 U6519 ( .A(mem[678]), .Y(n7238) );
  INVX1 U6520 ( .A(mem[1041]), .Y(n6875) );
  INVX1 U6521 ( .A(mem[942]), .Y(n6974) );
  INVX1 U6522 ( .A(mem[249]), .Y(n7667) );
  INVX1 U6523 ( .A(mem[150]), .Y(n7766) );
  INVX1 U6524 ( .A(mem[778]), .Y(n7138) );
  INVX1 U6525 ( .A(mem[679]), .Y(n7237) );
  INVX1 U6526 ( .A(mem[1042]), .Y(n6874) );
  INVX1 U6527 ( .A(mem[943]), .Y(n6973) );
  INVX1 U6528 ( .A(mem[250]), .Y(n7666) );
  INVX1 U6529 ( .A(mem[151]), .Y(n7765) );
  INVX1 U6530 ( .A(mem[779]), .Y(n7137) );
  INVX1 U6531 ( .A(mem[680]), .Y(n7236) );
  INVX1 U6532 ( .A(mem[1043]), .Y(n6873) );
  INVX1 U6533 ( .A(mem[944]), .Y(n6972) );
  INVX1 U6534 ( .A(mem[251]), .Y(n7665) );
  INVX1 U6535 ( .A(mem[152]), .Y(n7764) );
  INVX1 U6536 ( .A(mem[780]), .Y(n7136) );
  INVX1 U6537 ( .A(mem[681]), .Y(n7235) );
  INVX1 U6538 ( .A(mem[1044]), .Y(n6872) );
  INVX1 U6539 ( .A(mem[945]), .Y(n6971) );
  INVX1 U6540 ( .A(mem[252]), .Y(n7664) );
  INVX1 U6541 ( .A(mem[153]), .Y(n7763) );
  INVX1 U6542 ( .A(mem[781]), .Y(n7135) );
  INVX1 U6543 ( .A(mem[682]), .Y(n7234) );
  INVX1 U6544 ( .A(mem[1045]), .Y(n6871) );
  INVX1 U6545 ( .A(mem[946]), .Y(n6970) );
  INVX1 U6546 ( .A(mem[253]), .Y(n7663) );
  INVX1 U6547 ( .A(mem[154]), .Y(n7762) );
  INVX1 U6548 ( .A(mem[782]), .Y(n7134) );
  INVX1 U6549 ( .A(mem[683]), .Y(n7233) );
  INVX1 U6550 ( .A(mem[1046]), .Y(n6870) );
  INVX1 U6551 ( .A(mem[947]), .Y(n6969) );
  INVX1 U6552 ( .A(mem[254]), .Y(n7662) );
  INVX1 U6553 ( .A(mem[155]), .Y(n7761) );
  INVX1 U6554 ( .A(mem[783]), .Y(n7133) );
  INVX1 U6555 ( .A(mem[684]), .Y(n7232) );
  INVX1 U6556 ( .A(mem[1047]), .Y(n6869) );
  INVX1 U6557 ( .A(mem[948]), .Y(n6968) );
  INVX1 U6558 ( .A(mem[255]), .Y(n7661) );
  INVX1 U6559 ( .A(mem[156]), .Y(n7760) );
  INVX1 U6560 ( .A(mem[784]), .Y(n7132) );
  INVX1 U6561 ( .A(mem[685]), .Y(n7231) );
  INVX1 U6562 ( .A(mem[1048]), .Y(n6868) );
  INVX1 U6563 ( .A(mem[949]), .Y(n6967) );
  INVX1 U6564 ( .A(mem[256]), .Y(n7660) );
  INVX1 U6565 ( .A(mem[157]), .Y(n7759) );
  INVX1 U6566 ( .A(mem[785]), .Y(n7131) );
  INVX1 U6567 ( .A(mem[686]), .Y(n7230) );
  INVX1 U6568 ( .A(mem[1049]), .Y(n6867) );
  INVX1 U6569 ( .A(mem[950]), .Y(n6966) );
  INVX1 U6570 ( .A(mem[257]), .Y(n7659) );
  INVX1 U6571 ( .A(mem[158]), .Y(n7758) );
  INVX1 U6572 ( .A(mem[786]), .Y(n7130) );
  INVX1 U6573 ( .A(mem[687]), .Y(n7229) );
  INVX1 U6574 ( .A(mem[1050]), .Y(n6866) );
  INVX1 U6575 ( .A(mem[951]), .Y(n6965) );
  INVX1 U6576 ( .A(mem[258]), .Y(n7658) );
  INVX1 U6577 ( .A(mem[159]), .Y(n7757) );
  INVX1 U6578 ( .A(mem[787]), .Y(n7129) );
  INVX1 U6579 ( .A(mem[688]), .Y(n7228) );
  INVX1 U6580 ( .A(mem[1051]), .Y(n6865) );
  INVX1 U6581 ( .A(mem[952]), .Y(n6964) );
  INVX1 U6582 ( .A(mem[259]), .Y(n7657) );
  INVX1 U6583 ( .A(mem[160]), .Y(n7756) );
  INVX1 U6584 ( .A(mem[788]), .Y(n7128) );
  INVX1 U6585 ( .A(mem[689]), .Y(n7227) );
  INVX1 U6586 ( .A(mem[1052]), .Y(n6864) );
  INVX1 U6587 ( .A(mem[953]), .Y(n6963) );
  INVX1 U6588 ( .A(mem[260]), .Y(n7656) );
  INVX1 U6589 ( .A(mem[161]), .Y(n7755) );
  INVX1 U6590 ( .A(mem[789]), .Y(n7127) );
  INVX1 U6591 ( .A(mem[690]), .Y(n7226) );
  INVX1 U6592 ( .A(mem[1053]), .Y(n6863) );
  INVX1 U6593 ( .A(mem[954]), .Y(n6962) );
  INVX1 U6594 ( .A(mem[261]), .Y(n7655) );
  INVX1 U6595 ( .A(mem[162]), .Y(n7754) );
  INVX1 U6596 ( .A(mem[790]), .Y(n7126) );
  INVX1 U6597 ( .A(mem[691]), .Y(n7225) );
  INVX1 U6598 ( .A(mem[1054]), .Y(n6862) );
  INVX1 U6599 ( .A(mem[955]), .Y(n6961) );
  INVX1 U6600 ( .A(mem[262]), .Y(n7654) );
  INVX1 U6601 ( .A(mem[163]), .Y(n7753) );
  INVX1 U6602 ( .A(mem[791]), .Y(n7125) );
  INVX1 U6603 ( .A(mem[692]), .Y(n7224) );
  INVX1 U6604 ( .A(mem[1055]), .Y(n6861) );
  INVX1 U6605 ( .A(mem[956]), .Y(n6960) );
  INVX1 U6606 ( .A(mem[263]), .Y(n7653) );
  INVX1 U6607 ( .A(mem[164]), .Y(n7752) );
  INVX1 U6608 ( .A(mem[495]), .Y(n7421) );
  INVX1 U6609 ( .A(mem[396]), .Y(n7520) );
  INVX1 U6610 ( .A(mem[496]), .Y(n7420) );
  INVX1 U6611 ( .A(mem[397]), .Y(n7519) );
  INVX1 U6612 ( .A(mem[497]), .Y(n7419) );
  INVX1 U6613 ( .A(mem[398]), .Y(n7518) );
  INVX1 U6614 ( .A(mem[498]), .Y(n7418) );
  INVX1 U6615 ( .A(mem[399]), .Y(n7517) );
  INVX1 U6616 ( .A(mem[499]), .Y(n7417) );
  INVX1 U6617 ( .A(mem[400]), .Y(n7516) );
  INVX1 U6618 ( .A(mem[500]), .Y(n7416) );
  INVX1 U6619 ( .A(mem[401]), .Y(n7515) );
  INVX1 U6620 ( .A(mem[501]), .Y(n7415) );
  INVX1 U6621 ( .A(mem[402]), .Y(n7514) );
  INVX1 U6622 ( .A(mem[502]), .Y(n7414) );
  INVX1 U6623 ( .A(mem[403]), .Y(n7513) );
  INVX1 U6624 ( .A(mem[503]), .Y(n7413) );
  INVX1 U6625 ( .A(mem[404]), .Y(n7512) );
  INVX1 U6626 ( .A(mem[504]), .Y(n7412) );
  INVX1 U6627 ( .A(mem[405]), .Y(n7511) );
  INVX1 U6628 ( .A(mem[505]), .Y(n7411) );
  INVX1 U6629 ( .A(mem[406]), .Y(n7510) );
  INVX1 U6630 ( .A(mem[506]), .Y(n7410) );
  INVX1 U6631 ( .A(mem[407]), .Y(n7509) );
  INVX1 U6632 ( .A(mem[507]), .Y(n7409) );
  INVX1 U6633 ( .A(mem[408]), .Y(n7508) );
  INVX1 U6634 ( .A(mem[508]), .Y(n7408) );
  INVX1 U6635 ( .A(mem[409]), .Y(n7507) );
  INVX1 U6636 ( .A(mem[509]), .Y(n7407) );
  INVX1 U6637 ( .A(mem[410]), .Y(n7506) );
  INVX1 U6638 ( .A(mem[510]), .Y(n7406) );
  INVX1 U6639 ( .A(mem[411]), .Y(n7505) );
  INVX1 U6640 ( .A(mem[511]), .Y(n7405) );
  INVX1 U6641 ( .A(mem[412]), .Y(n7504) );
  INVX1 U6642 ( .A(mem[512]), .Y(n7404) );
  INVX1 U6643 ( .A(mem[413]), .Y(n7503) );
  INVX1 U6644 ( .A(mem[513]), .Y(n7403) );
  INVX1 U6645 ( .A(mem[414]), .Y(n7502) );
  INVX1 U6646 ( .A(mem[514]), .Y(n7402) );
  INVX1 U6647 ( .A(mem[415]), .Y(n7501) );
  INVX1 U6648 ( .A(mem[515]), .Y(n7401) );
  INVX1 U6649 ( .A(mem[416]), .Y(n7500) );
  INVX1 U6650 ( .A(mem[516]), .Y(n7400) );
  INVX1 U6651 ( .A(mem[417]), .Y(n7499) );
  INVX1 U6652 ( .A(mem[517]), .Y(n7399) );
  INVX1 U6653 ( .A(mem[418]), .Y(n7498) );
  INVX1 U6654 ( .A(mem[518]), .Y(n7398) );
  INVX1 U6655 ( .A(mem[419]), .Y(n7497) );
  INVX1 U6656 ( .A(mem[519]), .Y(n7397) );
  INVX1 U6657 ( .A(mem[420]), .Y(n7496) );
  INVX1 U6658 ( .A(mem[520]), .Y(n7396) );
  INVX1 U6659 ( .A(mem[421]), .Y(n7495) );
  INVX1 U6660 ( .A(mem[521]), .Y(n7395) );
  INVX1 U6661 ( .A(mem[422]), .Y(n7494) );
  INVX1 U6662 ( .A(mem[522]), .Y(n7394) );
  INVX1 U6663 ( .A(mem[423]), .Y(n7493) );
  INVX1 U6664 ( .A(mem[523]), .Y(n7393) );
  INVX1 U6665 ( .A(mem[424]), .Y(n7492) );
  INVX1 U6666 ( .A(mem[524]), .Y(n7392) );
  INVX1 U6667 ( .A(mem[425]), .Y(n7491) );
  INVX1 U6668 ( .A(mem[525]), .Y(n7391) );
  INVX1 U6669 ( .A(mem[426]), .Y(n7490) );
  INVX1 U6670 ( .A(mem[526]), .Y(n7390) );
  INVX1 U6671 ( .A(mem[427]), .Y(n7489) );
  INVX1 U6672 ( .A(mem[527]), .Y(n7389) );
  INVX1 U6673 ( .A(mem[428]), .Y(n7488) );
  INVX1 U6674 ( .A(n4454), .Y(n6847) );
  INVX1 U6675 ( .A(n3292), .Y(n6846) );
  AND2X1 U6676 ( .A(data_in[2]), .B(n6843), .Y(n3385) );
  AND2X1 U6677 ( .A(data_in[3]), .B(n6843), .Y(n3383) );
  AND2X1 U6678 ( .A(data_in[4]), .B(n6843), .Y(n3381) );
  AND2X1 U6679 ( .A(data_in[5]), .B(n6843), .Y(n3379) );
  AND2X1 U6680 ( .A(data_in[6]), .B(n6843), .Y(n3377) );
  AND2X1 U6681 ( .A(data_in[7]), .B(n6843), .Y(n3375) );
  AND2X1 U6682 ( .A(data_in[8]), .B(n6843), .Y(n3373) );
  AND2X1 U6683 ( .A(data_in[9]), .B(n6843), .Y(n3371) );
  AND2X1 U6684 ( .A(data_in[10]), .B(n6843), .Y(n3369) );
  AND2X1 U6685 ( .A(data_in[11]), .B(n6843), .Y(n3367) );
  AND2X1 U6686 ( .A(data_in[12]), .B(n6843), .Y(n3365) );
  AND2X1 U6687 ( .A(data_in[13]), .B(n6843), .Y(n3363) );
  AND2X1 U6688 ( .A(data_in[14]), .B(n6843), .Y(n3361) );
  AND2X1 U6689 ( .A(data_in[15]), .B(n6843), .Y(n3359) );
  AND2X1 U6690 ( .A(data_in[16]), .B(n6843), .Y(n3357) );
  AND2X1 U6691 ( .A(data_in[17]), .B(n6843), .Y(n3355) );
  AND2X1 U6692 ( .A(data_in[18]), .B(n6843), .Y(n3353) );
  AND2X1 U6693 ( .A(data_in[19]), .B(n6843), .Y(n3351) );
  AND2X1 U6694 ( .A(data_in[20]), .B(n6843), .Y(n3349) );
  AND2X1 U6695 ( .A(data_in[21]), .B(n6843), .Y(n3347) );
  AND2X1 U6696 ( .A(data_in[22]), .B(n6843), .Y(n3345) );
  AND2X1 U6697 ( .A(data_in[23]), .B(n6843), .Y(n3343) );
  AND2X1 U6698 ( .A(data_in[24]), .B(n6843), .Y(n3341) );
  AND2X1 U6699 ( .A(data_in[25]), .B(n6843), .Y(n3339) );
  AND2X1 U6700 ( .A(data_in[26]), .B(n6843), .Y(n3337) );
  AND2X1 U6701 ( .A(data_in[27]), .B(n6843), .Y(n3335) );
  AND2X1 U6702 ( .A(data_in[28]), .B(n6843), .Y(n3333) );
  AND2X1 U6703 ( .A(data_in[29]), .B(n6843), .Y(n3331) );
  AND2X1 U6704 ( .A(data_in[30]), .B(n6843), .Y(n3329) );
  AND2X1 U6705 ( .A(data_in[31]), .B(n6843), .Y(n3327) );
  AND2X1 U6706 ( .A(data_in[32]), .B(n6843), .Y(n3325) );
  AND2X1 U6707 ( .A(data_in[0]), .B(n6843), .Y(n3389) );
  AND2X1 U6708 ( .A(data_in[1]), .B(n6843), .Y(n3387) );
endmodule


module FIFO_DEPTH_P25_WIDTH41 ( clk, reset, data_in, put, get, data_out, 
        empty_bar, full_bar, fillcount );
  input [40:0] data_in;
  output [40:0] data_out;
  output [5:0] fillcount;
  input clk, reset, put, get;
  output empty_bar, full_bar;
  wire   n12, n13, n14, n15, n16, n5721, n1842, n1843, n1844, n1845, n1846,
         n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
         n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
         n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
         n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
         n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
         n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
         n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
         n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
         n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
         n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
         n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
         n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
         n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
         n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
         n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
         n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
         n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
         n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
         n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
         n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
         n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
         n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
         n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
         n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
         n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
         n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
         n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
         n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
         n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
         n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
         n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
         n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
         n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
         n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
         n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
         n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
         n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
         n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
         n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056,
         n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
         n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076,
         n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
         n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096,
         n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
         n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
         n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831;
  wire   [4:0] wr_ptr;
  wire   [1311:0] mem;
  assign full_bar = 1'b1;

  DFFPOSX1 wr_ptr_reg_0_ ( .D(n3163), .CLK(clk), .Q(wr_ptr[0]) );
  DFFPOSX1 rd_ptr_reg_4_ ( .D(n5723), .CLK(clk), .Q(n16) );
  DFFPOSX1 rd_ptr_reg_0_ ( .D(n3161), .CLK(clk), .Q(n12) );
  DFFPOSX1 rd_ptr_reg_1_ ( .D(n3160), .CLK(clk), .Q(n13) );
  DFFPOSX1 rd_ptr_reg_2_ ( .D(n3159), .CLK(clk), .Q(n14) );
  DFFPOSX1 rd_ptr_reg_3_ ( .D(n3158), .CLK(clk), .Q(n15) );
  DFFPOSX1 wr_ptr_reg_4_ ( .D(n3157), .CLK(clk), .Q(wr_ptr[4]) );
  DFFPOSX1 wr_ptr_reg_1_ ( .D(n3156), .CLK(clk), .Q(wr_ptr[1]) );
  DFFPOSX1 wr_ptr_reg_2_ ( .D(n3155), .CLK(clk), .Q(wr_ptr[2]) );
  DFFPOSX1 wr_ptr_reg_3_ ( .D(n3154), .CLK(clk), .Q(wr_ptr[3]) );
  DFFPOSX1 data_out_reg_40_ ( .D(n5737), .CLK(clk), .Q(data_out[40]) );
  DFFPOSX1 data_out_reg_39_ ( .D(n5758), .CLK(clk), .Q(data_out[39]) );
  DFFPOSX1 data_out_reg_38_ ( .D(n5744), .CLK(clk), .Q(data_out[38]) );
  DFFPOSX1 data_out_reg_37_ ( .D(n5736), .CLK(clk), .Q(data_out[37]) );
  DFFPOSX1 data_out_reg_36_ ( .D(n5757), .CLK(clk), .Q(data_out[36]) );
  DFFPOSX1 data_out_reg_35_ ( .D(n5756), .CLK(clk), .Q(data_out[35]) );
  DFFPOSX1 data_out_reg_34_ ( .D(n5755), .CLK(clk), .Q(data_out[34]) );
  DFFPOSX1 data_out_reg_33_ ( .D(n5754), .CLK(clk), .Q(data_out[33]) );
  DFFPOSX1 data_out_reg_32_ ( .D(n5753), .CLK(clk), .Q(data_out[32]) );
  DFFPOSX1 data_out_reg_31_ ( .D(n5752), .CLK(clk), .Q(data_out[31]) );
  DFFPOSX1 data_out_reg_30_ ( .D(n5751), .CLK(clk), .Q(data_out[30]) );
  DFFPOSX1 data_out_reg_29_ ( .D(n5750), .CLK(clk), .Q(data_out[29]) );
  DFFPOSX1 data_out_reg_28_ ( .D(n5749), .CLK(clk), .Q(data_out[28]) );
  DFFPOSX1 data_out_reg_27_ ( .D(n5748), .CLK(clk), .Q(data_out[27]) );
  DFFPOSX1 data_out_reg_26_ ( .D(n5747), .CLK(clk), .Q(data_out[26]) );
  DFFPOSX1 data_out_reg_25_ ( .D(n5746), .CLK(clk), .Q(data_out[25]) );
  DFFPOSX1 data_out_reg_24_ ( .D(n5745), .CLK(clk), .Q(data_out[24]) );
  DFFPOSX1 data_out_reg_23_ ( .D(n5735), .CLK(clk), .Q(data_out[23]) );
  DFFPOSX1 data_out_reg_22_ ( .D(n5734), .CLK(clk), .Q(data_out[22]) );
  DFFPOSX1 data_out_reg_21_ ( .D(n5733), .CLK(clk), .Q(data_out[21]) );
  DFFPOSX1 data_out_reg_20_ ( .D(n5732), .CLK(clk), .Q(data_out[20]) );
  DFFPOSX1 data_out_reg_19_ ( .D(n5731), .CLK(clk), .Q(data_out[19]) );
  DFFPOSX1 data_out_reg_18_ ( .D(n5730), .CLK(clk), .Q(data_out[18]) );
  DFFPOSX1 data_out_reg_17_ ( .D(n5729), .CLK(clk), .Q(data_out[17]) );
  DFFPOSX1 data_out_reg_16_ ( .D(n5728), .CLK(clk), .Q(data_out[16]) );
  DFFPOSX1 data_out_reg_15_ ( .D(n5727), .CLK(clk), .Q(data_out[15]) );
  DFFPOSX1 data_out_reg_14_ ( .D(n5726), .CLK(clk), .Q(data_out[14]) );
  DFFPOSX1 data_out_reg_13_ ( .D(n5725), .CLK(clk), .Q(data_out[13]) );
  DFFPOSX1 data_out_reg_12_ ( .D(n5724), .CLK(clk), .Q(data_out[12]) );
  DFFPOSX1 data_out_reg_11_ ( .D(n5764), .CLK(clk), .Q(data_out[11]) );
  DFFPOSX1 data_out_reg_10_ ( .D(n5743), .CLK(clk), .Q(data_out[10]) );
  DFFPOSX1 data_out_reg_9_ ( .D(n5763), .CLK(clk), .Q(data_out[9]) );
  DFFPOSX1 data_out_reg_8_ ( .D(n5742), .CLK(clk), .Q(data_out[8]) );
  DFFPOSX1 data_out_reg_7_ ( .D(n5762), .CLK(clk), .Q(data_out[7]) );
  DFFPOSX1 data_out_reg_6_ ( .D(n5741), .CLK(clk), .Q(data_out[6]) );
  DFFPOSX1 data_out_reg_5_ ( .D(n5761), .CLK(clk), .Q(data_out[5]) );
  DFFPOSX1 data_out_reg_4_ ( .D(n5740), .CLK(clk), .Q(data_out[4]) );
  DFFPOSX1 data_out_reg_3_ ( .D(n5760), .CLK(clk), .Q(data_out[3]) );
  DFFPOSX1 data_out_reg_2_ ( .D(n5739), .CLK(clk), .Q(data_out[2]) );
  DFFPOSX1 data_out_reg_1_ ( .D(n5759), .CLK(clk), .Q(data_out[1]) );
  DFFPOSX1 data_out_reg_0_ ( .D(n5738), .CLK(clk), .Q(data_out[0]) );
  DFFPOSX1 mem_reg_31__40_ ( .D(n3153), .CLK(clk), .Q(mem[1311]) );
  DFFPOSX1 mem_reg_31__39_ ( .D(n3152), .CLK(clk), .Q(mem[1310]) );
  DFFPOSX1 mem_reg_31__38_ ( .D(n3151), .CLK(clk), .Q(mem[1309]) );
  DFFPOSX1 mem_reg_31__37_ ( .D(n3150), .CLK(clk), .Q(mem[1308]) );
  DFFPOSX1 mem_reg_31__36_ ( .D(n3149), .CLK(clk), .Q(mem[1307]) );
  DFFPOSX1 mem_reg_31__35_ ( .D(n3148), .CLK(clk), .Q(mem[1306]) );
  DFFPOSX1 mem_reg_31__34_ ( .D(n3147), .CLK(clk), .Q(mem[1305]) );
  DFFPOSX1 mem_reg_31__33_ ( .D(n3146), .CLK(clk), .Q(mem[1304]) );
  DFFPOSX1 mem_reg_31__32_ ( .D(n3145), .CLK(clk), .Q(mem[1303]) );
  DFFPOSX1 mem_reg_31__31_ ( .D(n3144), .CLK(clk), .Q(mem[1302]) );
  DFFPOSX1 mem_reg_31__30_ ( .D(n3143), .CLK(clk), .Q(mem[1301]) );
  DFFPOSX1 mem_reg_31__29_ ( .D(n3142), .CLK(clk), .Q(mem[1300]) );
  DFFPOSX1 mem_reg_31__28_ ( .D(n3141), .CLK(clk), .Q(mem[1299]) );
  DFFPOSX1 mem_reg_31__27_ ( .D(n3140), .CLK(clk), .Q(mem[1298]) );
  DFFPOSX1 mem_reg_31__26_ ( .D(n3139), .CLK(clk), .Q(mem[1297]) );
  DFFPOSX1 mem_reg_31__25_ ( .D(n3138), .CLK(clk), .Q(mem[1296]) );
  DFFPOSX1 mem_reg_31__24_ ( .D(n3137), .CLK(clk), .Q(mem[1295]) );
  DFFPOSX1 mem_reg_31__23_ ( .D(n3136), .CLK(clk), .Q(mem[1294]) );
  DFFPOSX1 mem_reg_31__22_ ( .D(n3135), .CLK(clk), .Q(mem[1293]) );
  DFFPOSX1 mem_reg_31__21_ ( .D(n3134), .CLK(clk), .Q(mem[1292]) );
  DFFPOSX1 mem_reg_31__20_ ( .D(n3133), .CLK(clk), .Q(mem[1291]) );
  DFFPOSX1 mem_reg_31__19_ ( .D(n3132), .CLK(clk), .Q(mem[1290]) );
  DFFPOSX1 mem_reg_31__18_ ( .D(n3131), .CLK(clk), .Q(mem[1289]) );
  DFFPOSX1 mem_reg_31__17_ ( .D(n3130), .CLK(clk), .Q(mem[1288]) );
  DFFPOSX1 mem_reg_31__16_ ( .D(n3129), .CLK(clk), .Q(mem[1287]) );
  DFFPOSX1 mem_reg_31__15_ ( .D(n3128), .CLK(clk), .Q(mem[1286]) );
  DFFPOSX1 mem_reg_31__14_ ( .D(n3127), .CLK(clk), .Q(mem[1285]) );
  DFFPOSX1 mem_reg_31__13_ ( .D(n3126), .CLK(clk), .Q(mem[1284]) );
  DFFPOSX1 mem_reg_31__12_ ( .D(n3125), .CLK(clk), .Q(mem[1283]) );
  DFFPOSX1 mem_reg_31__11_ ( .D(n3124), .CLK(clk), .Q(mem[1282]) );
  DFFPOSX1 mem_reg_31__10_ ( .D(n3123), .CLK(clk), .Q(mem[1281]) );
  DFFPOSX1 mem_reg_31__9_ ( .D(n3122), .CLK(clk), .Q(mem[1280]) );
  DFFPOSX1 mem_reg_31__8_ ( .D(n3121), .CLK(clk), .Q(mem[1279]) );
  DFFPOSX1 mem_reg_31__7_ ( .D(n3120), .CLK(clk), .Q(mem[1278]) );
  DFFPOSX1 mem_reg_31__6_ ( .D(n3119), .CLK(clk), .Q(mem[1277]) );
  DFFPOSX1 mem_reg_31__5_ ( .D(n3118), .CLK(clk), .Q(mem[1276]) );
  DFFPOSX1 mem_reg_31__4_ ( .D(n3117), .CLK(clk), .Q(mem[1275]) );
  DFFPOSX1 mem_reg_31__3_ ( .D(n3116), .CLK(clk), .Q(mem[1274]) );
  DFFPOSX1 mem_reg_31__2_ ( .D(n3115), .CLK(clk), .Q(mem[1273]) );
  DFFPOSX1 mem_reg_31__1_ ( .D(n3114), .CLK(clk), .Q(mem[1272]) );
  DFFPOSX1 mem_reg_31__0_ ( .D(n3113), .CLK(clk), .Q(mem[1271]) );
  DFFPOSX1 mem_reg_30__40_ ( .D(n3112), .CLK(clk), .Q(mem[1270]) );
  DFFPOSX1 mem_reg_30__39_ ( .D(n3111), .CLK(clk), .Q(mem[1269]) );
  DFFPOSX1 mem_reg_30__38_ ( .D(n3110), .CLK(clk), .Q(mem[1268]) );
  DFFPOSX1 mem_reg_30__37_ ( .D(n3109), .CLK(clk), .Q(mem[1267]) );
  DFFPOSX1 mem_reg_30__36_ ( .D(n3108), .CLK(clk), .Q(mem[1266]) );
  DFFPOSX1 mem_reg_30__35_ ( .D(n3107), .CLK(clk), .Q(mem[1265]) );
  DFFPOSX1 mem_reg_30__34_ ( .D(n3106), .CLK(clk), .Q(mem[1264]) );
  DFFPOSX1 mem_reg_30__33_ ( .D(n3105), .CLK(clk), .Q(mem[1263]) );
  DFFPOSX1 mem_reg_30__32_ ( .D(n3104), .CLK(clk), .Q(mem[1262]) );
  DFFPOSX1 mem_reg_30__31_ ( .D(n3103), .CLK(clk), .Q(mem[1261]) );
  DFFPOSX1 mem_reg_30__30_ ( .D(n3102), .CLK(clk), .Q(mem[1260]) );
  DFFPOSX1 mem_reg_30__29_ ( .D(n3101), .CLK(clk), .Q(mem[1259]) );
  DFFPOSX1 mem_reg_30__28_ ( .D(n3100), .CLK(clk), .Q(mem[1258]) );
  DFFPOSX1 mem_reg_30__27_ ( .D(n3099), .CLK(clk), .Q(mem[1257]) );
  DFFPOSX1 mem_reg_30__26_ ( .D(n3098), .CLK(clk), .Q(mem[1256]) );
  DFFPOSX1 mem_reg_30__25_ ( .D(n3097), .CLK(clk), .Q(mem[1255]) );
  DFFPOSX1 mem_reg_30__24_ ( .D(n3096), .CLK(clk), .Q(mem[1254]) );
  DFFPOSX1 mem_reg_30__23_ ( .D(n3095), .CLK(clk), .Q(mem[1253]) );
  DFFPOSX1 mem_reg_30__22_ ( .D(n3094), .CLK(clk), .Q(mem[1252]) );
  DFFPOSX1 mem_reg_30__21_ ( .D(n3093), .CLK(clk), .Q(mem[1251]) );
  DFFPOSX1 mem_reg_30__20_ ( .D(n3092), .CLK(clk), .Q(mem[1250]) );
  DFFPOSX1 mem_reg_30__19_ ( .D(n3091), .CLK(clk), .Q(mem[1249]) );
  DFFPOSX1 mem_reg_30__18_ ( .D(n3090), .CLK(clk), .Q(mem[1248]) );
  DFFPOSX1 mem_reg_30__17_ ( .D(n3089), .CLK(clk), .Q(mem[1247]) );
  DFFPOSX1 mem_reg_30__16_ ( .D(n3088), .CLK(clk), .Q(mem[1246]) );
  DFFPOSX1 mem_reg_30__15_ ( .D(n3087), .CLK(clk), .Q(mem[1245]) );
  DFFPOSX1 mem_reg_30__14_ ( .D(n3086), .CLK(clk), .Q(mem[1244]) );
  DFFPOSX1 mem_reg_30__13_ ( .D(n3085), .CLK(clk), .Q(mem[1243]) );
  DFFPOSX1 mem_reg_30__12_ ( .D(n3084), .CLK(clk), .Q(mem[1242]) );
  DFFPOSX1 mem_reg_30__11_ ( .D(n3083), .CLK(clk), .Q(mem[1241]) );
  DFFPOSX1 mem_reg_30__10_ ( .D(n3082), .CLK(clk), .Q(mem[1240]) );
  DFFPOSX1 mem_reg_30__9_ ( .D(n3081), .CLK(clk), .Q(mem[1239]) );
  DFFPOSX1 mem_reg_30__8_ ( .D(n3080), .CLK(clk), .Q(mem[1238]) );
  DFFPOSX1 mem_reg_30__7_ ( .D(n3079), .CLK(clk), .Q(mem[1237]) );
  DFFPOSX1 mem_reg_30__6_ ( .D(n3078), .CLK(clk), .Q(mem[1236]) );
  DFFPOSX1 mem_reg_30__5_ ( .D(n3077), .CLK(clk), .Q(mem[1235]) );
  DFFPOSX1 mem_reg_30__4_ ( .D(n3076), .CLK(clk), .Q(mem[1234]) );
  DFFPOSX1 mem_reg_30__3_ ( .D(n3075), .CLK(clk), .Q(mem[1233]) );
  DFFPOSX1 mem_reg_30__2_ ( .D(n3074), .CLK(clk), .Q(mem[1232]) );
  DFFPOSX1 mem_reg_30__1_ ( .D(n3073), .CLK(clk), .Q(mem[1231]) );
  DFFPOSX1 mem_reg_30__0_ ( .D(n3072), .CLK(clk), .Q(mem[1230]) );
  DFFPOSX1 mem_reg_29__40_ ( .D(n3071), .CLK(clk), .Q(mem[1229]) );
  DFFPOSX1 mem_reg_29__39_ ( .D(n3070), .CLK(clk), .Q(mem[1228]) );
  DFFPOSX1 mem_reg_29__38_ ( .D(n3069), .CLK(clk), .Q(mem[1227]) );
  DFFPOSX1 mem_reg_29__37_ ( .D(n3068), .CLK(clk), .Q(mem[1226]) );
  DFFPOSX1 mem_reg_29__36_ ( .D(n3067), .CLK(clk), .Q(mem[1225]) );
  DFFPOSX1 mem_reg_29__35_ ( .D(n3066), .CLK(clk), .Q(mem[1224]) );
  DFFPOSX1 mem_reg_29__34_ ( .D(n3065), .CLK(clk), .Q(mem[1223]) );
  DFFPOSX1 mem_reg_29__33_ ( .D(n3064), .CLK(clk), .Q(mem[1222]) );
  DFFPOSX1 mem_reg_29__32_ ( .D(n3063), .CLK(clk), .Q(mem[1221]) );
  DFFPOSX1 mem_reg_29__31_ ( .D(n3062), .CLK(clk), .Q(mem[1220]) );
  DFFPOSX1 mem_reg_29__30_ ( .D(n3061), .CLK(clk), .Q(mem[1219]) );
  DFFPOSX1 mem_reg_29__29_ ( .D(n3060), .CLK(clk), .Q(mem[1218]) );
  DFFPOSX1 mem_reg_29__28_ ( .D(n3059), .CLK(clk), .Q(mem[1217]) );
  DFFPOSX1 mem_reg_29__27_ ( .D(n3058), .CLK(clk), .Q(mem[1216]) );
  DFFPOSX1 mem_reg_29__26_ ( .D(n3057), .CLK(clk), .Q(mem[1215]) );
  DFFPOSX1 mem_reg_29__25_ ( .D(n3056), .CLK(clk), .Q(mem[1214]) );
  DFFPOSX1 mem_reg_29__24_ ( .D(n3055), .CLK(clk), .Q(mem[1213]) );
  DFFPOSX1 mem_reg_29__23_ ( .D(n3054), .CLK(clk), .Q(mem[1212]) );
  DFFPOSX1 mem_reg_29__22_ ( .D(n3053), .CLK(clk), .Q(mem[1211]) );
  DFFPOSX1 mem_reg_29__21_ ( .D(n3052), .CLK(clk), .Q(mem[1210]) );
  DFFPOSX1 mem_reg_29__20_ ( .D(n3051), .CLK(clk), .Q(mem[1209]) );
  DFFPOSX1 mem_reg_29__19_ ( .D(n3050), .CLK(clk), .Q(mem[1208]) );
  DFFPOSX1 mem_reg_29__18_ ( .D(n3049), .CLK(clk), .Q(mem[1207]) );
  DFFPOSX1 mem_reg_29__17_ ( .D(n3048), .CLK(clk), .Q(mem[1206]) );
  DFFPOSX1 mem_reg_29__16_ ( .D(n3047), .CLK(clk), .Q(mem[1205]) );
  DFFPOSX1 mem_reg_29__15_ ( .D(n3046), .CLK(clk), .Q(mem[1204]) );
  DFFPOSX1 mem_reg_29__14_ ( .D(n3045), .CLK(clk), .Q(mem[1203]) );
  DFFPOSX1 mem_reg_29__13_ ( .D(n3044), .CLK(clk), .Q(mem[1202]) );
  DFFPOSX1 mem_reg_29__12_ ( .D(n3043), .CLK(clk), .Q(mem[1201]) );
  DFFPOSX1 mem_reg_29__11_ ( .D(n3042), .CLK(clk), .Q(mem[1200]) );
  DFFPOSX1 mem_reg_29__10_ ( .D(n3041), .CLK(clk), .Q(mem[1199]) );
  DFFPOSX1 mem_reg_29__9_ ( .D(n3040), .CLK(clk), .Q(mem[1198]) );
  DFFPOSX1 mem_reg_29__8_ ( .D(n3039), .CLK(clk), .Q(mem[1197]) );
  DFFPOSX1 mem_reg_29__7_ ( .D(n3038), .CLK(clk), .Q(mem[1196]) );
  DFFPOSX1 mem_reg_29__6_ ( .D(n3037), .CLK(clk), .Q(mem[1195]) );
  DFFPOSX1 mem_reg_29__5_ ( .D(n3036), .CLK(clk), .Q(mem[1194]) );
  DFFPOSX1 mem_reg_29__4_ ( .D(n3035), .CLK(clk), .Q(mem[1193]) );
  DFFPOSX1 mem_reg_29__3_ ( .D(n3034), .CLK(clk), .Q(mem[1192]) );
  DFFPOSX1 mem_reg_29__2_ ( .D(n3033), .CLK(clk), .Q(mem[1191]) );
  DFFPOSX1 mem_reg_29__1_ ( .D(n3032), .CLK(clk), .Q(mem[1190]) );
  DFFPOSX1 mem_reg_29__0_ ( .D(n3031), .CLK(clk), .Q(mem[1189]) );
  DFFPOSX1 mem_reg_28__40_ ( .D(n3030), .CLK(clk), .Q(mem[1188]) );
  DFFPOSX1 mem_reg_28__39_ ( .D(n3029), .CLK(clk), .Q(mem[1187]) );
  DFFPOSX1 mem_reg_28__38_ ( .D(n3028), .CLK(clk), .Q(mem[1186]) );
  DFFPOSX1 mem_reg_28__37_ ( .D(n3027), .CLK(clk), .Q(mem[1185]) );
  DFFPOSX1 mem_reg_28__36_ ( .D(n3026), .CLK(clk), .Q(mem[1184]) );
  DFFPOSX1 mem_reg_28__35_ ( .D(n3025), .CLK(clk), .Q(mem[1183]) );
  DFFPOSX1 mem_reg_28__34_ ( .D(n3024), .CLK(clk), .Q(mem[1182]) );
  DFFPOSX1 mem_reg_28__33_ ( .D(n3023), .CLK(clk), .Q(mem[1181]) );
  DFFPOSX1 mem_reg_28__32_ ( .D(n3022), .CLK(clk), .Q(mem[1180]) );
  DFFPOSX1 mem_reg_28__31_ ( .D(n3021), .CLK(clk), .Q(mem[1179]) );
  DFFPOSX1 mem_reg_28__30_ ( .D(n3020), .CLK(clk), .Q(mem[1178]) );
  DFFPOSX1 mem_reg_28__29_ ( .D(n3019), .CLK(clk), .Q(mem[1177]) );
  DFFPOSX1 mem_reg_28__28_ ( .D(n3018), .CLK(clk), .Q(mem[1176]) );
  DFFPOSX1 mem_reg_28__27_ ( .D(n3017), .CLK(clk), .Q(mem[1175]) );
  DFFPOSX1 mem_reg_28__26_ ( .D(n3016), .CLK(clk), .Q(mem[1174]) );
  DFFPOSX1 mem_reg_28__25_ ( .D(n3015), .CLK(clk), .Q(mem[1173]) );
  DFFPOSX1 mem_reg_28__24_ ( .D(n3014), .CLK(clk), .Q(mem[1172]) );
  DFFPOSX1 mem_reg_28__23_ ( .D(n3013), .CLK(clk), .Q(mem[1171]) );
  DFFPOSX1 mem_reg_28__22_ ( .D(n3012), .CLK(clk), .Q(mem[1170]) );
  DFFPOSX1 mem_reg_28__21_ ( .D(n3011), .CLK(clk), .Q(mem[1169]) );
  DFFPOSX1 mem_reg_28__20_ ( .D(n3010), .CLK(clk), .Q(mem[1168]) );
  DFFPOSX1 mem_reg_28__19_ ( .D(n3009), .CLK(clk), .Q(mem[1167]) );
  DFFPOSX1 mem_reg_28__18_ ( .D(n3008), .CLK(clk), .Q(mem[1166]) );
  DFFPOSX1 mem_reg_28__17_ ( .D(n3007), .CLK(clk), .Q(mem[1165]) );
  DFFPOSX1 mem_reg_28__16_ ( .D(n3006), .CLK(clk), .Q(mem[1164]) );
  DFFPOSX1 mem_reg_28__15_ ( .D(n3005), .CLK(clk), .Q(mem[1163]) );
  DFFPOSX1 mem_reg_28__14_ ( .D(n3004), .CLK(clk), .Q(mem[1162]) );
  DFFPOSX1 mem_reg_28__13_ ( .D(n3003), .CLK(clk), .Q(mem[1161]) );
  DFFPOSX1 mem_reg_28__12_ ( .D(n3002), .CLK(clk), .Q(mem[1160]) );
  DFFPOSX1 mem_reg_28__11_ ( .D(n3001), .CLK(clk), .Q(mem[1159]) );
  DFFPOSX1 mem_reg_28__10_ ( .D(n3000), .CLK(clk), .Q(mem[1158]) );
  DFFPOSX1 mem_reg_28__9_ ( .D(n2999), .CLK(clk), .Q(mem[1157]) );
  DFFPOSX1 mem_reg_28__8_ ( .D(n2998), .CLK(clk), .Q(mem[1156]) );
  DFFPOSX1 mem_reg_28__7_ ( .D(n2997), .CLK(clk), .Q(mem[1155]) );
  DFFPOSX1 mem_reg_28__6_ ( .D(n2996), .CLK(clk), .Q(mem[1154]) );
  DFFPOSX1 mem_reg_28__5_ ( .D(n2995), .CLK(clk), .Q(mem[1153]) );
  DFFPOSX1 mem_reg_28__4_ ( .D(n2994), .CLK(clk), .Q(mem[1152]) );
  DFFPOSX1 mem_reg_28__3_ ( .D(n2993), .CLK(clk), .Q(mem[1151]) );
  DFFPOSX1 mem_reg_28__2_ ( .D(n2992), .CLK(clk), .Q(mem[1150]) );
  DFFPOSX1 mem_reg_28__1_ ( .D(n2991), .CLK(clk), .Q(mem[1149]) );
  DFFPOSX1 mem_reg_28__0_ ( .D(n2990), .CLK(clk), .Q(mem[1148]) );
  DFFPOSX1 mem_reg_27__40_ ( .D(n2989), .CLK(clk), .Q(mem[1147]) );
  DFFPOSX1 mem_reg_27__39_ ( .D(n2988), .CLK(clk), .Q(mem[1146]) );
  DFFPOSX1 mem_reg_27__38_ ( .D(n2987), .CLK(clk), .Q(mem[1145]) );
  DFFPOSX1 mem_reg_27__37_ ( .D(n2986), .CLK(clk), .Q(mem[1144]) );
  DFFPOSX1 mem_reg_27__36_ ( .D(n2985), .CLK(clk), .Q(mem[1143]) );
  DFFPOSX1 mem_reg_27__35_ ( .D(n2984), .CLK(clk), .Q(mem[1142]) );
  DFFPOSX1 mem_reg_27__34_ ( .D(n2983), .CLK(clk), .Q(mem[1141]) );
  DFFPOSX1 mem_reg_27__33_ ( .D(n2982), .CLK(clk), .Q(mem[1140]) );
  DFFPOSX1 mem_reg_27__32_ ( .D(n2981), .CLK(clk), .Q(mem[1139]) );
  DFFPOSX1 mem_reg_27__31_ ( .D(n2980), .CLK(clk), .Q(mem[1138]) );
  DFFPOSX1 mem_reg_27__30_ ( .D(n2979), .CLK(clk), .Q(mem[1137]) );
  DFFPOSX1 mem_reg_27__29_ ( .D(n2978), .CLK(clk), .Q(mem[1136]) );
  DFFPOSX1 mem_reg_27__28_ ( .D(n2977), .CLK(clk), .Q(mem[1135]) );
  DFFPOSX1 mem_reg_27__27_ ( .D(n2976), .CLK(clk), .Q(mem[1134]) );
  DFFPOSX1 mem_reg_27__26_ ( .D(n2975), .CLK(clk), .Q(mem[1133]) );
  DFFPOSX1 mem_reg_27__25_ ( .D(n2974), .CLK(clk), .Q(mem[1132]) );
  DFFPOSX1 mem_reg_27__24_ ( .D(n2973), .CLK(clk), .Q(mem[1131]) );
  DFFPOSX1 mem_reg_27__23_ ( .D(n2972), .CLK(clk), .Q(mem[1130]) );
  DFFPOSX1 mem_reg_27__22_ ( .D(n2971), .CLK(clk), .Q(mem[1129]) );
  DFFPOSX1 mem_reg_27__21_ ( .D(n2970), .CLK(clk), .Q(mem[1128]) );
  DFFPOSX1 mem_reg_27__20_ ( .D(n2969), .CLK(clk), .Q(mem[1127]) );
  DFFPOSX1 mem_reg_27__19_ ( .D(n2968), .CLK(clk), .Q(mem[1126]) );
  DFFPOSX1 mem_reg_27__18_ ( .D(n2967), .CLK(clk), .Q(mem[1125]) );
  DFFPOSX1 mem_reg_27__17_ ( .D(n2966), .CLK(clk), .Q(mem[1124]) );
  DFFPOSX1 mem_reg_27__16_ ( .D(n2965), .CLK(clk), .Q(mem[1123]) );
  DFFPOSX1 mem_reg_27__15_ ( .D(n2964), .CLK(clk), .Q(mem[1122]) );
  DFFPOSX1 mem_reg_27__14_ ( .D(n2963), .CLK(clk), .Q(mem[1121]) );
  DFFPOSX1 mem_reg_27__13_ ( .D(n2962), .CLK(clk), .Q(mem[1120]) );
  DFFPOSX1 mem_reg_27__12_ ( .D(n2961), .CLK(clk), .Q(mem[1119]) );
  DFFPOSX1 mem_reg_27__11_ ( .D(n2960), .CLK(clk), .Q(mem[1118]) );
  DFFPOSX1 mem_reg_27__10_ ( .D(n2959), .CLK(clk), .Q(mem[1117]) );
  DFFPOSX1 mem_reg_27__9_ ( .D(n2958), .CLK(clk), .Q(mem[1116]) );
  DFFPOSX1 mem_reg_27__8_ ( .D(n2957), .CLK(clk), .Q(mem[1115]) );
  DFFPOSX1 mem_reg_27__7_ ( .D(n2956), .CLK(clk), .Q(mem[1114]) );
  DFFPOSX1 mem_reg_27__6_ ( .D(n2955), .CLK(clk), .Q(mem[1113]) );
  DFFPOSX1 mem_reg_27__5_ ( .D(n2954), .CLK(clk), .Q(mem[1112]) );
  DFFPOSX1 mem_reg_27__4_ ( .D(n2953), .CLK(clk), .Q(mem[1111]) );
  DFFPOSX1 mem_reg_27__3_ ( .D(n2952), .CLK(clk), .Q(mem[1110]) );
  DFFPOSX1 mem_reg_27__2_ ( .D(n2951), .CLK(clk), .Q(mem[1109]) );
  DFFPOSX1 mem_reg_27__1_ ( .D(n2950), .CLK(clk), .Q(mem[1108]) );
  DFFPOSX1 mem_reg_27__0_ ( .D(n2949), .CLK(clk), .Q(mem[1107]) );
  DFFPOSX1 mem_reg_26__40_ ( .D(n2948), .CLK(clk), .Q(mem[1106]) );
  DFFPOSX1 mem_reg_26__39_ ( .D(n2947), .CLK(clk), .Q(mem[1105]) );
  DFFPOSX1 mem_reg_26__38_ ( .D(n2946), .CLK(clk), .Q(mem[1104]) );
  DFFPOSX1 mem_reg_26__37_ ( .D(n2945), .CLK(clk), .Q(mem[1103]) );
  DFFPOSX1 mem_reg_26__36_ ( .D(n2944), .CLK(clk), .Q(mem[1102]) );
  DFFPOSX1 mem_reg_26__35_ ( .D(n2943), .CLK(clk), .Q(mem[1101]) );
  DFFPOSX1 mem_reg_26__34_ ( .D(n2942), .CLK(clk), .Q(mem[1100]) );
  DFFPOSX1 mem_reg_26__33_ ( .D(n2941), .CLK(clk), .Q(mem[1099]) );
  DFFPOSX1 mem_reg_26__32_ ( .D(n2940), .CLK(clk), .Q(mem[1098]) );
  DFFPOSX1 mem_reg_26__31_ ( .D(n2939), .CLK(clk), .Q(mem[1097]) );
  DFFPOSX1 mem_reg_26__30_ ( .D(n2938), .CLK(clk), .Q(mem[1096]) );
  DFFPOSX1 mem_reg_26__29_ ( .D(n2937), .CLK(clk), .Q(mem[1095]) );
  DFFPOSX1 mem_reg_26__28_ ( .D(n2936), .CLK(clk), .Q(mem[1094]) );
  DFFPOSX1 mem_reg_26__27_ ( .D(n2935), .CLK(clk), .Q(mem[1093]) );
  DFFPOSX1 mem_reg_26__26_ ( .D(n2934), .CLK(clk), .Q(mem[1092]) );
  DFFPOSX1 mem_reg_26__25_ ( .D(n2933), .CLK(clk), .Q(mem[1091]) );
  DFFPOSX1 mem_reg_26__24_ ( .D(n2932), .CLK(clk), .Q(mem[1090]) );
  DFFPOSX1 mem_reg_26__23_ ( .D(n2931), .CLK(clk), .Q(mem[1089]) );
  DFFPOSX1 mem_reg_26__22_ ( .D(n2930), .CLK(clk), .Q(mem[1088]) );
  DFFPOSX1 mem_reg_26__21_ ( .D(n2929), .CLK(clk), .Q(mem[1087]) );
  DFFPOSX1 mem_reg_26__20_ ( .D(n2928), .CLK(clk), .Q(mem[1086]) );
  DFFPOSX1 mem_reg_26__19_ ( .D(n2927), .CLK(clk), .Q(mem[1085]) );
  DFFPOSX1 mem_reg_26__18_ ( .D(n2926), .CLK(clk), .Q(mem[1084]) );
  DFFPOSX1 mem_reg_26__17_ ( .D(n2925), .CLK(clk), .Q(mem[1083]) );
  DFFPOSX1 mem_reg_26__16_ ( .D(n2924), .CLK(clk), .Q(mem[1082]) );
  DFFPOSX1 mem_reg_26__15_ ( .D(n2923), .CLK(clk), .Q(mem[1081]) );
  DFFPOSX1 mem_reg_26__14_ ( .D(n2922), .CLK(clk), .Q(mem[1080]) );
  DFFPOSX1 mem_reg_26__13_ ( .D(n2921), .CLK(clk), .Q(mem[1079]) );
  DFFPOSX1 mem_reg_26__12_ ( .D(n2920), .CLK(clk), .Q(mem[1078]) );
  DFFPOSX1 mem_reg_26__11_ ( .D(n2919), .CLK(clk), .Q(mem[1077]) );
  DFFPOSX1 mem_reg_26__10_ ( .D(n2918), .CLK(clk), .Q(mem[1076]) );
  DFFPOSX1 mem_reg_26__9_ ( .D(n2917), .CLK(clk), .Q(mem[1075]) );
  DFFPOSX1 mem_reg_26__8_ ( .D(n2916), .CLK(clk), .Q(mem[1074]) );
  DFFPOSX1 mem_reg_26__7_ ( .D(n2915), .CLK(clk), .Q(mem[1073]) );
  DFFPOSX1 mem_reg_26__6_ ( .D(n2914), .CLK(clk), .Q(mem[1072]) );
  DFFPOSX1 mem_reg_26__5_ ( .D(n2913), .CLK(clk), .Q(mem[1071]) );
  DFFPOSX1 mem_reg_26__4_ ( .D(n2912), .CLK(clk), .Q(mem[1070]) );
  DFFPOSX1 mem_reg_26__3_ ( .D(n2911), .CLK(clk), .Q(mem[1069]) );
  DFFPOSX1 mem_reg_26__2_ ( .D(n2910), .CLK(clk), .Q(mem[1068]) );
  DFFPOSX1 mem_reg_26__1_ ( .D(n2909), .CLK(clk), .Q(mem[1067]) );
  DFFPOSX1 mem_reg_26__0_ ( .D(n2908), .CLK(clk), .Q(mem[1066]) );
  DFFPOSX1 mem_reg_25__40_ ( .D(n2907), .CLK(clk), .Q(mem[1065]) );
  DFFPOSX1 mem_reg_25__39_ ( .D(n2906), .CLK(clk), .Q(mem[1064]) );
  DFFPOSX1 mem_reg_25__38_ ( .D(n2905), .CLK(clk), .Q(mem[1063]) );
  DFFPOSX1 mem_reg_25__37_ ( .D(n2904), .CLK(clk), .Q(mem[1062]) );
  DFFPOSX1 mem_reg_25__36_ ( .D(n2903), .CLK(clk), .Q(mem[1061]) );
  DFFPOSX1 mem_reg_25__35_ ( .D(n2902), .CLK(clk), .Q(mem[1060]) );
  DFFPOSX1 mem_reg_25__34_ ( .D(n2901), .CLK(clk), .Q(mem[1059]) );
  DFFPOSX1 mem_reg_25__33_ ( .D(n2900), .CLK(clk), .Q(mem[1058]) );
  DFFPOSX1 mem_reg_25__32_ ( .D(n2899), .CLK(clk), .Q(mem[1057]) );
  DFFPOSX1 mem_reg_25__31_ ( .D(n2898), .CLK(clk), .Q(mem[1056]) );
  DFFPOSX1 mem_reg_25__30_ ( .D(n2897), .CLK(clk), .Q(mem[1055]) );
  DFFPOSX1 mem_reg_25__29_ ( .D(n2896), .CLK(clk), .Q(mem[1054]) );
  DFFPOSX1 mem_reg_25__28_ ( .D(n2895), .CLK(clk), .Q(mem[1053]) );
  DFFPOSX1 mem_reg_25__27_ ( .D(n2894), .CLK(clk), .Q(mem[1052]) );
  DFFPOSX1 mem_reg_25__26_ ( .D(n2893), .CLK(clk), .Q(mem[1051]) );
  DFFPOSX1 mem_reg_25__25_ ( .D(n2892), .CLK(clk), .Q(mem[1050]) );
  DFFPOSX1 mem_reg_25__24_ ( .D(n2891), .CLK(clk), .Q(mem[1049]) );
  DFFPOSX1 mem_reg_25__23_ ( .D(n2890), .CLK(clk), .Q(mem[1048]) );
  DFFPOSX1 mem_reg_25__22_ ( .D(n2889), .CLK(clk), .Q(mem[1047]) );
  DFFPOSX1 mem_reg_25__21_ ( .D(n2888), .CLK(clk), .Q(mem[1046]) );
  DFFPOSX1 mem_reg_25__20_ ( .D(n2887), .CLK(clk), .Q(mem[1045]) );
  DFFPOSX1 mem_reg_25__19_ ( .D(n2886), .CLK(clk), .Q(mem[1044]) );
  DFFPOSX1 mem_reg_25__18_ ( .D(n2885), .CLK(clk), .Q(mem[1043]) );
  DFFPOSX1 mem_reg_25__17_ ( .D(n2884), .CLK(clk), .Q(mem[1042]) );
  DFFPOSX1 mem_reg_25__16_ ( .D(n2883), .CLK(clk), .Q(mem[1041]) );
  DFFPOSX1 mem_reg_25__15_ ( .D(n2882), .CLK(clk), .Q(mem[1040]) );
  DFFPOSX1 mem_reg_25__14_ ( .D(n2881), .CLK(clk), .Q(mem[1039]) );
  DFFPOSX1 mem_reg_25__13_ ( .D(n2880), .CLK(clk), .Q(mem[1038]) );
  DFFPOSX1 mem_reg_25__12_ ( .D(n2879), .CLK(clk), .Q(mem[1037]) );
  DFFPOSX1 mem_reg_25__11_ ( .D(n2878), .CLK(clk), .Q(mem[1036]) );
  DFFPOSX1 mem_reg_25__10_ ( .D(n2877), .CLK(clk), .Q(mem[1035]) );
  DFFPOSX1 mem_reg_25__9_ ( .D(n2876), .CLK(clk), .Q(mem[1034]) );
  DFFPOSX1 mem_reg_25__8_ ( .D(n2875), .CLK(clk), .Q(mem[1033]) );
  DFFPOSX1 mem_reg_25__7_ ( .D(n2874), .CLK(clk), .Q(mem[1032]) );
  DFFPOSX1 mem_reg_25__6_ ( .D(n2873), .CLK(clk), .Q(mem[1031]) );
  DFFPOSX1 mem_reg_25__5_ ( .D(n2872), .CLK(clk), .Q(mem[1030]) );
  DFFPOSX1 mem_reg_25__4_ ( .D(n2871), .CLK(clk), .Q(mem[1029]) );
  DFFPOSX1 mem_reg_25__3_ ( .D(n2870), .CLK(clk), .Q(mem[1028]) );
  DFFPOSX1 mem_reg_25__2_ ( .D(n2869), .CLK(clk), .Q(mem[1027]) );
  DFFPOSX1 mem_reg_25__1_ ( .D(n2868), .CLK(clk), .Q(mem[1026]) );
  DFFPOSX1 mem_reg_25__0_ ( .D(n2867), .CLK(clk), .Q(mem[1025]) );
  DFFPOSX1 mem_reg_24__40_ ( .D(n2866), .CLK(clk), .Q(mem[1024]) );
  DFFPOSX1 mem_reg_24__39_ ( .D(n2865), .CLK(clk), .Q(mem[1023]) );
  DFFPOSX1 mem_reg_24__38_ ( .D(n2864), .CLK(clk), .Q(mem[1022]) );
  DFFPOSX1 mem_reg_24__37_ ( .D(n2863), .CLK(clk), .Q(mem[1021]) );
  DFFPOSX1 mem_reg_24__36_ ( .D(n2862), .CLK(clk), .Q(mem[1020]) );
  DFFPOSX1 mem_reg_24__35_ ( .D(n2861), .CLK(clk), .Q(mem[1019]) );
  DFFPOSX1 mem_reg_24__34_ ( .D(n2860), .CLK(clk), .Q(mem[1018]) );
  DFFPOSX1 mem_reg_24__33_ ( .D(n2859), .CLK(clk), .Q(mem[1017]) );
  DFFPOSX1 mem_reg_24__32_ ( .D(n2858), .CLK(clk), .Q(mem[1016]) );
  DFFPOSX1 mem_reg_24__31_ ( .D(n2857), .CLK(clk), .Q(mem[1015]) );
  DFFPOSX1 mem_reg_24__30_ ( .D(n2856), .CLK(clk), .Q(mem[1014]) );
  DFFPOSX1 mem_reg_24__29_ ( .D(n2855), .CLK(clk), .Q(mem[1013]) );
  DFFPOSX1 mem_reg_24__28_ ( .D(n2854), .CLK(clk), .Q(mem[1012]) );
  DFFPOSX1 mem_reg_24__27_ ( .D(n2853), .CLK(clk), .Q(mem[1011]) );
  DFFPOSX1 mem_reg_24__26_ ( .D(n2852), .CLK(clk), .Q(mem[1010]) );
  DFFPOSX1 mem_reg_24__25_ ( .D(n2851), .CLK(clk), .Q(mem[1009]) );
  DFFPOSX1 mem_reg_24__24_ ( .D(n2850), .CLK(clk), .Q(mem[1008]) );
  DFFPOSX1 mem_reg_24__23_ ( .D(n2849), .CLK(clk), .Q(mem[1007]) );
  DFFPOSX1 mem_reg_24__22_ ( .D(n2848), .CLK(clk), .Q(mem[1006]) );
  DFFPOSX1 mem_reg_24__21_ ( .D(n2847), .CLK(clk), .Q(mem[1005]) );
  DFFPOSX1 mem_reg_24__20_ ( .D(n2846), .CLK(clk), .Q(mem[1004]) );
  DFFPOSX1 mem_reg_24__19_ ( .D(n2845), .CLK(clk), .Q(mem[1003]) );
  DFFPOSX1 mem_reg_24__18_ ( .D(n2844), .CLK(clk), .Q(mem[1002]) );
  DFFPOSX1 mem_reg_24__17_ ( .D(n2843), .CLK(clk), .Q(mem[1001]) );
  DFFPOSX1 mem_reg_24__16_ ( .D(n2842), .CLK(clk), .Q(mem[1000]) );
  DFFPOSX1 mem_reg_24__15_ ( .D(n2841), .CLK(clk), .Q(mem[999]) );
  DFFPOSX1 mem_reg_24__14_ ( .D(n2840), .CLK(clk), .Q(mem[998]) );
  DFFPOSX1 mem_reg_24__13_ ( .D(n2839), .CLK(clk), .Q(mem[997]) );
  DFFPOSX1 mem_reg_24__12_ ( .D(n2838), .CLK(clk), .Q(mem[996]) );
  DFFPOSX1 mem_reg_24__11_ ( .D(n2837), .CLK(clk), .Q(mem[995]) );
  DFFPOSX1 mem_reg_24__10_ ( .D(n2836), .CLK(clk), .Q(mem[994]) );
  DFFPOSX1 mem_reg_24__9_ ( .D(n2835), .CLK(clk), .Q(mem[993]) );
  DFFPOSX1 mem_reg_24__8_ ( .D(n2834), .CLK(clk), .Q(mem[992]) );
  DFFPOSX1 mem_reg_24__7_ ( .D(n2833), .CLK(clk), .Q(mem[991]) );
  DFFPOSX1 mem_reg_24__6_ ( .D(n2832), .CLK(clk), .Q(mem[990]) );
  DFFPOSX1 mem_reg_24__5_ ( .D(n2831), .CLK(clk), .Q(mem[989]) );
  DFFPOSX1 mem_reg_24__4_ ( .D(n2830), .CLK(clk), .Q(mem[988]) );
  DFFPOSX1 mem_reg_24__3_ ( .D(n2829), .CLK(clk), .Q(mem[987]) );
  DFFPOSX1 mem_reg_24__2_ ( .D(n2828), .CLK(clk), .Q(mem[986]) );
  DFFPOSX1 mem_reg_24__1_ ( .D(n2827), .CLK(clk), .Q(mem[985]) );
  DFFPOSX1 mem_reg_24__0_ ( .D(n2826), .CLK(clk), .Q(mem[984]) );
  DFFPOSX1 mem_reg_23__40_ ( .D(n2825), .CLK(clk), .Q(mem[983]) );
  DFFPOSX1 mem_reg_23__39_ ( .D(n2824), .CLK(clk), .Q(mem[982]) );
  DFFPOSX1 mem_reg_23__38_ ( .D(n2823), .CLK(clk), .Q(mem[981]) );
  DFFPOSX1 mem_reg_23__37_ ( .D(n2822), .CLK(clk), .Q(mem[980]) );
  DFFPOSX1 mem_reg_23__36_ ( .D(n2821), .CLK(clk), .Q(mem[979]) );
  DFFPOSX1 mem_reg_23__35_ ( .D(n2820), .CLK(clk), .Q(mem[978]) );
  DFFPOSX1 mem_reg_23__34_ ( .D(n2819), .CLK(clk), .Q(mem[977]) );
  DFFPOSX1 mem_reg_23__33_ ( .D(n2818), .CLK(clk), .Q(mem[976]) );
  DFFPOSX1 mem_reg_23__32_ ( .D(n2817), .CLK(clk), .Q(mem[975]) );
  DFFPOSX1 mem_reg_23__31_ ( .D(n2816), .CLK(clk), .Q(mem[974]) );
  DFFPOSX1 mem_reg_23__30_ ( .D(n2815), .CLK(clk), .Q(mem[973]) );
  DFFPOSX1 mem_reg_23__29_ ( .D(n2814), .CLK(clk), .Q(mem[972]) );
  DFFPOSX1 mem_reg_23__28_ ( .D(n2813), .CLK(clk), .Q(mem[971]) );
  DFFPOSX1 mem_reg_23__27_ ( .D(n2812), .CLK(clk), .Q(mem[970]) );
  DFFPOSX1 mem_reg_23__26_ ( .D(n2811), .CLK(clk), .Q(mem[969]) );
  DFFPOSX1 mem_reg_23__25_ ( .D(n2810), .CLK(clk), .Q(mem[968]) );
  DFFPOSX1 mem_reg_23__24_ ( .D(n2809), .CLK(clk), .Q(mem[967]) );
  DFFPOSX1 mem_reg_23__23_ ( .D(n2808), .CLK(clk), .Q(mem[966]) );
  DFFPOSX1 mem_reg_23__22_ ( .D(n2807), .CLK(clk), .Q(mem[965]) );
  DFFPOSX1 mem_reg_23__21_ ( .D(n2806), .CLK(clk), .Q(mem[964]) );
  DFFPOSX1 mem_reg_23__20_ ( .D(n2805), .CLK(clk), .Q(mem[963]) );
  DFFPOSX1 mem_reg_23__19_ ( .D(n2804), .CLK(clk), .Q(mem[962]) );
  DFFPOSX1 mem_reg_23__18_ ( .D(n2803), .CLK(clk), .Q(mem[961]) );
  DFFPOSX1 mem_reg_23__17_ ( .D(n2802), .CLK(clk), .Q(mem[960]) );
  DFFPOSX1 mem_reg_23__16_ ( .D(n2801), .CLK(clk), .Q(mem[959]) );
  DFFPOSX1 mem_reg_23__15_ ( .D(n2800), .CLK(clk), .Q(mem[958]) );
  DFFPOSX1 mem_reg_23__14_ ( .D(n2799), .CLK(clk), .Q(mem[957]) );
  DFFPOSX1 mem_reg_23__13_ ( .D(n2798), .CLK(clk), .Q(mem[956]) );
  DFFPOSX1 mem_reg_23__12_ ( .D(n2797), .CLK(clk), .Q(mem[955]) );
  DFFPOSX1 mem_reg_23__11_ ( .D(n2796), .CLK(clk), .Q(mem[954]) );
  DFFPOSX1 mem_reg_23__10_ ( .D(n2795), .CLK(clk), .Q(mem[953]) );
  DFFPOSX1 mem_reg_23__9_ ( .D(n2794), .CLK(clk), .Q(mem[952]) );
  DFFPOSX1 mem_reg_23__8_ ( .D(n2793), .CLK(clk), .Q(mem[951]) );
  DFFPOSX1 mem_reg_23__7_ ( .D(n2792), .CLK(clk), .Q(mem[950]) );
  DFFPOSX1 mem_reg_23__6_ ( .D(n2791), .CLK(clk), .Q(mem[949]) );
  DFFPOSX1 mem_reg_23__5_ ( .D(n2790), .CLK(clk), .Q(mem[948]) );
  DFFPOSX1 mem_reg_23__4_ ( .D(n2789), .CLK(clk), .Q(mem[947]) );
  DFFPOSX1 mem_reg_23__3_ ( .D(n2788), .CLK(clk), .Q(mem[946]) );
  DFFPOSX1 mem_reg_23__2_ ( .D(n2787), .CLK(clk), .Q(mem[945]) );
  DFFPOSX1 mem_reg_23__1_ ( .D(n2786), .CLK(clk), .Q(mem[944]) );
  DFFPOSX1 mem_reg_23__0_ ( .D(n2785), .CLK(clk), .Q(mem[943]) );
  DFFPOSX1 mem_reg_22__40_ ( .D(n2784), .CLK(clk), .Q(mem[942]) );
  DFFPOSX1 mem_reg_22__39_ ( .D(n2783), .CLK(clk), .Q(mem[941]) );
  DFFPOSX1 mem_reg_22__38_ ( .D(n2782), .CLK(clk), .Q(mem[940]) );
  DFFPOSX1 mem_reg_22__37_ ( .D(n2781), .CLK(clk), .Q(mem[939]) );
  DFFPOSX1 mem_reg_22__36_ ( .D(n2780), .CLK(clk), .Q(mem[938]) );
  DFFPOSX1 mem_reg_22__35_ ( .D(n2779), .CLK(clk), .Q(mem[937]) );
  DFFPOSX1 mem_reg_22__34_ ( .D(n2778), .CLK(clk), .Q(mem[936]) );
  DFFPOSX1 mem_reg_22__33_ ( .D(n2777), .CLK(clk), .Q(mem[935]) );
  DFFPOSX1 mem_reg_22__32_ ( .D(n2776), .CLK(clk), .Q(mem[934]) );
  DFFPOSX1 mem_reg_22__31_ ( .D(n2775), .CLK(clk), .Q(mem[933]) );
  DFFPOSX1 mem_reg_22__30_ ( .D(n2774), .CLK(clk), .Q(mem[932]) );
  DFFPOSX1 mem_reg_22__29_ ( .D(n2773), .CLK(clk), .Q(mem[931]) );
  DFFPOSX1 mem_reg_22__28_ ( .D(n2772), .CLK(clk), .Q(mem[930]) );
  DFFPOSX1 mem_reg_22__27_ ( .D(n2771), .CLK(clk), .Q(mem[929]) );
  DFFPOSX1 mem_reg_22__26_ ( .D(n2770), .CLK(clk), .Q(mem[928]) );
  DFFPOSX1 mem_reg_22__25_ ( .D(n2769), .CLK(clk), .Q(mem[927]) );
  DFFPOSX1 mem_reg_22__24_ ( .D(n2768), .CLK(clk), .Q(mem[926]) );
  DFFPOSX1 mem_reg_22__23_ ( .D(n2767), .CLK(clk), .Q(mem[925]) );
  DFFPOSX1 mem_reg_22__22_ ( .D(n2766), .CLK(clk), .Q(mem[924]) );
  DFFPOSX1 mem_reg_22__21_ ( .D(n2765), .CLK(clk), .Q(mem[923]) );
  DFFPOSX1 mem_reg_22__20_ ( .D(n2764), .CLK(clk), .Q(mem[922]) );
  DFFPOSX1 mem_reg_22__19_ ( .D(n2763), .CLK(clk), .Q(mem[921]) );
  DFFPOSX1 mem_reg_22__18_ ( .D(n2762), .CLK(clk), .Q(mem[920]) );
  DFFPOSX1 mem_reg_22__17_ ( .D(n2761), .CLK(clk), .Q(mem[919]) );
  DFFPOSX1 mem_reg_22__16_ ( .D(n2760), .CLK(clk), .Q(mem[918]) );
  DFFPOSX1 mem_reg_22__15_ ( .D(n2759), .CLK(clk), .Q(mem[917]) );
  DFFPOSX1 mem_reg_22__14_ ( .D(n2758), .CLK(clk), .Q(mem[916]) );
  DFFPOSX1 mem_reg_22__13_ ( .D(n2757), .CLK(clk), .Q(mem[915]) );
  DFFPOSX1 mem_reg_22__12_ ( .D(n2756), .CLK(clk), .Q(mem[914]) );
  DFFPOSX1 mem_reg_22__11_ ( .D(n2755), .CLK(clk), .Q(mem[913]) );
  DFFPOSX1 mem_reg_22__10_ ( .D(n2754), .CLK(clk), .Q(mem[912]) );
  DFFPOSX1 mem_reg_22__9_ ( .D(n2753), .CLK(clk), .Q(mem[911]) );
  DFFPOSX1 mem_reg_22__8_ ( .D(n2752), .CLK(clk), .Q(mem[910]) );
  DFFPOSX1 mem_reg_22__7_ ( .D(n2751), .CLK(clk), .Q(mem[909]) );
  DFFPOSX1 mem_reg_22__6_ ( .D(n2750), .CLK(clk), .Q(mem[908]) );
  DFFPOSX1 mem_reg_22__5_ ( .D(n2749), .CLK(clk), .Q(mem[907]) );
  DFFPOSX1 mem_reg_22__4_ ( .D(n2748), .CLK(clk), .Q(mem[906]) );
  DFFPOSX1 mem_reg_22__3_ ( .D(n2747), .CLK(clk), .Q(mem[905]) );
  DFFPOSX1 mem_reg_22__2_ ( .D(n2746), .CLK(clk), .Q(mem[904]) );
  DFFPOSX1 mem_reg_22__1_ ( .D(n2745), .CLK(clk), .Q(mem[903]) );
  DFFPOSX1 mem_reg_22__0_ ( .D(n2744), .CLK(clk), .Q(mem[902]) );
  DFFPOSX1 mem_reg_21__40_ ( .D(n2743), .CLK(clk), .Q(mem[901]) );
  DFFPOSX1 mem_reg_21__39_ ( .D(n2742), .CLK(clk), .Q(mem[900]) );
  DFFPOSX1 mem_reg_21__38_ ( .D(n2741), .CLK(clk), .Q(mem[899]) );
  DFFPOSX1 mem_reg_21__37_ ( .D(n2740), .CLK(clk), .Q(mem[898]) );
  DFFPOSX1 mem_reg_21__36_ ( .D(n2739), .CLK(clk), .Q(mem[897]) );
  DFFPOSX1 mem_reg_21__35_ ( .D(n2738), .CLK(clk), .Q(mem[896]) );
  DFFPOSX1 mem_reg_21__34_ ( .D(n2737), .CLK(clk), .Q(mem[895]) );
  DFFPOSX1 mem_reg_21__33_ ( .D(n2736), .CLK(clk), .Q(mem[894]) );
  DFFPOSX1 mem_reg_21__32_ ( .D(n2735), .CLK(clk), .Q(mem[893]) );
  DFFPOSX1 mem_reg_21__31_ ( .D(n2734), .CLK(clk), .Q(mem[892]) );
  DFFPOSX1 mem_reg_21__30_ ( .D(n2733), .CLK(clk), .Q(mem[891]) );
  DFFPOSX1 mem_reg_21__29_ ( .D(n2732), .CLK(clk), .Q(mem[890]) );
  DFFPOSX1 mem_reg_21__28_ ( .D(n2731), .CLK(clk), .Q(mem[889]) );
  DFFPOSX1 mem_reg_21__27_ ( .D(n2730), .CLK(clk), .Q(mem[888]) );
  DFFPOSX1 mem_reg_21__26_ ( .D(n2729), .CLK(clk), .Q(mem[887]) );
  DFFPOSX1 mem_reg_21__25_ ( .D(n2728), .CLK(clk), .Q(mem[886]) );
  DFFPOSX1 mem_reg_21__24_ ( .D(n2727), .CLK(clk), .Q(mem[885]) );
  DFFPOSX1 mem_reg_21__23_ ( .D(n2726), .CLK(clk), .Q(mem[884]) );
  DFFPOSX1 mem_reg_21__22_ ( .D(n2725), .CLK(clk), .Q(mem[883]) );
  DFFPOSX1 mem_reg_21__21_ ( .D(n2724), .CLK(clk), .Q(mem[882]) );
  DFFPOSX1 mem_reg_21__20_ ( .D(n2723), .CLK(clk), .Q(mem[881]) );
  DFFPOSX1 mem_reg_21__19_ ( .D(n2722), .CLK(clk), .Q(mem[880]) );
  DFFPOSX1 mem_reg_21__18_ ( .D(n2721), .CLK(clk), .Q(mem[879]) );
  DFFPOSX1 mem_reg_21__17_ ( .D(n2720), .CLK(clk), .Q(mem[878]) );
  DFFPOSX1 mem_reg_21__16_ ( .D(n2719), .CLK(clk), .Q(mem[877]) );
  DFFPOSX1 mem_reg_21__15_ ( .D(n2718), .CLK(clk), .Q(mem[876]) );
  DFFPOSX1 mem_reg_21__14_ ( .D(n2717), .CLK(clk), .Q(mem[875]) );
  DFFPOSX1 mem_reg_21__13_ ( .D(n2716), .CLK(clk), .Q(mem[874]) );
  DFFPOSX1 mem_reg_21__12_ ( .D(n2715), .CLK(clk), .Q(mem[873]) );
  DFFPOSX1 mem_reg_21__11_ ( .D(n2714), .CLK(clk), .Q(mem[872]) );
  DFFPOSX1 mem_reg_21__10_ ( .D(n2713), .CLK(clk), .Q(mem[871]) );
  DFFPOSX1 mem_reg_21__9_ ( .D(n2712), .CLK(clk), .Q(mem[870]) );
  DFFPOSX1 mem_reg_21__8_ ( .D(n2711), .CLK(clk), .Q(mem[869]) );
  DFFPOSX1 mem_reg_21__7_ ( .D(n2710), .CLK(clk), .Q(mem[868]) );
  DFFPOSX1 mem_reg_21__6_ ( .D(n2709), .CLK(clk), .Q(mem[867]) );
  DFFPOSX1 mem_reg_21__5_ ( .D(n2708), .CLK(clk), .Q(mem[866]) );
  DFFPOSX1 mem_reg_21__4_ ( .D(n2707), .CLK(clk), .Q(mem[865]) );
  DFFPOSX1 mem_reg_21__3_ ( .D(n2706), .CLK(clk), .Q(mem[864]) );
  DFFPOSX1 mem_reg_21__2_ ( .D(n2705), .CLK(clk), .Q(mem[863]) );
  DFFPOSX1 mem_reg_21__1_ ( .D(n2704), .CLK(clk), .Q(mem[862]) );
  DFFPOSX1 mem_reg_21__0_ ( .D(n2703), .CLK(clk), .Q(mem[861]) );
  DFFPOSX1 mem_reg_20__40_ ( .D(n2702), .CLK(clk), .Q(mem[860]) );
  DFFPOSX1 mem_reg_20__39_ ( .D(n2701), .CLK(clk), .Q(mem[859]) );
  DFFPOSX1 mem_reg_20__38_ ( .D(n2700), .CLK(clk), .Q(mem[858]) );
  DFFPOSX1 mem_reg_20__37_ ( .D(n2699), .CLK(clk), .Q(mem[857]) );
  DFFPOSX1 mem_reg_20__36_ ( .D(n2698), .CLK(clk), .Q(mem[856]) );
  DFFPOSX1 mem_reg_20__35_ ( .D(n2697), .CLK(clk), .Q(mem[855]) );
  DFFPOSX1 mem_reg_20__34_ ( .D(n2696), .CLK(clk), .Q(mem[854]) );
  DFFPOSX1 mem_reg_20__33_ ( .D(n2695), .CLK(clk), .Q(mem[853]) );
  DFFPOSX1 mem_reg_20__32_ ( .D(n2694), .CLK(clk), .Q(mem[852]) );
  DFFPOSX1 mem_reg_20__31_ ( .D(n2693), .CLK(clk), .Q(mem[851]) );
  DFFPOSX1 mem_reg_20__30_ ( .D(n2692), .CLK(clk), .Q(mem[850]) );
  DFFPOSX1 mem_reg_20__29_ ( .D(n2691), .CLK(clk), .Q(mem[849]) );
  DFFPOSX1 mem_reg_20__28_ ( .D(n2690), .CLK(clk), .Q(mem[848]) );
  DFFPOSX1 mem_reg_20__27_ ( .D(n2689), .CLK(clk), .Q(mem[847]) );
  DFFPOSX1 mem_reg_20__26_ ( .D(n2688), .CLK(clk), .Q(mem[846]) );
  DFFPOSX1 mem_reg_20__25_ ( .D(n2687), .CLK(clk), .Q(mem[845]) );
  DFFPOSX1 mem_reg_20__24_ ( .D(n2686), .CLK(clk), .Q(mem[844]) );
  DFFPOSX1 mem_reg_20__23_ ( .D(n2685), .CLK(clk), .Q(mem[843]) );
  DFFPOSX1 mem_reg_20__22_ ( .D(n2684), .CLK(clk), .Q(mem[842]) );
  DFFPOSX1 mem_reg_20__21_ ( .D(n2683), .CLK(clk), .Q(mem[841]) );
  DFFPOSX1 mem_reg_20__20_ ( .D(n2682), .CLK(clk), .Q(mem[840]) );
  DFFPOSX1 mem_reg_20__19_ ( .D(n2681), .CLK(clk), .Q(mem[839]) );
  DFFPOSX1 mem_reg_20__18_ ( .D(n2680), .CLK(clk), .Q(mem[838]) );
  DFFPOSX1 mem_reg_20__17_ ( .D(n2679), .CLK(clk), .Q(mem[837]) );
  DFFPOSX1 mem_reg_20__16_ ( .D(n2678), .CLK(clk), .Q(mem[836]) );
  DFFPOSX1 mem_reg_20__15_ ( .D(n2677), .CLK(clk), .Q(mem[835]) );
  DFFPOSX1 mem_reg_20__14_ ( .D(n2676), .CLK(clk), .Q(mem[834]) );
  DFFPOSX1 mem_reg_20__13_ ( .D(n2675), .CLK(clk), .Q(mem[833]) );
  DFFPOSX1 mem_reg_20__12_ ( .D(n2674), .CLK(clk), .Q(mem[832]) );
  DFFPOSX1 mem_reg_20__11_ ( .D(n2673), .CLK(clk), .Q(mem[831]) );
  DFFPOSX1 mem_reg_20__10_ ( .D(n2672), .CLK(clk), .Q(mem[830]) );
  DFFPOSX1 mem_reg_20__9_ ( .D(n2671), .CLK(clk), .Q(mem[829]) );
  DFFPOSX1 mem_reg_20__8_ ( .D(n2670), .CLK(clk), .Q(mem[828]) );
  DFFPOSX1 mem_reg_20__7_ ( .D(n2669), .CLK(clk), .Q(mem[827]) );
  DFFPOSX1 mem_reg_20__6_ ( .D(n2668), .CLK(clk), .Q(mem[826]) );
  DFFPOSX1 mem_reg_20__5_ ( .D(n2667), .CLK(clk), .Q(mem[825]) );
  DFFPOSX1 mem_reg_20__4_ ( .D(n2666), .CLK(clk), .Q(mem[824]) );
  DFFPOSX1 mem_reg_20__3_ ( .D(n2665), .CLK(clk), .Q(mem[823]) );
  DFFPOSX1 mem_reg_20__2_ ( .D(n2664), .CLK(clk), .Q(mem[822]) );
  DFFPOSX1 mem_reg_20__1_ ( .D(n2663), .CLK(clk), .Q(mem[821]) );
  DFFPOSX1 mem_reg_20__0_ ( .D(n2662), .CLK(clk), .Q(mem[820]) );
  DFFPOSX1 mem_reg_19__40_ ( .D(n2661), .CLK(clk), .Q(mem[819]) );
  DFFPOSX1 mem_reg_19__39_ ( .D(n2660), .CLK(clk), .Q(mem[818]) );
  DFFPOSX1 mem_reg_19__38_ ( .D(n2659), .CLK(clk), .Q(mem[817]) );
  DFFPOSX1 mem_reg_19__37_ ( .D(n2658), .CLK(clk), .Q(mem[816]) );
  DFFPOSX1 mem_reg_19__36_ ( .D(n2657), .CLK(clk), .Q(mem[815]) );
  DFFPOSX1 mem_reg_19__35_ ( .D(n2656), .CLK(clk), .Q(mem[814]) );
  DFFPOSX1 mem_reg_19__34_ ( .D(n2655), .CLK(clk), .Q(mem[813]) );
  DFFPOSX1 mem_reg_19__33_ ( .D(n2654), .CLK(clk), .Q(mem[812]) );
  DFFPOSX1 mem_reg_19__32_ ( .D(n2653), .CLK(clk), .Q(mem[811]) );
  DFFPOSX1 mem_reg_19__31_ ( .D(n2652), .CLK(clk), .Q(mem[810]) );
  DFFPOSX1 mem_reg_19__30_ ( .D(n2651), .CLK(clk), .Q(mem[809]) );
  DFFPOSX1 mem_reg_19__29_ ( .D(n2650), .CLK(clk), .Q(mem[808]) );
  DFFPOSX1 mem_reg_19__28_ ( .D(n2649), .CLK(clk), .Q(mem[807]) );
  DFFPOSX1 mem_reg_19__27_ ( .D(n2648), .CLK(clk), .Q(mem[806]) );
  DFFPOSX1 mem_reg_19__26_ ( .D(n2647), .CLK(clk), .Q(mem[805]) );
  DFFPOSX1 mem_reg_19__25_ ( .D(n2646), .CLK(clk), .Q(mem[804]) );
  DFFPOSX1 mem_reg_19__24_ ( .D(n2645), .CLK(clk), .Q(mem[803]) );
  DFFPOSX1 mem_reg_19__23_ ( .D(n2644), .CLK(clk), .Q(mem[802]) );
  DFFPOSX1 mem_reg_19__22_ ( .D(n2643), .CLK(clk), .Q(mem[801]) );
  DFFPOSX1 mem_reg_19__21_ ( .D(n2642), .CLK(clk), .Q(mem[800]) );
  DFFPOSX1 mem_reg_19__20_ ( .D(n2641), .CLK(clk), .Q(mem[799]) );
  DFFPOSX1 mem_reg_19__19_ ( .D(n2640), .CLK(clk), .Q(mem[798]) );
  DFFPOSX1 mem_reg_19__18_ ( .D(n2639), .CLK(clk), .Q(mem[797]) );
  DFFPOSX1 mem_reg_19__17_ ( .D(n2638), .CLK(clk), .Q(mem[796]) );
  DFFPOSX1 mem_reg_19__16_ ( .D(n2637), .CLK(clk), .Q(mem[795]) );
  DFFPOSX1 mem_reg_19__15_ ( .D(n2636), .CLK(clk), .Q(mem[794]) );
  DFFPOSX1 mem_reg_19__14_ ( .D(n2635), .CLK(clk), .Q(mem[793]) );
  DFFPOSX1 mem_reg_19__13_ ( .D(n2634), .CLK(clk), .Q(mem[792]) );
  DFFPOSX1 mem_reg_19__12_ ( .D(n2633), .CLK(clk), .Q(mem[791]) );
  DFFPOSX1 mem_reg_19__11_ ( .D(n2632), .CLK(clk), .Q(mem[790]) );
  DFFPOSX1 mem_reg_19__10_ ( .D(n2631), .CLK(clk), .Q(mem[789]) );
  DFFPOSX1 mem_reg_19__9_ ( .D(n2630), .CLK(clk), .Q(mem[788]) );
  DFFPOSX1 mem_reg_19__8_ ( .D(n2629), .CLK(clk), .Q(mem[787]) );
  DFFPOSX1 mem_reg_19__7_ ( .D(n2628), .CLK(clk), .Q(mem[786]) );
  DFFPOSX1 mem_reg_19__6_ ( .D(n2627), .CLK(clk), .Q(mem[785]) );
  DFFPOSX1 mem_reg_19__5_ ( .D(n2626), .CLK(clk), .Q(mem[784]) );
  DFFPOSX1 mem_reg_19__4_ ( .D(n2625), .CLK(clk), .Q(mem[783]) );
  DFFPOSX1 mem_reg_19__3_ ( .D(n2624), .CLK(clk), .Q(mem[782]) );
  DFFPOSX1 mem_reg_19__2_ ( .D(n2623), .CLK(clk), .Q(mem[781]) );
  DFFPOSX1 mem_reg_19__1_ ( .D(n2622), .CLK(clk), .Q(mem[780]) );
  DFFPOSX1 mem_reg_19__0_ ( .D(n2621), .CLK(clk), .Q(mem[779]) );
  DFFPOSX1 mem_reg_18__40_ ( .D(n2620), .CLK(clk), .Q(mem[778]) );
  DFFPOSX1 mem_reg_18__39_ ( .D(n2619), .CLK(clk), .Q(mem[777]) );
  DFFPOSX1 mem_reg_18__38_ ( .D(n2618), .CLK(clk), .Q(mem[776]) );
  DFFPOSX1 mem_reg_18__37_ ( .D(n2617), .CLK(clk), .Q(mem[775]) );
  DFFPOSX1 mem_reg_18__36_ ( .D(n2616), .CLK(clk), .Q(mem[774]) );
  DFFPOSX1 mem_reg_18__35_ ( .D(n2615), .CLK(clk), .Q(mem[773]) );
  DFFPOSX1 mem_reg_18__34_ ( .D(n2614), .CLK(clk), .Q(mem[772]) );
  DFFPOSX1 mem_reg_18__33_ ( .D(n2613), .CLK(clk), .Q(mem[771]) );
  DFFPOSX1 mem_reg_18__32_ ( .D(n2612), .CLK(clk), .Q(mem[770]) );
  DFFPOSX1 mem_reg_18__31_ ( .D(n2611), .CLK(clk), .Q(mem[769]) );
  DFFPOSX1 mem_reg_18__30_ ( .D(n2610), .CLK(clk), .Q(mem[768]) );
  DFFPOSX1 mem_reg_18__29_ ( .D(n2609), .CLK(clk), .Q(mem[767]) );
  DFFPOSX1 mem_reg_18__28_ ( .D(n2608), .CLK(clk), .Q(mem[766]) );
  DFFPOSX1 mem_reg_18__27_ ( .D(n2607), .CLK(clk), .Q(mem[765]) );
  DFFPOSX1 mem_reg_18__26_ ( .D(n2606), .CLK(clk), .Q(mem[764]) );
  DFFPOSX1 mem_reg_18__25_ ( .D(n2605), .CLK(clk), .Q(mem[763]) );
  DFFPOSX1 mem_reg_18__24_ ( .D(n2604), .CLK(clk), .Q(mem[762]) );
  DFFPOSX1 mem_reg_18__23_ ( .D(n2603), .CLK(clk), .Q(mem[761]) );
  DFFPOSX1 mem_reg_18__22_ ( .D(n2602), .CLK(clk), .Q(mem[760]) );
  DFFPOSX1 mem_reg_18__21_ ( .D(n2601), .CLK(clk), .Q(mem[759]) );
  DFFPOSX1 mem_reg_18__20_ ( .D(n2600), .CLK(clk), .Q(mem[758]) );
  DFFPOSX1 mem_reg_18__19_ ( .D(n2599), .CLK(clk), .Q(mem[757]) );
  DFFPOSX1 mem_reg_18__18_ ( .D(n2598), .CLK(clk), .Q(mem[756]) );
  DFFPOSX1 mem_reg_18__17_ ( .D(n2597), .CLK(clk), .Q(mem[755]) );
  DFFPOSX1 mem_reg_18__16_ ( .D(n2596), .CLK(clk), .Q(mem[754]) );
  DFFPOSX1 mem_reg_18__15_ ( .D(n2595), .CLK(clk), .Q(mem[753]) );
  DFFPOSX1 mem_reg_18__14_ ( .D(n2594), .CLK(clk), .Q(mem[752]) );
  DFFPOSX1 mem_reg_18__13_ ( .D(n2593), .CLK(clk), .Q(mem[751]) );
  DFFPOSX1 mem_reg_18__12_ ( .D(n2592), .CLK(clk), .Q(mem[750]) );
  DFFPOSX1 mem_reg_18__11_ ( .D(n2591), .CLK(clk), .Q(mem[749]) );
  DFFPOSX1 mem_reg_18__10_ ( .D(n2590), .CLK(clk), .Q(mem[748]) );
  DFFPOSX1 mem_reg_18__9_ ( .D(n2589), .CLK(clk), .Q(mem[747]) );
  DFFPOSX1 mem_reg_18__8_ ( .D(n2588), .CLK(clk), .Q(mem[746]) );
  DFFPOSX1 mem_reg_18__7_ ( .D(n2587), .CLK(clk), .Q(mem[745]) );
  DFFPOSX1 mem_reg_18__6_ ( .D(n2586), .CLK(clk), .Q(mem[744]) );
  DFFPOSX1 mem_reg_18__5_ ( .D(n2585), .CLK(clk), .Q(mem[743]) );
  DFFPOSX1 mem_reg_18__4_ ( .D(n2584), .CLK(clk), .Q(mem[742]) );
  DFFPOSX1 mem_reg_18__3_ ( .D(n2583), .CLK(clk), .Q(mem[741]) );
  DFFPOSX1 mem_reg_18__2_ ( .D(n2582), .CLK(clk), .Q(mem[740]) );
  DFFPOSX1 mem_reg_18__1_ ( .D(n2581), .CLK(clk), .Q(mem[739]) );
  DFFPOSX1 mem_reg_18__0_ ( .D(n2580), .CLK(clk), .Q(mem[738]) );
  DFFPOSX1 mem_reg_17__40_ ( .D(n2579), .CLK(clk), .Q(mem[737]) );
  DFFPOSX1 mem_reg_17__39_ ( .D(n2578), .CLK(clk), .Q(mem[736]) );
  DFFPOSX1 mem_reg_17__38_ ( .D(n2577), .CLK(clk), .Q(mem[735]) );
  DFFPOSX1 mem_reg_17__37_ ( .D(n2576), .CLK(clk), .Q(mem[734]) );
  DFFPOSX1 mem_reg_17__36_ ( .D(n2575), .CLK(clk), .Q(mem[733]) );
  DFFPOSX1 mem_reg_17__35_ ( .D(n2574), .CLK(clk), .Q(mem[732]) );
  DFFPOSX1 mem_reg_17__34_ ( .D(n2573), .CLK(clk), .Q(mem[731]) );
  DFFPOSX1 mem_reg_17__33_ ( .D(n2572), .CLK(clk), .Q(mem[730]) );
  DFFPOSX1 mem_reg_17__32_ ( .D(n2571), .CLK(clk), .Q(mem[729]) );
  DFFPOSX1 mem_reg_17__31_ ( .D(n2570), .CLK(clk), .Q(mem[728]) );
  DFFPOSX1 mem_reg_17__30_ ( .D(n2569), .CLK(clk), .Q(mem[727]) );
  DFFPOSX1 mem_reg_17__29_ ( .D(n2568), .CLK(clk), .Q(mem[726]) );
  DFFPOSX1 mem_reg_17__28_ ( .D(n2567), .CLK(clk), .Q(mem[725]) );
  DFFPOSX1 mem_reg_17__27_ ( .D(n2566), .CLK(clk), .Q(mem[724]) );
  DFFPOSX1 mem_reg_17__26_ ( .D(n2565), .CLK(clk), .Q(mem[723]) );
  DFFPOSX1 mem_reg_17__25_ ( .D(n2564), .CLK(clk), .Q(mem[722]) );
  DFFPOSX1 mem_reg_17__24_ ( .D(n2563), .CLK(clk), .Q(mem[721]) );
  DFFPOSX1 mem_reg_17__23_ ( .D(n2562), .CLK(clk), .Q(mem[720]) );
  DFFPOSX1 mem_reg_17__22_ ( .D(n2561), .CLK(clk), .Q(mem[719]) );
  DFFPOSX1 mem_reg_17__21_ ( .D(n2560), .CLK(clk), .Q(mem[718]) );
  DFFPOSX1 mem_reg_17__20_ ( .D(n2559), .CLK(clk), .Q(mem[717]) );
  DFFPOSX1 mem_reg_17__19_ ( .D(n2558), .CLK(clk), .Q(mem[716]) );
  DFFPOSX1 mem_reg_17__18_ ( .D(n2557), .CLK(clk), .Q(mem[715]) );
  DFFPOSX1 mem_reg_17__17_ ( .D(n2556), .CLK(clk), .Q(mem[714]) );
  DFFPOSX1 mem_reg_17__16_ ( .D(n2555), .CLK(clk), .Q(mem[713]) );
  DFFPOSX1 mem_reg_17__15_ ( .D(n2554), .CLK(clk), .Q(mem[712]) );
  DFFPOSX1 mem_reg_17__14_ ( .D(n2553), .CLK(clk), .Q(mem[711]) );
  DFFPOSX1 mem_reg_17__13_ ( .D(n2552), .CLK(clk), .Q(mem[710]) );
  DFFPOSX1 mem_reg_17__12_ ( .D(n2551), .CLK(clk), .Q(mem[709]) );
  DFFPOSX1 mem_reg_17__11_ ( .D(n2550), .CLK(clk), .Q(mem[708]) );
  DFFPOSX1 mem_reg_17__10_ ( .D(n2549), .CLK(clk), .Q(mem[707]) );
  DFFPOSX1 mem_reg_17__9_ ( .D(n2548), .CLK(clk), .Q(mem[706]) );
  DFFPOSX1 mem_reg_17__8_ ( .D(n2547), .CLK(clk), .Q(mem[705]) );
  DFFPOSX1 mem_reg_17__7_ ( .D(n2546), .CLK(clk), .Q(mem[704]) );
  DFFPOSX1 mem_reg_17__6_ ( .D(n2545), .CLK(clk), .Q(mem[703]) );
  DFFPOSX1 mem_reg_17__5_ ( .D(n2544), .CLK(clk), .Q(mem[702]) );
  DFFPOSX1 mem_reg_17__4_ ( .D(n2543), .CLK(clk), .Q(mem[701]) );
  DFFPOSX1 mem_reg_17__3_ ( .D(n2542), .CLK(clk), .Q(mem[700]) );
  DFFPOSX1 mem_reg_17__2_ ( .D(n2541), .CLK(clk), .Q(mem[699]) );
  DFFPOSX1 mem_reg_17__1_ ( .D(n2540), .CLK(clk), .Q(mem[698]) );
  DFFPOSX1 mem_reg_17__0_ ( .D(n2539), .CLK(clk), .Q(mem[697]) );
  DFFPOSX1 mem_reg_16__40_ ( .D(n2538), .CLK(clk), .Q(mem[696]) );
  DFFPOSX1 mem_reg_16__39_ ( .D(n2537), .CLK(clk), .Q(mem[695]) );
  DFFPOSX1 mem_reg_16__38_ ( .D(n2536), .CLK(clk), .Q(mem[694]) );
  DFFPOSX1 mem_reg_16__37_ ( .D(n2535), .CLK(clk), .Q(mem[693]) );
  DFFPOSX1 mem_reg_16__36_ ( .D(n2534), .CLK(clk), .Q(mem[692]) );
  DFFPOSX1 mem_reg_16__35_ ( .D(n2533), .CLK(clk), .Q(mem[691]) );
  DFFPOSX1 mem_reg_16__34_ ( .D(n2532), .CLK(clk), .Q(mem[690]) );
  DFFPOSX1 mem_reg_16__33_ ( .D(n2531), .CLK(clk), .Q(mem[689]) );
  DFFPOSX1 mem_reg_16__32_ ( .D(n2530), .CLK(clk), .Q(mem[688]) );
  DFFPOSX1 mem_reg_16__31_ ( .D(n2529), .CLK(clk), .Q(mem[687]) );
  DFFPOSX1 mem_reg_16__30_ ( .D(n2528), .CLK(clk), .Q(mem[686]) );
  DFFPOSX1 mem_reg_16__29_ ( .D(n2527), .CLK(clk), .Q(mem[685]) );
  DFFPOSX1 mem_reg_16__28_ ( .D(n2526), .CLK(clk), .Q(mem[684]) );
  DFFPOSX1 mem_reg_16__27_ ( .D(n2525), .CLK(clk), .Q(mem[683]) );
  DFFPOSX1 mem_reg_16__26_ ( .D(n2524), .CLK(clk), .Q(mem[682]) );
  DFFPOSX1 mem_reg_16__25_ ( .D(n2523), .CLK(clk), .Q(mem[681]) );
  DFFPOSX1 mem_reg_16__24_ ( .D(n2522), .CLK(clk), .Q(mem[680]) );
  DFFPOSX1 mem_reg_16__23_ ( .D(n2521), .CLK(clk), .Q(mem[679]) );
  DFFPOSX1 mem_reg_16__22_ ( .D(n2520), .CLK(clk), .Q(mem[678]) );
  DFFPOSX1 mem_reg_16__21_ ( .D(n2519), .CLK(clk), .Q(mem[677]) );
  DFFPOSX1 mem_reg_16__20_ ( .D(n2518), .CLK(clk), .Q(mem[676]) );
  DFFPOSX1 mem_reg_16__19_ ( .D(n2517), .CLK(clk), .Q(mem[675]) );
  DFFPOSX1 mem_reg_16__18_ ( .D(n2516), .CLK(clk), .Q(mem[674]) );
  DFFPOSX1 mem_reg_16__17_ ( .D(n2515), .CLK(clk), .Q(mem[673]) );
  DFFPOSX1 mem_reg_16__16_ ( .D(n2514), .CLK(clk), .Q(mem[672]) );
  DFFPOSX1 mem_reg_16__15_ ( .D(n2513), .CLK(clk), .Q(mem[671]) );
  DFFPOSX1 mem_reg_16__14_ ( .D(n2512), .CLK(clk), .Q(mem[670]) );
  DFFPOSX1 mem_reg_16__13_ ( .D(n2511), .CLK(clk), .Q(mem[669]) );
  DFFPOSX1 mem_reg_16__12_ ( .D(n2510), .CLK(clk), .Q(mem[668]) );
  DFFPOSX1 mem_reg_16__11_ ( .D(n2509), .CLK(clk), .Q(mem[667]) );
  DFFPOSX1 mem_reg_16__10_ ( .D(n2508), .CLK(clk), .Q(mem[666]) );
  DFFPOSX1 mem_reg_16__9_ ( .D(n2507), .CLK(clk), .Q(mem[665]) );
  DFFPOSX1 mem_reg_16__8_ ( .D(n2506), .CLK(clk), .Q(mem[664]) );
  DFFPOSX1 mem_reg_16__7_ ( .D(n2505), .CLK(clk), .Q(mem[663]) );
  DFFPOSX1 mem_reg_16__6_ ( .D(n2504), .CLK(clk), .Q(mem[662]) );
  DFFPOSX1 mem_reg_16__5_ ( .D(n2503), .CLK(clk), .Q(mem[661]) );
  DFFPOSX1 mem_reg_16__4_ ( .D(n2502), .CLK(clk), .Q(mem[660]) );
  DFFPOSX1 mem_reg_16__3_ ( .D(n2501), .CLK(clk), .Q(mem[659]) );
  DFFPOSX1 mem_reg_16__2_ ( .D(n2500), .CLK(clk), .Q(mem[658]) );
  DFFPOSX1 mem_reg_16__1_ ( .D(n2499), .CLK(clk), .Q(mem[657]) );
  DFFPOSX1 mem_reg_16__0_ ( .D(n2498), .CLK(clk), .Q(mem[656]) );
  DFFPOSX1 mem_reg_15__40_ ( .D(n2497), .CLK(clk), .Q(mem[655]) );
  DFFPOSX1 mem_reg_15__39_ ( .D(n2496), .CLK(clk), .Q(mem[654]) );
  DFFPOSX1 mem_reg_15__38_ ( .D(n2495), .CLK(clk), .Q(mem[653]) );
  DFFPOSX1 mem_reg_15__37_ ( .D(n2494), .CLK(clk), .Q(mem[652]) );
  DFFPOSX1 mem_reg_15__36_ ( .D(n2493), .CLK(clk), .Q(mem[651]) );
  DFFPOSX1 mem_reg_15__35_ ( .D(n2492), .CLK(clk), .Q(mem[650]) );
  DFFPOSX1 mem_reg_15__34_ ( .D(n2491), .CLK(clk), .Q(mem[649]) );
  DFFPOSX1 mem_reg_15__33_ ( .D(n2490), .CLK(clk), .Q(mem[648]) );
  DFFPOSX1 mem_reg_15__32_ ( .D(n2489), .CLK(clk), .Q(mem[647]) );
  DFFPOSX1 mem_reg_15__31_ ( .D(n2488), .CLK(clk), .Q(mem[646]) );
  DFFPOSX1 mem_reg_15__30_ ( .D(n2487), .CLK(clk), .Q(mem[645]) );
  DFFPOSX1 mem_reg_15__29_ ( .D(n2486), .CLK(clk), .Q(mem[644]) );
  DFFPOSX1 mem_reg_15__28_ ( .D(n2485), .CLK(clk), .Q(mem[643]) );
  DFFPOSX1 mem_reg_15__27_ ( .D(n2484), .CLK(clk), .Q(mem[642]) );
  DFFPOSX1 mem_reg_15__26_ ( .D(n2483), .CLK(clk), .Q(mem[641]) );
  DFFPOSX1 mem_reg_15__25_ ( .D(n2482), .CLK(clk), .Q(mem[640]) );
  DFFPOSX1 mem_reg_15__24_ ( .D(n2481), .CLK(clk), .Q(mem[639]) );
  DFFPOSX1 mem_reg_15__23_ ( .D(n2480), .CLK(clk), .Q(mem[638]) );
  DFFPOSX1 mem_reg_15__22_ ( .D(n2479), .CLK(clk), .Q(mem[637]) );
  DFFPOSX1 mem_reg_15__21_ ( .D(n2478), .CLK(clk), .Q(mem[636]) );
  DFFPOSX1 mem_reg_15__20_ ( .D(n2477), .CLK(clk), .Q(mem[635]) );
  DFFPOSX1 mem_reg_15__19_ ( .D(n2476), .CLK(clk), .Q(mem[634]) );
  DFFPOSX1 mem_reg_15__18_ ( .D(n2475), .CLK(clk), .Q(mem[633]) );
  DFFPOSX1 mem_reg_15__17_ ( .D(n2474), .CLK(clk), .Q(mem[632]) );
  DFFPOSX1 mem_reg_15__16_ ( .D(n2473), .CLK(clk), .Q(mem[631]) );
  DFFPOSX1 mem_reg_15__15_ ( .D(n2472), .CLK(clk), .Q(mem[630]) );
  DFFPOSX1 mem_reg_15__14_ ( .D(n2471), .CLK(clk), .Q(mem[629]) );
  DFFPOSX1 mem_reg_15__13_ ( .D(n2470), .CLK(clk), .Q(mem[628]) );
  DFFPOSX1 mem_reg_15__12_ ( .D(n2469), .CLK(clk), .Q(mem[627]) );
  DFFPOSX1 mem_reg_15__11_ ( .D(n2468), .CLK(clk), .Q(mem[626]) );
  DFFPOSX1 mem_reg_15__10_ ( .D(n2467), .CLK(clk), .Q(mem[625]) );
  DFFPOSX1 mem_reg_15__9_ ( .D(n2466), .CLK(clk), .Q(mem[624]) );
  DFFPOSX1 mem_reg_15__8_ ( .D(n2465), .CLK(clk), .Q(mem[623]) );
  DFFPOSX1 mem_reg_15__7_ ( .D(n2464), .CLK(clk), .Q(mem[622]) );
  DFFPOSX1 mem_reg_15__6_ ( .D(n2463), .CLK(clk), .Q(mem[621]) );
  DFFPOSX1 mem_reg_15__5_ ( .D(n2462), .CLK(clk), .Q(mem[620]) );
  DFFPOSX1 mem_reg_15__4_ ( .D(n2461), .CLK(clk), .Q(mem[619]) );
  DFFPOSX1 mem_reg_15__3_ ( .D(n2460), .CLK(clk), .Q(mem[618]) );
  DFFPOSX1 mem_reg_15__2_ ( .D(n2459), .CLK(clk), .Q(mem[617]) );
  DFFPOSX1 mem_reg_15__1_ ( .D(n2458), .CLK(clk), .Q(mem[616]) );
  DFFPOSX1 mem_reg_15__0_ ( .D(n2457), .CLK(clk), .Q(mem[615]) );
  DFFPOSX1 mem_reg_14__40_ ( .D(n2456), .CLK(clk), .Q(mem[614]) );
  DFFPOSX1 mem_reg_14__39_ ( .D(n2455), .CLK(clk), .Q(mem[613]) );
  DFFPOSX1 mem_reg_14__38_ ( .D(n2454), .CLK(clk), .Q(mem[612]) );
  DFFPOSX1 mem_reg_14__37_ ( .D(n2453), .CLK(clk), .Q(mem[611]) );
  DFFPOSX1 mem_reg_14__36_ ( .D(n2452), .CLK(clk), .Q(mem[610]) );
  DFFPOSX1 mem_reg_14__35_ ( .D(n2451), .CLK(clk), .Q(mem[609]) );
  DFFPOSX1 mem_reg_14__34_ ( .D(n2450), .CLK(clk), .Q(mem[608]) );
  DFFPOSX1 mem_reg_14__33_ ( .D(n2449), .CLK(clk), .Q(mem[607]) );
  DFFPOSX1 mem_reg_14__32_ ( .D(n2448), .CLK(clk), .Q(mem[606]) );
  DFFPOSX1 mem_reg_14__31_ ( .D(n2447), .CLK(clk), .Q(mem[605]) );
  DFFPOSX1 mem_reg_14__30_ ( .D(n2446), .CLK(clk), .Q(mem[604]) );
  DFFPOSX1 mem_reg_14__29_ ( .D(n2445), .CLK(clk), .Q(mem[603]) );
  DFFPOSX1 mem_reg_14__28_ ( .D(n2444), .CLK(clk), .Q(mem[602]) );
  DFFPOSX1 mem_reg_14__27_ ( .D(n2443), .CLK(clk), .Q(mem[601]) );
  DFFPOSX1 mem_reg_14__26_ ( .D(n2442), .CLK(clk), .Q(mem[600]) );
  DFFPOSX1 mem_reg_14__25_ ( .D(n2441), .CLK(clk), .Q(mem[599]) );
  DFFPOSX1 mem_reg_14__24_ ( .D(n2440), .CLK(clk), .Q(mem[598]) );
  DFFPOSX1 mem_reg_14__23_ ( .D(n2439), .CLK(clk), .Q(mem[597]) );
  DFFPOSX1 mem_reg_14__22_ ( .D(n2438), .CLK(clk), .Q(mem[596]) );
  DFFPOSX1 mem_reg_14__21_ ( .D(n2437), .CLK(clk), .Q(mem[595]) );
  DFFPOSX1 mem_reg_14__20_ ( .D(n2436), .CLK(clk), .Q(mem[594]) );
  DFFPOSX1 mem_reg_14__19_ ( .D(n2435), .CLK(clk), .Q(mem[593]) );
  DFFPOSX1 mem_reg_14__18_ ( .D(n2434), .CLK(clk), .Q(mem[592]) );
  DFFPOSX1 mem_reg_14__17_ ( .D(n2433), .CLK(clk), .Q(mem[591]) );
  DFFPOSX1 mem_reg_14__16_ ( .D(n2432), .CLK(clk), .Q(mem[590]) );
  DFFPOSX1 mem_reg_14__15_ ( .D(n2431), .CLK(clk), .Q(mem[589]) );
  DFFPOSX1 mem_reg_14__14_ ( .D(n2430), .CLK(clk), .Q(mem[588]) );
  DFFPOSX1 mem_reg_14__13_ ( .D(n2429), .CLK(clk), .Q(mem[587]) );
  DFFPOSX1 mem_reg_14__12_ ( .D(n2428), .CLK(clk), .Q(mem[586]) );
  DFFPOSX1 mem_reg_14__11_ ( .D(n2427), .CLK(clk), .Q(mem[585]) );
  DFFPOSX1 mem_reg_14__10_ ( .D(n2426), .CLK(clk), .Q(mem[584]) );
  DFFPOSX1 mem_reg_14__9_ ( .D(n2425), .CLK(clk), .Q(mem[583]) );
  DFFPOSX1 mem_reg_14__8_ ( .D(n2424), .CLK(clk), .Q(mem[582]) );
  DFFPOSX1 mem_reg_14__7_ ( .D(n2423), .CLK(clk), .Q(mem[581]) );
  DFFPOSX1 mem_reg_14__6_ ( .D(n2422), .CLK(clk), .Q(mem[580]) );
  DFFPOSX1 mem_reg_14__5_ ( .D(n2421), .CLK(clk), .Q(mem[579]) );
  DFFPOSX1 mem_reg_14__4_ ( .D(n2420), .CLK(clk), .Q(mem[578]) );
  DFFPOSX1 mem_reg_14__3_ ( .D(n2419), .CLK(clk), .Q(mem[577]) );
  DFFPOSX1 mem_reg_14__2_ ( .D(n2418), .CLK(clk), .Q(mem[576]) );
  DFFPOSX1 mem_reg_14__1_ ( .D(n2417), .CLK(clk), .Q(mem[575]) );
  DFFPOSX1 mem_reg_14__0_ ( .D(n2416), .CLK(clk), .Q(mem[574]) );
  DFFPOSX1 mem_reg_13__40_ ( .D(n2415), .CLK(clk), .Q(mem[573]) );
  DFFPOSX1 mem_reg_13__39_ ( .D(n2414), .CLK(clk), .Q(mem[572]) );
  DFFPOSX1 mem_reg_13__38_ ( .D(n2413), .CLK(clk), .Q(mem[571]) );
  DFFPOSX1 mem_reg_13__37_ ( .D(n2412), .CLK(clk), .Q(mem[570]) );
  DFFPOSX1 mem_reg_13__36_ ( .D(n2411), .CLK(clk), .Q(mem[569]) );
  DFFPOSX1 mem_reg_13__35_ ( .D(n2410), .CLK(clk), .Q(mem[568]) );
  DFFPOSX1 mem_reg_13__34_ ( .D(n2409), .CLK(clk), .Q(mem[567]) );
  DFFPOSX1 mem_reg_13__33_ ( .D(n2408), .CLK(clk), .Q(mem[566]) );
  DFFPOSX1 mem_reg_13__32_ ( .D(n2407), .CLK(clk), .Q(mem[565]) );
  DFFPOSX1 mem_reg_13__31_ ( .D(n2406), .CLK(clk), .Q(mem[564]) );
  DFFPOSX1 mem_reg_13__30_ ( .D(n2405), .CLK(clk), .Q(mem[563]) );
  DFFPOSX1 mem_reg_13__29_ ( .D(n2404), .CLK(clk), .Q(mem[562]) );
  DFFPOSX1 mem_reg_13__28_ ( .D(n2403), .CLK(clk), .Q(mem[561]) );
  DFFPOSX1 mem_reg_13__27_ ( .D(n2402), .CLK(clk), .Q(mem[560]) );
  DFFPOSX1 mem_reg_13__26_ ( .D(n2401), .CLK(clk), .Q(mem[559]) );
  DFFPOSX1 mem_reg_13__25_ ( .D(n2400), .CLK(clk), .Q(mem[558]) );
  DFFPOSX1 mem_reg_13__24_ ( .D(n2399), .CLK(clk), .Q(mem[557]) );
  DFFPOSX1 mem_reg_13__23_ ( .D(n2398), .CLK(clk), .Q(mem[556]) );
  DFFPOSX1 mem_reg_13__22_ ( .D(n2397), .CLK(clk), .Q(mem[555]) );
  DFFPOSX1 mem_reg_13__21_ ( .D(n2396), .CLK(clk), .Q(mem[554]) );
  DFFPOSX1 mem_reg_13__20_ ( .D(n2395), .CLK(clk), .Q(mem[553]) );
  DFFPOSX1 mem_reg_13__19_ ( .D(n2394), .CLK(clk), .Q(mem[552]) );
  DFFPOSX1 mem_reg_13__18_ ( .D(n2393), .CLK(clk), .Q(mem[551]) );
  DFFPOSX1 mem_reg_13__17_ ( .D(n2392), .CLK(clk), .Q(mem[550]) );
  DFFPOSX1 mem_reg_13__16_ ( .D(n2391), .CLK(clk), .Q(mem[549]) );
  DFFPOSX1 mem_reg_13__15_ ( .D(n2390), .CLK(clk), .Q(mem[548]) );
  DFFPOSX1 mem_reg_13__14_ ( .D(n2389), .CLK(clk), .Q(mem[547]) );
  DFFPOSX1 mem_reg_13__13_ ( .D(n2388), .CLK(clk), .Q(mem[546]) );
  DFFPOSX1 mem_reg_13__12_ ( .D(n2387), .CLK(clk), .Q(mem[545]) );
  DFFPOSX1 mem_reg_13__11_ ( .D(n2386), .CLK(clk), .Q(mem[544]) );
  DFFPOSX1 mem_reg_13__10_ ( .D(n2385), .CLK(clk), .Q(mem[543]) );
  DFFPOSX1 mem_reg_13__9_ ( .D(n2384), .CLK(clk), .Q(mem[542]) );
  DFFPOSX1 mem_reg_13__8_ ( .D(n2383), .CLK(clk), .Q(mem[541]) );
  DFFPOSX1 mem_reg_13__7_ ( .D(n2382), .CLK(clk), .Q(mem[540]) );
  DFFPOSX1 mem_reg_13__6_ ( .D(n2381), .CLK(clk), .Q(mem[539]) );
  DFFPOSX1 mem_reg_13__5_ ( .D(n2380), .CLK(clk), .Q(mem[538]) );
  DFFPOSX1 mem_reg_13__4_ ( .D(n2379), .CLK(clk), .Q(mem[537]) );
  DFFPOSX1 mem_reg_13__3_ ( .D(n2378), .CLK(clk), .Q(mem[536]) );
  DFFPOSX1 mem_reg_13__2_ ( .D(n2377), .CLK(clk), .Q(mem[535]) );
  DFFPOSX1 mem_reg_13__1_ ( .D(n2376), .CLK(clk), .Q(mem[534]) );
  DFFPOSX1 mem_reg_13__0_ ( .D(n2375), .CLK(clk), .Q(mem[533]) );
  DFFPOSX1 mem_reg_12__40_ ( .D(n2374), .CLK(clk), .Q(mem[532]) );
  DFFPOSX1 mem_reg_12__39_ ( .D(n2373), .CLK(clk), .Q(mem[531]) );
  DFFPOSX1 mem_reg_12__38_ ( .D(n2372), .CLK(clk), .Q(mem[530]) );
  DFFPOSX1 mem_reg_12__37_ ( .D(n2371), .CLK(clk), .Q(mem[529]) );
  DFFPOSX1 mem_reg_12__36_ ( .D(n2370), .CLK(clk), .Q(mem[528]) );
  DFFPOSX1 mem_reg_12__35_ ( .D(n2369), .CLK(clk), .Q(mem[527]) );
  DFFPOSX1 mem_reg_12__34_ ( .D(n2368), .CLK(clk), .Q(mem[526]) );
  DFFPOSX1 mem_reg_12__33_ ( .D(n2367), .CLK(clk), .Q(mem[525]) );
  DFFPOSX1 mem_reg_12__32_ ( .D(n2366), .CLK(clk), .Q(mem[524]) );
  DFFPOSX1 mem_reg_12__31_ ( .D(n2365), .CLK(clk), .Q(mem[523]) );
  DFFPOSX1 mem_reg_12__30_ ( .D(n2364), .CLK(clk), .Q(mem[522]) );
  DFFPOSX1 mem_reg_12__29_ ( .D(n2363), .CLK(clk), .Q(mem[521]) );
  DFFPOSX1 mem_reg_12__28_ ( .D(n2362), .CLK(clk), .Q(mem[520]) );
  DFFPOSX1 mem_reg_12__27_ ( .D(n2361), .CLK(clk), .Q(mem[519]) );
  DFFPOSX1 mem_reg_12__26_ ( .D(n2360), .CLK(clk), .Q(mem[518]) );
  DFFPOSX1 mem_reg_12__25_ ( .D(n2359), .CLK(clk), .Q(mem[517]) );
  DFFPOSX1 mem_reg_12__24_ ( .D(n2358), .CLK(clk), .Q(mem[516]) );
  DFFPOSX1 mem_reg_12__23_ ( .D(n2357), .CLK(clk), .Q(mem[515]) );
  DFFPOSX1 mem_reg_12__22_ ( .D(n2356), .CLK(clk), .Q(mem[514]) );
  DFFPOSX1 mem_reg_12__21_ ( .D(n2355), .CLK(clk), .Q(mem[513]) );
  DFFPOSX1 mem_reg_12__20_ ( .D(n2354), .CLK(clk), .Q(mem[512]) );
  DFFPOSX1 mem_reg_12__19_ ( .D(n2353), .CLK(clk), .Q(mem[511]) );
  DFFPOSX1 mem_reg_12__18_ ( .D(n2352), .CLK(clk), .Q(mem[510]) );
  DFFPOSX1 mem_reg_12__17_ ( .D(n2351), .CLK(clk), .Q(mem[509]) );
  DFFPOSX1 mem_reg_12__16_ ( .D(n2350), .CLK(clk), .Q(mem[508]) );
  DFFPOSX1 mem_reg_12__15_ ( .D(n2349), .CLK(clk), .Q(mem[507]) );
  DFFPOSX1 mem_reg_12__14_ ( .D(n2348), .CLK(clk), .Q(mem[506]) );
  DFFPOSX1 mem_reg_12__13_ ( .D(n2347), .CLK(clk), .Q(mem[505]) );
  DFFPOSX1 mem_reg_12__12_ ( .D(n2346), .CLK(clk), .Q(mem[504]) );
  DFFPOSX1 mem_reg_12__11_ ( .D(n2345), .CLK(clk), .Q(mem[503]) );
  DFFPOSX1 mem_reg_12__10_ ( .D(n2344), .CLK(clk), .Q(mem[502]) );
  DFFPOSX1 mem_reg_12__9_ ( .D(n2343), .CLK(clk), .Q(mem[501]) );
  DFFPOSX1 mem_reg_12__8_ ( .D(n2342), .CLK(clk), .Q(mem[500]) );
  DFFPOSX1 mem_reg_12__7_ ( .D(n2341), .CLK(clk), .Q(mem[499]) );
  DFFPOSX1 mem_reg_12__6_ ( .D(n2340), .CLK(clk), .Q(mem[498]) );
  DFFPOSX1 mem_reg_12__5_ ( .D(n2339), .CLK(clk), .Q(mem[497]) );
  DFFPOSX1 mem_reg_12__4_ ( .D(n2338), .CLK(clk), .Q(mem[496]) );
  DFFPOSX1 mem_reg_12__3_ ( .D(n2337), .CLK(clk), .Q(mem[495]) );
  DFFPOSX1 mem_reg_12__2_ ( .D(n2336), .CLK(clk), .Q(mem[494]) );
  DFFPOSX1 mem_reg_12__1_ ( .D(n2335), .CLK(clk), .Q(mem[493]) );
  DFFPOSX1 mem_reg_12__0_ ( .D(n2334), .CLK(clk), .Q(mem[492]) );
  DFFPOSX1 mem_reg_11__40_ ( .D(n2333), .CLK(clk), .Q(mem[491]) );
  DFFPOSX1 mem_reg_11__39_ ( .D(n2332), .CLK(clk), .Q(mem[490]) );
  DFFPOSX1 mem_reg_11__38_ ( .D(n2331), .CLK(clk), .Q(mem[489]) );
  DFFPOSX1 mem_reg_11__37_ ( .D(n2330), .CLK(clk), .Q(mem[488]) );
  DFFPOSX1 mem_reg_11__36_ ( .D(n2329), .CLK(clk), .Q(mem[487]) );
  DFFPOSX1 mem_reg_11__35_ ( .D(n2328), .CLK(clk), .Q(mem[486]) );
  DFFPOSX1 mem_reg_11__34_ ( .D(n2327), .CLK(clk), .Q(mem[485]) );
  DFFPOSX1 mem_reg_11__33_ ( .D(n2326), .CLK(clk), .Q(mem[484]) );
  DFFPOSX1 mem_reg_11__32_ ( .D(n2325), .CLK(clk), .Q(mem[483]) );
  DFFPOSX1 mem_reg_11__31_ ( .D(n2324), .CLK(clk), .Q(mem[482]) );
  DFFPOSX1 mem_reg_11__30_ ( .D(n2323), .CLK(clk), .Q(mem[481]) );
  DFFPOSX1 mem_reg_11__29_ ( .D(n2322), .CLK(clk), .Q(mem[480]) );
  DFFPOSX1 mem_reg_11__28_ ( .D(n2321), .CLK(clk), .Q(mem[479]) );
  DFFPOSX1 mem_reg_11__27_ ( .D(n2320), .CLK(clk), .Q(mem[478]) );
  DFFPOSX1 mem_reg_11__26_ ( .D(n2319), .CLK(clk), .Q(mem[477]) );
  DFFPOSX1 mem_reg_11__25_ ( .D(n2318), .CLK(clk), .Q(mem[476]) );
  DFFPOSX1 mem_reg_11__24_ ( .D(n2317), .CLK(clk), .Q(mem[475]) );
  DFFPOSX1 mem_reg_11__23_ ( .D(n2316), .CLK(clk), .Q(mem[474]) );
  DFFPOSX1 mem_reg_11__22_ ( .D(n2315), .CLK(clk), .Q(mem[473]) );
  DFFPOSX1 mem_reg_11__21_ ( .D(n2314), .CLK(clk), .Q(mem[472]) );
  DFFPOSX1 mem_reg_11__20_ ( .D(n2313), .CLK(clk), .Q(mem[471]) );
  DFFPOSX1 mem_reg_11__19_ ( .D(n2312), .CLK(clk), .Q(mem[470]) );
  DFFPOSX1 mem_reg_11__18_ ( .D(n2311), .CLK(clk), .Q(mem[469]) );
  DFFPOSX1 mem_reg_11__17_ ( .D(n2310), .CLK(clk), .Q(mem[468]) );
  DFFPOSX1 mem_reg_11__16_ ( .D(n2309), .CLK(clk), .Q(mem[467]) );
  DFFPOSX1 mem_reg_11__15_ ( .D(n2308), .CLK(clk), .Q(mem[466]) );
  DFFPOSX1 mem_reg_11__14_ ( .D(n2307), .CLK(clk), .Q(mem[465]) );
  DFFPOSX1 mem_reg_11__13_ ( .D(n2306), .CLK(clk), .Q(mem[464]) );
  DFFPOSX1 mem_reg_11__12_ ( .D(n2305), .CLK(clk), .Q(mem[463]) );
  DFFPOSX1 mem_reg_11__11_ ( .D(n2304), .CLK(clk), .Q(mem[462]) );
  DFFPOSX1 mem_reg_11__10_ ( .D(n2303), .CLK(clk), .Q(mem[461]) );
  DFFPOSX1 mem_reg_11__9_ ( .D(n2302), .CLK(clk), .Q(mem[460]) );
  DFFPOSX1 mem_reg_11__8_ ( .D(n2301), .CLK(clk), .Q(mem[459]) );
  DFFPOSX1 mem_reg_11__7_ ( .D(n2300), .CLK(clk), .Q(mem[458]) );
  DFFPOSX1 mem_reg_11__6_ ( .D(n2299), .CLK(clk), .Q(mem[457]) );
  DFFPOSX1 mem_reg_11__5_ ( .D(n2298), .CLK(clk), .Q(mem[456]) );
  DFFPOSX1 mem_reg_11__4_ ( .D(n2297), .CLK(clk), .Q(mem[455]) );
  DFFPOSX1 mem_reg_11__3_ ( .D(n2296), .CLK(clk), .Q(mem[454]) );
  DFFPOSX1 mem_reg_11__2_ ( .D(n2295), .CLK(clk), .Q(mem[453]) );
  DFFPOSX1 mem_reg_11__1_ ( .D(n2294), .CLK(clk), .Q(mem[452]) );
  DFFPOSX1 mem_reg_11__0_ ( .D(n2293), .CLK(clk), .Q(mem[451]) );
  DFFPOSX1 mem_reg_10__40_ ( .D(n2292), .CLK(clk), .Q(mem[450]) );
  DFFPOSX1 mem_reg_10__39_ ( .D(n2291), .CLK(clk), .Q(mem[449]) );
  DFFPOSX1 mem_reg_10__38_ ( .D(n2290), .CLK(clk), .Q(mem[448]) );
  DFFPOSX1 mem_reg_10__37_ ( .D(n2289), .CLK(clk), .Q(mem[447]) );
  DFFPOSX1 mem_reg_10__36_ ( .D(n2288), .CLK(clk), .Q(mem[446]) );
  DFFPOSX1 mem_reg_10__35_ ( .D(n2287), .CLK(clk), .Q(mem[445]) );
  DFFPOSX1 mem_reg_10__34_ ( .D(n2286), .CLK(clk), .Q(mem[444]) );
  DFFPOSX1 mem_reg_10__33_ ( .D(n2285), .CLK(clk), .Q(mem[443]) );
  DFFPOSX1 mem_reg_10__32_ ( .D(n2284), .CLK(clk), .Q(mem[442]) );
  DFFPOSX1 mem_reg_10__31_ ( .D(n2283), .CLK(clk), .Q(mem[441]) );
  DFFPOSX1 mem_reg_10__30_ ( .D(n2282), .CLK(clk), .Q(mem[440]) );
  DFFPOSX1 mem_reg_10__29_ ( .D(n2281), .CLK(clk), .Q(mem[439]) );
  DFFPOSX1 mem_reg_10__28_ ( .D(n2280), .CLK(clk), .Q(mem[438]) );
  DFFPOSX1 mem_reg_10__27_ ( .D(n2279), .CLK(clk), .Q(mem[437]) );
  DFFPOSX1 mem_reg_10__26_ ( .D(n2278), .CLK(clk), .Q(mem[436]) );
  DFFPOSX1 mem_reg_10__25_ ( .D(n2277), .CLK(clk), .Q(mem[435]) );
  DFFPOSX1 mem_reg_10__24_ ( .D(n2276), .CLK(clk), .Q(mem[434]) );
  DFFPOSX1 mem_reg_10__23_ ( .D(n2275), .CLK(clk), .Q(mem[433]) );
  DFFPOSX1 mem_reg_10__22_ ( .D(n2274), .CLK(clk), .Q(mem[432]) );
  DFFPOSX1 mem_reg_10__21_ ( .D(n2273), .CLK(clk), .Q(mem[431]) );
  DFFPOSX1 mem_reg_10__20_ ( .D(n2272), .CLK(clk), .Q(mem[430]) );
  DFFPOSX1 mem_reg_10__19_ ( .D(n2271), .CLK(clk), .Q(mem[429]) );
  DFFPOSX1 mem_reg_10__18_ ( .D(n2270), .CLK(clk), .Q(mem[428]) );
  DFFPOSX1 mem_reg_10__17_ ( .D(n2269), .CLK(clk), .Q(mem[427]) );
  DFFPOSX1 mem_reg_10__16_ ( .D(n2268), .CLK(clk), .Q(mem[426]) );
  DFFPOSX1 mem_reg_10__15_ ( .D(n2267), .CLK(clk), .Q(mem[425]) );
  DFFPOSX1 mem_reg_10__14_ ( .D(n2266), .CLK(clk), .Q(mem[424]) );
  DFFPOSX1 mem_reg_10__13_ ( .D(n2265), .CLK(clk), .Q(mem[423]) );
  DFFPOSX1 mem_reg_10__12_ ( .D(n2264), .CLK(clk), .Q(mem[422]) );
  DFFPOSX1 mem_reg_10__11_ ( .D(n2263), .CLK(clk), .Q(mem[421]) );
  DFFPOSX1 mem_reg_10__10_ ( .D(n2262), .CLK(clk), .Q(mem[420]) );
  DFFPOSX1 mem_reg_10__9_ ( .D(n2261), .CLK(clk), .Q(mem[419]) );
  DFFPOSX1 mem_reg_10__8_ ( .D(n2260), .CLK(clk), .Q(mem[418]) );
  DFFPOSX1 mem_reg_10__7_ ( .D(n2259), .CLK(clk), .Q(mem[417]) );
  DFFPOSX1 mem_reg_10__6_ ( .D(n2258), .CLK(clk), .Q(mem[416]) );
  DFFPOSX1 mem_reg_10__5_ ( .D(n2257), .CLK(clk), .Q(mem[415]) );
  DFFPOSX1 mem_reg_10__4_ ( .D(n2256), .CLK(clk), .Q(mem[414]) );
  DFFPOSX1 mem_reg_10__3_ ( .D(n2255), .CLK(clk), .Q(mem[413]) );
  DFFPOSX1 mem_reg_10__2_ ( .D(n2254), .CLK(clk), .Q(mem[412]) );
  DFFPOSX1 mem_reg_10__1_ ( .D(n2253), .CLK(clk), .Q(mem[411]) );
  DFFPOSX1 mem_reg_10__0_ ( .D(n2252), .CLK(clk), .Q(mem[410]) );
  DFFPOSX1 mem_reg_9__40_ ( .D(n2251), .CLK(clk), .Q(mem[409]) );
  DFFPOSX1 mem_reg_9__39_ ( .D(n2250), .CLK(clk), .Q(mem[408]) );
  DFFPOSX1 mem_reg_9__38_ ( .D(n2249), .CLK(clk), .Q(mem[407]) );
  DFFPOSX1 mem_reg_9__37_ ( .D(n2248), .CLK(clk), .Q(mem[406]) );
  DFFPOSX1 mem_reg_9__36_ ( .D(n2247), .CLK(clk), .Q(mem[405]) );
  DFFPOSX1 mem_reg_9__35_ ( .D(n2246), .CLK(clk), .Q(mem[404]) );
  DFFPOSX1 mem_reg_9__34_ ( .D(n2245), .CLK(clk), .Q(mem[403]) );
  DFFPOSX1 mem_reg_9__33_ ( .D(n2244), .CLK(clk), .Q(mem[402]) );
  DFFPOSX1 mem_reg_9__32_ ( .D(n2243), .CLK(clk), .Q(mem[401]) );
  DFFPOSX1 mem_reg_9__31_ ( .D(n2242), .CLK(clk), .Q(mem[400]) );
  DFFPOSX1 mem_reg_9__30_ ( .D(n2241), .CLK(clk), .Q(mem[399]) );
  DFFPOSX1 mem_reg_9__29_ ( .D(n2240), .CLK(clk), .Q(mem[398]) );
  DFFPOSX1 mem_reg_9__28_ ( .D(n2239), .CLK(clk), .Q(mem[397]) );
  DFFPOSX1 mem_reg_9__27_ ( .D(n2238), .CLK(clk), .Q(mem[396]) );
  DFFPOSX1 mem_reg_9__26_ ( .D(n2237), .CLK(clk), .Q(mem[395]) );
  DFFPOSX1 mem_reg_9__25_ ( .D(n2236), .CLK(clk), .Q(mem[394]) );
  DFFPOSX1 mem_reg_9__24_ ( .D(n2235), .CLK(clk), .Q(mem[393]) );
  DFFPOSX1 mem_reg_9__23_ ( .D(n2234), .CLK(clk), .Q(mem[392]) );
  DFFPOSX1 mem_reg_9__22_ ( .D(n2233), .CLK(clk), .Q(mem[391]) );
  DFFPOSX1 mem_reg_9__21_ ( .D(n2232), .CLK(clk), .Q(mem[390]) );
  DFFPOSX1 mem_reg_9__20_ ( .D(n2231), .CLK(clk), .Q(mem[389]) );
  DFFPOSX1 mem_reg_9__19_ ( .D(n2230), .CLK(clk), .Q(mem[388]) );
  DFFPOSX1 mem_reg_9__18_ ( .D(n2229), .CLK(clk), .Q(mem[387]) );
  DFFPOSX1 mem_reg_9__17_ ( .D(n2228), .CLK(clk), .Q(mem[386]) );
  DFFPOSX1 mem_reg_9__16_ ( .D(n2227), .CLK(clk), .Q(mem[385]) );
  DFFPOSX1 mem_reg_9__15_ ( .D(n2226), .CLK(clk), .Q(mem[384]) );
  DFFPOSX1 mem_reg_9__14_ ( .D(n2225), .CLK(clk), .Q(mem[383]) );
  DFFPOSX1 mem_reg_9__13_ ( .D(n2224), .CLK(clk), .Q(mem[382]) );
  DFFPOSX1 mem_reg_9__12_ ( .D(n2223), .CLK(clk), .Q(mem[381]) );
  DFFPOSX1 mem_reg_9__11_ ( .D(n2222), .CLK(clk), .Q(mem[380]) );
  DFFPOSX1 mem_reg_9__10_ ( .D(n2221), .CLK(clk), .Q(mem[379]) );
  DFFPOSX1 mem_reg_9__9_ ( .D(n2220), .CLK(clk), .Q(mem[378]) );
  DFFPOSX1 mem_reg_9__8_ ( .D(n2219), .CLK(clk), .Q(mem[377]) );
  DFFPOSX1 mem_reg_9__7_ ( .D(n2218), .CLK(clk), .Q(mem[376]) );
  DFFPOSX1 mem_reg_9__6_ ( .D(n2217), .CLK(clk), .Q(mem[375]) );
  DFFPOSX1 mem_reg_9__5_ ( .D(n2216), .CLK(clk), .Q(mem[374]) );
  DFFPOSX1 mem_reg_9__4_ ( .D(n2215), .CLK(clk), .Q(mem[373]) );
  DFFPOSX1 mem_reg_9__3_ ( .D(n2214), .CLK(clk), .Q(mem[372]) );
  DFFPOSX1 mem_reg_9__2_ ( .D(n2213), .CLK(clk), .Q(mem[371]) );
  DFFPOSX1 mem_reg_9__1_ ( .D(n2212), .CLK(clk), .Q(mem[370]) );
  DFFPOSX1 mem_reg_9__0_ ( .D(n2211), .CLK(clk), .Q(mem[369]) );
  DFFPOSX1 mem_reg_8__40_ ( .D(n2210), .CLK(clk), .Q(mem[368]) );
  DFFPOSX1 mem_reg_8__39_ ( .D(n2209), .CLK(clk), .Q(mem[367]) );
  DFFPOSX1 mem_reg_8__38_ ( .D(n2208), .CLK(clk), .Q(mem[366]) );
  DFFPOSX1 mem_reg_8__37_ ( .D(n2207), .CLK(clk), .Q(mem[365]) );
  DFFPOSX1 mem_reg_8__36_ ( .D(n2206), .CLK(clk), .Q(mem[364]) );
  DFFPOSX1 mem_reg_8__35_ ( .D(n2205), .CLK(clk), .Q(mem[363]) );
  DFFPOSX1 mem_reg_8__34_ ( .D(n2204), .CLK(clk), .Q(mem[362]) );
  DFFPOSX1 mem_reg_8__33_ ( .D(n2203), .CLK(clk), .Q(mem[361]) );
  DFFPOSX1 mem_reg_8__32_ ( .D(n2202), .CLK(clk), .Q(mem[360]) );
  DFFPOSX1 mem_reg_8__31_ ( .D(n2201), .CLK(clk), .Q(mem[359]) );
  DFFPOSX1 mem_reg_8__30_ ( .D(n2200), .CLK(clk), .Q(mem[358]) );
  DFFPOSX1 mem_reg_8__29_ ( .D(n2199), .CLK(clk), .Q(mem[357]) );
  DFFPOSX1 mem_reg_8__28_ ( .D(n2198), .CLK(clk), .Q(mem[356]) );
  DFFPOSX1 mem_reg_8__27_ ( .D(n2197), .CLK(clk), .Q(mem[355]) );
  DFFPOSX1 mem_reg_8__26_ ( .D(n2196), .CLK(clk), .Q(mem[354]) );
  DFFPOSX1 mem_reg_8__25_ ( .D(n2195), .CLK(clk), .Q(mem[353]) );
  DFFPOSX1 mem_reg_8__24_ ( .D(n2194), .CLK(clk), .Q(mem[352]) );
  DFFPOSX1 mem_reg_8__23_ ( .D(n2193), .CLK(clk), .Q(mem[351]) );
  DFFPOSX1 mem_reg_8__22_ ( .D(n2192), .CLK(clk), .Q(mem[350]) );
  DFFPOSX1 mem_reg_8__21_ ( .D(n2191), .CLK(clk), .Q(mem[349]) );
  DFFPOSX1 mem_reg_8__20_ ( .D(n2190), .CLK(clk), .Q(mem[348]) );
  DFFPOSX1 mem_reg_8__19_ ( .D(n2189), .CLK(clk), .Q(mem[347]) );
  DFFPOSX1 mem_reg_8__18_ ( .D(n2188), .CLK(clk), .Q(mem[346]) );
  DFFPOSX1 mem_reg_8__17_ ( .D(n2187), .CLK(clk), .Q(mem[345]) );
  DFFPOSX1 mem_reg_8__16_ ( .D(n2186), .CLK(clk), .Q(mem[344]) );
  DFFPOSX1 mem_reg_8__15_ ( .D(n2185), .CLK(clk), .Q(mem[343]) );
  DFFPOSX1 mem_reg_8__14_ ( .D(n2184), .CLK(clk), .Q(mem[342]) );
  DFFPOSX1 mem_reg_8__13_ ( .D(n2183), .CLK(clk), .Q(mem[341]) );
  DFFPOSX1 mem_reg_8__12_ ( .D(n2182), .CLK(clk), .Q(mem[340]) );
  DFFPOSX1 mem_reg_8__11_ ( .D(n2181), .CLK(clk), .Q(mem[339]) );
  DFFPOSX1 mem_reg_8__10_ ( .D(n2180), .CLK(clk), .Q(mem[338]) );
  DFFPOSX1 mem_reg_8__9_ ( .D(n2179), .CLK(clk), .Q(mem[337]) );
  DFFPOSX1 mem_reg_8__8_ ( .D(n2178), .CLK(clk), .Q(mem[336]) );
  DFFPOSX1 mem_reg_8__7_ ( .D(n2177), .CLK(clk), .Q(mem[335]) );
  DFFPOSX1 mem_reg_8__6_ ( .D(n2176), .CLK(clk), .Q(mem[334]) );
  DFFPOSX1 mem_reg_8__5_ ( .D(n2175), .CLK(clk), .Q(mem[333]) );
  DFFPOSX1 mem_reg_8__4_ ( .D(n2174), .CLK(clk), .Q(mem[332]) );
  DFFPOSX1 mem_reg_8__3_ ( .D(n2173), .CLK(clk), .Q(mem[331]) );
  DFFPOSX1 mem_reg_8__2_ ( .D(n2172), .CLK(clk), .Q(mem[330]) );
  DFFPOSX1 mem_reg_8__1_ ( .D(n2171), .CLK(clk), .Q(mem[329]) );
  DFFPOSX1 mem_reg_8__0_ ( .D(n2170), .CLK(clk), .Q(mem[328]) );
  DFFPOSX1 mem_reg_7__40_ ( .D(n2169), .CLK(clk), .Q(mem[327]) );
  DFFPOSX1 mem_reg_7__39_ ( .D(n2168), .CLK(clk), .Q(mem[326]) );
  DFFPOSX1 mem_reg_7__38_ ( .D(n2167), .CLK(clk), .Q(mem[325]) );
  DFFPOSX1 mem_reg_7__37_ ( .D(n2166), .CLK(clk), .Q(mem[324]) );
  DFFPOSX1 mem_reg_7__36_ ( .D(n2165), .CLK(clk), .Q(mem[323]) );
  DFFPOSX1 mem_reg_7__35_ ( .D(n2164), .CLK(clk), .Q(mem[322]) );
  DFFPOSX1 mem_reg_7__34_ ( .D(n2163), .CLK(clk), .Q(mem[321]) );
  DFFPOSX1 mem_reg_7__33_ ( .D(n2162), .CLK(clk), .Q(mem[320]) );
  DFFPOSX1 mem_reg_7__32_ ( .D(n2161), .CLK(clk), .Q(mem[319]) );
  DFFPOSX1 mem_reg_7__31_ ( .D(n2160), .CLK(clk), .Q(mem[318]) );
  DFFPOSX1 mem_reg_7__30_ ( .D(n2159), .CLK(clk), .Q(mem[317]) );
  DFFPOSX1 mem_reg_7__29_ ( .D(n2158), .CLK(clk), .Q(mem[316]) );
  DFFPOSX1 mem_reg_7__28_ ( .D(n2157), .CLK(clk), .Q(mem[315]) );
  DFFPOSX1 mem_reg_7__27_ ( .D(n2156), .CLK(clk), .Q(mem[314]) );
  DFFPOSX1 mem_reg_7__26_ ( .D(n2155), .CLK(clk), .Q(mem[313]) );
  DFFPOSX1 mem_reg_7__25_ ( .D(n2154), .CLK(clk), .Q(mem[312]) );
  DFFPOSX1 mem_reg_7__24_ ( .D(n2153), .CLK(clk), .Q(mem[311]) );
  DFFPOSX1 mem_reg_7__23_ ( .D(n2152), .CLK(clk), .Q(mem[310]) );
  DFFPOSX1 mem_reg_7__22_ ( .D(n2151), .CLK(clk), .Q(mem[309]) );
  DFFPOSX1 mem_reg_7__21_ ( .D(n2150), .CLK(clk), .Q(mem[308]) );
  DFFPOSX1 mem_reg_7__20_ ( .D(n2149), .CLK(clk), .Q(mem[307]) );
  DFFPOSX1 mem_reg_7__19_ ( .D(n2148), .CLK(clk), .Q(mem[306]) );
  DFFPOSX1 mem_reg_7__18_ ( .D(n2147), .CLK(clk), .Q(mem[305]) );
  DFFPOSX1 mem_reg_7__17_ ( .D(n2146), .CLK(clk), .Q(mem[304]) );
  DFFPOSX1 mem_reg_7__16_ ( .D(n2145), .CLK(clk), .Q(mem[303]) );
  DFFPOSX1 mem_reg_7__15_ ( .D(n2144), .CLK(clk), .Q(mem[302]) );
  DFFPOSX1 mem_reg_7__14_ ( .D(n2143), .CLK(clk), .Q(mem[301]) );
  DFFPOSX1 mem_reg_7__13_ ( .D(n2142), .CLK(clk), .Q(mem[300]) );
  DFFPOSX1 mem_reg_7__12_ ( .D(n2141), .CLK(clk), .Q(mem[299]) );
  DFFPOSX1 mem_reg_7__11_ ( .D(n2140), .CLK(clk), .Q(mem[298]) );
  DFFPOSX1 mem_reg_7__10_ ( .D(n2139), .CLK(clk), .Q(mem[297]) );
  DFFPOSX1 mem_reg_7__9_ ( .D(n2138), .CLK(clk), .Q(mem[296]) );
  DFFPOSX1 mem_reg_7__8_ ( .D(n2137), .CLK(clk), .Q(mem[295]) );
  DFFPOSX1 mem_reg_7__7_ ( .D(n2136), .CLK(clk), .Q(mem[294]) );
  DFFPOSX1 mem_reg_7__6_ ( .D(n2135), .CLK(clk), .Q(mem[293]) );
  DFFPOSX1 mem_reg_7__5_ ( .D(n2134), .CLK(clk), .Q(mem[292]) );
  DFFPOSX1 mem_reg_7__4_ ( .D(n2133), .CLK(clk), .Q(mem[291]) );
  DFFPOSX1 mem_reg_7__3_ ( .D(n2132), .CLK(clk), .Q(mem[290]) );
  DFFPOSX1 mem_reg_7__2_ ( .D(n2131), .CLK(clk), .Q(mem[289]) );
  DFFPOSX1 mem_reg_7__1_ ( .D(n2130), .CLK(clk), .Q(mem[288]) );
  DFFPOSX1 mem_reg_7__0_ ( .D(n2129), .CLK(clk), .Q(mem[287]) );
  DFFPOSX1 mem_reg_6__40_ ( .D(n2128), .CLK(clk), .Q(mem[286]) );
  DFFPOSX1 mem_reg_6__39_ ( .D(n2127), .CLK(clk), .Q(mem[285]) );
  DFFPOSX1 mem_reg_6__38_ ( .D(n2126), .CLK(clk), .Q(mem[284]) );
  DFFPOSX1 mem_reg_6__37_ ( .D(n2125), .CLK(clk), .Q(mem[283]) );
  DFFPOSX1 mem_reg_6__36_ ( .D(n2124), .CLK(clk), .Q(mem[282]) );
  DFFPOSX1 mem_reg_6__35_ ( .D(n2123), .CLK(clk), .Q(mem[281]) );
  DFFPOSX1 mem_reg_6__34_ ( .D(n2122), .CLK(clk), .Q(mem[280]) );
  DFFPOSX1 mem_reg_6__33_ ( .D(n2121), .CLK(clk), .Q(mem[279]) );
  DFFPOSX1 mem_reg_6__32_ ( .D(n2120), .CLK(clk), .Q(mem[278]) );
  DFFPOSX1 mem_reg_6__31_ ( .D(n2119), .CLK(clk), .Q(mem[277]) );
  DFFPOSX1 mem_reg_6__30_ ( .D(n2118), .CLK(clk), .Q(mem[276]) );
  DFFPOSX1 mem_reg_6__29_ ( .D(n2117), .CLK(clk), .Q(mem[275]) );
  DFFPOSX1 mem_reg_6__28_ ( .D(n2116), .CLK(clk), .Q(mem[274]) );
  DFFPOSX1 mem_reg_6__27_ ( .D(n2115), .CLK(clk), .Q(mem[273]) );
  DFFPOSX1 mem_reg_6__26_ ( .D(n2114), .CLK(clk), .Q(mem[272]) );
  DFFPOSX1 mem_reg_6__25_ ( .D(n2113), .CLK(clk), .Q(mem[271]) );
  DFFPOSX1 mem_reg_6__24_ ( .D(n2112), .CLK(clk), .Q(mem[270]) );
  DFFPOSX1 mem_reg_6__23_ ( .D(n2111), .CLK(clk), .Q(mem[269]) );
  DFFPOSX1 mem_reg_6__22_ ( .D(n2110), .CLK(clk), .Q(mem[268]) );
  DFFPOSX1 mem_reg_6__21_ ( .D(n2109), .CLK(clk), .Q(mem[267]) );
  DFFPOSX1 mem_reg_6__20_ ( .D(n2108), .CLK(clk), .Q(mem[266]) );
  DFFPOSX1 mem_reg_6__19_ ( .D(n2107), .CLK(clk), .Q(mem[265]) );
  DFFPOSX1 mem_reg_6__18_ ( .D(n2106), .CLK(clk), .Q(mem[264]) );
  DFFPOSX1 mem_reg_6__17_ ( .D(n2105), .CLK(clk), .Q(mem[263]) );
  DFFPOSX1 mem_reg_6__16_ ( .D(n2104), .CLK(clk), .Q(mem[262]) );
  DFFPOSX1 mem_reg_6__15_ ( .D(n2103), .CLK(clk), .Q(mem[261]) );
  DFFPOSX1 mem_reg_6__14_ ( .D(n2102), .CLK(clk), .Q(mem[260]) );
  DFFPOSX1 mem_reg_6__13_ ( .D(n2101), .CLK(clk), .Q(mem[259]) );
  DFFPOSX1 mem_reg_6__12_ ( .D(n2100), .CLK(clk), .Q(mem[258]) );
  DFFPOSX1 mem_reg_6__11_ ( .D(n2099), .CLK(clk), .Q(mem[257]) );
  DFFPOSX1 mem_reg_6__10_ ( .D(n2098), .CLK(clk), .Q(mem[256]) );
  DFFPOSX1 mem_reg_6__9_ ( .D(n2097), .CLK(clk), .Q(mem[255]) );
  DFFPOSX1 mem_reg_6__8_ ( .D(n2096), .CLK(clk), .Q(mem[254]) );
  DFFPOSX1 mem_reg_6__7_ ( .D(n2095), .CLK(clk), .Q(mem[253]) );
  DFFPOSX1 mem_reg_6__6_ ( .D(n2094), .CLK(clk), .Q(mem[252]) );
  DFFPOSX1 mem_reg_6__5_ ( .D(n2093), .CLK(clk), .Q(mem[251]) );
  DFFPOSX1 mem_reg_6__4_ ( .D(n2092), .CLK(clk), .Q(mem[250]) );
  DFFPOSX1 mem_reg_6__3_ ( .D(n2091), .CLK(clk), .Q(mem[249]) );
  DFFPOSX1 mem_reg_6__2_ ( .D(n2090), .CLK(clk), .Q(mem[248]) );
  DFFPOSX1 mem_reg_6__1_ ( .D(n2089), .CLK(clk), .Q(mem[247]) );
  DFFPOSX1 mem_reg_6__0_ ( .D(n2088), .CLK(clk), .Q(mem[246]) );
  DFFPOSX1 mem_reg_5__40_ ( .D(n2087), .CLK(clk), .Q(mem[245]) );
  DFFPOSX1 mem_reg_5__39_ ( .D(n2086), .CLK(clk), .Q(mem[244]) );
  DFFPOSX1 mem_reg_5__38_ ( .D(n2085), .CLK(clk), .Q(mem[243]) );
  DFFPOSX1 mem_reg_5__37_ ( .D(n2084), .CLK(clk), .Q(mem[242]) );
  DFFPOSX1 mem_reg_5__36_ ( .D(n2083), .CLK(clk), .Q(mem[241]) );
  DFFPOSX1 mem_reg_5__35_ ( .D(n2082), .CLK(clk), .Q(mem[240]) );
  DFFPOSX1 mem_reg_5__34_ ( .D(n2081), .CLK(clk), .Q(mem[239]) );
  DFFPOSX1 mem_reg_5__33_ ( .D(n2080), .CLK(clk), .Q(mem[238]) );
  DFFPOSX1 mem_reg_5__32_ ( .D(n2079), .CLK(clk), .Q(mem[237]) );
  DFFPOSX1 mem_reg_5__31_ ( .D(n2078), .CLK(clk), .Q(mem[236]) );
  DFFPOSX1 mem_reg_5__30_ ( .D(n2077), .CLK(clk), .Q(mem[235]) );
  DFFPOSX1 mem_reg_5__29_ ( .D(n2076), .CLK(clk), .Q(mem[234]) );
  DFFPOSX1 mem_reg_5__28_ ( .D(n2075), .CLK(clk), .Q(mem[233]) );
  DFFPOSX1 mem_reg_5__27_ ( .D(n2074), .CLK(clk), .Q(mem[232]) );
  DFFPOSX1 mem_reg_5__26_ ( .D(n2073), .CLK(clk), .Q(mem[231]) );
  DFFPOSX1 mem_reg_5__25_ ( .D(n2072), .CLK(clk), .Q(mem[230]) );
  DFFPOSX1 mem_reg_5__24_ ( .D(n2071), .CLK(clk), .Q(mem[229]) );
  DFFPOSX1 mem_reg_5__23_ ( .D(n2070), .CLK(clk), .Q(mem[228]) );
  DFFPOSX1 mem_reg_5__22_ ( .D(n2069), .CLK(clk), .Q(mem[227]) );
  DFFPOSX1 mem_reg_5__21_ ( .D(n2068), .CLK(clk), .Q(mem[226]) );
  DFFPOSX1 mem_reg_5__20_ ( .D(n2067), .CLK(clk), .Q(mem[225]) );
  DFFPOSX1 mem_reg_5__19_ ( .D(n2066), .CLK(clk), .Q(mem[224]) );
  DFFPOSX1 mem_reg_5__18_ ( .D(n2065), .CLK(clk), .Q(mem[223]) );
  DFFPOSX1 mem_reg_5__17_ ( .D(n2064), .CLK(clk), .Q(mem[222]) );
  DFFPOSX1 mem_reg_5__16_ ( .D(n2063), .CLK(clk), .Q(mem[221]) );
  DFFPOSX1 mem_reg_5__15_ ( .D(n2062), .CLK(clk), .Q(mem[220]) );
  DFFPOSX1 mem_reg_5__14_ ( .D(n2061), .CLK(clk), .Q(mem[219]) );
  DFFPOSX1 mem_reg_5__13_ ( .D(n2060), .CLK(clk), .Q(mem[218]) );
  DFFPOSX1 mem_reg_5__12_ ( .D(n2059), .CLK(clk), .Q(mem[217]) );
  DFFPOSX1 mem_reg_5__11_ ( .D(n2058), .CLK(clk), .Q(mem[216]) );
  DFFPOSX1 mem_reg_5__10_ ( .D(n2057), .CLK(clk), .Q(mem[215]) );
  DFFPOSX1 mem_reg_5__9_ ( .D(n2056), .CLK(clk), .Q(mem[214]) );
  DFFPOSX1 mem_reg_5__8_ ( .D(n2055), .CLK(clk), .Q(mem[213]) );
  DFFPOSX1 mem_reg_5__7_ ( .D(n2054), .CLK(clk), .Q(mem[212]) );
  DFFPOSX1 mem_reg_5__6_ ( .D(n2053), .CLK(clk), .Q(mem[211]) );
  DFFPOSX1 mem_reg_5__5_ ( .D(n2052), .CLK(clk), .Q(mem[210]) );
  DFFPOSX1 mem_reg_5__4_ ( .D(n2051), .CLK(clk), .Q(mem[209]) );
  DFFPOSX1 mem_reg_5__3_ ( .D(n2050), .CLK(clk), .Q(mem[208]) );
  DFFPOSX1 mem_reg_5__2_ ( .D(n2049), .CLK(clk), .Q(mem[207]) );
  DFFPOSX1 mem_reg_5__1_ ( .D(n2048), .CLK(clk), .Q(mem[206]) );
  DFFPOSX1 mem_reg_5__0_ ( .D(n2047), .CLK(clk), .Q(mem[205]) );
  DFFPOSX1 mem_reg_4__40_ ( .D(n2046), .CLK(clk), .Q(mem[204]) );
  DFFPOSX1 mem_reg_4__39_ ( .D(n2045), .CLK(clk), .Q(mem[203]) );
  DFFPOSX1 mem_reg_4__38_ ( .D(n2044), .CLK(clk), .Q(mem[202]) );
  DFFPOSX1 mem_reg_4__37_ ( .D(n2043), .CLK(clk), .Q(mem[201]) );
  DFFPOSX1 mem_reg_4__36_ ( .D(n2042), .CLK(clk), .Q(mem[200]) );
  DFFPOSX1 mem_reg_4__35_ ( .D(n2041), .CLK(clk), .Q(mem[199]) );
  DFFPOSX1 mem_reg_4__34_ ( .D(n2040), .CLK(clk), .Q(mem[198]) );
  DFFPOSX1 mem_reg_4__33_ ( .D(n2039), .CLK(clk), .Q(mem[197]) );
  DFFPOSX1 mem_reg_4__32_ ( .D(n2038), .CLK(clk), .Q(mem[196]) );
  DFFPOSX1 mem_reg_4__31_ ( .D(n2037), .CLK(clk), .Q(mem[195]) );
  DFFPOSX1 mem_reg_4__30_ ( .D(n2036), .CLK(clk), .Q(mem[194]) );
  DFFPOSX1 mem_reg_4__29_ ( .D(n2035), .CLK(clk), .Q(mem[193]) );
  DFFPOSX1 mem_reg_4__28_ ( .D(n2034), .CLK(clk), .Q(mem[192]) );
  DFFPOSX1 mem_reg_4__27_ ( .D(n2033), .CLK(clk), .Q(mem[191]) );
  DFFPOSX1 mem_reg_4__26_ ( .D(n2032), .CLK(clk), .Q(mem[190]) );
  DFFPOSX1 mem_reg_4__25_ ( .D(n2031), .CLK(clk), .Q(mem[189]) );
  DFFPOSX1 mem_reg_4__24_ ( .D(n2030), .CLK(clk), .Q(mem[188]) );
  DFFPOSX1 mem_reg_4__23_ ( .D(n2029), .CLK(clk), .Q(mem[187]) );
  DFFPOSX1 mem_reg_4__22_ ( .D(n2028), .CLK(clk), .Q(mem[186]) );
  DFFPOSX1 mem_reg_4__21_ ( .D(n2027), .CLK(clk), .Q(mem[185]) );
  DFFPOSX1 mem_reg_4__20_ ( .D(n2026), .CLK(clk), .Q(mem[184]) );
  DFFPOSX1 mem_reg_4__19_ ( .D(n2025), .CLK(clk), .Q(mem[183]) );
  DFFPOSX1 mem_reg_4__18_ ( .D(n2024), .CLK(clk), .Q(mem[182]) );
  DFFPOSX1 mem_reg_4__17_ ( .D(n2023), .CLK(clk), .Q(mem[181]) );
  DFFPOSX1 mem_reg_4__16_ ( .D(n2022), .CLK(clk), .Q(mem[180]) );
  DFFPOSX1 mem_reg_4__15_ ( .D(n2021), .CLK(clk), .Q(mem[179]) );
  DFFPOSX1 mem_reg_4__14_ ( .D(n2020), .CLK(clk), .Q(mem[178]) );
  DFFPOSX1 mem_reg_4__13_ ( .D(n2019), .CLK(clk), .Q(mem[177]) );
  DFFPOSX1 mem_reg_4__12_ ( .D(n2018), .CLK(clk), .Q(mem[176]) );
  DFFPOSX1 mem_reg_4__11_ ( .D(n2017), .CLK(clk), .Q(mem[175]) );
  DFFPOSX1 mem_reg_4__10_ ( .D(n2016), .CLK(clk), .Q(mem[174]) );
  DFFPOSX1 mem_reg_4__9_ ( .D(n2015), .CLK(clk), .Q(mem[173]) );
  DFFPOSX1 mem_reg_4__8_ ( .D(n2014), .CLK(clk), .Q(mem[172]) );
  DFFPOSX1 mem_reg_4__7_ ( .D(n2013), .CLK(clk), .Q(mem[171]) );
  DFFPOSX1 mem_reg_4__6_ ( .D(n2012), .CLK(clk), .Q(mem[170]) );
  DFFPOSX1 mem_reg_4__5_ ( .D(n2011), .CLK(clk), .Q(mem[169]) );
  DFFPOSX1 mem_reg_4__4_ ( .D(n2010), .CLK(clk), .Q(mem[168]) );
  DFFPOSX1 mem_reg_4__3_ ( .D(n2009), .CLK(clk), .Q(mem[167]) );
  DFFPOSX1 mem_reg_4__2_ ( .D(n2008), .CLK(clk), .Q(mem[166]) );
  DFFPOSX1 mem_reg_4__1_ ( .D(n2007), .CLK(clk), .Q(mem[165]) );
  DFFPOSX1 mem_reg_4__0_ ( .D(n2006), .CLK(clk), .Q(mem[164]) );
  DFFPOSX1 mem_reg_3__40_ ( .D(n2005), .CLK(clk), .Q(mem[163]) );
  DFFPOSX1 mem_reg_3__39_ ( .D(n2004), .CLK(clk), .Q(mem[162]) );
  DFFPOSX1 mem_reg_3__38_ ( .D(n2003), .CLK(clk), .Q(mem[161]) );
  DFFPOSX1 mem_reg_3__37_ ( .D(n2002), .CLK(clk), .Q(mem[160]) );
  DFFPOSX1 mem_reg_3__36_ ( .D(n2001), .CLK(clk), .Q(mem[159]) );
  DFFPOSX1 mem_reg_3__35_ ( .D(n2000), .CLK(clk), .Q(mem[158]) );
  DFFPOSX1 mem_reg_3__34_ ( .D(n1999), .CLK(clk), .Q(mem[157]) );
  DFFPOSX1 mem_reg_3__33_ ( .D(n1998), .CLK(clk), .Q(mem[156]) );
  DFFPOSX1 mem_reg_3__32_ ( .D(n1997), .CLK(clk), .Q(mem[155]) );
  DFFPOSX1 mem_reg_3__31_ ( .D(n1996), .CLK(clk), .Q(mem[154]) );
  DFFPOSX1 mem_reg_3__30_ ( .D(n1995), .CLK(clk), .Q(mem[153]) );
  DFFPOSX1 mem_reg_3__29_ ( .D(n1994), .CLK(clk), .Q(mem[152]) );
  DFFPOSX1 mem_reg_3__28_ ( .D(n1993), .CLK(clk), .Q(mem[151]) );
  DFFPOSX1 mem_reg_3__27_ ( .D(n1992), .CLK(clk), .Q(mem[150]) );
  DFFPOSX1 mem_reg_3__26_ ( .D(n1991), .CLK(clk), .Q(mem[149]) );
  DFFPOSX1 mem_reg_3__25_ ( .D(n1990), .CLK(clk), .Q(mem[148]) );
  DFFPOSX1 mem_reg_3__24_ ( .D(n1989), .CLK(clk), .Q(mem[147]) );
  DFFPOSX1 mem_reg_3__23_ ( .D(n1988), .CLK(clk), .Q(mem[146]) );
  DFFPOSX1 mem_reg_3__22_ ( .D(n1987), .CLK(clk), .Q(mem[145]) );
  DFFPOSX1 mem_reg_3__21_ ( .D(n1986), .CLK(clk), .Q(mem[144]) );
  DFFPOSX1 mem_reg_3__20_ ( .D(n1985), .CLK(clk), .Q(mem[143]) );
  DFFPOSX1 mem_reg_3__19_ ( .D(n1984), .CLK(clk), .Q(mem[142]) );
  DFFPOSX1 mem_reg_3__18_ ( .D(n1983), .CLK(clk), .Q(mem[141]) );
  DFFPOSX1 mem_reg_3__17_ ( .D(n1982), .CLK(clk), .Q(mem[140]) );
  DFFPOSX1 mem_reg_3__16_ ( .D(n1981), .CLK(clk), .Q(mem[139]) );
  DFFPOSX1 mem_reg_3__15_ ( .D(n1980), .CLK(clk), .Q(mem[138]) );
  DFFPOSX1 mem_reg_3__14_ ( .D(n1979), .CLK(clk), .Q(mem[137]) );
  DFFPOSX1 mem_reg_3__13_ ( .D(n1978), .CLK(clk), .Q(mem[136]) );
  DFFPOSX1 mem_reg_3__12_ ( .D(n1977), .CLK(clk), .Q(mem[135]) );
  DFFPOSX1 mem_reg_3__11_ ( .D(n1976), .CLK(clk), .Q(mem[134]) );
  DFFPOSX1 mem_reg_3__10_ ( .D(n1975), .CLK(clk), .Q(mem[133]) );
  DFFPOSX1 mem_reg_3__9_ ( .D(n1974), .CLK(clk), .Q(mem[132]) );
  DFFPOSX1 mem_reg_3__8_ ( .D(n1973), .CLK(clk), .Q(mem[131]) );
  DFFPOSX1 mem_reg_3__7_ ( .D(n1972), .CLK(clk), .Q(mem[130]) );
  DFFPOSX1 mem_reg_3__6_ ( .D(n1971), .CLK(clk), .Q(mem[129]) );
  DFFPOSX1 mem_reg_3__5_ ( .D(n1970), .CLK(clk), .Q(mem[128]) );
  DFFPOSX1 mem_reg_3__4_ ( .D(n1969), .CLK(clk), .Q(mem[127]) );
  DFFPOSX1 mem_reg_3__3_ ( .D(n1968), .CLK(clk), .Q(mem[126]) );
  DFFPOSX1 mem_reg_3__2_ ( .D(n1967), .CLK(clk), .Q(mem[125]) );
  DFFPOSX1 mem_reg_3__1_ ( .D(n1966), .CLK(clk), .Q(mem[124]) );
  DFFPOSX1 mem_reg_3__0_ ( .D(n1965), .CLK(clk), .Q(mem[123]) );
  DFFPOSX1 mem_reg_2__40_ ( .D(n1964), .CLK(clk), .Q(mem[122]) );
  DFFPOSX1 mem_reg_2__39_ ( .D(n1963), .CLK(clk), .Q(mem[121]) );
  DFFPOSX1 mem_reg_2__38_ ( .D(n1962), .CLK(clk), .Q(mem[120]) );
  DFFPOSX1 mem_reg_2__37_ ( .D(n1961), .CLK(clk), .Q(mem[119]) );
  DFFPOSX1 mem_reg_2__36_ ( .D(n1960), .CLK(clk), .Q(mem[118]) );
  DFFPOSX1 mem_reg_2__35_ ( .D(n1959), .CLK(clk), .Q(mem[117]) );
  DFFPOSX1 mem_reg_2__34_ ( .D(n1958), .CLK(clk), .Q(mem[116]) );
  DFFPOSX1 mem_reg_2__33_ ( .D(n1957), .CLK(clk), .Q(mem[115]) );
  DFFPOSX1 mem_reg_2__32_ ( .D(n1956), .CLK(clk), .Q(mem[114]) );
  DFFPOSX1 mem_reg_2__31_ ( .D(n1955), .CLK(clk), .Q(mem[113]) );
  DFFPOSX1 mem_reg_2__30_ ( .D(n1954), .CLK(clk), .Q(mem[112]) );
  DFFPOSX1 mem_reg_2__29_ ( .D(n1953), .CLK(clk), .Q(mem[111]) );
  DFFPOSX1 mem_reg_2__28_ ( .D(n1952), .CLK(clk), .Q(mem[110]) );
  DFFPOSX1 mem_reg_2__27_ ( .D(n1951), .CLK(clk), .Q(mem[109]) );
  DFFPOSX1 mem_reg_2__26_ ( .D(n1950), .CLK(clk), .Q(mem[108]) );
  DFFPOSX1 mem_reg_2__25_ ( .D(n1949), .CLK(clk), .Q(mem[107]) );
  DFFPOSX1 mem_reg_2__24_ ( .D(n1948), .CLK(clk), .Q(mem[106]) );
  DFFPOSX1 mem_reg_2__23_ ( .D(n1947), .CLK(clk), .Q(mem[105]) );
  DFFPOSX1 mem_reg_2__22_ ( .D(n1946), .CLK(clk), .Q(mem[104]) );
  DFFPOSX1 mem_reg_2__21_ ( .D(n1945), .CLK(clk), .Q(mem[103]) );
  DFFPOSX1 mem_reg_2__20_ ( .D(n1944), .CLK(clk), .Q(mem[102]) );
  DFFPOSX1 mem_reg_2__19_ ( .D(n1943), .CLK(clk), .Q(mem[101]) );
  DFFPOSX1 mem_reg_2__18_ ( .D(n1942), .CLK(clk), .Q(mem[100]) );
  DFFPOSX1 mem_reg_2__17_ ( .D(n1941), .CLK(clk), .Q(mem[99]) );
  DFFPOSX1 mem_reg_2__16_ ( .D(n1940), .CLK(clk), .Q(mem[98]) );
  DFFPOSX1 mem_reg_2__15_ ( .D(n1939), .CLK(clk), .Q(mem[97]) );
  DFFPOSX1 mem_reg_2__14_ ( .D(n1938), .CLK(clk), .Q(mem[96]) );
  DFFPOSX1 mem_reg_2__13_ ( .D(n1937), .CLK(clk), .Q(mem[95]) );
  DFFPOSX1 mem_reg_2__12_ ( .D(n1936), .CLK(clk), .Q(mem[94]) );
  DFFPOSX1 mem_reg_2__11_ ( .D(n1935), .CLK(clk), .Q(mem[93]) );
  DFFPOSX1 mem_reg_2__10_ ( .D(n1934), .CLK(clk), .Q(mem[92]) );
  DFFPOSX1 mem_reg_2__9_ ( .D(n1933), .CLK(clk), .Q(mem[91]) );
  DFFPOSX1 mem_reg_2__8_ ( .D(n1932), .CLK(clk), .Q(mem[90]) );
  DFFPOSX1 mem_reg_2__7_ ( .D(n1931), .CLK(clk), .Q(mem[89]) );
  DFFPOSX1 mem_reg_2__6_ ( .D(n1930), .CLK(clk), .Q(mem[88]) );
  DFFPOSX1 mem_reg_2__5_ ( .D(n1929), .CLK(clk), .Q(mem[87]) );
  DFFPOSX1 mem_reg_2__4_ ( .D(n1928), .CLK(clk), .Q(mem[86]) );
  DFFPOSX1 mem_reg_2__3_ ( .D(n1927), .CLK(clk), .Q(mem[85]) );
  DFFPOSX1 mem_reg_2__2_ ( .D(n1926), .CLK(clk), .Q(mem[84]) );
  DFFPOSX1 mem_reg_2__1_ ( .D(n1925), .CLK(clk), .Q(mem[83]) );
  DFFPOSX1 mem_reg_2__0_ ( .D(n1924), .CLK(clk), .Q(mem[82]) );
  DFFPOSX1 mem_reg_1__40_ ( .D(n1923), .CLK(clk), .Q(mem[81]) );
  DFFPOSX1 mem_reg_1__39_ ( .D(n1922), .CLK(clk), .Q(mem[80]) );
  DFFPOSX1 mem_reg_1__38_ ( .D(n1921), .CLK(clk), .Q(mem[79]) );
  DFFPOSX1 mem_reg_1__37_ ( .D(n1920), .CLK(clk), .Q(mem[78]) );
  DFFPOSX1 mem_reg_1__36_ ( .D(n1919), .CLK(clk), .Q(mem[77]) );
  DFFPOSX1 mem_reg_1__35_ ( .D(n1918), .CLK(clk), .Q(mem[76]) );
  DFFPOSX1 mem_reg_1__34_ ( .D(n1917), .CLK(clk), .Q(mem[75]) );
  DFFPOSX1 mem_reg_1__33_ ( .D(n1916), .CLK(clk), .Q(mem[74]) );
  DFFPOSX1 mem_reg_1__32_ ( .D(n1915), .CLK(clk), .Q(mem[73]) );
  DFFPOSX1 mem_reg_1__31_ ( .D(n1914), .CLK(clk), .Q(mem[72]) );
  DFFPOSX1 mem_reg_1__30_ ( .D(n1913), .CLK(clk), .Q(mem[71]) );
  DFFPOSX1 mem_reg_1__29_ ( .D(n1912), .CLK(clk), .Q(mem[70]) );
  DFFPOSX1 mem_reg_1__28_ ( .D(n1911), .CLK(clk), .Q(mem[69]) );
  DFFPOSX1 mem_reg_1__27_ ( .D(n1910), .CLK(clk), .Q(mem[68]) );
  DFFPOSX1 mem_reg_1__26_ ( .D(n1909), .CLK(clk), .Q(mem[67]) );
  DFFPOSX1 mem_reg_1__25_ ( .D(n1908), .CLK(clk), .Q(mem[66]) );
  DFFPOSX1 mem_reg_1__24_ ( .D(n1907), .CLK(clk), .Q(mem[65]) );
  DFFPOSX1 mem_reg_1__23_ ( .D(n1906), .CLK(clk), .Q(mem[64]) );
  DFFPOSX1 mem_reg_1__22_ ( .D(n1905), .CLK(clk), .Q(mem[63]) );
  DFFPOSX1 mem_reg_1__21_ ( .D(n1904), .CLK(clk), .Q(mem[62]) );
  DFFPOSX1 mem_reg_1__20_ ( .D(n1903), .CLK(clk), .Q(mem[61]) );
  DFFPOSX1 mem_reg_1__19_ ( .D(n1902), .CLK(clk), .Q(mem[60]) );
  DFFPOSX1 mem_reg_1__18_ ( .D(n1901), .CLK(clk), .Q(mem[59]) );
  DFFPOSX1 mem_reg_1__17_ ( .D(n1900), .CLK(clk), .Q(mem[58]) );
  DFFPOSX1 mem_reg_1__16_ ( .D(n1899), .CLK(clk), .Q(mem[57]) );
  DFFPOSX1 mem_reg_1__15_ ( .D(n1898), .CLK(clk), .Q(mem[56]) );
  DFFPOSX1 mem_reg_1__14_ ( .D(n1897), .CLK(clk), .Q(mem[55]) );
  DFFPOSX1 mem_reg_1__13_ ( .D(n1896), .CLK(clk), .Q(mem[54]) );
  DFFPOSX1 mem_reg_1__12_ ( .D(n1895), .CLK(clk), .Q(mem[53]) );
  DFFPOSX1 mem_reg_1__11_ ( .D(n1894), .CLK(clk), .Q(mem[52]) );
  DFFPOSX1 mem_reg_1__10_ ( .D(n1893), .CLK(clk), .Q(mem[51]) );
  DFFPOSX1 mem_reg_1__9_ ( .D(n1892), .CLK(clk), .Q(mem[50]) );
  DFFPOSX1 mem_reg_1__8_ ( .D(n1891), .CLK(clk), .Q(mem[49]) );
  DFFPOSX1 mem_reg_1__7_ ( .D(n1890), .CLK(clk), .Q(mem[48]) );
  DFFPOSX1 mem_reg_1__6_ ( .D(n1889), .CLK(clk), .Q(mem[47]) );
  DFFPOSX1 mem_reg_1__5_ ( .D(n1888), .CLK(clk), .Q(mem[46]) );
  DFFPOSX1 mem_reg_1__4_ ( .D(n1887), .CLK(clk), .Q(mem[45]) );
  DFFPOSX1 mem_reg_1__3_ ( .D(n1886), .CLK(clk), .Q(mem[44]) );
  DFFPOSX1 mem_reg_1__2_ ( .D(n1885), .CLK(clk), .Q(mem[43]) );
  DFFPOSX1 mem_reg_1__1_ ( .D(n1884), .CLK(clk), .Q(mem[42]) );
  DFFPOSX1 mem_reg_1__0_ ( .D(n1883), .CLK(clk), .Q(mem[41]) );
  DFFPOSX1 mem_reg_0__40_ ( .D(n1882), .CLK(clk), .Q(mem[40]) );
  DFFPOSX1 mem_reg_0__39_ ( .D(n1881), .CLK(clk), .Q(mem[39]) );
  DFFPOSX1 mem_reg_0__38_ ( .D(n1880), .CLK(clk), .Q(mem[38]) );
  DFFPOSX1 mem_reg_0__37_ ( .D(n1879), .CLK(clk), .Q(mem[37]) );
  DFFPOSX1 mem_reg_0__36_ ( .D(n1878), .CLK(clk), .Q(mem[36]) );
  DFFPOSX1 mem_reg_0__35_ ( .D(n1877), .CLK(clk), .Q(mem[35]) );
  DFFPOSX1 mem_reg_0__34_ ( .D(n1876), .CLK(clk), .Q(mem[34]) );
  DFFPOSX1 mem_reg_0__33_ ( .D(n1875), .CLK(clk), .Q(mem[33]) );
  DFFPOSX1 mem_reg_0__32_ ( .D(n1874), .CLK(clk), .Q(mem[32]) );
  DFFPOSX1 mem_reg_0__31_ ( .D(n1873), .CLK(clk), .Q(mem[31]) );
  DFFPOSX1 mem_reg_0__30_ ( .D(n1872), .CLK(clk), .Q(mem[30]) );
  DFFPOSX1 mem_reg_0__29_ ( .D(n1871), .CLK(clk), .Q(mem[29]) );
  DFFPOSX1 mem_reg_0__28_ ( .D(n1870), .CLK(clk), .Q(mem[28]) );
  DFFPOSX1 mem_reg_0__27_ ( .D(n1869), .CLK(clk), .Q(mem[27]) );
  DFFPOSX1 mem_reg_0__26_ ( .D(n1868), .CLK(clk), .Q(mem[26]) );
  DFFPOSX1 mem_reg_0__25_ ( .D(n1867), .CLK(clk), .Q(mem[25]) );
  DFFPOSX1 mem_reg_0__24_ ( .D(n1866), .CLK(clk), .Q(mem[24]) );
  DFFPOSX1 mem_reg_0__23_ ( .D(n1865), .CLK(clk), .Q(mem[23]) );
  DFFPOSX1 mem_reg_0__22_ ( .D(n1864), .CLK(clk), .Q(mem[22]) );
  DFFPOSX1 mem_reg_0__21_ ( .D(n1863), .CLK(clk), .Q(mem[21]) );
  DFFPOSX1 mem_reg_0__20_ ( .D(n1862), .CLK(clk), .Q(mem[20]) );
  DFFPOSX1 mem_reg_0__19_ ( .D(n1861), .CLK(clk), .Q(mem[19]) );
  DFFPOSX1 mem_reg_0__18_ ( .D(n1860), .CLK(clk), .Q(mem[18]) );
  DFFPOSX1 mem_reg_0__17_ ( .D(n1859), .CLK(clk), .Q(mem[17]) );
  DFFPOSX1 mem_reg_0__16_ ( .D(n1858), .CLK(clk), .Q(mem[16]) );
  DFFPOSX1 mem_reg_0__15_ ( .D(n1857), .CLK(clk), .Q(mem[15]) );
  DFFPOSX1 mem_reg_0__14_ ( .D(n1856), .CLK(clk), .Q(mem[14]) );
  DFFPOSX1 mem_reg_0__13_ ( .D(n1855), .CLK(clk), .Q(mem[13]) );
  DFFPOSX1 mem_reg_0__12_ ( .D(n1854), .CLK(clk), .Q(mem[12]) );
  DFFPOSX1 mem_reg_0__11_ ( .D(n1853), .CLK(clk), .Q(mem[11]) );
  DFFPOSX1 mem_reg_0__10_ ( .D(n1852), .CLK(clk), .Q(mem[10]) );
  DFFPOSX1 mem_reg_0__9_ ( .D(n1851), .CLK(clk), .Q(mem[9]) );
  DFFPOSX1 mem_reg_0__8_ ( .D(n1850), .CLK(clk), .Q(mem[8]) );
  DFFPOSX1 mem_reg_0__7_ ( .D(n1849), .CLK(clk), .Q(mem[7]) );
  DFFPOSX1 mem_reg_0__6_ ( .D(n1848), .CLK(clk), .Q(mem[6]) );
  DFFPOSX1 mem_reg_0__5_ ( .D(n1847), .CLK(clk), .Q(mem[5]) );
  DFFPOSX1 mem_reg_0__4_ ( .D(n1846), .CLK(clk), .Q(mem[4]) );
  DFFPOSX1 mem_reg_0__3_ ( .D(n1845), .CLK(clk), .Q(mem[3]) );
  DFFPOSX1 mem_reg_0__2_ ( .D(n1844), .CLK(clk), .Q(mem[2]) );
  DFFPOSX1 mem_reg_0__1_ ( .D(n1843), .CLK(clk), .Q(mem[1]) );
  DFFPOSX1 mem_reg_0__0_ ( .D(n1842), .CLK(clk), .Q(mem[0]) );
  OAI21X1 U1433 ( .A(n8503), .B(n8510), .C(n1342), .Y(fillcount[5]) );
  OAI21X1 U1434 ( .A(n7115), .B(n16), .C(n8515), .Y(n1342) );
  NAND3X1 U1435 ( .A(n6333), .B(n1345), .C(n1346), .Y(n5507) );
  NOR3X1 U1436 ( .A(n7032), .B(n7073), .C(n7114), .Y(n1346) );
  NAND3X1 U1438 ( .A(n4046), .B(n6662), .C(n6991), .Y(n1351) );
  AOI22X1 U1439 ( .A(n1354), .B(n9040), .C(n8490), .D(n8917), .Y(n1353) );
  NAND3X1 U1441 ( .A(n6291), .B(n6661), .C(n6990), .Y(n1350) );
  AOI22X1 U1442 ( .A(n1359), .B(n9122), .C(n1360), .D(n8958), .Y(n1358) );
  AOI22X1 U1444 ( .A(n1362), .B(n9163), .C(n1363), .D(n9081), .Y(n1356) );
  NAND3X1 U1446 ( .A(n1366), .B(n6660), .C(n6989), .Y(n1365) );
  AOI22X1 U1447 ( .A(n1354), .B(n8712), .C(n8485), .D(n8589), .Y(n1368) );
  NAND3X1 U1449 ( .A(n6290), .B(n6659), .C(n6988), .Y(n1364) );
  AOI22X1 U1450 ( .A(n1359), .B(n8794), .C(n1360), .D(n8630), .Y(n1371) );
  AOI22X1 U1452 ( .A(n1362), .B(n8835), .C(n1363), .D(n8753), .Y(n1369) );
  NAND3X1 U1454 ( .A(n1374), .B(n6658), .C(n6987), .Y(n1373) );
  AOI22X1 U1455 ( .A(n1354), .B(n9696), .C(n8483), .D(n9573), .Y(n1376) );
  NAND3X1 U1457 ( .A(n6289), .B(n6657), .C(n6986), .Y(n1372) );
  AOI22X1 U1458 ( .A(n1359), .B(n9778), .C(n1360), .D(n9614), .Y(n1379) );
  AOI22X1 U1460 ( .A(n1362), .B(n9819), .C(n1363), .D(n9737), .Y(n1377) );
  NAND3X1 U1461 ( .A(n1382), .B(n6656), .C(n6985), .Y(n1381) );
  AOI22X1 U1462 ( .A(n1354), .B(n9368), .C(n8487), .D(n9245), .Y(n1384) );
  NAND3X1 U1464 ( .A(n6288), .B(n6655), .C(n6984), .Y(n1380) );
  AOI22X1 U1465 ( .A(n1359), .B(n9450), .C(n1360), .D(n9286), .Y(n1387) );
  AOI22X1 U1467 ( .A(n1362), .B(n9491), .C(n1363), .D(n9409), .Y(n1385) );
  NAND3X1 U1469 ( .A(n6332), .B(n1389), .C(n1390), .Y(n5508) );
  NOR3X1 U1470 ( .A(n7031), .B(n7072), .C(n7113), .Y(n1390) );
  NAND3X1 U1472 ( .A(n4046), .B(n6654), .C(n6983), .Y(n1395) );
  AOI22X1 U1473 ( .A(n1354), .B(n9042), .C(n8486), .D(n8919), .Y(n1397) );
  NAND3X1 U1475 ( .A(n6287), .B(n6653), .C(n6982), .Y(n1394) );
  AOI22X1 U1476 ( .A(n1359), .B(n9124), .C(n1360), .D(n8960), .Y(n1400) );
  AOI22X1 U1478 ( .A(n1362), .B(n9165), .C(n1363), .D(n9083), .Y(n1398) );
  NAND3X1 U1480 ( .A(n1366), .B(n6652), .C(n6981), .Y(n1402) );
  AOI22X1 U1481 ( .A(n1354), .B(n8714), .C(n8486), .D(n8591), .Y(n1404) );
  NAND3X1 U1483 ( .A(n6286), .B(n6651), .C(n6980), .Y(n1401) );
  AOI22X1 U1484 ( .A(n1359), .B(n8796), .C(n1360), .D(n8632), .Y(n1407) );
  AOI22X1 U1486 ( .A(n1362), .B(n8837), .C(n1363), .D(n8755), .Y(n1405) );
  NAND3X1 U1488 ( .A(n1374), .B(n6650), .C(n6979), .Y(n1409) );
  AOI22X1 U1489 ( .A(n1354), .B(n9698), .C(n8484), .D(n9575), .Y(n1411) );
  NAND3X1 U1491 ( .A(n6285), .B(n6649), .C(n6978), .Y(n1408) );
  AOI22X1 U1492 ( .A(n1359), .B(n9780), .C(n1360), .D(n9616), .Y(n1414) );
  AOI22X1 U1494 ( .A(n1362), .B(n9821), .C(n1363), .D(n9739), .Y(n1412) );
  NAND3X1 U1495 ( .A(n1382), .B(n6648), .C(n6977), .Y(n1416) );
  AOI22X1 U1496 ( .A(n1354), .B(n9370), .C(n8488), .D(n9247), .Y(n1418) );
  NAND3X1 U1498 ( .A(n6284), .B(n6647), .C(n6976), .Y(n1415) );
  AOI22X1 U1499 ( .A(n1359), .B(n9452), .C(n1360), .D(n9288), .Y(n1421) );
  AOI22X1 U1501 ( .A(n1362), .B(n9493), .C(n1363), .D(n9411), .Y(n1419) );
  NAND3X1 U1503 ( .A(n6331), .B(n1423), .C(n1424), .Y(n5509) );
  NOR3X1 U1504 ( .A(n7030), .B(n7071), .C(n7112), .Y(n1424) );
  NAND3X1 U1506 ( .A(n4046), .B(n6646), .C(n6975), .Y(n1429) );
  AOI22X1 U1507 ( .A(n1354), .B(n9044), .C(n8491), .D(n8921), .Y(n1431) );
  NAND3X1 U1509 ( .A(n6283), .B(n6645), .C(n6974), .Y(n1428) );
  AOI22X1 U1510 ( .A(n1359), .B(n9126), .C(n1360), .D(n8962), .Y(n1434) );
  AOI22X1 U1512 ( .A(n1362), .B(n9167), .C(n1363), .D(n9085), .Y(n1432) );
  NAND3X1 U1514 ( .A(n1366), .B(n6644), .C(n6973), .Y(n1436) );
  AOI22X1 U1515 ( .A(n1354), .B(n8716), .C(n8487), .D(n8593), .Y(n1438) );
  NAND3X1 U1517 ( .A(n6282), .B(n6643), .C(n6972), .Y(n1435) );
  AOI22X1 U1518 ( .A(n1359), .B(n8798), .C(n1360), .D(n8634), .Y(n1441) );
  AOI22X1 U1520 ( .A(n1362), .B(n8839), .C(n1363), .D(n8757), .Y(n1439) );
  NAND3X1 U1522 ( .A(n1374), .B(n6642), .C(n6971), .Y(n1443) );
  AOI22X1 U1523 ( .A(n1354), .B(n9700), .C(n8483), .D(n9577), .Y(n1445) );
  NAND3X1 U1525 ( .A(n6281), .B(n6641), .C(n6970), .Y(n1442) );
  AOI22X1 U1526 ( .A(n1359), .B(n9782), .C(n1360), .D(n9618), .Y(n1448) );
  AOI22X1 U1528 ( .A(n1362), .B(n9823), .C(n1363), .D(n9741), .Y(n1446) );
  NAND3X1 U1529 ( .A(n1382), .B(n6640), .C(n6969), .Y(n1450) );
  AOI22X1 U1530 ( .A(n1354), .B(n9372), .C(n8490), .D(n9249), .Y(n1452) );
  NAND3X1 U1532 ( .A(n6280), .B(n6639), .C(n6968), .Y(n1449) );
  AOI22X1 U1533 ( .A(n1359), .B(n9454), .C(n1360), .D(n9290), .Y(n1455) );
  AOI22X1 U1535 ( .A(n1362), .B(n9495), .C(n1363), .D(n9413), .Y(n1453) );
  NAND3X1 U1537 ( .A(n6330), .B(n1457), .C(n1458), .Y(n5510) );
  NOR3X1 U1538 ( .A(n7029), .B(n7070), .C(n7111), .Y(n1458) );
  NAND3X1 U1540 ( .A(n4046), .B(n6638), .C(n6967), .Y(n1463) );
  AOI22X1 U1541 ( .A(n1354), .B(n9046), .C(n8485), .D(n8923), .Y(n1465) );
  NAND3X1 U1543 ( .A(n6279), .B(n6637), .C(n6966), .Y(n1462) );
  AOI22X1 U1544 ( .A(n1359), .B(n9128), .C(n1360), .D(n8964), .Y(n1468) );
  AOI22X1 U1546 ( .A(n1362), .B(n9169), .C(n1363), .D(n9087), .Y(n1466) );
  NAND3X1 U1548 ( .A(n1366), .B(n6636), .C(n6965), .Y(n1470) );
  AOI22X1 U1549 ( .A(n1354), .B(n8718), .C(n8489), .D(n8595), .Y(n1472) );
  NAND3X1 U1551 ( .A(n6278), .B(n6635), .C(n6964), .Y(n1469) );
  AOI22X1 U1552 ( .A(n1359), .B(n8800), .C(n1360), .D(n8636), .Y(n1475) );
  AOI22X1 U1554 ( .A(n1362), .B(n8841), .C(n1363), .D(n8759), .Y(n1473) );
  NAND3X1 U1556 ( .A(n1374), .B(n6634), .C(n6963), .Y(n1477) );
  AOI22X1 U1557 ( .A(n1354), .B(n9702), .C(n8483), .D(n9579), .Y(n1479) );
  NAND3X1 U1559 ( .A(n6277), .B(n6633), .C(n6962), .Y(n1476) );
  AOI22X1 U1560 ( .A(n1359), .B(n9784), .C(n1360), .D(n9620), .Y(n1482) );
  AOI22X1 U1562 ( .A(n1362), .B(n9825), .C(n1363), .D(n9743), .Y(n1480) );
  NAND3X1 U1563 ( .A(n1382), .B(n6632), .C(n6961), .Y(n1484) );
  AOI22X1 U1564 ( .A(n1354), .B(n9374), .C(n8491), .D(n9251), .Y(n1486) );
  NAND3X1 U1566 ( .A(n6276), .B(n6631), .C(n6960), .Y(n1483) );
  AOI22X1 U1567 ( .A(n1359), .B(n9456), .C(n1360), .D(n9292), .Y(n1489) );
  AOI22X1 U1569 ( .A(n1362), .B(n9497), .C(n1363), .D(n9415), .Y(n1487) );
  NAND3X1 U1571 ( .A(n6329), .B(n1491), .C(n1492), .Y(n5511) );
  NOR3X1 U1572 ( .A(n7028), .B(n7069), .C(n7110), .Y(n1492) );
  NAND3X1 U1574 ( .A(n4046), .B(n6630), .C(n6959), .Y(n1497) );
  AOI22X1 U1575 ( .A(n1354), .B(n9048), .C(n8486), .D(n8925), .Y(n1499) );
  NAND3X1 U1577 ( .A(n6275), .B(n6629), .C(n6958), .Y(n1496) );
  AOI22X1 U1578 ( .A(n1359), .B(n9130), .C(n1360), .D(n8966), .Y(n1502) );
  AOI22X1 U1580 ( .A(n1362), .B(n9171), .C(n1363), .D(n9089), .Y(n1500) );
  NAND3X1 U1582 ( .A(n1366), .B(n6628), .C(n6957), .Y(n1504) );
  AOI22X1 U1583 ( .A(n1354), .B(n8720), .C(n8488), .D(n8597), .Y(n1506) );
  NAND3X1 U1585 ( .A(n6274), .B(n6627), .C(n6956), .Y(n1503) );
  AOI22X1 U1586 ( .A(n1359), .B(n8802), .C(n1360), .D(n8638), .Y(n1509) );
  AOI22X1 U1588 ( .A(n1362), .B(n8843), .C(n1363), .D(n8761), .Y(n1507) );
  NAND3X1 U1590 ( .A(n1374), .B(n6626), .C(n6955), .Y(n1511) );
  AOI22X1 U1591 ( .A(n1354), .B(n9704), .C(n8483), .D(n9581), .Y(n1513) );
  NAND3X1 U1593 ( .A(n6273), .B(n6625), .C(n6954), .Y(n1510) );
  AOI22X1 U1594 ( .A(n1359), .B(n9786), .C(n1360), .D(n9622), .Y(n1516) );
  AOI22X1 U1596 ( .A(n1362), .B(n9827), .C(n1363), .D(n9745), .Y(n1514) );
  NAND3X1 U1597 ( .A(n1382), .B(n6624), .C(n6953), .Y(n1518) );
  AOI22X1 U1598 ( .A(n1354), .B(n9376), .C(n1355), .D(n9253), .Y(n1520) );
  NAND3X1 U1600 ( .A(n6272), .B(n6623), .C(n6952), .Y(n1517) );
  AOI22X1 U1601 ( .A(n1359), .B(n9458), .C(n1360), .D(n9294), .Y(n1523) );
  AOI22X1 U1603 ( .A(n1362), .B(n9499), .C(n1363), .D(n9417), .Y(n1521) );
  NAND3X1 U1605 ( .A(n6328), .B(n1525), .C(n1526), .Y(n5512) );
  NOR3X1 U1606 ( .A(n7027), .B(n7068), .C(n7109), .Y(n1526) );
  NAND3X1 U1608 ( .A(n4046), .B(n6622), .C(n6951), .Y(n1531) );
  AOI22X1 U1609 ( .A(n1354), .B(n9050), .C(n8490), .D(n8927), .Y(n1533) );
  NAND3X1 U1611 ( .A(n6271), .B(n6621), .C(n6950), .Y(n1530) );
  AOI22X1 U1612 ( .A(n1359), .B(n9132), .C(n1360), .D(n8968), .Y(n1536) );
  AOI22X1 U1614 ( .A(n1362), .B(n9173), .C(n1363), .D(n9091), .Y(n1534) );
  NAND3X1 U1616 ( .A(n1366), .B(n6620), .C(n6949), .Y(n1538) );
  AOI22X1 U1617 ( .A(n1354), .B(n8722), .C(n8491), .D(n8599), .Y(n1540) );
  NAND3X1 U1619 ( .A(n6270), .B(n6619), .C(n6948), .Y(n1537) );
  AOI22X1 U1620 ( .A(n1359), .B(n8804), .C(n1360), .D(n8640), .Y(n1543) );
  AOI22X1 U1622 ( .A(n1362), .B(n8845), .C(n1363), .D(n8763), .Y(n1541) );
  NAND3X1 U1624 ( .A(n1374), .B(n6618), .C(n6947), .Y(n1545) );
  AOI22X1 U1625 ( .A(n1354), .B(n9706), .C(n8484), .D(n9583), .Y(n1547) );
  NAND3X1 U1627 ( .A(n6269), .B(n6617), .C(n6946), .Y(n1544) );
  AOI22X1 U1628 ( .A(n1359), .B(n9788), .C(n1360), .D(n9624), .Y(n1550) );
  AOI22X1 U1630 ( .A(n1362), .B(n9829), .C(n1363), .D(n9747), .Y(n1548) );
  NAND3X1 U1631 ( .A(n1382), .B(n6616), .C(n6945), .Y(n1552) );
  AOI22X1 U1632 ( .A(n1354), .B(n9378), .C(n1355), .D(n9255), .Y(n1554) );
  NAND3X1 U1634 ( .A(n6268), .B(n6615), .C(n6944), .Y(n1551) );
  AOI22X1 U1635 ( .A(n1359), .B(n9460), .C(n1360), .D(n9296), .Y(n1557) );
  AOI22X1 U1637 ( .A(n1362), .B(n9501), .C(n1363), .D(n9419), .Y(n1555) );
  NAND3X1 U1639 ( .A(n6327), .B(n1559), .C(n1560), .Y(n5513) );
  NOR3X1 U1640 ( .A(n7026), .B(n7067), .C(n7108), .Y(n1560) );
  NAND3X1 U1642 ( .A(n4046), .B(n6614), .C(n6943), .Y(n1565) );
  AOI22X1 U1643 ( .A(n1354), .B(n9012), .C(n8487), .D(n8889), .Y(n1567) );
  NAND3X1 U1645 ( .A(n6267), .B(n6613), .C(n6942), .Y(n1564) );
  AOI22X1 U1646 ( .A(n1359), .B(n9094), .C(n1360), .D(n8930), .Y(n1570) );
  AOI22X1 U1648 ( .A(n1362), .B(n9135), .C(n1363), .D(n9053), .Y(n1568) );
  NAND3X1 U1650 ( .A(n1366), .B(n6612), .C(n6941), .Y(n1572) );
  AOI22X1 U1651 ( .A(n1354), .B(n8684), .C(n8486), .D(n8561), .Y(n1574) );
  NAND3X1 U1653 ( .A(n6266), .B(n6611), .C(n6940), .Y(n1571) );
  AOI22X1 U1654 ( .A(n1359), .B(n8766), .C(n1360), .D(n8602), .Y(n1577) );
  AOI22X1 U1656 ( .A(n1362), .B(n8807), .C(n1363), .D(n8725), .Y(n1575) );
  NAND3X1 U1658 ( .A(n1374), .B(n6610), .C(n6939), .Y(n1579) );
  AOI22X1 U1659 ( .A(n1354), .B(n9668), .C(n8489), .D(n9545), .Y(n1581) );
  NAND3X1 U1661 ( .A(n6265), .B(n6609), .C(n6938), .Y(n1578) );
  AOI22X1 U1662 ( .A(n1359), .B(n9750), .C(n1360), .D(n9586), .Y(n1584) );
  AOI22X1 U1664 ( .A(n1362), .B(n9791), .C(n1363), .D(n9709), .Y(n1582) );
  NAND3X1 U1665 ( .A(n1382), .B(n6608), .C(n6937), .Y(n1586) );
  AOI22X1 U1666 ( .A(n1354), .B(n9340), .C(n1355), .D(n9217), .Y(n1588) );
  NAND3X1 U1668 ( .A(n6264), .B(n6607), .C(n6936), .Y(n1585) );
  AOI22X1 U1669 ( .A(n1359), .B(n9422), .C(n1360), .D(n9258), .Y(n1591) );
  AOI22X1 U1671 ( .A(n1362), .B(n9463), .C(n1363), .D(n9381), .Y(n1589) );
  NAND3X1 U1673 ( .A(n6326), .B(n1593), .C(n1594), .Y(n5514) );
  NOR3X1 U1674 ( .A(n7025), .B(n7066), .C(n7107), .Y(n1594) );
  NAND3X1 U1676 ( .A(n4046), .B(n6606), .C(n6935), .Y(n1599) );
  AOI22X1 U1677 ( .A(n1354), .B(n9015), .C(n8485), .D(n8892), .Y(n1601) );
  NAND3X1 U1679 ( .A(n6263), .B(n6605), .C(n6934), .Y(n1598) );
  AOI22X1 U1680 ( .A(n1359), .B(n9097), .C(n1360), .D(n8933), .Y(n1604) );
  AOI22X1 U1682 ( .A(n1362), .B(n9138), .C(n1363), .D(n9056), .Y(n1602) );
  NAND3X1 U1684 ( .A(n1366), .B(n6604), .C(n6933), .Y(n1606) );
  AOI22X1 U1685 ( .A(n1354), .B(n8687), .C(n8491), .D(n8564), .Y(n1608) );
  NAND3X1 U1687 ( .A(n6262), .B(n6603), .C(n6932), .Y(n1605) );
  AOI22X1 U1688 ( .A(n1359), .B(n8769), .C(n1360), .D(n8605), .Y(n1611) );
  AOI22X1 U1690 ( .A(n1362), .B(n8810), .C(n1363), .D(n8728), .Y(n1609) );
  NAND3X1 U1692 ( .A(n1374), .B(n6602), .C(n6931), .Y(n1613) );
  AOI22X1 U1693 ( .A(n1354), .B(n9671), .C(n8488), .D(n9548), .Y(n1615) );
  NAND3X1 U1695 ( .A(n6261), .B(n6601), .C(n6930), .Y(n1612) );
  AOI22X1 U1696 ( .A(n1359), .B(n9753), .C(n1360), .D(n9589), .Y(n1618) );
  AOI22X1 U1698 ( .A(n1362), .B(n9794), .C(n1363), .D(n9712), .Y(n1616) );
  NAND3X1 U1699 ( .A(n1382), .B(n6600), .C(n6929), .Y(n1620) );
  AOI22X1 U1700 ( .A(n1354), .B(n9343), .C(n1355), .D(n9220), .Y(n1622) );
  NAND3X1 U1702 ( .A(n6260), .B(n6599), .C(n6928), .Y(n1619) );
  AOI22X1 U1703 ( .A(n1359), .B(n9425), .C(n1360), .D(n9261), .Y(n1625) );
  AOI22X1 U1705 ( .A(n1362), .B(n9466), .C(n1363), .D(n9384), .Y(n1623) );
  NAND3X1 U1707 ( .A(n6325), .B(n1627), .C(n1628), .Y(n5515) );
  NOR3X1 U1708 ( .A(n7024), .B(n7065), .C(n7106), .Y(n1628) );
  NAND3X1 U1710 ( .A(n4046), .B(n6598), .C(n6927), .Y(n1633) );
  AOI22X1 U1711 ( .A(n1354), .B(n9016), .C(n8490), .D(n8893), .Y(n1635) );
  NAND3X1 U1713 ( .A(n6259), .B(n6597), .C(n6926), .Y(n1632) );
  AOI22X1 U1714 ( .A(n1359), .B(n9098), .C(n1360), .D(n8934), .Y(n1638) );
  AOI22X1 U1716 ( .A(n1362), .B(n9139), .C(n1363), .D(n9057), .Y(n1636) );
  NAND3X1 U1718 ( .A(n1366), .B(n6596), .C(n6925), .Y(n1640) );
  AOI22X1 U1719 ( .A(n1354), .B(n8688), .C(n8491), .D(n8565), .Y(n1642) );
  NAND3X1 U1721 ( .A(n6258), .B(n6595), .C(n6924), .Y(n1639) );
  AOI22X1 U1722 ( .A(n1359), .B(n8770), .C(n1360), .D(n8606), .Y(n1645) );
  AOI22X1 U1724 ( .A(n1362), .B(n8811), .C(n1363), .D(n8729), .Y(n1643) );
  NAND3X1 U1726 ( .A(n1374), .B(n6594), .C(n6923), .Y(n1647) );
  AOI22X1 U1727 ( .A(n1354), .B(n9672), .C(n8489), .D(n9549), .Y(n1649) );
  NAND3X1 U1729 ( .A(n6257), .B(n6593), .C(n6922), .Y(n1646) );
  AOI22X1 U1730 ( .A(n1359), .B(n9754), .C(n1360), .D(n9590), .Y(n1652) );
  AOI22X1 U1732 ( .A(n1362), .B(n9795), .C(n1363), .D(n9713), .Y(n1650) );
  NAND3X1 U1733 ( .A(n1382), .B(n6592), .C(n6921), .Y(n1654) );
  AOI22X1 U1734 ( .A(n1354), .B(n9344), .C(n8486), .D(n9221), .Y(n1656) );
  NAND3X1 U1736 ( .A(n6256), .B(n6591), .C(n6920), .Y(n1653) );
  AOI22X1 U1737 ( .A(n1359), .B(n9426), .C(n1360), .D(n9262), .Y(n1659) );
  AOI22X1 U1739 ( .A(n1362), .B(n9467), .C(n1363), .D(n9385), .Y(n1657) );
  NAND3X1 U1741 ( .A(n6324), .B(n1661), .C(n1662), .Y(n5516) );
  NOR3X1 U1742 ( .A(n7023), .B(n7064), .C(n7105), .Y(n1662) );
  NAND3X1 U1744 ( .A(n4046), .B(n6590), .C(n6919), .Y(n1667) );
  AOI22X1 U1745 ( .A(n1354), .B(n9017), .C(n8491), .D(n8894), .Y(n1669) );
  NAND3X1 U1747 ( .A(n6255), .B(n6589), .C(n6918), .Y(n1666) );
  AOI22X1 U1748 ( .A(n1359), .B(n9099), .C(n8469), .D(n8935), .Y(n1672) );
  AOI22X1 U1750 ( .A(n1362), .B(n9140), .C(n8437), .D(n9058), .Y(n1670) );
  NAND3X1 U1752 ( .A(n1366), .B(n6588), .C(n6917), .Y(n1674) );
  AOI22X1 U1753 ( .A(n1354), .B(n8689), .C(n8489), .D(n8566), .Y(n1676) );
  NAND3X1 U1755 ( .A(n6254), .B(n6587), .C(n6916), .Y(n1673) );
  AOI22X1 U1756 ( .A(n1359), .B(n8771), .C(n8468), .D(n8607), .Y(n1679) );
  AOI22X1 U1758 ( .A(n1362), .B(n8812), .C(n8439), .D(n8730), .Y(n1677) );
  NAND3X1 U1760 ( .A(n1374), .B(n6586), .C(n6915), .Y(n1681) );
  AOI22X1 U1761 ( .A(n1354), .B(n9673), .C(n8488), .D(n9550), .Y(n1683) );
  NAND3X1 U1763 ( .A(n6253), .B(n6585), .C(n6914), .Y(n1680) );
  AOI22X1 U1764 ( .A(n1359), .B(n9755), .C(n1360), .D(n9591), .Y(n1686) );
  AOI22X1 U1766 ( .A(n1362), .B(n9796), .C(n1363), .D(n9714), .Y(n1684) );
  NAND3X1 U1767 ( .A(n1382), .B(n6584), .C(n6913), .Y(n1688) );
  AOI22X1 U1768 ( .A(n8492), .B(n9345), .C(n8484), .D(n9222), .Y(n1690) );
  NAND3X1 U1770 ( .A(n6252), .B(n6583), .C(n6912), .Y(n1687) );
  AOI22X1 U1771 ( .A(n8477), .B(n9427), .C(n8465), .D(n9263), .Y(n1693) );
  AOI22X1 U1773 ( .A(n8446), .B(n9468), .C(n8438), .D(n9386), .Y(n1691) );
  NAND3X1 U1775 ( .A(n6323), .B(n1695), .C(n1696), .Y(n5517) );
  NOR3X1 U1776 ( .A(n7022), .B(n7063), .C(n7104), .Y(n1696) );
  NAND3X1 U1778 ( .A(n4046), .B(n6582), .C(n6911), .Y(n1701) );
  AOI22X1 U1779 ( .A(n8496), .B(n9018), .C(n8485), .D(n8895), .Y(n1703) );
  NAND3X1 U1781 ( .A(n6251), .B(n6581), .C(n6910), .Y(n1700) );
  AOI22X1 U1782 ( .A(n8479), .B(n9100), .C(n8470), .D(n8936), .Y(n1706) );
  AOI22X1 U1784 ( .A(n8451), .B(n9141), .C(n8442), .D(n9059), .Y(n1704) );
  NAND3X1 U1786 ( .A(n1366), .B(n6580), .C(n6909), .Y(n1708) );
  AOI22X1 U1787 ( .A(n8498), .B(n8690), .C(n8488), .D(n8567), .Y(n1710) );
  NAND3X1 U1789 ( .A(n6250), .B(n6579), .C(n6908), .Y(n1707) );
  AOI22X1 U1790 ( .A(n8478), .B(n8772), .C(n8472), .D(n8608), .Y(n1713) );
  AOI22X1 U1792 ( .A(n8447), .B(n8813), .C(n8435), .D(n8731), .Y(n1711) );
  NAND3X1 U1794 ( .A(n1374), .B(n6578), .C(n6907), .Y(n1715) );
  AOI22X1 U1795 ( .A(n8495), .B(n9674), .C(n8490), .D(n9551), .Y(n1717) );
  NAND3X1 U1797 ( .A(n6249), .B(n6577), .C(n6906), .Y(n1714) );
  AOI22X1 U1798 ( .A(n8474), .B(n9756), .C(n8467), .D(n9592), .Y(n1720) );
  AOI22X1 U1800 ( .A(n8449), .B(n9797), .C(n8438), .D(n9715), .Y(n1718) );
  NAND3X1 U1801 ( .A(n1382), .B(n6576), .C(n6905), .Y(n1722) );
  AOI22X1 U1802 ( .A(n8493), .B(n9346), .C(n8487), .D(n9223), .Y(n1724) );
  NAND3X1 U1804 ( .A(n6248), .B(n6575), .C(n6904), .Y(n1721) );
  AOI22X1 U1805 ( .A(n8476), .B(n9428), .C(n8467), .D(n9264), .Y(n1727) );
  AOI22X1 U1807 ( .A(n8445), .B(n9469), .C(n8440), .D(n9387), .Y(n1725) );
  NAND3X1 U1809 ( .A(n6322), .B(n1729), .C(n1730), .Y(n5518) );
  NOR3X1 U1810 ( .A(n7021), .B(n7062), .C(n7103), .Y(n1730) );
  NAND3X1 U1812 ( .A(n4046), .B(n6574), .C(n6903), .Y(n1735) );
  AOI22X1 U1813 ( .A(n8494), .B(n9019), .C(n8491), .D(n8896), .Y(n1737) );
  NAND3X1 U1815 ( .A(n6247), .B(n6573), .C(n6902), .Y(n1734) );
  AOI22X1 U1816 ( .A(n8480), .B(n9101), .C(n8471), .D(n8937), .Y(n1740) );
  AOI22X1 U1818 ( .A(n8452), .B(n9142), .C(n8443), .D(n9060), .Y(n1738) );
  NAND3X1 U1820 ( .A(n1366), .B(n6572), .C(n6901), .Y(n1742) );
  AOI22X1 U1821 ( .A(n8497), .B(n8691), .C(n8491), .D(n8568), .Y(n1744) );
  NAND3X1 U1823 ( .A(n6246), .B(n6571), .C(n6900), .Y(n1741) );
  AOI22X1 U1824 ( .A(n8477), .B(n8773), .C(n8465), .D(n8609), .Y(n1747) );
  AOI22X1 U1826 ( .A(n8446), .B(n8814), .C(n8436), .D(n8732), .Y(n1745) );
  NAND3X1 U1828 ( .A(n1374), .B(n6570), .C(n6899), .Y(n1749) );
  AOI22X1 U1829 ( .A(n8492), .B(n9675), .C(n8491), .D(n9552), .Y(n1751) );
  NAND3X1 U1831 ( .A(n6245), .B(n6569), .C(n6898), .Y(n1748) );
  AOI22X1 U1832 ( .A(n8475), .B(n9757), .C(n8466), .D(n9593), .Y(n1754) );
  AOI22X1 U1834 ( .A(n8448), .B(n9798), .C(n8440), .D(n9716), .Y(n1752) );
  NAND3X1 U1835 ( .A(n1382), .B(n6568), .C(n6897), .Y(n1756) );
  AOI22X1 U1836 ( .A(n8498), .B(n9347), .C(n8491), .D(n9224), .Y(n1758) );
  NAND3X1 U1838 ( .A(n6244), .B(n6567), .C(n6896), .Y(n1755) );
  AOI22X1 U1839 ( .A(n8474), .B(n9429), .C(n8466), .D(n9265), .Y(n1761) );
  AOI22X1 U1841 ( .A(n8449), .B(n9470), .C(n8441), .D(n9388), .Y(n1759) );
  NAND3X1 U1843 ( .A(n6321), .B(n1763), .C(n1764), .Y(n5519) );
  NOR3X1 U1844 ( .A(n7020), .B(n7061), .C(n7102), .Y(n1764) );
  NAND3X1 U1846 ( .A(n4046), .B(n6566), .C(n6895), .Y(n1769) );
  AOI22X1 U1847 ( .A(n8495), .B(n9020), .C(n8491), .D(n8897), .Y(n1771) );
  NAND3X1 U1849 ( .A(n6243), .B(n6565), .C(n6894), .Y(n1768) );
  AOI22X1 U1850 ( .A(n8474), .B(n9102), .C(n8464), .D(n8938), .Y(n1774) );
  AOI22X1 U1852 ( .A(n8450), .B(n9143), .C(n8435), .D(n9061), .Y(n1772) );
  NAND3X1 U1854 ( .A(n1366), .B(n6564), .C(n6893), .Y(n1776) );
  AOI22X1 U1855 ( .A(n8496), .B(n8692), .C(n8491), .D(n8569), .Y(n1778) );
  NAND3X1 U1857 ( .A(n6242), .B(n6563), .C(n6892), .Y(n1775) );
  AOI22X1 U1858 ( .A(n8476), .B(n8774), .C(n8464), .D(n8610), .Y(n1781) );
  AOI22X1 U1860 ( .A(n8445), .B(n8815), .C(n8435), .D(n8733), .Y(n1779) );
  NAND3X1 U1862 ( .A(n1374), .B(n6562), .C(n6891), .Y(n1783) );
  AOI22X1 U1863 ( .A(n8493), .B(n9676), .C(n8491), .D(n9553), .Y(n1785) );
  NAND3X1 U1865 ( .A(n6241), .B(n6561), .C(n6890), .Y(n1782) );
  AOI22X1 U1866 ( .A(n1359), .B(n9758), .C(n8464), .D(n9594), .Y(n1788) );
  AOI22X1 U1868 ( .A(n1362), .B(n9799), .C(n8435), .D(n9717), .Y(n1786) );
  NAND3X1 U1869 ( .A(n1382), .B(n6560), .C(n6889), .Y(n1790) );
  AOI22X1 U1870 ( .A(n8497), .B(n9348), .C(n8491), .D(n9225), .Y(n1792) );
  NAND3X1 U1872 ( .A(n6240), .B(n6559), .C(n6888), .Y(n1789) );
  AOI22X1 U1873 ( .A(n8475), .B(n9430), .C(n8464), .D(n9266), .Y(n1795) );
  AOI22X1 U1875 ( .A(n8448), .B(n9471), .C(n8435), .D(n9389), .Y(n1793) );
  NAND3X1 U1877 ( .A(n6320), .B(n1797), .C(n1798), .Y(n5520) );
  NOR3X1 U1878 ( .A(n7019), .B(n7060), .C(n7101), .Y(n1798) );
  NAND3X1 U1880 ( .A(n4046), .B(n6558), .C(n6887), .Y(n1803) );
  AOI22X1 U1881 ( .A(n8492), .B(n9021), .C(n8491), .D(n8898), .Y(n1805) );
  NAND3X1 U1883 ( .A(n6239), .B(n6557), .C(n6886), .Y(n1802) );
  AOI22X1 U1884 ( .A(n8474), .B(n9103), .C(n8464), .D(n8939), .Y(n1808) );
  AOI22X1 U1886 ( .A(n8445), .B(n9144), .C(n8435), .D(n9062), .Y(n1806) );
  NAND3X1 U1888 ( .A(n1366), .B(n6556), .C(n6885), .Y(n1810) );
  AOI22X1 U1889 ( .A(n8492), .B(n8693), .C(n8491), .D(n8570), .Y(n1812) );
  NAND3X1 U1891 ( .A(n6238), .B(n6555), .C(n6884), .Y(n1809) );
  AOI22X1 U1892 ( .A(n8474), .B(n8775), .C(n8464), .D(n8611), .Y(n1815) );
  AOI22X1 U1894 ( .A(n8445), .B(n8816), .C(n8435), .D(n8734), .Y(n1813) );
  NAND3X1 U1896 ( .A(n1374), .B(n6554), .C(n6883), .Y(n1817) );
  AOI22X1 U1897 ( .A(n8492), .B(n9677), .C(n8491), .D(n9554), .Y(n1819) );
  NAND3X1 U1899 ( .A(n6237), .B(n6553), .C(n6882), .Y(n1816) );
  AOI22X1 U1900 ( .A(n8474), .B(n9759), .C(n8464), .D(n9595), .Y(n1822) );
  AOI22X1 U1902 ( .A(n8445), .B(n9800), .C(n8435), .D(n9718), .Y(n1820) );
  NAND3X1 U1903 ( .A(n1382), .B(n6552), .C(n6881), .Y(n1824) );
  AOI22X1 U1904 ( .A(n8492), .B(n9349), .C(n8491), .D(n9226), .Y(n1826) );
  NAND3X1 U1906 ( .A(n6236), .B(n6551), .C(n6880), .Y(n1823) );
  AOI22X1 U1907 ( .A(n8474), .B(n9431), .C(n8464), .D(n9267), .Y(n1829) );
  AOI22X1 U1909 ( .A(n8445), .B(n9472), .C(n8435), .D(n9390), .Y(n1827) );
  NAND3X1 U1911 ( .A(n6319), .B(n1831), .C(n1832), .Y(n5521) );
  NOR3X1 U1912 ( .A(n7018), .B(n7059), .C(n7100), .Y(n1832) );
  NAND3X1 U1914 ( .A(n4046), .B(n6550), .C(n6879), .Y(n1837) );
  AOI22X1 U1915 ( .A(n8492), .B(n9022), .C(n8490), .D(n8899), .Y(n1839) );
  NAND3X1 U1917 ( .A(n6235), .B(n6549), .C(n6878), .Y(n1836) );
  AOI22X1 U1918 ( .A(n8474), .B(n9104), .C(n8464), .D(n8940), .Y(n3164) );
  AOI22X1 U1920 ( .A(n8445), .B(n9145), .C(n8435), .D(n9063), .Y(n1840) );
  NAND3X1 U1922 ( .A(n1366), .B(n6548), .C(n6877), .Y(n3166) );
  AOI22X1 U1923 ( .A(n8492), .B(n8694), .C(n8490), .D(n8571), .Y(n3168) );
  NAND3X1 U1925 ( .A(n6234), .B(n6547), .C(n6876), .Y(n3165) );
  AOI22X1 U1926 ( .A(n8474), .B(n8776), .C(n8464), .D(n8612), .Y(n3171) );
  AOI22X1 U1928 ( .A(n8445), .B(n8817), .C(n8435), .D(n8735), .Y(n3169) );
  NAND3X1 U1930 ( .A(n1374), .B(n6546), .C(n6875), .Y(n3173) );
  AOI22X1 U1931 ( .A(n8492), .B(n9678), .C(n8490), .D(n9555), .Y(n3175) );
  NAND3X1 U1933 ( .A(n6233), .B(n6545), .C(n6874), .Y(n3172) );
  AOI22X1 U1934 ( .A(n8474), .B(n9760), .C(n8464), .D(n9596), .Y(n3178) );
  AOI22X1 U1936 ( .A(n8445), .B(n9801), .C(n8435), .D(n9719), .Y(n3176) );
  NAND3X1 U1937 ( .A(n1382), .B(n6544), .C(n6873), .Y(n3180) );
  AOI22X1 U1938 ( .A(n8492), .B(n9350), .C(n8490), .D(n9227), .Y(n3182) );
  NAND3X1 U1940 ( .A(n6232), .B(n6543), .C(n6872), .Y(n3179) );
  AOI22X1 U1941 ( .A(n8474), .B(n9432), .C(n8464), .D(n9268), .Y(n3185) );
  AOI22X1 U1943 ( .A(n8445), .B(n9473), .C(n8435), .D(n9391), .Y(n3183) );
  NAND3X1 U1945 ( .A(n6318), .B(n3187), .C(n3188), .Y(n5522) );
  NOR3X1 U1946 ( .A(n7017), .B(n7058), .C(n7099), .Y(n3188) );
  NAND3X1 U1948 ( .A(n4046), .B(n6542), .C(n6871), .Y(n3193) );
  AOI22X1 U1949 ( .A(n8492), .B(n9023), .C(n8490), .D(n8900), .Y(n3195) );
  NAND3X1 U1951 ( .A(n6231), .B(n6541), .C(n6870), .Y(n3192) );
  AOI22X1 U1952 ( .A(n8474), .B(n9105), .C(n8465), .D(n8941), .Y(n3198) );
  AOI22X1 U1954 ( .A(n8445), .B(n9146), .C(n8436), .D(n9064), .Y(n3196) );
  NAND3X1 U1956 ( .A(n1366), .B(n6540), .C(n6869), .Y(n3200) );
  AOI22X1 U1957 ( .A(n8492), .B(n8695), .C(n8490), .D(n8572), .Y(n3202) );
  NAND3X1 U1959 ( .A(n6230), .B(n6539), .C(n6868), .Y(n3199) );
  AOI22X1 U1960 ( .A(n8474), .B(n8777), .C(n8465), .D(n8613), .Y(n3205) );
  AOI22X1 U1962 ( .A(n8445), .B(n8818), .C(n8436), .D(n8736), .Y(n3203) );
  NAND3X1 U1964 ( .A(n1374), .B(n6538), .C(n6867), .Y(n3207) );
  AOI22X1 U1965 ( .A(n8492), .B(n9679), .C(n8490), .D(n9556), .Y(n3209) );
  NAND3X1 U1967 ( .A(n6229), .B(n6537), .C(n6866), .Y(n3206) );
  AOI22X1 U1968 ( .A(n8474), .B(n9761), .C(n8465), .D(n9597), .Y(n3212) );
  AOI22X1 U1970 ( .A(n8445), .B(n9802), .C(n8436), .D(n9720), .Y(n3210) );
  NAND3X1 U1971 ( .A(n1382), .B(n6536), .C(n6865), .Y(n3214) );
  AOI22X1 U1972 ( .A(n8492), .B(n9351), .C(n8490), .D(n9228), .Y(n3216) );
  NAND3X1 U1974 ( .A(n6228), .B(n6535), .C(n6864), .Y(n3213) );
  AOI22X1 U1975 ( .A(n8474), .B(n9433), .C(n8465), .D(n9269), .Y(n3219) );
  AOI22X1 U1977 ( .A(n8445), .B(n9474), .C(n8436), .D(n9392), .Y(n3217) );
  NAND3X1 U1979 ( .A(n6317), .B(n3221), .C(n3222), .Y(n5523) );
  NOR3X1 U1980 ( .A(n7016), .B(n7057), .C(n7098), .Y(n3222) );
  NAND3X1 U1982 ( .A(n4046), .B(n6534), .C(n6863), .Y(n3227) );
  AOI22X1 U1983 ( .A(n8492), .B(n9024), .C(n8490), .D(n8901), .Y(n3229) );
  NAND3X1 U1985 ( .A(n6227), .B(n6533), .C(n6862), .Y(n3226) );
  AOI22X1 U1986 ( .A(n8474), .B(n9106), .C(n8465), .D(n8942), .Y(n3232) );
  AOI22X1 U1988 ( .A(n8445), .B(n9147), .C(n8436), .D(n9065), .Y(n3230) );
  NAND3X1 U1990 ( .A(n1366), .B(n6532), .C(n6861), .Y(n3234) );
  AOI22X1 U1991 ( .A(n8493), .B(n8696), .C(n8490), .D(n8573), .Y(n3236) );
  NAND3X1 U1993 ( .A(n6226), .B(n6531), .C(n6860), .Y(n3233) );
  AOI22X1 U1994 ( .A(n8475), .B(n8778), .C(n8465), .D(n8614), .Y(n3239) );
  AOI22X1 U1996 ( .A(n8446), .B(n8819), .C(n8436), .D(n8737), .Y(n3237) );
  NAND3X1 U1998 ( .A(n1374), .B(n6530), .C(n6859), .Y(n3241) );
  AOI22X1 U1999 ( .A(n8493), .B(n9680), .C(n8490), .D(n9557), .Y(n3243) );
  NAND3X1 U2001 ( .A(n6225), .B(n6529), .C(n6858), .Y(n3240) );
  AOI22X1 U2002 ( .A(n8475), .B(n9762), .C(n8465), .D(n9598), .Y(n3246) );
  AOI22X1 U2004 ( .A(n8446), .B(n9803), .C(n8436), .D(n9721), .Y(n3244) );
  NAND3X1 U2005 ( .A(n1382), .B(n6528), .C(n6857), .Y(n3248) );
  AOI22X1 U2006 ( .A(n8493), .B(n9352), .C(n8490), .D(n9229), .Y(n3250) );
  NAND3X1 U2008 ( .A(n6224), .B(n6527), .C(n6856), .Y(n3247) );
  AOI22X1 U2009 ( .A(n8475), .B(n9434), .C(n8465), .D(n9270), .Y(n3253) );
  AOI22X1 U2011 ( .A(n8446), .B(n9475), .C(n8436), .D(n9393), .Y(n3251) );
  NAND3X1 U2013 ( .A(n6316), .B(n3255), .C(n3256), .Y(n5524) );
  NOR3X1 U2014 ( .A(n7015), .B(n7056), .C(n7097), .Y(n3256) );
  NAND3X1 U2016 ( .A(n4046), .B(n6526), .C(n6855), .Y(n3261) );
  AOI22X1 U2017 ( .A(n8493), .B(n9025), .C(n8489), .D(n8902), .Y(n3263) );
  NAND3X1 U2019 ( .A(n6223), .B(n6525), .C(n6854), .Y(n3260) );
  AOI22X1 U2020 ( .A(n8475), .B(n9107), .C(n8465), .D(n8943), .Y(n3266) );
  AOI22X1 U2022 ( .A(n8446), .B(n9148), .C(n8436), .D(n9066), .Y(n3264) );
  NAND3X1 U2024 ( .A(n1366), .B(n6524), .C(n6853), .Y(n3268) );
  AOI22X1 U2025 ( .A(n8493), .B(n8697), .C(n8489), .D(n8574), .Y(n3270) );
  NAND3X1 U2027 ( .A(n6222), .B(n6523), .C(n6852), .Y(n3267) );
  AOI22X1 U2028 ( .A(n8475), .B(n8779), .C(n8465), .D(n8615), .Y(n3273) );
  AOI22X1 U2030 ( .A(n8446), .B(n8820), .C(n8436), .D(n8738), .Y(n3271) );
  NAND3X1 U2032 ( .A(n1374), .B(n6522), .C(n6851), .Y(n3275) );
  AOI22X1 U2033 ( .A(n8493), .B(n9681), .C(n8489), .D(n9558), .Y(n3277) );
  NAND3X1 U2035 ( .A(n6221), .B(n6521), .C(n6850), .Y(n3274) );
  AOI22X1 U2036 ( .A(n8475), .B(n9763), .C(n8465), .D(n9599), .Y(n3280) );
  AOI22X1 U2038 ( .A(n8446), .B(n9804), .C(n8436), .D(n9722), .Y(n3278) );
  NAND3X1 U2039 ( .A(n1382), .B(n6520), .C(n6849), .Y(n3282) );
  AOI22X1 U2040 ( .A(n8493), .B(n9353), .C(n8489), .D(n9230), .Y(n3284) );
  NAND3X1 U2042 ( .A(n6220), .B(n6519), .C(n6848), .Y(n3281) );
  AOI22X1 U2043 ( .A(n8475), .B(n9435), .C(n8465), .D(n9271), .Y(n3287) );
  AOI22X1 U2045 ( .A(n8446), .B(n9476), .C(n8436), .D(n9394), .Y(n3285) );
  NAND3X1 U2047 ( .A(n6315), .B(n3289), .C(n3290), .Y(n5525) );
  NOR3X1 U2048 ( .A(n7014), .B(n7055), .C(n7096), .Y(n3290) );
  NAND3X1 U2050 ( .A(n4046), .B(n6518), .C(n6847), .Y(n3295) );
  AOI22X1 U2051 ( .A(n8493), .B(n9026), .C(n8489), .D(n8903), .Y(n3297) );
  NAND3X1 U2053 ( .A(n6219), .B(n6517), .C(n6846), .Y(n3294) );
  AOI22X1 U2054 ( .A(n8475), .B(n9108), .C(n8466), .D(n8944), .Y(n3300) );
  AOI22X1 U2056 ( .A(n8446), .B(n9149), .C(n8437), .D(n9067), .Y(n3298) );
  NAND3X1 U2058 ( .A(n1366), .B(n6516), .C(n6845), .Y(n3302) );
  AOI22X1 U2059 ( .A(n8493), .B(n8698), .C(n8489), .D(n8575), .Y(n3304) );
  NAND3X1 U2061 ( .A(n6218), .B(n6515), .C(n6844), .Y(n3301) );
  AOI22X1 U2062 ( .A(n8475), .B(n8780), .C(n8466), .D(n8616), .Y(n3307) );
  AOI22X1 U2064 ( .A(n8446), .B(n8821), .C(n8437), .D(n8739), .Y(n3305) );
  NAND3X1 U2066 ( .A(n1374), .B(n6514), .C(n6843), .Y(n3309) );
  AOI22X1 U2067 ( .A(n8493), .B(n9682), .C(n8489), .D(n9559), .Y(n3311) );
  NAND3X1 U2069 ( .A(n6217), .B(n6513), .C(n6842), .Y(n3308) );
  AOI22X1 U2070 ( .A(n8475), .B(n9764), .C(n8466), .D(n9600), .Y(n3314) );
  AOI22X1 U2072 ( .A(n8446), .B(n9805), .C(n8437), .D(n9723), .Y(n3312) );
  NAND3X1 U2073 ( .A(n1382), .B(n6512), .C(n6841), .Y(n3316) );
  AOI22X1 U2074 ( .A(n8493), .B(n9354), .C(n8489), .D(n9231), .Y(n3318) );
  NAND3X1 U2076 ( .A(n6216), .B(n6511), .C(n6840), .Y(n3315) );
  AOI22X1 U2077 ( .A(n8475), .B(n9436), .C(n8466), .D(n9272), .Y(n3321) );
  AOI22X1 U2079 ( .A(n8446), .B(n9477), .C(n8437), .D(n9395), .Y(n3319) );
  NAND3X1 U2081 ( .A(n6314), .B(n3323), .C(n3324), .Y(n5526) );
  NOR3X1 U2082 ( .A(n7013), .B(n7054), .C(n7095), .Y(n3324) );
  NAND3X1 U2084 ( .A(n4046), .B(n6510), .C(n6839), .Y(n3329) );
  AOI22X1 U2085 ( .A(n8493), .B(n9027), .C(n8489), .D(n8904), .Y(n3331) );
  NAND3X1 U2087 ( .A(n6215), .B(n6509), .C(n6838), .Y(n3328) );
  AOI22X1 U2088 ( .A(n8475), .B(n9109), .C(n8466), .D(n8945), .Y(n3334) );
  AOI22X1 U2090 ( .A(n8446), .B(n9150), .C(n8437), .D(n9068), .Y(n3332) );
  NAND3X1 U2092 ( .A(n1366), .B(n6508), .C(n6837), .Y(n3336) );
  AOI22X1 U2093 ( .A(n8493), .B(n8699), .C(n8489), .D(n8576), .Y(n3338) );
  NAND3X1 U2095 ( .A(n6214), .B(n6507), .C(n6836), .Y(n3335) );
  AOI22X1 U2096 ( .A(n8475), .B(n8781), .C(n8466), .D(n8617), .Y(n3341) );
  AOI22X1 U2098 ( .A(n8446), .B(n8822), .C(n8437), .D(n8740), .Y(n3339) );
  NAND3X1 U2100 ( .A(n1374), .B(n6506), .C(n6835), .Y(n3343) );
  AOI22X1 U2101 ( .A(n8496), .B(n9683), .C(n8489), .D(n9560), .Y(n3345) );
  NAND3X1 U2103 ( .A(n6213), .B(n6505), .C(n6834), .Y(n3342) );
  AOI22X1 U2104 ( .A(n8476), .B(n9765), .C(n8466), .D(n9601), .Y(n3348) );
  AOI22X1 U2106 ( .A(n8447), .B(n9806), .C(n8437), .D(n9724), .Y(n3346) );
  NAND3X1 U2107 ( .A(n1382), .B(n6504), .C(n6833), .Y(n3350) );
  AOI22X1 U2108 ( .A(n8498), .B(n9355), .C(n8489), .D(n9232), .Y(n3352) );
  NAND3X1 U2110 ( .A(n6212), .B(n6503), .C(n6832), .Y(n3349) );
  AOI22X1 U2111 ( .A(n8476), .B(n9437), .C(n8466), .D(n9273), .Y(n3355) );
  AOI22X1 U2113 ( .A(n8447), .B(n9478), .C(n8437), .D(n9396), .Y(n3353) );
  NAND3X1 U2115 ( .A(n6313), .B(n3357), .C(n3358), .Y(n5527) );
  NOR3X1 U2116 ( .A(n7012), .B(n7053), .C(n7094), .Y(n3358) );
  NAND3X1 U2118 ( .A(n4046), .B(n6502), .C(n6831), .Y(n3363) );
  AOI22X1 U2119 ( .A(n8494), .B(n9013), .C(n8488), .D(n8890), .Y(n3365) );
  NAND3X1 U2121 ( .A(n6211), .B(n6501), .C(n6830), .Y(n3362) );
  AOI22X1 U2122 ( .A(n8476), .B(n9095), .C(n8466), .D(n8931), .Y(n3368) );
  AOI22X1 U2124 ( .A(n8447), .B(n9136), .C(n8437), .D(n9054), .Y(n3366) );
  NAND3X1 U2126 ( .A(n1366), .B(n6500), .C(n6829), .Y(n3370) );
  AOI22X1 U2127 ( .A(n8493), .B(n8685), .C(n8488), .D(n8562), .Y(n3372) );
  NAND3X1 U2129 ( .A(n6210), .B(n6499), .C(n6828), .Y(n3369) );
  AOI22X1 U2130 ( .A(n8476), .B(n8767), .C(n8466), .D(n8603), .Y(n3375) );
  AOI22X1 U2132 ( .A(n8447), .B(n8808), .C(n8437), .D(n8726), .Y(n3373) );
  NAND3X1 U2134 ( .A(n1374), .B(n6498), .C(n6827), .Y(n3377) );
  AOI22X1 U2135 ( .A(n8494), .B(n9669), .C(n8488), .D(n9546), .Y(n3379) );
  NAND3X1 U2137 ( .A(n6209), .B(n6497), .C(n6826), .Y(n3376) );
  AOI22X1 U2138 ( .A(n8476), .B(n9751), .C(n8466), .D(n9587), .Y(n3382) );
  AOI22X1 U2140 ( .A(n8447), .B(n9792), .C(n8437), .D(n9710), .Y(n3380) );
  NAND3X1 U2141 ( .A(n1382), .B(n6496), .C(n6825), .Y(n3384) );
  AOI22X1 U2142 ( .A(n8497), .B(n9341), .C(n8488), .D(n9218), .Y(n3386) );
  NAND3X1 U2144 ( .A(n6208), .B(n6495), .C(n6824), .Y(n3383) );
  AOI22X1 U2145 ( .A(n8476), .B(n9423), .C(n8466), .D(n9259), .Y(n3389) );
  AOI22X1 U2147 ( .A(n8447), .B(n9464), .C(n8437), .D(n9382), .Y(n3387) );
  NAND3X1 U2149 ( .A(n6312), .B(n3391), .C(n3392), .Y(n5528) );
  NOR3X1 U2150 ( .A(n7011), .B(n7052), .C(n7093), .Y(n3392) );
  NAND3X1 U2152 ( .A(n4046), .B(n6494), .C(n6823), .Y(n3397) );
  AOI22X1 U2153 ( .A(n8495), .B(n9041), .C(n8488), .D(n8918), .Y(n3399) );
  NAND3X1 U2155 ( .A(n6207), .B(n6493), .C(n6822), .Y(n3396) );
  AOI22X1 U2156 ( .A(n8476), .B(n9123), .C(n8467), .D(n8959), .Y(n3402) );
  AOI22X1 U2158 ( .A(n8447), .B(n9164), .C(n8438), .D(n9082), .Y(n3400) );
  NAND3X1 U2160 ( .A(n1366), .B(n6492), .C(n6821), .Y(n3404) );
  AOI22X1 U2161 ( .A(n8498), .B(n8713), .C(n8488), .D(n8590), .Y(n3406) );
  NAND3X1 U2163 ( .A(n6206), .B(n6491), .C(n6820), .Y(n3403) );
  AOI22X1 U2164 ( .A(n8476), .B(n8795), .C(n8467), .D(n8631), .Y(n3409) );
  AOI22X1 U2166 ( .A(n8447), .B(n8836), .C(n8438), .D(n8754), .Y(n3407) );
  NAND3X1 U2168 ( .A(n1374), .B(n6490), .C(n6819), .Y(n3411) );
  AOI22X1 U2169 ( .A(n8495), .B(n9697), .C(n8488), .D(n9574), .Y(n3413) );
  NAND3X1 U2171 ( .A(n6205), .B(n6489), .C(n6818), .Y(n3410) );
  AOI22X1 U2172 ( .A(n8476), .B(n9779), .C(n8467), .D(n9615), .Y(n3416) );
  AOI22X1 U2174 ( .A(n8447), .B(n9820), .C(n8438), .D(n9738), .Y(n3414) );
  NAND3X1 U2175 ( .A(n1382), .B(n6488), .C(n6817), .Y(n3418) );
  AOI22X1 U2176 ( .A(n8496), .B(n9369), .C(n8488), .D(n9246), .Y(n3420) );
  NAND3X1 U2178 ( .A(n6204), .B(n6487), .C(n6816), .Y(n3417) );
  AOI22X1 U2179 ( .A(n8476), .B(n9451), .C(n8467), .D(n9287), .Y(n3423) );
  AOI22X1 U2181 ( .A(n8447), .B(n9492), .C(n8438), .D(n9410), .Y(n3421) );
  NAND3X1 U2183 ( .A(n6311), .B(n3425), .C(n3426), .Y(n5529) );
  NOR3X1 U2184 ( .A(n7010), .B(n7051), .C(n7092), .Y(n3426) );
  NAND3X1 U2186 ( .A(n4046), .B(n6486), .C(n6815), .Y(n3431) );
  AOI22X1 U2187 ( .A(n8492), .B(n9043), .C(n8488), .D(n8920), .Y(n3433) );
  NAND3X1 U2189 ( .A(n6203), .B(n6485), .C(n6814), .Y(n3430) );
  AOI22X1 U2190 ( .A(n8476), .B(n9125), .C(n8467), .D(n8961), .Y(n3436) );
  AOI22X1 U2192 ( .A(n8447), .B(n9166), .C(n8438), .D(n9084), .Y(n3434) );
  NAND3X1 U2194 ( .A(n1366), .B(n6484), .C(n6813), .Y(n3438) );
  AOI22X1 U2195 ( .A(n8497), .B(n8715), .C(n8488), .D(n8592), .Y(n3440) );
  NAND3X1 U2197 ( .A(n6202), .B(n6483), .C(n6812), .Y(n3437) );
  AOI22X1 U2198 ( .A(n8476), .B(n8797), .C(n8467), .D(n8633), .Y(n3443) );
  AOI22X1 U2200 ( .A(n8447), .B(n8838), .C(n8438), .D(n8756), .Y(n3441) );
  NAND3X1 U2202 ( .A(n1374), .B(n6482), .C(n6811), .Y(n3445) );
  AOI22X1 U2203 ( .A(n8494), .B(n9699), .C(n8488), .D(n9576), .Y(n3447) );
  NAND3X1 U2205 ( .A(n6201), .B(n6481), .C(n6810), .Y(n3444) );
  AOI22X1 U2206 ( .A(n8476), .B(n9781), .C(n8467), .D(n9617), .Y(n3450) );
  AOI22X1 U2208 ( .A(n8447), .B(n9822), .C(n8438), .D(n9740), .Y(n3448) );
  NAND3X1 U2209 ( .A(n1382), .B(n6480), .C(n6809), .Y(n3452) );
  AOI22X1 U2210 ( .A(n8494), .B(n9371), .C(n8488), .D(n9248), .Y(n3454) );
  NAND3X1 U2212 ( .A(n6200), .B(n6479), .C(n6808), .Y(n3451) );
  AOI22X1 U2213 ( .A(n8477), .B(n9453), .C(n8467), .D(n9289), .Y(n3457) );
  AOI22X1 U2215 ( .A(n8448), .B(n9494), .C(n8438), .D(n9412), .Y(n3455) );
  NAND3X1 U2217 ( .A(n6310), .B(n3459), .C(n3460), .Y(n5530) );
  NOR3X1 U2218 ( .A(n7009), .B(n7050), .C(n7091), .Y(n3460) );
  NAND3X1 U2220 ( .A(n4046), .B(n6478), .C(n6807), .Y(n3465) );
  AOI22X1 U2221 ( .A(n8494), .B(n9045), .C(n8484), .D(n8922), .Y(n3467) );
  NAND3X1 U2223 ( .A(n6199), .B(n6477), .C(n6806), .Y(n3464) );
  AOI22X1 U2224 ( .A(n8477), .B(n9127), .C(n8467), .D(n8963), .Y(n3470) );
  AOI22X1 U2226 ( .A(n8448), .B(n9168), .C(n8438), .D(n9086), .Y(n3468) );
  NAND3X1 U2228 ( .A(n1366), .B(n6476), .C(n6805), .Y(n3472) );
  AOI22X1 U2229 ( .A(n8494), .B(n8717), .C(n8485), .D(n8594), .Y(n3474) );
  NAND3X1 U2231 ( .A(n6198), .B(n6475), .C(n6804), .Y(n3471) );
  AOI22X1 U2232 ( .A(n8477), .B(n8799), .C(n8467), .D(n8635), .Y(n3477) );
  AOI22X1 U2234 ( .A(n8448), .B(n8840), .C(n8438), .D(n8758), .Y(n3475) );
  NAND3X1 U2236 ( .A(n1374), .B(n6474), .C(n6803), .Y(n3479) );
  AOI22X1 U2237 ( .A(n8494), .B(n9701), .C(n8484), .D(n9578), .Y(n3481) );
  NAND3X1 U2239 ( .A(n6197), .B(n6473), .C(n6802), .Y(n3478) );
  AOI22X1 U2240 ( .A(n8477), .B(n9783), .C(n8467), .D(n9619), .Y(n3484) );
  AOI22X1 U2242 ( .A(n8448), .B(n9824), .C(n8438), .D(n9742), .Y(n3482) );
  NAND3X1 U2243 ( .A(n1382), .B(n6472), .C(n6801), .Y(n3486) );
  AOI22X1 U2244 ( .A(n8494), .B(n9373), .C(n8490), .D(n9250), .Y(n3488) );
  NAND3X1 U2246 ( .A(n6196), .B(n6471), .C(n6800), .Y(n3485) );
  AOI22X1 U2247 ( .A(n8477), .B(n9455), .C(n8467), .D(n9291), .Y(n3491) );
  AOI22X1 U2249 ( .A(n8448), .B(n9496), .C(n8438), .D(n9414), .Y(n3489) );
  NAND3X1 U2251 ( .A(n6309), .B(n3493), .C(n3494), .Y(n5531) );
  NOR3X1 U2252 ( .A(n7008), .B(n7049), .C(n7090), .Y(n3494) );
  NAND3X1 U2254 ( .A(n4046), .B(n6470), .C(n6799), .Y(n3499) );
  AOI22X1 U2255 ( .A(n8494), .B(n9047), .C(n1355), .D(n8924), .Y(n3501) );
  NAND3X1 U2257 ( .A(n6195), .B(n6469), .C(n6798), .Y(n3498) );
  AOI22X1 U2258 ( .A(n8477), .B(n9129), .C(n8468), .D(n8965), .Y(n3504) );
  AOI22X1 U2260 ( .A(n8448), .B(n9170), .C(n8439), .D(n9088), .Y(n3502) );
  NAND3X1 U2262 ( .A(n1366), .B(n6468), .C(n6797), .Y(n3506) );
  AOI22X1 U2263 ( .A(n8494), .B(n8719), .C(n8486), .D(n8596), .Y(n3508) );
  NAND3X1 U2265 ( .A(n6194), .B(n6467), .C(n6796), .Y(n3505) );
  AOI22X1 U2266 ( .A(n8477), .B(n8801), .C(n8468), .D(n8637), .Y(n3511) );
  AOI22X1 U2268 ( .A(n8448), .B(n8842), .C(n8439), .D(n8760), .Y(n3509) );
  NAND3X1 U2270 ( .A(n1374), .B(n6466), .C(n6795), .Y(n3513) );
  AOI22X1 U2271 ( .A(n8494), .B(n9703), .C(n8490), .D(n9580), .Y(n3515) );
  NAND3X1 U2273 ( .A(n6193), .B(n6465), .C(n6794), .Y(n3512) );
  AOI22X1 U2274 ( .A(n8477), .B(n9785), .C(n8468), .D(n9621), .Y(n3518) );
  AOI22X1 U2276 ( .A(n8448), .B(n9826), .C(n8439), .D(n9744), .Y(n3516) );
  NAND3X1 U2277 ( .A(n8431), .B(n6464), .C(n6793), .Y(n3520) );
  AOI22X1 U2278 ( .A(n8494), .B(n9375), .C(n8487), .D(n9252), .Y(n3522) );
  NAND3X1 U2280 ( .A(n6192), .B(n6463), .C(n6792), .Y(n3519) );
  AOI22X1 U2281 ( .A(n8477), .B(n9457), .C(n8468), .D(n9293), .Y(n3525) );
  AOI22X1 U2283 ( .A(n8448), .B(n9498), .C(n8439), .D(n9416), .Y(n3523) );
  NAND3X1 U2285 ( .A(n6308), .B(n3527), .C(n3528), .Y(n5532) );
  NOR3X1 U2286 ( .A(n7007), .B(n7048), .C(n7089), .Y(n3528) );
  NAND3X1 U2288 ( .A(n4046), .B(n6462), .C(n6791), .Y(n3533) );
  AOI22X1 U2289 ( .A(n8494), .B(n9049), .C(n8489), .D(n8926), .Y(n3535) );
  NAND3X1 U2291 ( .A(n6191), .B(n6461), .C(n6790), .Y(n3532) );
  AOI22X1 U2292 ( .A(n8477), .B(n9131), .C(n8468), .D(n8967), .Y(n3538) );
  AOI22X1 U2294 ( .A(n8448), .B(n9172), .C(n8439), .D(n9090), .Y(n3536) );
  NAND3X1 U2296 ( .A(n1366), .B(n6460), .C(n6789), .Y(n3540) );
  AOI22X1 U2297 ( .A(n8494), .B(n8721), .C(n8483), .D(n8598), .Y(n3542) );
  NAND3X1 U2299 ( .A(n6190), .B(n6459), .C(n6788), .Y(n3539) );
  AOI22X1 U2300 ( .A(n8477), .B(n8803), .C(n8468), .D(n8639), .Y(n3545) );
  AOI22X1 U2302 ( .A(n8448), .B(n8844), .C(n8439), .D(n8762), .Y(n3543) );
  NAND3X1 U2304 ( .A(n1374), .B(n6458), .C(n6787), .Y(n3547) );
  AOI22X1 U2305 ( .A(n8494), .B(n9705), .C(n8487), .D(n9582), .Y(n3549) );
  NAND3X1 U2307 ( .A(n6189), .B(n6457), .C(n6786), .Y(n3546) );
  AOI22X1 U2308 ( .A(n8477), .B(n9787), .C(n8468), .D(n9623), .Y(n3552) );
  AOI22X1 U2310 ( .A(n8448), .B(n9828), .C(n8439), .D(n9746), .Y(n3550) );
  NAND3X1 U2311 ( .A(n8431), .B(n6456), .C(n6785), .Y(n3554) );
  AOI22X1 U2312 ( .A(n8494), .B(n9377), .C(n8485), .D(n9254), .Y(n3556) );
  NAND3X1 U2314 ( .A(n6188), .B(n6455), .C(n6784), .Y(n3553) );
  AOI22X1 U2315 ( .A(n8477), .B(n9459), .C(n8468), .D(n9295), .Y(n3559) );
  AOI22X1 U2317 ( .A(n8448), .B(n9500), .C(n8439), .D(n9418), .Y(n3557) );
  NAND3X1 U2319 ( .A(n6307), .B(n3561), .C(n3562), .Y(n5533) );
  NOR3X1 U2320 ( .A(n7006), .B(n7047), .C(n7088), .Y(n3562) );
  NAND3X1 U2322 ( .A(n4046), .B(n6454), .C(n6783), .Y(n3567) );
  AOI22X1 U2323 ( .A(n8495), .B(n9051), .C(n8487), .D(n8928), .Y(n3569) );
  NAND3X1 U2325 ( .A(n6187), .B(n6453), .C(n6782), .Y(n3566) );
  AOI22X1 U2326 ( .A(n8478), .B(n9133), .C(n8468), .D(n8969), .Y(n3572) );
  AOI22X1 U2328 ( .A(n8449), .B(n9174), .C(n8439), .D(n9092), .Y(n3570) );
  NAND3X1 U2330 ( .A(n1366), .B(n6452), .C(n6781), .Y(n3574) );
  AOI22X1 U2331 ( .A(n8495), .B(n8723), .C(n8487), .D(n8600), .Y(n3576) );
  NAND3X1 U2333 ( .A(n6186), .B(n6451), .C(n6780), .Y(n3573) );
  AOI22X1 U2334 ( .A(n8478), .B(n8805), .C(n8468), .D(n8641), .Y(n3579) );
  AOI22X1 U2336 ( .A(n8449), .B(n8846), .C(n8439), .D(n8764), .Y(n3577) );
  NAND3X1 U2338 ( .A(n1374), .B(n6450), .C(n6779), .Y(n3581) );
  AOI22X1 U2339 ( .A(n8495), .B(n9707), .C(n8487), .D(n9584), .Y(n3583) );
  NAND3X1 U2341 ( .A(n6185), .B(n6449), .C(n6778), .Y(n3580) );
  AOI22X1 U2342 ( .A(n8478), .B(n9789), .C(n8468), .D(n9625), .Y(n3586) );
  AOI22X1 U2344 ( .A(n8449), .B(n9830), .C(n8439), .D(n9748), .Y(n3584) );
  NAND3X1 U2345 ( .A(n8431), .B(n6448), .C(n6777), .Y(n3588) );
  AOI22X1 U2346 ( .A(n8495), .B(n9379), .C(n8487), .D(n9256), .Y(n3590) );
  NAND3X1 U2348 ( .A(n6184), .B(n6447), .C(n6776), .Y(n3587) );
  AOI22X1 U2349 ( .A(n8478), .B(n9461), .C(n8468), .D(n9297), .Y(n3593) );
  AOI22X1 U2351 ( .A(n8449), .B(n9502), .C(n8439), .D(n9420), .Y(n3591) );
  NAND3X1 U2353 ( .A(n6306), .B(n3595), .C(n3596), .Y(n5534) );
  NOR3X1 U2354 ( .A(n7005), .B(n7046), .C(n7087), .Y(n3596) );
  NAND3X1 U2356 ( .A(n4046), .B(n6446), .C(n6775), .Y(n3601) );
  AOI22X1 U2357 ( .A(n8495), .B(n9011), .C(n8487), .D(n8888), .Y(n3603) );
  NAND3X1 U2359 ( .A(n6183), .B(n6445), .C(n6774), .Y(n3600) );
  AOI22X1 U2360 ( .A(n8478), .B(n9093), .C(n8469), .D(n8929), .Y(n3606) );
  AOI22X1 U2362 ( .A(n8449), .B(n9134), .C(n8440), .D(n9052), .Y(n3604) );
  NAND3X1 U2364 ( .A(n1366), .B(n6444), .C(n6773), .Y(n3608) );
  AOI22X1 U2365 ( .A(n8495), .B(n8683), .C(n8487), .D(n8560), .Y(n3610) );
  NAND3X1 U2367 ( .A(n6182), .B(n6443), .C(n6772), .Y(n3607) );
  AOI22X1 U2368 ( .A(n8478), .B(n8765), .C(n8469), .D(n8601), .Y(n3613) );
  AOI22X1 U2370 ( .A(n8449), .B(n8806), .C(n8440), .D(n8724), .Y(n3611) );
  NAND3X1 U2372 ( .A(n1374), .B(n6442), .C(n6771), .Y(n3615) );
  AOI22X1 U2373 ( .A(n8495), .B(n9667), .C(n8487), .D(n9544), .Y(n3617) );
  NAND3X1 U2375 ( .A(n6181), .B(n6441), .C(n6770), .Y(n3614) );
  AOI22X1 U2376 ( .A(n8478), .B(n9749), .C(n8469), .D(n9585), .Y(n3620) );
  AOI22X1 U2378 ( .A(n8449), .B(n9790), .C(n8440), .D(n9708), .Y(n3618) );
  NAND3X1 U2379 ( .A(n8431), .B(n6440), .C(n6769), .Y(n3622) );
  AOI22X1 U2380 ( .A(n8495), .B(n9339), .C(n8487), .D(n9216), .Y(n3624) );
  NAND3X1 U2382 ( .A(n6180), .B(n6439), .C(n6768), .Y(n3621) );
  AOI22X1 U2383 ( .A(n8478), .B(n9421), .C(n8469), .D(n9257), .Y(n3627) );
  AOI22X1 U2385 ( .A(n8449), .B(n9462), .C(n8440), .D(n9380), .Y(n3625) );
  NAND3X1 U2387 ( .A(n6305), .B(n3629), .C(n3630), .Y(n5535) );
  NOR3X1 U2388 ( .A(n7004), .B(n7045), .C(n7086), .Y(n3630) );
  NAND3X1 U2390 ( .A(n4046), .B(n6438), .C(n6767), .Y(n3635) );
  AOI22X1 U2391 ( .A(n8495), .B(n9014), .C(n8487), .D(n8891), .Y(n3637) );
  NAND3X1 U2393 ( .A(n6179), .B(n6437), .C(n6766), .Y(n3634) );
  AOI22X1 U2394 ( .A(n8478), .B(n9096), .C(n8469), .D(n8932), .Y(n3640) );
  AOI22X1 U2396 ( .A(n8449), .B(n9137), .C(n8440), .D(n9055), .Y(n3638) );
  NAND3X1 U2398 ( .A(n1366), .B(n6436), .C(n6765), .Y(n3642) );
  AOI22X1 U2399 ( .A(n8495), .B(n8686), .C(n8487), .D(n8563), .Y(n3644) );
  NAND3X1 U2401 ( .A(n6178), .B(n6435), .C(n6764), .Y(n3641) );
  AOI22X1 U2402 ( .A(n8478), .B(n8768), .C(n8469), .D(n8604), .Y(n3647) );
  AOI22X1 U2404 ( .A(n8449), .B(n8809), .C(n8440), .D(n8727), .Y(n3645) );
  NAND3X1 U2406 ( .A(n1374), .B(n6434), .C(n6763), .Y(n3649) );
  AOI22X1 U2407 ( .A(n8495), .B(n9670), .C(n8487), .D(n9547), .Y(n3651) );
  NAND3X1 U2409 ( .A(n6177), .B(n6433), .C(n6762), .Y(n3648) );
  AOI22X1 U2410 ( .A(n8478), .B(n9752), .C(n8469), .D(n9588), .Y(n3654) );
  AOI22X1 U2412 ( .A(n8449), .B(n9793), .C(n8440), .D(n9711), .Y(n3652) );
  NAND3X1 U2413 ( .A(n8431), .B(n6432), .C(n6761), .Y(n3656) );
  AOI22X1 U2414 ( .A(n8495), .B(n9342), .C(n8487), .D(n9219), .Y(n3658) );
  NAND3X1 U2416 ( .A(n6176), .B(n6431), .C(n6760), .Y(n3655) );
  AOI22X1 U2417 ( .A(n8478), .B(n9424), .C(n8469), .D(n9260), .Y(n3661) );
  AOI22X1 U2419 ( .A(n8449), .B(n9465), .C(n8440), .D(n9383), .Y(n3659) );
  NAND3X1 U2421 ( .A(n6304), .B(n3663), .C(n3664), .Y(n5536) );
  NOR3X1 U2422 ( .A(n7003), .B(n7044), .C(n7085), .Y(n3664) );
  NAND3X1 U2424 ( .A(n4046), .B(n6430), .C(n6759), .Y(n3669) );
  AOI22X1 U2425 ( .A(n8495), .B(n9028), .C(n8486), .D(n8905), .Y(n3671) );
  NAND3X1 U2427 ( .A(n6175), .B(n6429), .C(n6758), .Y(n3668) );
  AOI22X1 U2428 ( .A(n8478), .B(n9110), .C(n8469), .D(n8946), .Y(n3674) );
  AOI22X1 U2430 ( .A(n8449), .B(n9151), .C(n8440), .D(n9069), .Y(n3672) );
  NAND3X1 U2432 ( .A(n1366), .B(n6428), .C(n6757), .Y(n3676) );
  AOI22X1 U2433 ( .A(n8496), .B(n8700), .C(n8486), .D(n8577), .Y(n3678) );
  NAND3X1 U2435 ( .A(n6174), .B(n6427), .C(n6756), .Y(n3675) );
  AOI22X1 U2436 ( .A(n8475), .B(n8782), .C(n8469), .D(n8618), .Y(n3681) );
  AOI22X1 U2438 ( .A(n8450), .B(n8823), .C(n8440), .D(n8741), .Y(n3679) );
  NAND3X1 U2440 ( .A(n8433), .B(n6426), .C(n6755), .Y(n3683) );
  AOI22X1 U2441 ( .A(n8496), .B(n9684), .C(n8486), .D(n9561), .Y(n3685) );
  NAND3X1 U2443 ( .A(n6173), .B(n6425), .C(n6754), .Y(n3682) );
  AOI22X1 U2444 ( .A(n8479), .B(n9766), .C(n8469), .D(n9602), .Y(n3688) );
  AOI22X1 U2446 ( .A(n8450), .B(n9807), .C(n8440), .D(n9725), .Y(n3686) );
  NAND3X1 U2447 ( .A(n8431), .B(n6424), .C(n6753), .Y(n3690) );
  AOI22X1 U2448 ( .A(n8496), .B(n9356), .C(n8486), .D(n9233), .Y(n3692) );
  NAND3X1 U2450 ( .A(n6172), .B(n6423), .C(n6752), .Y(n3689) );
  AOI22X1 U2451 ( .A(n8475), .B(n9438), .C(n8469), .D(n9274), .Y(n3695) );
  AOI22X1 U2453 ( .A(n8450), .B(n9479), .C(n8440), .D(n9397), .Y(n3693) );
  NAND3X1 U2455 ( .A(n6303), .B(n3697), .C(n3698), .Y(n5537) );
  NOR3X1 U2456 ( .A(n7002), .B(n7043), .C(n7084), .Y(n3698) );
  NAND3X1 U2458 ( .A(n4046), .B(n6422), .C(n6751), .Y(n3703) );
  AOI22X1 U2459 ( .A(n8496), .B(n9029), .C(n8486), .D(n8906), .Y(n3705) );
  NAND3X1 U2461 ( .A(n6171), .B(n6421), .C(n6750), .Y(n3702) );
  AOI22X1 U2462 ( .A(n8478), .B(n9111), .C(n8470), .D(n8947), .Y(n3708) );
  AOI22X1 U2464 ( .A(n8450), .B(n9152), .C(n8441), .D(n9070), .Y(n3706) );
  NAND3X1 U2466 ( .A(n1366), .B(n6420), .C(n6749), .Y(n3710) );
  AOI22X1 U2467 ( .A(n8496), .B(n8701), .C(n8486), .D(n8578), .Y(n3712) );
  NAND3X1 U2469 ( .A(n6170), .B(n6419), .C(n6748), .Y(n3709) );
  AOI22X1 U2470 ( .A(n8479), .B(n8783), .C(n8470), .D(n8619), .Y(n3715) );
  AOI22X1 U2472 ( .A(n8450), .B(n8824), .C(n8441), .D(n8742), .Y(n3713) );
  NAND3X1 U2474 ( .A(n8433), .B(n6418), .C(n6747), .Y(n3717) );
  AOI22X1 U2475 ( .A(n8496), .B(n9685), .C(n8486), .D(n9562), .Y(n3719) );
  NAND3X1 U2477 ( .A(n6169), .B(n6417), .C(n6746), .Y(n3716) );
  AOI22X1 U2478 ( .A(n8480), .B(n9767), .C(n8470), .D(n9603), .Y(n3722) );
  AOI22X1 U2480 ( .A(n8450), .B(n9808), .C(n8441), .D(n9726), .Y(n3720) );
  NAND3X1 U2481 ( .A(n8431), .B(n6416), .C(n6745), .Y(n3724) );
  AOI22X1 U2482 ( .A(n8496), .B(n9357), .C(n8486), .D(n9234), .Y(n3726) );
  NAND3X1 U2484 ( .A(n6168), .B(n6415), .C(n6744), .Y(n3723) );
  AOI22X1 U2485 ( .A(n8479), .B(n9439), .C(n8470), .D(n9275), .Y(n3729) );
  AOI22X1 U2487 ( .A(n8450), .B(n9480), .C(n8441), .D(n9398), .Y(n3727) );
  NAND3X1 U2489 ( .A(n6302), .B(n3731), .C(n3732), .Y(n5538) );
  NOR3X1 U2490 ( .A(n7001), .B(n7042), .C(n7083), .Y(n3732) );
  NAND3X1 U2492 ( .A(n4046), .B(n6414), .C(n6743), .Y(n3737) );
  AOI22X1 U2493 ( .A(n8496), .B(n9030), .C(n8486), .D(n8907), .Y(n3739) );
  NAND3X1 U2495 ( .A(n6167), .B(n6413), .C(n6742), .Y(n3736) );
  AOI22X1 U2496 ( .A(n8477), .B(n9112), .C(n8470), .D(n8948), .Y(n3742) );
  AOI22X1 U2498 ( .A(n8450), .B(n9153), .C(n8441), .D(n9071), .Y(n3740) );
  NAND3X1 U2500 ( .A(n1366), .B(n6412), .C(n6741), .Y(n3744) );
  AOI22X1 U2501 ( .A(n8496), .B(n8702), .C(n8486), .D(n8579), .Y(n3746) );
  NAND3X1 U2503 ( .A(n6166), .B(n6411), .C(n6740), .Y(n3743) );
  AOI22X1 U2504 ( .A(n8480), .B(n8784), .C(n8470), .D(n8620), .Y(n3749) );
  AOI22X1 U2506 ( .A(n8450), .B(n8825), .C(n8441), .D(n8743), .Y(n3747) );
  NAND3X1 U2508 ( .A(n8433), .B(n6410), .C(n6739), .Y(n3751) );
  AOI22X1 U2509 ( .A(n8496), .B(n9686), .C(n8486), .D(n9563), .Y(n3753) );
  NAND3X1 U2511 ( .A(n6165), .B(n6409), .C(n6738), .Y(n3750) );
  AOI22X1 U2512 ( .A(n8478), .B(n9768), .C(n8470), .D(n9604), .Y(n3756) );
  AOI22X1 U2514 ( .A(n8450), .B(n9809), .C(n8441), .D(n9727), .Y(n3754) );
  NAND3X1 U2515 ( .A(n8431), .B(n6408), .C(n6737), .Y(n3758) );
  AOI22X1 U2516 ( .A(n8496), .B(n9358), .C(n8486), .D(n9235), .Y(n3760) );
  NAND3X1 U2518 ( .A(n6164), .B(n6407), .C(n6736), .Y(n3757) );
  AOI22X1 U2519 ( .A(n8480), .B(n9440), .C(n8470), .D(n9276), .Y(n3763) );
  AOI22X1 U2521 ( .A(n8450), .B(n9481), .C(n8441), .D(n9399), .Y(n3761) );
  NAND3X1 U2523 ( .A(n6301), .B(n3765), .C(n3766), .Y(n5539) );
  NOR3X1 U2524 ( .A(n7000), .B(n7041), .C(n7082), .Y(n3766) );
  NAND3X1 U2526 ( .A(n4046), .B(n6406), .C(n6735), .Y(n3771) );
  AOI22X1 U2527 ( .A(n8496), .B(n9031), .C(n8485), .D(n8908), .Y(n3773) );
  NAND3X1 U2529 ( .A(n6163), .B(n6405), .C(n6734), .Y(n3770) );
  AOI22X1 U2530 ( .A(n8476), .B(n9113), .C(n8470), .D(n8949), .Y(n3776) );
  AOI22X1 U2532 ( .A(n8450), .B(n9154), .C(n8441), .D(n9072), .Y(n3774) );
  NAND3X1 U2534 ( .A(n1366), .B(n6404), .C(n6733), .Y(n3778) );
  AOI22X1 U2535 ( .A(n8496), .B(n8703), .C(n8485), .D(n8580), .Y(n3780) );
  NAND3X1 U2537 ( .A(n6162), .B(n6403), .C(n6732), .Y(n3777) );
  AOI22X1 U2538 ( .A(n8478), .B(n8785), .C(n8470), .D(n8621), .Y(n3783) );
  AOI22X1 U2540 ( .A(n8450), .B(n8826), .C(n8441), .D(n8744), .Y(n3781) );
  NAND3X1 U2542 ( .A(n8433), .B(n6402), .C(n6731), .Y(n3785) );
  AOI22X1 U2543 ( .A(n8497), .B(n9687), .C(n8485), .D(n9564), .Y(n3787) );
  NAND3X1 U2545 ( .A(n6161), .B(n6401), .C(n6730), .Y(n3784) );
  AOI22X1 U2546 ( .A(n8479), .B(n9769), .C(n8470), .D(n9605), .Y(n3790) );
  AOI22X1 U2548 ( .A(n8451), .B(n9810), .C(n8441), .D(n9728), .Y(n3788) );
  NAND3X1 U2549 ( .A(n8431), .B(n6400), .C(n6729), .Y(n3792) );
  AOI22X1 U2550 ( .A(n8497), .B(n9359), .C(n8485), .D(n9236), .Y(n3794) );
  NAND3X1 U2552 ( .A(n6160), .B(n6399), .C(n6728), .Y(n3791) );
  AOI22X1 U2553 ( .A(n8479), .B(n9441), .C(n8470), .D(n9277), .Y(n3797) );
  AOI22X1 U2555 ( .A(n8451), .B(n9482), .C(n8441), .D(n9400), .Y(n3795) );
  NAND3X1 U2557 ( .A(n6300), .B(n3799), .C(n3800), .Y(n5540) );
  NOR3X1 U2558 ( .A(n6999), .B(n7040), .C(n7081), .Y(n3800) );
  NAND3X1 U2560 ( .A(n4046), .B(n6398), .C(n6727), .Y(n3805) );
  AOI22X1 U2561 ( .A(n8497), .B(n9032), .C(n8485), .D(n8909), .Y(n3807) );
  NAND3X1 U2563 ( .A(n6159), .B(n6397), .C(n6726), .Y(n3804) );
  AOI22X1 U2564 ( .A(n8479), .B(n9114), .C(n8471), .D(n8950), .Y(n3810) );
  AOI22X1 U2566 ( .A(n8451), .B(n9155), .C(n8442), .D(n9073), .Y(n3808) );
  NAND3X1 U2568 ( .A(n1366), .B(n6396), .C(n6725), .Y(n3812) );
  AOI22X1 U2569 ( .A(n8497), .B(n8704), .C(n8485), .D(n8581), .Y(n3814) );
  NAND3X1 U2571 ( .A(n6158), .B(n6395), .C(n6724), .Y(n3811) );
  AOI22X1 U2572 ( .A(n8479), .B(n8786), .C(n8471), .D(n8622), .Y(n3817) );
  AOI22X1 U2574 ( .A(n8451), .B(n8827), .C(n8442), .D(n8745), .Y(n3815) );
  NAND3X1 U2576 ( .A(n8433), .B(n6394), .C(n6723), .Y(n3819) );
  AOI22X1 U2577 ( .A(n8497), .B(n9688), .C(n8485), .D(n9565), .Y(n3821) );
  NAND3X1 U2579 ( .A(n6157), .B(n6393), .C(n6722), .Y(n3818) );
  AOI22X1 U2580 ( .A(n8479), .B(n9770), .C(n8471), .D(n9606), .Y(n3824) );
  AOI22X1 U2582 ( .A(n8451), .B(n9811), .C(n8442), .D(n9729), .Y(n3822) );
  NAND3X1 U2583 ( .A(n8431), .B(n6392), .C(n6721), .Y(n3826) );
  AOI22X1 U2584 ( .A(n8497), .B(n9360), .C(n8485), .D(n9237), .Y(n3828) );
  NAND3X1 U2586 ( .A(n6156), .B(n6391), .C(n6720), .Y(n3825) );
  AOI22X1 U2587 ( .A(n8479), .B(n9442), .C(n8471), .D(n9278), .Y(n3831) );
  AOI22X1 U2589 ( .A(n8451), .B(n9483), .C(n8442), .D(n9401), .Y(n3829) );
  NAND3X1 U2591 ( .A(n6299), .B(n3833), .C(n3834), .Y(n5541) );
  NOR3X1 U2592 ( .A(n6998), .B(n7039), .C(n7080), .Y(n3834) );
  NAND3X1 U2594 ( .A(n4046), .B(n6390), .C(n6719), .Y(n3839) );
  AOI22X1 U2595 ( .A(n8497), .B(n9033), .C(n8485), .D(n8910), .Y(n3841) );
  NAND3X1 U2597 ( .A(n6155), .B(n6389), .C(n6718), .Y(n3838) );
  AOI22X1 U2598 ( .A(n8479), .B(n9115), .C(n8471), .D(n8951), .Y(n3844) );
  AOI22X1 U2600 ( .A(n8451), .B(n9156), .C(n8442), .D(n9074), .Y(n3842) );
  NAND3X1 U2602 ( .A(n1366), .B(n6388), .C(n6717), .Y(n3846) );
  AOI22X1 U2603 ( .A(n8497), .B(n8705), .C(n8485), .D(n8582), .Y(n3848) );
  NAND3X1 U2605 ( .A(n6154), .B(n6387), .C(n6716), .Y(n3845) );
  AOI22X1 U2606 ( .A(n8479), .B(n8787), .C(n8471), .D(n8623), .Y(n3851) );
  AOI22X1 U2608 ( .A(n8451), .B(n8828), .C(n8442), .D(n8746), .Y(n3849) );
  NAND3X1 U2610 ( .A(n8433), .B(n6386), .C(n6715), .Y(n3853) );
  AOI22X1 U2611 ( .A(n8497), .B(n9689), .C(n8485), .D(n9566), .Y(n3855) );
  NAND3X1 U2613 ( .A(n6153), .B(n6385), .C(n6714), .Y(n3852) );
  AOI22X1 U2614 ( .A(n8479), .B(n9771), .C(n8471), .D(n9607), .Y(n3858) );
  AOI22X1 U2616 ( .A(n8451), .B(n9812), .C(n8442), .D(n9730), .Y(n3856) );
  NAND3X1 U2617 ( .A(n8431), .B(n6384), .C(n6713), .Y(n3860) );
  AOI22X1 U2618 ( .A(n8497), .B(n9361), .C(n8485), .D(n9238), .Y(n3862) );
  NAND3X1 U2620 ( .A(n6152), .B(n6383), .C(n6712), .Y(n3859) );
  AOI22X1 U2621 ( .A(n8479), .B(n9443), .C(n8471), .D(n9279), .Y(n3865) );
  AOI22X1 U2623 ( .A(n8451), .B(n9484), .C(n8442), .D(n9402), .Y(n3863) );
  NAND3X1 U2625 ( .A(n6298), .B(n3867), .C(n3868), .Y(n5542) );
  NOR3X1 U2626 ( .A(n6997), .B(n7038), .C(n7079), .Y(n3868) );
  NAND3X1 U2628 ( .A(n4046), .B(n6382), .C(n6711), .Y(n3873) );
  AOI22X1 U2629 ( .A(n8497), .B(n9034), .C(n8484), .D(n8911), .Y(n3875) );
  NAND3X1 U2631 ( .A(n6151), .B(n6381), .C(n6710), .Y(n3872) );
  AOI22X1 U2632 ( .A(n8479), .B(n9116), .C(n8471), .D(n8952), .Y(n3878) );
  AOI22X1 U2634 ( .A(n8451), .B(n9157), .C(n8442), .D(n9075), .Y(n3876) );
  NAND3X1 U2636 ( .A(n1366), .B(n6380), .C(n6709), .Y(n3880) );
  AOI22X1 U2637 ( .A(n8497), .B(n8706), .C(n8484), .D(n8583), .Y(n3882) );
  NAND3X1 U2639 ( .A(n6150), .B(n6379), .C(n6708), .Y(n3879) );
  AOI22X1 U2640 ( .A(n8479), .B(n8788), .C(n8471), .D(n8624), .Y(n3885) );
  AOI22X1 U2642 ( .A(n8451), .B(n8829), .C(n8442), .D(n8747), .Y(n3883) );
  NAND3X1 U2644 ( .A(n8433), .B(n6378), .C(n6707), .Y(n3887) );
  AOI22X1 U2645 ( .A(n8497), .B(n9690), .C(n8484), .D(n9567), .Y(n3889) );
  NAND3X1 U2647 ( .A(n6149), .B(n6377), .C(n6706), .Y(n3886) );
  AOI22X1 U2648 ( .A(n8479), .B(n9772), .C(n8471), .D(n9608), .Y(n3892) );
  AOI22X1 U2650 ( .A(n8451), .B(n9813), .C(n8442), .D(n9731), .Y(n3890) );
  NAND3X1 U2651 ( .A(n8431), .B(n6376), .C(n6705), .Y(n3894) );
  AOI22X1 U2652 ( .A(n8498), .B(n9362), .C(n8484), .D(n9239), .Y(n3896) );
  NAND3X1 U2654 ( .A(n6148), .B(n6375), .C(n6704), .Y(n3893) );
  AOI22X1 U2655 ( .A(n8480), .B(n9444), .C(n8471), .D(n9280), .Y(n3899) );
  AOI22X1 U2657 ( .A(n8452), .B(n9485), .C(n8442), .D(n9403), .Y(n3897) );
  NAND3X1 U2659 ( .A(n6297), .B(n3901), .C(n3902), .Y(n5543) );
  NOR3X1 U2660 ( .A(n6996), .B(n7037), .C(n7078), .Y(n3902) );
  NAND3X1 U2662 ( .A(n4046), .B(n6374), .C(n6703), .Y(n3907) );
  AOI22X1 U2663 ( .A(n8498), .B(n9035), .C(n8484), .D(n8912), .Y(n3909) );
  NAND3X1 U2665 ( .A(n6147), .B(n6373), .C(n6702), .Y(n3906) );
  AOI22X1 U2666 ( .A(n8480), .B(n9117), .C(n8472), .D(n8953), .Y(n3912) );
  AOI22X1 U2668 ( .A(n8452), .B(n9158), .C(n8443), .D(n9076), .Y(n3910) );
  NAND3X1 U2670 ( .A(n1366), .B(n6372), .C(n6701), .Y(n3914) );
  AOI22X1 U2671 ( .A(n8498), .B(n8707), .C(n8484), .D(n8584), .Y(n3916) );
  NAND3X1 U2673 ( .A(n6146), .B(n6371), .C(n6700), .Y(n3913) );
  AOI22X1 U2674 ( .A(n8480), .B(n8789), .C(n8472), .D(n8625), .Y(n3919) );
  AOI22X1 U2676 ( .A(n8452), .B(n8830), .C(n8443), .D(n8748), .Y(n3917) );
  NAND3X1 U2678 ( .A(n8433), .B(n6370), .C(n6699), .Y(n3921) );
  AOI22X1 U2679 ( .A(n8498), .B(n9691), .C(n8484), .D(n9568), .Y(n3923) );
  NAND3X1 U2681 ( .A(n6145), .B(n6369), .C(n6698), .Y(n3920) );
  AOI22X1 U2682 ( .A(n8480), .B(n9773), .C(n8472), .D(n9609), .Y(n3926) );
  AOI22X1 U2684 ( .A(n8452), .B(n9814), .C(n8443), .D(n9732), .Y(n3924) );
  NAND3X1 U2685 ( .A(n1382), .B(n6368), .C(n6697), .Y(n3928) );
  AOI22X1 U2686 ( .A(n8498), .B(n9363), .C(n8484), .D(n9240), .Y(n3930) );
  NAND3X1 U2688 ( .A(n6144), .B(n6367), .C(n6696), .Y(n3927) );
  AOI22X1 U2689 ( .A(n8480), .B(n9445), .C(n8472), .D(n9281), .Y(n3933) );
  AOI22X1 U2691 ( .A(n8452), .B(n9486), .C(n8443), .D(n9404), .Y(n3931) );
  NAND3X1 U2693 ( .A(n6296), .B(n3935), .C(n3936), .Y(n5544) );
  NOR3X1 U2694 ( .A(n6995), .B(n7036), .C(n7077), .Y(n3936) );
  NAND3X1 U2696 ( .A(n4046), .B(n6366), .C(n6695), .Y(n3941) );
  AOI22X1 U2697 ( .A(n8498), .B(n9036), .C(n8484), .D(n8913), .Y(n3943) );
  NAND3X1 U2699 ( .A(n6143), .B(n6365), .C(n6694), .Y(n3940) );
  AOI22X1 U2700 ( .A(n8480), .B(n9118), .C(n8472), .D(n8954), .Y(n3946) );
  AOI22X1 U2702 ( .A(n8452), .B(n9159), .C(n8443), .D(n9077), .Y(n3944) );
  NAND3X1 U2704 ( .A(n1366), .B(n6364), .C(n6693), .Y(n3948) );
  AOI22X1 U2705 ( .A(n8498), .B(n8708), .C(n8484), .D(n8585), .Y(n3950) );
  NAND3X1 U2707 ( .A(n6142), .B(n6363), .C(n6692), .Y(n3947) );
  AOI22X1 U2708 ( .A(n8480), .B(n8790), .C(n8472), .D(n8626), .Y(n3953) );
  AOI22X1 U2710 ( .A(n8452), .B(n8831), .C(n8443), .D(n8749), .Y(n3951) );
  NAND3X1 U2712 ( .A(n8433), .B(n6362), .C(n6691), .Y(n3955) );
  AOI22X1 U2713 ( .A(n8498), .B(n9692), .C(n8484), .D(n9569), .Y(n3957) );
  NAND3X1 U2715 ( .A(n6141), .B(n6361), .C(n6690), .Y(n3954) );
  AOI22X1 U2716 ( .A(n8480), .B(n9774), .C(n8472), .D(n9610), .Y(n3960) );
  AOI22X1 U2718 ( .A(n8452), .B(n9815), .C(n8443), .D(n9733), .Y(n3958) );
  NAND3X1 U2719 ( .A(n1382), .B(n6360), .C(n6689), .Y(n3962) );
  AOI22X1 U2720 ( .A(n8498), .B(n9364), .C(n8484), .D(n9241), .Y(n3964) );
  NAND3X1 U2722 ( .A(n6140), .B(n6359), .C(n6688), .Y(n3961) );
  AOI22X1 U2723 ( .A(n8480), .B(n9446), .C(n8472), .D(n9282), .Y(n3967) );
  AOI22X1 U2725 ( .A(n8452), .B(n9487), .C(n8443), .D(n9405), .Y(n3965) );
  NAND3X1 U2727 ( .A(n6295), .B(n3969), .C(n3970), .Y(n5545) );
  NOR3X1 U2728 ( .A(n6994), .B(n7035), .C(n7076), .Y(n3970) );
  NAND3X1 U2730 ( .A(n4046), .B(n6358), .C(n6687), .Y(n3975) );
  AOI22X1 U2731 ( .A(n8498), .B(n9037), .C(n8483), .D(n8914), .Y(n3977) );
  NAND3X1 U2733 ( .A(n6139), .B(n6357), .C(n6686), .Y(n3974) );
  AOI22X1 U2734 ( .A(n8480), .B(n9119), .C(n8472), .D(n8955), .Y(n3980) );
  AOI22X1 U2736 ( .A(n8452), .B(n9160), .C(n8443), .D(n9078), .Y(n3978) );
  NAND3X1 U2738 ( .A(n1366), .B(n6356), .C(n6685), .Y(n3982) );
  AOI22X1 U2739 ( .A(n8498), .B(n8709), .C(n8483), .D(n8586), .Y(n3984) );
  NAND3X1 U2741 ( .A(n6138), .B(n6355), .C(n6684), .Y(n3981) );
  AOI22X1 U2742 ( .A(n8480), .B(n8791), .C(n8472), .D(n8627), .Y(n3987) );
  AOI22X1 U2744 ( .A(n8452), .B(n8832), .C(n8443), .D(n8750), .Y(n3985) );
  NAND3X1 U2746 ( .A(n8433), .B(n6354), .C(n6683), .Y(n3989) );
  AOI22X1 U2747 ( .A(n8498), .B(n9693), .C(n8483), .D(n9570), .Y(n3991) );
  NAND3X1 U2749 ( .A(n6137), .B(n6353), .C(n6682), .Y(n3988) );
  AOI22X1 U2750 ( .A(n8480), .B(n9775), .C(n8472), .D(n9611), .Y(n3994) );
  AOI22X1 U2752 ( .A(n8452), .B(n9816), .C(n8443), .D(n9734), .Y(n3992) );
  NAND3X1 U2753 ( .A(n1382), .B(n6352), .C(n6681), .Y(n3996) );
  AOI22X1 U2754 ( .A(n8498), .B(n9365), .C(n8483), .D(n9242), .Y(n3998) );
  NAND3X1 U2756 ( .A(n6136), .B(n6351), .C(n6680), .Y(n3995) );
  AOI22X1 U2757 ( .A(n8480), .B(n9447), .C(n8472), .D(n9283), .Y(n4001) );
  AOI22X1 U2759 ( .A(n8452), .B(n9488), .C(n8443), .D(n9406), .Y(n3999) );
  NAND3X1 U2761 ( .A(n6294), .B(n4003), .C(n4004), .Y(n5546) );
  NOR3X1 U2762 ( .A(n6993), .B(n7034), .C(n7075), .Y(n4004) );
  NAND3X1 U2764 ( .A(n4046), .B(n6350), .C(n6679), .Y(n4009) );
  AOI22X1 U2765 ( .A(n1354), .B(n9038), .C(n8483), .D(n8915), .Y(n4011) );
  NAND3X1 U2767 ( .A(n6135), .B(n6349), .C(n6678), .Y(n4008) );
  AOI22X1 U2768 ( .A(n1359), .B(n9120), .C(n1360), .D(n8956), .Y(n4014) );
  AOI22X1 U2770 ( .A(n1362), .B(n9161), .C(n1363), .D(n9079), .Y(n4012) );
  NAND3X1 U2772 ( .A(n1366), .B(n6348), .C(n6677), .Y(n4016) );
  AOI22X1 U2773 ( .A(n1354), .B(n8710), .C(n8483), .D(n8587), .Y(n4018) );
  NAND3X1 U2775 ( .A(n6134), .B(n6347), .C(n6676), .Y(n4015) );
  AOI22X1 U2776 ( .A(n1359), .B(n8792), .C(n1360), .D(n8628), .Y(n4021) );
  AOI22X1 U2778 ( .A(n1362), .B(n8833), .C(n1363), .D(n8751), .Y(n4019) );
  NAND3X1 U2780 ( .A(n8433), .B(n6346), .C(n6675), .Y(n4023) );
  AOI22X1 U2781 ( .A(n1354), .B(n9694), .C(n8483), .D(n9571), .Y(n4025) );
  NAND3X1 U2783 ( .A(n6133), .B(n6345), .C(n6674), .Y(n4022) );
  AOI22X1 U2784 ( .A(n1359), .B(n9776), .C(n1360), .D(n9612), .Y(n4028) );
  AOI22X1 U2786 ( .A(n1362), .B(n9817), .C(n1363), .D(n9735), .Y(n4026) );
  NAND3X1 U2787 ( .A(n1382), .B(n6344), .C(n6673), .Y(n4030) );
  AOI22X1 U2788 ( .A(n1354), .B(n9366), .C(n8483), .D(n9243), .Y(n4032) );
  NAND3X1 U2790 ( .A(n6132), .B(n6343), .C(n6672), .Y(n4029) );
  AOI22X1 U2791 ( .A(n1359), .B(n9448), .C(n1360), .D(n9284), .Y(n4035) );
  AOI22X1 U2793 ( .A(n1362), .B(n9489), .C(n1363), .D(n9407), .Y(n4033) );
  NAND3X1 U2795 ( .A(n6293), .B(n4037), .C(n4038), .Y(n5547) );
  NOR3X1 U2796 ( .A(n6992), .B(n7033), .C(n7074), .Y(n4038) );
  NAND3X1 U2798 ( .A(n4046), .B(n6342), .C(n6671), .Y(n4043) );
  AOI22X1 U2799 ( .A(n1354), .B(n9039), .C(n8483), .D(n8916), .Y(n4045) );
  NAND3X1 U2801 ( .A(n6131), .B(n6341), .C(n6670), .Y(n4042) );
  AOI22X1 U2802 ( .A(n1359), .B(n9121), .C(n1360), .D(n8957), .Y(n4049) );
  AOI22X1 U2804 ( .A(n1362), .B(n9162), .C(n1363), .D(n9080), .Y(n4047) );
  NAND3X1 U2806 ( .A(n1366), .B(n6340), .C(n6669), .Y(n4051) );
  AOI22X1 U2807 ( .A(n1354), .B(n8711), .C(n8483), .D(n8588), .Y(n4053) );
  NAND3X1 U2809 ( .A(n6130), .B(n6339), .C(n6668), .Y(n4050) );
  AOI22X1 U2810 ( .A(n1359), .B(n8793), .C(n1360), .D(n8629), .Y(n4057) );
  AOI22X1 U2812 ( .A(n1362), .B(n8834), .C(n1363), .D(n8752), .Y(n4055) );
  NAND3X1 U2814 ( .A(n8433), .B(n6338), .C(n6667), .Y(n4059) );
  AOI22X1 U2815 ( .A(n1354), .B(n9695), .C(n8483), .D(n9572), .Y(n4061) );
  NOR3X1 U2817 ( .A(n15), .B(n16), .C(n8241), .Y(n1374) );
  NAND3X1 U2818 ( .A(n6129), .B(n6337), .C(n6666), .Y(n4058) );
  AOI22X1 U2819 ( .A(n1359), .B(n9777), .C(n1360), .D(n9613), .Y(n4065) );
  AOI22X1 U2821 ( .A(n1362), .B(n9818), .C(n1363), .D(n9736), .Y(n4063) );
  NAND3X1 U2822 ( .A(n1382), .B(n6336), .C(n6665), .Y(n4067) );
  AOI22X1 U2823 ( .A(n1354), .B(n9367), .C(n8483), .D(n9244), .Y(n4069) );
  NOR3X1 U2824 ( .A(n8512), .B(n12), .C(n8513), .Y(n1355) );
  NAND3X1 U2826 ( .A(n6128), .B(n6335), .C(n6664), .Y(n4066) );
  AOI22X1 U2827 ( .A(n1359), .B(n9449), .C(n1360), .D(n9285), .Y(n4072) );
  AOI22X1 U2829 ( .A(n1362), .B(n9490), .C(n1363), .D(n9408), .Y(n4070) );
  OAI21X1 U2832 ( .A(wr_ptr[0]), .B(n8424), .C(n4077), .Y(n3163) );
  NAND3X1 U2833 ( .A(n6292), .B(n8422), .C(n6663), .Y(n3162) );
  AOI22X1 U2834 ( .A(n4054), .B(n8331), .C(n4082), .D(n16), .Y(n4080) );
  NOR3X1 U2837 ( .A(n8514), .B(n16), .C(n8241), .Y(n1382) );
  OAI21X1 U2838 ( .A(n8511), .B(n8149), .C(n7971), .Y(n3161) );
  OAI21X1 U2840 ( .A(n7116), .B(n8512), .C(n5766), .Y(n3160) );
  NAND3X1 U2841 ( .A(n12), .B(n8512), .C(n4062), .Y(n4085) );
  OAI21X1 U2842 ( .A(n7116), .B(n8513), .C(n4086), .Y(n3159) );
  OAI21X1 U2843 ( .A(n1354), .B(n4073), .C(n4062), .Y(n4086) );
  AOI21X1 U2844 ( .A(n8511), .B(n4062), .C(n4082), .Y(n4084) );
  OAI21X1 U2845 ( .A(n6334), .B(n8514), .C(n5765), .Y(n3158) );
  NAND3X1 U2846 ( .A(n4062), .B(n8514), .C(n8427), .Y(n4088) );
  AOI21X1 U2847 ( .A(n4062), .B(n8331), .C(n4082), .Y(n4087) );
  NAND3X1 U2848 ( .A(n13), .B(n12), .C(n14), .Y(n4081) );
  NAND3X1 U2852 ( .A(n4090), .B(n4091), .C(n4092), .Y(n5721) );
  NOR3X1 U2853 ( .A(n4093), .B(fillcount[0]), .C(n4094), .Y(n4092) );
  OAI21X1 U2854 ( .A(n8058), .B(n8515), .C(n8057), .Y(n3157) );
  NAND3X1 U2855 ( .A(n8509), .B(n4076), .C(n8059), .Y(n4096) );
  AOI21X1 U2857 ( .A(n4076), .B(n8518), .C(n4098), .Y(n4095) );
  OAI21X1 U2858 ( .A(n8507), .B(n8516), .C(n7709), .Y(n3156) );
  NAND3X1 U2859 ( .A(wr_ptr[0]), .B(n8516), .C(n4076), .Y(n4099) );
  OAI21X1 U2860 ( .A(n7795), .B(n8517), .C(n4102), .Y(n3155) );
  AOI21X1 U2861 ( .A(n4076), .B(n8516), .C(n4100), .Y(n4101) );
  OAI21X1 U2862 ( .A(wr_ptr[0]), .B(n8424), .C(n8332), .Y(n4100) );
  OAI21X1 U2863 ( .A(n8508), .B(n8518), .C(n7968), .Y(n3154) );
  NAND3X1 U2864 ( .A(n4076), .B(n8518), .C(n8509), .Y(n4104) );
  OAI21X1 U2865 ( .A(n8509), .B(n8424), .C(n8332), .Y(n4098) );
  OAI21X1 U2868 ( .A(n4106), .B(n8519), .C(n8154), .Y(n3153) );
  OAI21X1 U2870 ( .A(n4106), .B(n8520), .C(n7972), .Y(n3152) );
  OAI21X1 U2872 ( .A(n4106), .B(n8521), .C(n7883), .Y(n3151) );
  OAI21X1 U2874 ( .A(n4106), .B(n8522), .C(n7796), .Y(n3150) );
  OAI21X1 U2876 ( .A(n4106), .B(n8523), .C(n7710), .Y(n3149) );
  OAI21X1 U2878 ( .A(n4106), .B(n8524), .C(n5798), .Y(n3148) );
  OAI21X1 U2880 ( .A(n4106), .B(n8525), .C(n7973), .Y(n3147) );
  OAI21X1 U2882 ( .A(n4106), .B(n8526), .C(n7884), .Y(n3146) );
  OAI21X1 U2884 ( .A(n4106), .B(n8527), .C(n7797), .Y(n3145) );
  OAI21X1 U2886 ( .A(n4106), .B(n8528), .C(n7711), .Y(n3144) );
  OAI21X1 U2888 ( .A(n4106), .B(n8529), .C(n7263), .Y(n3143) );
  OAI21X1 U2890 ( .A(n4106), .B(n8530), .C(n7190), .Y(n3142) );
  OAI21X1 U2892 ( .A(n4106), .B(n8531), .C(n7117), .Y(n3141) );
  OAI21X1 U2894 ( .A(n4106), .B(n8532), .C(n7634), .Y(n3140) );
  OAI21X1 U2896 ( .A(n4106), .B(n8533), .C(n7559), .Y(n3139) );
  OAI21X1 U2898 ( .A(n4106), .B(n8534), .C(n7484), .Y(n3138) );
  OAI21X1 U2900 ( .A(n4106), .B(n8535), .C(n7409), .Y(n3137) );
  OAI21X1 U2902 ( .A(n4106), .B(n8536), .C(n8335), .Y(n3136) );
  OAI21X1 U2904 ( .A(n4106), .B(n8537), .C(n8244), .Y(n3135) );
  OAI21X1 U2906 ( .A(n4106), .B(n8538), .C(n8155), .Y(n3134) );
  OAI21X1 U2908 ( .A(n4106), .B(n8539), .C(n8062), .Y(n3133) );
  OAI21X1 U2910 ( .A(n4106), .B(n8540), .C(n7336), .Y(n3132) );
  OAI21X1 U2912 ( .A(n4106), .B(n8541), .C(n7264), .Y(n3131) );
  OAI21X1 U2914 ( .A(n4106), .B(n8542), .C(n7191), .Y(n3130) );
  OAI21X1 U2916 ( .A(n4106), .B(n8543), .C(n7118), .Y(n3129) );
  OAI21X1 U2918 ( .A(n4106), .B(n8544), .C(n7635), .Y(n3128) );
  OAI21X1 U2920 ( .A(n4106), .B(n8545), .C(n7560), .Y(n3127) );
  OAI21X1 U2922 ( .A(n4106), .B(n8546), .C(n7485), .Y(n3126) );
  OAI21X1 U2924 ( .A(n4106), .B(n8547), .C(n7410), .Y(n3125) );
  OAI21X1 U2926 ( .A(n4106), .B(n8548), .C(n8336), .Y(n3124) );
  OAI21X1 U2928 ( .A(n4106), .B(n8549), .C(n8245), .Y(n3123) );
  OAI21X1 U2930 ( .A(n4106), .B(n8550), .C(n8156), .Y(n3122) );
  OAI21X1 U2932 ( .A(n4106), .B(n8551), .C(n8063), .Y(n3121) );
  OAI21X1 U2934 ( .A(n4106), .B(n8552), .C(n7337), .Y(n3120) );
  OAI21X1 U2936 ( .A(n4106), .B(n8553), .C(n7265), .Y(n3119) );
  OAI21X1 U2938 ( .A(n4106), .B(n8554), .C(n7192), .Y(n3118) );
  OAI21X1 U2940 ( .A(n4106), .B(n8555), .C(n7119), .Y(n3117) );
  OAI21X1 U2942 ( .A(n4106), .B(n8556), .C(n7636), .Y(n3116) );
  OAI21X1 U2944 ( .A(n4106), .B(n8557), .C(n7561), .Y(n3115) );
  OAI21X1 U2946 ( .A(n4106), .B(n8558), .C(n7486), .Y(n3114) );
  OAI21X1 U2948 ( .A(n4106), .B(n8559), .C(n7411), .Y(n3113) );
  OAI21X1 U2950 ( .A(n8153), .B(n8425), .C(n8501), .Y(n4106) );
  OAI21X1 U2951 ( .A(n4190), .B(n8560), .C(n8064), .Y(n3112) );
  OAI21X1 U2953 ( .A(n4190), .B(n8561), .C(n7885), .Y(n3111) );
  OAI21X1 U2955 ( .A(n4190), .B(n8562), .C(n7974), .Y(n3110) );
  OAI21X1 U2957 ( .A(n4190), .B(n8563), .C(n7712), .Y(n3109) );
  OAI21X1 U2959 ( .A(n4190), .B(n8564), .C(n7798), .Y(n3108) );
  OAI21X1 U2961 ( .A(n4190), .B(n8565), .C(n5797), .Y(n3107) );
  OAI21X1 U2963 ( .A(n4190), .B(n8566), .C(n7886), .Y(n3106) );
  OAI21X1 U2965 ( .A(n4190), .B(n8567), .C(n7975), .Y(n3105) );
  OAI21X1 U2967 ( .A(n4190), .B(n8568), .C(n7713), .Y(n3104) );
  OAI21X1 U2969 ( .A(n4190), .B(n8569), .C(n7799), .Y(n3103) );
  OAI21X1 U2971 ( .A(n4190), .B(n8570), .C(n7338), .Y(n3102) );
  OAI21X1 U2973 ( .A(n4190), .B(n8571), .C(n7120), .Y(n3101) );
  OAI21X1 U2975 ( .A(n4190), .B(n8572), .C(n7193), .Y(n3100) );
  OAI21X1 U2977 ( .A(n4190), .B(n8573), .C(n7562), .Y(n3099) );
  OAI21X1 U2979 ( .A(n4190), .B(n8574), .C(n7637), .Y(n3098) );
  OAI21X1 U2981 ( .A(n4190), .B(n8575), .C(n7412), .Y(n3097) );
  OAI21X1 U2983 ( .A(n4190), .B(n8576), .C(n7487), .Y(n3096) );
  OAI21X1 U2985 ( .A(n4190), .B(n8577), .C(n8246), .Y(n3095) );
  OAI21X1 U2987 ( .A(n4190), .B(n8578), .C(n8337), .Y(n3094) );
  OAI21X1 U2989 ( .A(n4190), .B(n8579), .C(n8065), .Y(n3093) );
  OAI21X1 U2991 ( .A(n4190), .B(n8580), .C(n8157), .Y(n3092) );
  OAI21X1 U2993 ( .A(n4190), .B(n8581), .C(n7266), .Y(n3091) );
  OAI21X1 U2995 ( .A(n4190), .B(n8582), .C(n7339), .Y(n3090) );
  OAI21X1 U2997 ( .A(n4190), .B(n8583), .C(n7121), .Y(n3089) );
  OAI21X1 U2999 ( .A(n4190), .B(n8584), .C(n7194), .Y(n3088) );
  OAI21X1 U3001 ( .A(n4190), .B(n8585), .C(n7563), .Y(n3087) );
  OAI21X1 U3003 ( .A(n4190), .B(n8586), .C(n7638), .Y(n3086) );
  OAI21X1 U3005 ( .A(n4190), .B(n8587), .C(n7413), .Y(n3085) );
  OAI21X1 U3007 ( .A(n4190), .B(n8588), .C(n7488), .Y(n3084) );
  OAI21X1 U3009 ( .A(n4190), .B(n8589), .C(n8247), .Y(n3083) );
  OAI21X1 U3011 ( .A(n4190), .B(n8590), .C(n8338), .Y(n3082) );
  OAI21X1 U3013 ( .A(n4190), .B(n8591), .C(n8066), .Y(n3081) );
  OAI21X1 U3015 ( .A(n4190), .B(n8592), .C(n8158), .Y(n3080) );
  OAI21X1 U3017 ( .A(n4190), .B(n8593), .C(n7267), .Y(n3079) );
  OAI21X1 U3019 ( .A(n4190), .B(n8594), .C(n7340), .Y(n3078) );
  OAI21X1 U3021 ( .A(n4190), .B(n8595), .C(n7122), .Y(n3077) );
  OAI21X1 U3023 ( .A(n4190), .B(n8596), .C(n7195), .Y(n3076) );
  OAI21X1 U3025 ( .A(n4190), .B(n8597), .C(n7564), .Y(n3075) );
  OAI21X1 U3027 ( .A(n4190), .B(n8598), .C(n7639), .Y(n3074) );
  OAI21X1 U3029 ( .A(n4190), .B(n8599), .C(n7414), .Y(n3073) );
  OAI21X1 U3031 ( .A(n4190), .B(n8600), .C(n7489), .Y(n3072) );
  OAI21X1 U3033 ( .A(n8425), .B(n8060), .C(n8501), .Y(n4190) );
  OAI21X1 U3034 ( .A(n4233), .B(n8601), .C(n8339), .Y(n3071) );
  OAI21X1 U3036 ( .A(n4233), .B(n8602), .C(n7800), .Y(n3070) );
  OAI21X1 U3038 ( .A(n4233), .B(n8603), .C(n7714), .Y(n3069) );
  OAI21X1 U3040 ( .A(n4233), .B(n8604), .C(n7976), .Y(n3068) );
  OAI21X1 U3042 ( .A(n4233), .B(n8605), .C(n7887), .Y(n3067) );
  OAI21X1 U3044 ( .A(n4233), .B(n8606), .C(n5796), .Y(n3066) );
  OAI21X1 U3046 ( .A(n4233), .B(n8607), .C(n7801), .Y(n3065) );
  OAI21X1 U3048 ( .A(n4233), .B(n8608), .C(n7715), .Y(n3064) );
  OAI21X1 U3050 ( .A(n4233), .B(n8609), .C(n7977), .Y(n3063) );
  OAI21X1 U3052 ( .A(n4233), .B(n8610), .C(n7888), .Y(n3062) );
  OAI21X1 U3054 ( .A(n4233), .B(n8611), .C(n7123), .Y(n3061) );
  OAI21X1 U3056 ( .A(n4233), .B(n8612), .C(n7341), .Y(n3060) );
  OAI21X1 U3058 ( .A(n4233), .B(n8613), .C(n7268), .Y(n3059) );
  OAI21X1 U3060 ( .A(n4233), .B(n8614), .C(n7490), .Y(n3058) );
  OAI21X1 U3062 ( .A(n4233), .B(n8615), .C(n7415), .Y(n3057) );
  OAI21X1 U3064 ( .A(n4233), .B(n8616), .C(n7640), .Y(n3056) );
  OAI21X1 U3066 ( .A(n4233), .B(n8617), .C(n7565), .Y(n3055) );
  OAI21X1 U3068 ( .A(n4233), .B(n8618), .C(n8159), .Y(n3054) );
  OAI21X1 U3070 ( .A(n4233), .B(n8619), .C(n8067), .Y(n3053) );
  OAI21X1 U3072 ( .A(n4233), .B(n8620), .C(n8340), .Y(n3052) );
  OAI21X1 U3074 ( .A(n4233), .B(n8621), .C(n8248), .Y(n3051) );
  OAI21X1 U3076 ( .A(n4233), .B(n8622), .C(n7196), .Y(n3050) );
  OAI21X1 U3078 ( .A(n4233), .B(n8623), .C(n7124), .Y(n3049) );
  OAI21X1 U3080 ( .A(n4233), .B(n8624), .C(n7342), .Y(n3048) );
  OAI21X1 U3082 ( .A(n4233), .B(n8625), .C(n7269), .Y(n3047) );
  OAI21X1 U3084 ( .A(n4233), .B(n8626), .C(n7491), .Y(n3046) );
  OAI21X1 U3086 ( .A(n4233), .B(n8627), .C(n7416), .Y(n3045) );
  OAI21X1 U3088 ( .A(n4233), .B(n8628), .C(n7641), .Y(n3044) );
  OAI21X1 U3090 ( .A(n4233), .B(n8629), .C(n7566), .Y(n3043) );
  OAI21X1 U3092 ( .A(n4233), .B(n8630), .C(n8160), .Y(n3042) );
  OAI21X1 U3094 ( .A(n4233), .B(n8631), .C(n8068), .Y(n3041) );
  OAI21X1 U3096 ( .A(n4233), .B(n8632), .C(n8341), .Y(n3040) );
  OAI21X1 U3098 ( .A(n4233), .B(n8633), .C(n8249), .Y(n3039) );
  OAI21X1 U3100 ( .A(n4233), .B(n8634), .C(n7197), .Y(n3038) );
  OAI21X1 U3102 ( .A(n4233), .B(n8635), .C(n7125), .Y(n3037) );
  OAI21X1 U3104 ( .A(n4233), .B(n8636), .C(n7343), .Y(n3036) );
  OAI21X1 U3106 ( .A(n4233), .B(n8637), .C(n7270), .Y(n3035) );
  OAI21X1 U3108 ( .A(n4233), .B(n8638), .C(n7492), .Y(n3034) );
  OAI21X1 U3110 ( .A(n4233), .B(n8639), .C(n7417), .Y(n3033) );
  OAI21X1 U3112 ( .A(n4233), .B(n8640), .C(n7642), .Y(n3032) );
  OAI21X1 U3114 ( .A(n4233), .B(n8641), .C(n7567), .Y(n3031) );
  OAI21X1 U3116 ( .A(n8425), .B(n7969), .C(n8501), .Y(n4233) );
  OAI21X1 U3117 ( .A(n4276), .B(n8642), .C(n8250), .Y(n3030) );
  OAI21X1 U3119 ( .A(n4276), .B(n8643), .C(n7716), .Y(n3029) );
  OAI21X1 U3121 ( .A(n4276), .B(n8644), .C(n7802), .Y(n3028) );
  OAI21X1 U3123 ( .A(n4276), .B(n8645), .C(n7889), .Y(n3027) );
  OAI21X1 U3125 ( .A(n4276), .B(n8646), .C(n7978), .Y(n3026) );
  OAI21X1 U3127 ( .A(n4276), .B(n8647), .C(n5795), .Y(n3025) );
  OAI21X1 U3129 ( .A(n4276), .B(n8648), .C(n7717), .Y(n3024) );
  OAI21X1 U3131 ( .A(n4276), .B(n8649), .C(n7803), .Y(n3023) );
  OAI21X1 U3133 ( .A(n4276), .B(n8650), .C(n7890), .Y(n3022) );
  OAI21X1 U3135 ( .A(n4276), .B(n8651), .C(n7979), .Y(n3021) );
  OAI21X1 U3137 ( .A(n4276), .B(n8652), .C(n7198), .Y(n3020) );
  OAI21X1 U3139 ( .A(n4276), .B(n8653), .C(n7271), .Y(n3019) );
  OAI21X1 U3141 ( .A(n4276), .B(n8654), .C(n7344), .Y(n3018) );
  OAI21X1 U3143 ( .A(n4276), .B(n8655), .C(n7418), .Y(n3017) );
  OAI21X1 U3145 ( .A(n4276), .B(n8656), .C(n7493), .Y(n3016) );
  OAI21X1 U3147 ( .A(n4276), .B(n8657), .C(n7568), .Y(n3015) );
  OAI21X1 U3149 ( .A(n4276), .B(n8658), .C(n7643), .Y(n3014) );
  OAI21X1 U3151 ( .A(n4276), .B(n8659), .C(n8069), .Y(n3013) );
  OAI21X1 U3153 ( .A(n4276), .B(n8660), .C(n8161), .Y(n3012) );
  OAI21X1 U3155 ( .A(n4276), .B(n8661), .C(n8251), .Y(n3011) );
  OAI21X1 U3157 ( .A(n4276), .B(n8662), .C(n8342), .Y(n3010) );
  OAI21X1 U3159 ( .A(n4276), .B(n8663), .C(n7126), .Y(n3009) );
  OAI21X1 U3161 ( .A(n4276), .B(n8664), .C(n7199), .Y(n3008) );
  OAI21X1 U3163 ( .A(n4276), .B(n8665), .C(n7272), .Y(n3007) );
  OAI21X1 U3165 ( .A(n4276), .B(n8666), .C(n7345), .Y(n3006) );
  OAI21X1 U3167 ( .A(n4276), .B(n8667), .C(n7419), .Y(n3005) );
  OAI21X1 U3169 ( .A(n4276), .B(n8668), .C(n7494), .Y(n3004) );
  OAI21X1 U3171 ( .A(n4276), .B(n8669), .C(n7569), .Y(n3003) );
  OAI21X1 U3173 ( .A(n4276), .B(n8670), .C(n7644), .Y(n3002) );
  OAI21X1 U3175 ( .A(n4276), .B(n8671), .C(n8070), .Y(n3001) );
  OAI21X1 U3177 ( .A(n4276), .B(n8672), .C(n8162), .Y(n3000) );
  OAI21X1 U3179 ( .A(n4276), .B(n8673), .C(n8252), .Y(n2999) );
  OAI21X1 U3181 ( .A(n4276), .B(n8674), .C(n8343), .Y(n2998) );
  OAI21X1 U3183 ( .A(n4276), .B(n8675), .C(n7127), .Y(n2997) );
  OAI21X1 U3185 ( .A(n4276), .B(n8676), .C(n7200), .Y(n2996) );
  OAI21X1 U3187 ( .A(n4276), .B(n8677), .C(n7273), .Y(n2995) );
  OAI21X1 U3189 ( .A(n4276), .B(n8678), .C(n7346), .Y(n2994) );
  OAI21X1 U3191 ( .A(n4276), .B(n8679), .C(n7420), .Y(n2993) );
  OAI21X1 U3193 ( .A(n4276), .B(n8680), .C(n7495), .Y(n2992) );
  OAI21X1 U3195 ( .A(n4276), .B(n8681), .C(n7570), .Y(n2991) );
  OAI21X1 U3197 ( .A(n4276), .B(n8682), .C(n7645), .Y(n2990) );
  OAI21X1 U3199 ( .A(n8425), .B(n8242), .C(n8501), .Y(n4276) );
  OAI21X1 U3200 ( .A(n4319), .B(n8683), .C(n7201), .Y(n2989) );
  OAI21X1 U3202 ( .A(n4319), .B(n8684), .C(n7646), .Y(n2988) );
  OAI21X1 U3204 ( .A(n4319), .B(n8685), .C(n7571), .Y(n2987) );
  OAI21X1 U3206 ( .A(n4319), .B(n8686), .C(n7496), .Y(n2986) );
  OAI21X1 U3208 ( .A(n4319), .B(n8687), .C(n7421), .Y(n2985) );
  OAI21X1 U3210 ( .A(n4319), .B(n8688), .C(n5794), .Y(n2984) );
  OAI21X1 U3212 ( .A(n4319), .B(n8689), .C(n7647), .Y(n2983) );
  OAI21X1 U3214 ( .A(n4319), .B(n8690), .C(n7572), .Y(n2982) );
  OAI21X1 U3216 ( .A(n4319), .B(n8691), .C(n7497), .Y(n2981) );
  OAI21X1 U3218 ( .A(n4319), .B(n8692), .C(n7422), .Y(n2980) );
  OAI21X1 U3220 ( .A(n4319), .B(n8693), .C(n8253), .Y(n2979) );
  OAI21X1 U3222 ( .A(n4319), .B(n8694), .C(n8163), .Y(n2978) );
  OAI21X1 U3224 ( .A(n4319), .B(n8695), .C(n8071), .Y(n2977) );
  OAI21X1 U3226 ( .A(n4319), .B(n8696), .C(n7980), .Y(n2976) );
  OAI21X1 U3228 ( .A(n4319), .B(n8697), .C(n7891), .Y(n2975) );
  OAI21X1 U3230 ( .A(n4319), .B(n8698), .C(n7804), .Y(n2974) );
  OAI21X1 U3232 ( .A(n4319), .B(n8699), .C(n7718), .Y(n2973) );
  OAI21X1 U3234 ( .A(n4319), .B(n8700), .C(n7347), .Y(n2972) );
  OAI21X1 U3236 ( .A(n4319), .B(n8701), .C(n7274), .Y(n2971) );
  OAI21X1 U3238 ( .A(n4319), .B(n8702), .C(n7202), .Y(n2970) );
  OAI21X1 U3240 ( .A(n4319), .B(n8703), .C(n7128), .Y(n2969) );
  OAI21X1 U3242 ( .A(n4319), .B(n8704), .C(n8344), .Y(n2968) );
  OAI21X1 U3244 ( .A(n4319), .B(n8705), .C(n8254), .Y(n2967) );
  OAI21X1 U3246 ( .A(n4319), .B(n8706), .C(n8164), .Y(n2966) );
  OAI21X1 U3248 ( .A(n4319), .B(n8707), .C(n8072), .Y(n2965) );
  OAI21X1 U3250 ( .A(n4319), .B(n8708), .C(n7981), .Y(n2964) );
  OAI21X1 U3252 ( .A(n4319), .B(n8709), .C(n7892), .Y(n2963) );
  OAI21X1 U3254 ( .A(n4319), .B(n8710), .C(n7805), .Y(n2962) );
  OAI21X1 U3256 ( .A(n4319), .B(n8711), .C(n7719), .Y(n2961) );
  OAI21X1 U3258 ( .A(n4319), .B(n8712), .C(n7348), .Y(n2960) );
  OAI21X1 U3260 ( .A(n4319), .B(n8713), .C(n7275), .Y(n2959) );
  OAI21X1 U3262 ( .A(n4319), .B(n8714), .C(n7203), .Y(n2958) );
  OAI21X1 U3264 ( .A(n4319), .B(n8715), .C(n7129), .Y(n2957) );
  OAI21X1 U3266 ( .A(n4319), .B(n8716), .C(n8345), .Y(n2956) );
  OAI21X1 U3268 ( .A(n4319), .B(n8717), .C(n8255), .Y(n2955) );
  OAI21X1 U3270 ( .A(n4319), .B(n8718), .C(n8165), .Y(n2954) );
  OAI21X1 U3272 ( .A(n4319), .B(n8719), .C(n8073), .Y(n2953) );
  OAI21X1 U3274 ( .A(n4319), .B(n8720), .C(n7982), .Y(n2952) );
  OAI21X1 U3276 ( .A(n4319), .B(n8721), .C(n7893), .Y(n2951) );
  OAI21X1 U3278 ( .A(n4319), .B(n8722), .C(n7806), .Y(n2950) );
  OAI21X1 U3280 ( .A(n4319), .B(n8723), .C(n7720), .Y(n2949) );
  OAI21X1 U3282 ( .A(n8243), .B(n8425), .C(n8501), .Y(n4319) );
  OAI21X1 U3283 ( .A(n4361), .B(n8724), .C(n7130), .Y(n2948) );
  OAI21X1 U3285 ( .A(n4361), .B(n8725), .C(n7573), .Y(n2947) );
  OAI21X1 U3287 ( .A(n4361), .B(n8726), .C(n7648), .Y(n2946) );
  OAI21X1 U3289 ( .A(n4361), .B(n8727), .C(n7423), .Y(n2945) );
  OAI21X1 U3291 ( .A(n4361), .B(n8728), .C(n7498), .Y(n2944) );
  OAI21X1 U3293 ( .A(n4361), .B(n8729), .C(n5793), .Y(n2943) );
  OAI21X1 U3295 ( .A(n4361), .B(n8730), .C(n7574), .Y(n2942) );
  OAI21X1 U3297 ( .A(n4361), .B(n8731), .C(n7649), .Y(n2941) );
  OAI21X1 U3299 ( .A(n4361), .B(n8732), .C(n7424), .Y(n2940) );
  OAI21X1 U3301 ( .A(n4361), .B(n8733), .C(n7499), .Y(n2939) );
  OAI21X1 U3303 ( .A(n4361), .B(n8734), .C(n8346), .Y(n2938) );
  OAI21X1 U3305 ( .A(n4361), .B(n8735), .C(n8074), .Y(n2937) );
  OAI21X1 U3307 ( .A(n4361), .B(n8736), .C(n8166), .Y(n2936) );
  OAI21X1 U3309 ( .A(n4361), .B(n8737), .C(n7894), .Y(n2935) );
  OAI21X1 U3311 ( .A(n4361), .B(n8738), .C(n7983), .Y(n2934) );
  OAI21X1 U3313 ( .A(n4361), .B(n8739), .C(n7721), .Y(n2933) );
  OAI21X1 U3315 ( .A(n4361), .B(n8740), .C(n7807), .Y(n2932) );
  OAI21X1 U3317 ( .A(n4361), .B(n8741), .C(n7276), .Y(n2931) );
  OAI21X1 U3319 ( .A(n4361), .B(n8742), .C(n7349), .Y(n2930) );
  OAI21X1 U3321 ( .A(n4361), .B(n8743), .C(n7131), .Y(n2929) );
  OAI21X1 U3323 ( .A(n4361), .B(n8744), .C(n7204), .Y(n2928) );
  OAI21X1 U3325 ( .A(n4361), .B(n8745), .C(n8256), .Y(n2927) );
  OAI21X1 U3327 ( .A(n4361), .B(n8746), .C(n8347), .Y(n2926) );
  OAI21X1 U3329 ( .A(n4361), .B(n8747), .C(n8075), .Y(n2925) );
  OAI21X1 U3331 ( .A(n4361), .B(n8748), .C(n8167), .Y(n2924) );
  OAI21X1 U3333 ( .A(n4361), .B(n8749), .C(n7895), .Y(n2923) );
  OAI21X1 U3335 ( .A(n4361), .B(n8750), .C(n7984), .Y(n2922) );
  OAI21X1 U3337 ( .A(n4361), .B(n8751), .C(n7722), .Y(n2921) );
  OAI21X1 U3339 ( .A(n4361), .B(n8752), .C(n7808), .Y(n2920) );
  OAI21X1 U3341 ( .A(n4361), .B(n8753), .C(n7277), .Y(n2919) );
  OAI21X1 U3343 ( .A(n4361), .B(n8754), .C(n7350), .Y(n2918) );
  OAI21X1 U3345 ( .A(n4361), .B(n8755), .C(n7132), .Y(n2917) );
  OAI21X1 U3347 ( .A(n4361), .B(n8756), .C(n7205), .Y(n2916) );
  OAI21X1 U3349 ( .A(n4361), .B(n8757), .C(n8257), .Y(n2915) );
  OAI21X1 U3351 ( .A(n4361), .B(n8758), .C(n8348), .Y(n2914) );
  OAI21X1 U3353 ( .A(n4361), .B(n8759), .C(n8076), .Y(n2913) );
  OAI21X1 U3355 ( .A(n4361), .B(n8760), .C(n8168), .Y(n2912) );
  OAI21X1 U3357 ( .A(n4361), .B(n8761), .C(n7896), .Y(n2911) );
  OAI21X1 U3359 ( .A(n4361), .B(n8762), .C(n7985), .Y(n2910) );
  OAI21X1 U3361 ( .A(n4361), .B(n8763), .C(n7723), .Y(n2909) );
  OAI21X1 U3363 ( .A(n4361), .B(n8764), .C(n7809), .Y(n2908) );
  OAI21X1 U3365 ( .A(n8425), .B(n7970), .C(n8501), .Y(n4361) );
  OAI21X1 U3366 ( .A(n4404), .B(n8765), .C(n7351), .Y(n2907) );
  OAI21X1 U3368 ( .A(n4404), .B(n8766), .C(n7500), .Y(n2906) );
  OAI21X1 U3370 ( .A(n4404), .B(n8767), .C(n7425), .Y(n2905) );
  OAI21X1 U3372 ( .A(n4404), .B(n8768), .C(n7650), .Y(n2904) );
  OAI21X1 U3374 ( .A(n4404), .B(n8769), .C(n7575), .Y(n2903) );
  OAI21X1 U3376 ( .A(n4404), .B(n8770), .C(n5792), .Y(n2902) );
  OAI21X1 U3378 ( .A(n4404), .B(n8771), .C(n7501), .Y(n2901) );
  OAI21X1 U3380 ( .A(n4404), .B(n8772), .C(n7426), .Y(n2900) );
  OAI21X1 U3382 ( .A(n4404), .B(n8773), .C(n7651), .Y(n2899) );
  OAI21X1 U3384 ( .A(n4404), .B(n8774), .C(n7576), .Y(n2898) );
  OAI21X1 U3386 ( .A(n4404), .B(n8775), .C(n8077), .Y(n2897) );
  OAI21X1 U3388 ( .A(n4404), .B(n8776), .C(n8349), .Y(n2896) );
  OAI21X1 U3390 ( .A(n4404), .B(n8777), .C(n8258), .Y(n2895) );
  OAI21X1 U3392 ( .A(n4404), .B(n8778), .C(n7810), .Y(n2894) );
  OAI21X1 U3394 ( .A(n4404), .B(n8779), .C(n7724), .Y(n2893) );
  OAI21X1 U3396 ( .A(n4404), .B(n8780), .C(n7986), .Y(n2892) );
  OAI21X1 U3398 ( .A(n4404), .B(n8781), .C(n7897), .Y(n2891) );
  OAI21X1 U3400 ( .A(n4404), .B(n8782), .C(n7206), .Y(n2890) );
  OAI21X1 U3402 ( .A(n4404), .B(n8783), .C(n7133), .Y(n2889) );
  OAI21X1 U3404 ( .A(n4404), .B(n8784), .C(n7352), .Y(n2888) );
  OAI21X1 U3406 ( .A(n4404), .B(n8785), .C(n7278), .Y(n2887) );
  OAI21X1 U3408 ( .A(n4404), .B(n8786), .C(n8169), .Y(n2886) );
  OAI21X1 U3410 ( .A(n4404), .B(n8787), .C(n8078), .Y(n2885) );
  OAI21X1 U3412 ( .A(n4404), .B(n8788), .C(n8350), .Y(n2884) );
  OAI21X1 U3414 ( .A(n4404), .B(n8789), .C(n8259), .Y(n2883) );
  OAI21X1 U3416 ( .A(n4404), .B(n8790), .C(n7811), .Y(n2882) );
  OAI21X1 U3418 ( .A(n4404), .B(n8791), .C(n7725), .Y(n2881) );
  OAI21X1 U3420 ( .A(n4404), .B(n8792), .C(n7987), .Y(n2880) );
  OAI21X1 U3422 ( .A(n4404), .B(n8793), .C(n7898), .Y(n2879) );
  OAI21X1 U3424 ( .A(n4404), .B(n8794), .C(n7207), .Y(n2878) );
  OAI21X1 U3426 ( .A(n4404), .B(n8795), .C(n7134), .Y(n2877) );
  OAI21X1 U3428 ( .A(n4404), .B(n8796), .C(n7353), .Y(n2876) );
  OAI21X1 U3430 ( .A(n4404), .B(n8797), .C(n7279), .Y(n2875) );
  OAI21X1 U3432 ( .A(n4404), .B(n8798), .C(n8170), .Y(n2874) );
  OAI21X1 U3434 ( .A(n4404), .B(n8799), .C(n8079), .Y(n2873) );
  OAI21X1 U3436 ( .A(n4404), .B(n8800), .C(n8351), .Y(n2872) );
  OAI21X1 U3438 ( .A(n4404), .B(n8801), .C(n8260), .Y(n2871) );
  OAI21X1 U3440 ( .A(n4404), .B(n8802), .C(n7812), .Y(n2870) );
  OAI21X1 U3442 ( .A(n4404), .B(n8803), .C(n7726), .Y(n2869) );
  OAI21X1 U3444 ( .A(n4404), .B(n8804), .C(n7988), .Y(n2868) );
  OAI21X1 U3446 ( .A(n4404), .B(n8805), .C(n7899), .Y(n2867) );
  OAI21X1 U3448 ( .A(n8425), .B(n8061), .C(n8501), .Y(n4404) );
  OAI21X1 U3449 ( .A(n4447), .B(n8806), .C(n7280), .Y(n2866) );
  OAI21X1 U3451 ( .A(n4447), .B(n8807), .C(n7427), .Y(n2865) );
  OAI21X1 U3453 ( .A(n4447), .B(n8808), .C(n7502), .Y(n2864) );
  OAI21X1 U3455 ( .A(n4447), .B(n8809), .C(n7577), .Y(n2863) );
  OAI21X1 U3457 ( .A(n4447), .B(n8810), .C(n7652), .Y(n2862) );
  OAI21X1 U3459 ( .A(n4447), .B(n8811), .C(n5791), .Y(n2861) );
  OAI21X1 U3461 ( .A(n4447), .B(n8812), .C(n7428), .Y(n2860) );
  OAI21X1 U3463 ( .A(n4447), .B(n8813), .C(n7503), .Y(n2859) );
  OAI21X1 U3465 ( .A(n4447), .B(n8814), .C(n7578), .Y(n2858) );
  OAI21X1 U3467 ( .A(n4447), .B(n8815), .C(n7653), .Y(n2857) );
  OAI21X1 U3469 ( .A(n4447), .B(n8816), .C(n8171), .Y(n2856) );
  OAI21X1 U3471 ( .A(n4447), .B(n8817), .C(n8261), .Y(n2855) );
  OAI21X1 U3473 ( .A(n4447), .B(n8818), .C(n8352), .Y(n2854) );
  OAI21X1 U3475 ( .A(n4447), .B(n8819), .C(n7727), .Y(n2853) );
  OAI21X1 U3477 ( .A(n4447), .B(n8820), .C(n7813), .Y(n2852) );
  OAI21X1 U3479 ( .A(n4447), .B(n8821), .C(n7900), .Y(n2851) );
  OAI21X1 U3481 ( .A(n4447), .B(n8822), .C(n7989), .Y(n2850) );
  OAI21X1 U3483 ( .A(n4447), .B(n8823), .C(n7135), .Y(n2849) );
  OAI21X1 U3485 ( .A(n4447), .B(n8824), .C(n7208), .Y(n2848) );
  OAI21X1 U3487 ( .A(n4447), .B(n8825), .C(n7281), .Y(n2847) );
  OAI21X1 U3489 ( .A(n4447), .B(n8826), .C(n7354), .Y(n2846) );
  OAI21X1 U3491 ( .A(n4447), .B(n8827), .C(n8080), .Y(n2845) );
  OAI21X1 U3493 ( .A(n4447), .B(n8828), .C(n8172), .Y(n2844) );
  OAI21X1 U3495 ( .A(n4447), .B(n8829), .C(n8262), .Y(n2843) );
  OAI21X1 U3497 ( .A(n4447), .B(n8830), .C(n8353), .Y(n2842) );
  OAI21X1 U3499 ( .A(n4447), .B(n8831), .C(n7728), .Y(n2841) );
  OAI21X1 U3501 ( .A(n4447), .B(n8832), .C(n7814), .Y(n2840) );
  OAI21X1 U3503 ( .A(n4447), .B(n8833), .C(n7901), .Y(n2839) );
  OAI21X1 U3505 ( .A(n4447), .B(n8834), .C(n7990), .Y(n2838) );
  OAI21X1 U3507 ( .A(n4447), .B(n8835), .C(n7136), .Y(n2837) );
  OAI21X1 U3509 ( .A(n4447), .B(n8836), .C(n7209), .Y(n2836) );
  OAI21X1 U3511 ( .A(n4447), .B(n8837), .C(n7282), .Y(n2835) );
  OAI21X1 U3513 ( .A(n4447), .B(n8838), .C(n7355), .Y(n2834) );
  OAI21X1 U3515 ( .A(n4447), .B(n8839), .C(n8081), .Y(n2833) );
  OAI21X1 U3517 ( .A(n4447), .B(n8840), .C(n8173), .Y(n2832) );
  OAI21X1 U3519 ( .A(n4447), .B(n8841), .C(n8263), .Y(n2831) );
  OAI21X1 U3521 ( .A(n4447), .B(n8842), .C(n8354), .Y(n2830) );
  OAI21X1 U3523 ( .A(n4447), .B(n8843), .C(n7729), .Y(n2829) );
  OAI21X1 U3525 ( .A(n4447), .B(n8844), .C(n7815), .Y(n2828) );
  OAI21X1 U3527 ( .A(n4447), .B(n8845), .C(n7902), .Y(n2827) );
  OAI21X1 U3529 ( .A(n4447), .B(n8846), .C(n7991), .Y(n2826) );
  OAI21X1 U3531 ( .A(n8425), .B(n8152), .C(n8501), .Y(n4447) );
  NAND3X1 U3532 ( .A(wr_ptr[4]), .B(wr_ptr[3]), .C(put), .Y(n4189) );
  OAI21X1 U3533 ( .A(n4490), .B(n8847), .C(n7504), .Y(n2825) );
  OAI21X1 U3535 ( .A(n4490), .B(n8848), .C(n7356), .Y(n2824) );
  OAI21X1 U3537 ( .A(n4490), .B(n8849), .C(n7283), .Y(n2823) );
  OAI21X1 U3539 ( .A(n4490), .B(n8850), .C(n7210), .Y(n2822) );
  OAI21X1 U3541 ( .A(n4490), .B(n8851), .C(n7137), .Y(n2821) );
  OAI21X1 U3543 ( .A(n4490), .B(n8852), .C(n5790), .Y(n2820) );
  OAI21X1 U3545 ( .A(n4490), .B(n8853), .C(n7357), .Y(n2819) );
  OAI21X1 U3547 ( .A(n4490), .B(n8854), .C(n7284), .Y(n2818) );
  OAI21X1 U3549 ( .A(n4490), .B(n8855), .C(n7211), .Y(n2817) );
  OAI21X1 U3551 ( .A(n4490), .B(n8856), .C(n7138), .Y(n2816) );
  OAI21X1 U3553 ( .A(n4490), .B(n8857), .C(n7903), .Y(n2815) );
  OAI21X1 U3555 ( .A(n4490), .B(n8858), .C(n7816), .Y(n2814) );
  OAI21X1 U3557 ( .A(n4490), .B(n8859), .C(n7730), .Y(n2813) );
  OAI21X1 U3559 ( .A(n4490), .B(n8860), .C(n8355), .Y(n2812) );
  OAI21X1 U3561 ( .A(n4490), .B(n8861), .C(n8264), .Y(n2811) );
  OAI21X1 U3563 ( .A(n4490), .B(n8862), .C(n8174), .Y(n2810) );
  OAI21X1 U3565 ( .A(n4490), .B(n8863), .C(n8082), .Y(n2809) );
  OAI21X1 U3567 ( .A(n4490), .B(n8864), .C(n7654), .Y(n2808) );
  OAI21X1 U3569 ( .A(n4490), .B(n8865), .C(n7579), .Y(n2807) );
  OAI21X1 U3571 ( .A(n4490), .B(n8866), .C(n7505), .Y(n2806) );
  OAI21X1 U3573 ( .A(n4490), .B(n8867), .C(n7429), .Y(n2805) );
  OAI21X1 U3575 ( .A(n4490), .B(n8868), .C(n7992), .Y(n2804) );
  OAI21X1 U3577 ( .A(n4490), .B(n8869), .C(n7904), .Y(n2803) );
  OAI21X1 U3579 ( .A(n4490), .B(n8870), .C(n7817), .Y(n2802) );
  OAI21X1 U3581 ( .A(n4490), .B(n8871), .C(n7731), .Y(n2801) );
  OAI21X1 U3583 ( .A(n4490), .B(n8872), .C(n8356), .Y(n2800) );
  OAI21X1 U3585 ( .A(n4490), .B(n8873), .C(n8265), .Y(n2799) );
  OAI21X1 U3587 ( .A(n4490), .B(n8874), .C(n8175), .Y(n2798) );
  OAI21X1 U3589 ( .A(n4490), .B(n8875), .C(n8083), .Y(n2797) );
  OAI21X1 U3591 ( .A(n4490), .B(n8876), .C(n7655), .Y(n2796) );
  OAI21X1 U3593 ( .A(n4490), .B(n8877), .C(n7580), .Y(n2795) );
  OAI21X1 U3595 ( .A(n4490), .B(n8878), .C(n7506), .Y(n2794) );
  OAI21X1 U3597 ( .A(n4490), .B(n8879), .C(n7430), .Y(n2793) );
  OAI21X1 U3599 ( .A(n4490), .B(n8880), .C(n7993), .Y(n2792) );
  OAI21X1 U3601 ( .A(n4490), .B(n8881), .C(n7905), .Y(n2791) );
  OAI21X1 U3603 ( .A(n4490), .B(n8882), .C(n7818), .Y(n2790) );
  OAI21X1 U3605 ( .A(n4490), .B(n8883), .C(n7732), .Y(n2789) );
  OAI21X1 U3607 ( .A(n4490), .B(n8884), .C(n8357), .Y(n2788) );
  OAI21X1 U3609 ( .A(n4490), .B(n8885), .C(n8266), .Y(n2787) );
  OAI21X1 U3611 ( .A(n4490), .B(n8886), .C(n8176), .Y(n2786) );
  OAI21X1 U3613 ( .A(n4490), .B(n8887), .C(n8084), .Y(n2785) );
  OAI21X1 U3615 ( .A(n8153), .B(n8333), .C(n8500), .Y(n4490) );
  OAI21X1 U3616 ( .A(n4533), .B(n8888), .C(n7431), .Y(n2784) );
  OAI21X1 U3618 ( .A(n4533), .B(n8889), .C(n7285), .Y(n2783) );
  OAI21X1 U3620 ( .A(n4533), .B(n8890), .C(n7358), .Y(n2782) );
  OAI21X1 U3622 ( .A(n4533), .B(n8891), .C(n7139), .Y(n2781) );
  OAI21X1 U3624 ( .A(n4533), .B(n8892), .C(n7212), .Y(n2780) );
  OAI21X1 U3626 ( .A(n4533), .B(n8893), .C(n5789), .Y(n2779) );
  OAI21X1 U3628 ( .A(n4533), .B(n8894), .C(n7286), .Y(n2778) );
  OAI21X1 U3630 ( .A(n4533), .B(n8895), .C(n7359), .Y(n2777) );
  OAI21X1 U3632 ( .A(n4533), .B(n8896), .C(n7140), .Y(n2776) );
  OAI21X1 U3634 ( .A(n4533), .B(n8897), .C(n7213), .Y(n2775) );
  OAI21X1 U3636 ( .A(n4533), .B(n8898), .C(n7994), .Y(n2774) );
  OAI21X1 U3638 ( .A(n4533), .B(n8899), .C(n7733), .Y(n2773) );
  OAI21X1 U3640 ( .A(n4533), .B(n8900), .C(n7819), .Y(n2772) );
  OAI21X1 U3642 ( .A(n4533), .B(n8901), .C(n8267), .Y(n2771) );
  OAI21X1 U3644 ( .A(n4533), .B(n8902), .C(n8358), .Y(n2770) );
  OAI21X1 U3646 ( .A(n4533), .B(n8903), .C(n8085), .Y(n2769) );
  OAI21X1 U3648 ( .A(n4533), .B(n8904), .C(n8177), .Y(n2768) );
  OAI21X1 U3650 ( .A(n4533), .B(n8905), .C(n7581), .Y(n2767) );
  OAI21X1 U3652 ( .A(n4533), .B(n8906), .C(n7656), .Y(n2766) );
  OAI21X1 U3654 ( .A(n4533), .B(n8907), .C(n7432), .Y(n2765) );
  OAI21X1 U3656 ( .A(n4533), .B(n8908), .C(n7507), .Y(n2764) );
  OAI21X1 U3658 ( .A(n4533), .B(n8909), .C(n7906), .Y(n2763) );
  OAI21X1 U3660 ( .A(n4533), .B(n8910), .C(n7995), .Y(n2762) );
  OAI21X1 U3662 ( .A(n4533), .B(n8911), .C(n7734), .Y(n2761) );
  OAI21X1 U3664 ( .A(n4533), .B(n8912), .C(n7820), .Y(n2760) );
  OAI21X1 U3666 ( .A(n4533), .B(n8913), .C(n8268), .Y(n2759) );
  OAI21X1 U3668 ( .A(n4533), .B(n8914), .C(n8359), .Y(n2758) );
  OAI21X1 U3670 ( .A(n4533), .B(n8915), .C(n8086), .Y(n2757) );
  OAI21X1 U3672 ( .A(n4533), .B(n8916), .C(n8178), .Y(n2756) );
  OAI21X1 U3674 ( .A(n4533), .B(n8917), .C(n7582), .Y(n2755) );
  OAI21X1 U3676 ( .A(n4533), .B(n8918), .C(n7657), .Y(n2754) );
  OAI21X1 U3678 ( .A(n4533), .B(n8919), .C(n7433), .Y(n2753) );
  OAI21X1 U3680 ( .A(n4533), .B(n8920), .C(n7508), .Y(n2752) );
  OAI21X1 U3682 ( .A(n4533), .B(n8921), .C(n7907), .Y(n2751) );
  OAI21X1 U3684 ( .A(n4533), .B(n8922), .C(n7996), .Y(n2750) );
  OAI21X1 U3686 ( .A(n4533), .B(n8923), .C(n7735), .Y(n2749) );
  OAI21X1 U3688 ( .A(n4533), .B(n8924), .C(n7821), .Y(n2748) );
  OAI21X1 U3690 ( .A(n4533), .B(n8925), .C(n8269), .Y(n2747) );
  OAI21X1 U3692 ( .A(n4533), .B(n8926), .C(n8360), .Y(n2746) );
  OAI21X1 U3694 ( .A(n4533), .B(n8927), .C(n8087), .Y(n2745) );
  OAI21X1 U3696 ( .A(n4533), .B(n8928), .C(n8179), .Y(n2744) );
  OAI21X1 U3698 ( .A(n8060), .B(n8333), .C(n8501), .Y(n4533) );
  OAI21X1 U3699 ( .A(n4575), .B(n8929), .C(n7658), .Y(n2743) );
  OAI21X1 U3701 ( .A(n4575), .B(n8930), .C(n7214), .Y(n2742) );
  OAI21X1 U3703 ( .A(n4575), .B(n8931), .C(n7141), .Y(n2741) );
  OAI21X1 U3705 ( .A(n4575), .B(n8932), .C(n7360), .Y(n2740) );
  OAI21X1 U3707 ( .A(n4575), .B(n8933), .C(n7287), .Y(n2739) );
  OAI21X1 U3709 ( .A(n4575), .B(n8934), .C(n5788), .Y(n2738) );
  OAI21X1 U3711 ( .A(n4575), .B(n8935), .C(n7215), .Y(n2737) );
  OAI21X1 U3713 ( .A(n4575), .B(n8936), .C(n7142), .Y(n2736) );
  OAI21X1 U3715 ( .A(n4575), .B(n8937), .C(n7361), .Y(n2735) );
  OAI21X1 U3717 ( .A(n4575), .B(n8938), .C(n7288), .Y(n2734) );
  OAI21X1 U3719 ( .A(n4575), .B(n8939), .C(n7736), .Y(n2733) );
  OAI21X1 U3721 ( .A(n4575), .B(n8940), .C(n7997), .Y(n2732) );
  OAI21X1 U3723 ( .A(n4575), .B(n8941), .C(n7908), .Y(n2731) );
  OAI21X1 U3725 ( .A(n4575), .B(n8942), .C(n8180), .Y(n2730) );
  OAI21X1 U3727 ( .A(n4575), .B(n8943), .C(n8088), .Y(n2729) );
  OAI21X1 U3729 ( .A(n4575), .B(n8944), .C(n8361), .Y(n2728) );
  OAI21X1 U3731 ( .A(n4575), .B(n8945), .C(n8270), .Y(n2727) );
  OAI21X1 U3733 ( .A(n4575), .B(n8946), .C(n7509), .Y(n2726) );
  OAI21X1 U3735 ( .A(n4575), .B(n8947), .C(n7434), .Y(n2725) );
  OAI21X1 U3737 ( .A(n4575), .B(n8948), .C(n7659), .Y(n2724) );
  OAI21X1 U3739 ( .A(n4575), .B(n8949), .C(n7583), .Y(n2723) );
  OAI21X1 U3741 ( .A(n4575), .B(n8950), .C(n7822), .Y(n2722) );
  OAI21X1 U3743 ( .A(n4575), .B(n8951), .C(n7737), .Y(n2721) );
  OAI21X1 U3745 ( .A(n4575), .B(n8952), .C(n7998), .Y(n2720) );
  OAI21X1 U3747 ( .A(n4575), .B(n8953), .C(n7909), .Y(n2719) );
  OAI21X1 U3749 ( .A(n4575), .B(n8954), .C(n8181), .Y(n2718) );
  OAI21X1 U3751 ( .A(n4575), .B(n8955), .C(n8089), .Y(n2717) );
  OAI21X1 U3753 ( .A(n4575), .B(n8956), .C(n8362), .Y(n2716) );
  OAI21X1 U3755 ( .A(n4575), .B(n8957), .C(n8271), .Y(n2715) );
  OAI21X1 U3757 ( .A(n4575), .B(n8958), .C(n7510), .Y(n2714) );
  OAI21X1 U3759 ( .A(n4575), .B(n8959), .C(n7435), .Y(n2713) );
  OAI21X1 U3761 ( .A(n4575), .B(n8960), .C(n7660), .Y(n2712) );
  OAI21X1 U3763 ( .A(n4575), .B(n8961), .C(n7584), .Y(n2711) );
  OAI21X1 U3765 ( .A(n4575), .B(n8962), .C(n7823), .Y(n2710) );
  OAI21X1 U3767 ( .A(n4575), .B(n8963), .C(n7738), .Y(n2709) );
  OAI21X1 U3769 ( .A(n4575), .B(n8964), .C(n7999), .Y(n2708) );
  OAI21X1 U3771 ( .A(n4575), .B(n8965), .C(n7910), .Y(n2707) );
  OAI21X1 U3773 ( .A(n4575), .B(n8966), .C(n8182), .Y(n2706) );
  OAI21X1 U3775 ( .A(n4575), .B(n8967), .C(n8090), .Y(n2705) );
  OAI21X1 U3777 ( .A(n4575), .B(n8968), .C(n8363), .Y(n2704) );
  OAI21X1 U3779 ( .A(n4575), .B(n8969), .C(n8272), .Y(n2703) );
  OAI21X1 U3781 ( .A(n7969), .B(n8333), .C(n8500), .Y(n4575) );
  OAI21X1 U3782 ( .A(n4617), .B(n8970), .C(n7585), .Y(n2702) );
  OAI21X1 U3784 ( .A(n4617), .B(n8971), .C(n7143), .Y(n2701) );
  OAI21X1 U3786 ( .A(n4617), .B(n8972), .C(n7216), .Y(n2700) );
  OAI21X1 U3788 ( .A(n4617), .B(n8973), .C(n7289), .Y(n2699) );
  OAI21X1 U3790 ( .A(n4617), .B(n8974), .C(n7362), .Y(n2698) );
  OAI21X1 U3792 ( .A(n4617), .B(n8975), .C(n5787), .Y(n2697) );
  OAI21X1 U3794 ( .A(n4617), .B(n8976), .C(n7144), .Y(n2696) );
  OAI21X1 U3796 ( .A(n4617), .B(n8977), .C(n7217), .Y(n2695) );
  OAI21X1 U3798 ( .A(n4617), .B(n8978), .C(n7290), .Y(n2694) );
  OAI21X1 U3800 ( .A(n4617), .B(n8979), .C(n7363), .Y(n2693) );
  OAI21X1 U3802 ( .A(n4617), .B(n8980), .C(n7824), .Y(n2692) );
  OAI21X1 U3804 ( .A(n4617), .B(n8981), .C(n7911), .Y(n2691) );
  OAI21X1 U3806 ( .A(n4617), .B(n8982), .C(n8000), .Y(n2690) );
  OAI21X1 U3808 ( .A(n4617), .B(n8983), .C(n8091), .Y(n2689) );
  OAI21X1 U3810 ( .A(n4617), .B(n8984), .C(n8183), .Y(n2688) );
  OAI21X1 U3812 ( .A(n4617), .B(n8985), .C(n8273), .Y(n2687) );
  OAI21X1 U3814 ( .A(n4617), .B(n8986), .C(n8364), .Y(n2686) );
  OAI21X1 U3816 ( .A(n4617), .B(n8987), .C(n7436), .Y(n2685) );
  OAI21X1 U3818 ( .A(n4617), .B(n8988), .C(n7511), .Y(n2684) );
  OAI21X1 U3820 ( .A(n4617), .B(n8989), .C(n7586), .Y(n2683) );
  OAI21X1 U3822 ( .A(n4617), .B(n8990), .C(n7661), .Y(n2682) );
  OAI21X1 U3824 ( .A(n4617), .B(n8991), .C(n7739), .Y(n2681) );
  OAI21X1 U3826 ( .A(n4617), .B(n8992), .C(n7825), .Y(n2680) );
  OAI21X1 U3828 ( .A(n4617), .B(n8993), .C(n7912), .Y(n2679) );
  OAI21X1 U3830 ( .A(n4617), .B(n8994), .C(n8001), .Y(n2678) );
  OAI21X1 U3832 ( .A(n4617), .B(n8995), .C(n8092), .Y(n2677) );
  OAI21X1 U3834 ( .A(n4617), .B(n8996), .C(n8184), .Y(n2676) );
  OAI21X1 U3836 ( .A(n4617), .B(n8997), .C(n8274), .Y(n2675) );
  OAI21X1 U3838 ( .A(n4617), .B(n8998), .C(n8365), .Y(n2674) );
  OAI21X1 U3840 ( .A(n4617), .B(n8999), .C(n7437), .Y(n2673) );
  OAI21X1 U3842 ( .A(n4617), .B(n9000), .C(n7512), .Y(n2672) );
  OAI21X1 U3844 ( .A(n4617), .B(n9001), .C(n7587), .Y(n2671) );
  OAI21X1 U3846 ( .A(n4617), .B(n9002), .C(n7662), .Y(n2670) );
  OAI21X1 U3848 ( .A(n4617), .B(n9003), .C(n7740), .Y(n2669) );
  OAI21X1 U3850 ( .A(n4617), .B(n9004), .C(n7826), .Y(n2668) );
  OAI21X1 U3852 ( .A(n4617), .B(n9005), .C(n7913), .Y(n2667) );
  OAI21X1 U3854 ( .A(n4617), .B(n9006), .C(n8002), .Y(n2666) );
  OAI21X1 U3856 ( .A(n4617), .B(n9007), .C(n8093), .Y(n2665) );
  OAI21X1 U3858 ( .A(n4617), .B(n9008), .C(n8185), .Y(n2664) );
  OAI21X1 U3860 ( .A(n4617), .B(n9009), .C(n8275), .Y(n2663) );
  OAI21X1 U3862 ( .A(n4617), .B(n9010), .C(n8366), .Y(n2662) );
  OAI21X1 U3864 ( .A(n8242), .B(n8333), .C(n8501), .Y(n4617) );
  OAI21X1 U3865 ( .A(n4659), .B(n9011), .C(n8186), .Y(n2661) );
  OAI21X1 U3867 ( .A(n4659), .B(n9012), .C(n8003), .Y(n2660) );
  OAI21X1 U3869 ( .A(n4659), .B(n9013), .C(n7914), .Y(n2659) );
  OAI21X1 U3871 ( .A(n4659), .B(n9014), .C(n7827), .Y(n2658) );
  OAI21X1 U3873 ( .A(n4659), .B(n9015), .C(n7741), .Y(n2657) );
  OAI21X1 U3875 ( .A(n4659), .B(n9016), .C(n5786), .Y(n2656) );
  OAI21X1 U3877 ( .A(n4659), .B(n9017), .C(n8004), .Y(n2655) );
  OAI21X1 U3879 ( .A(n4659), .B(n9018), .C(n7915), .Y(n2654) );
  OAI21X1 U3881 ( .A(n4659), .B(n9019), .C(n7828), .Y(n2653) );
  OAI21X1 U3883 ( .A(n4659), .B(n9020), .C(n7742), .Y(n2652) );
  OAI21X1 U3885 ( .A(n4659), .B(n9021), .C(n7291), .Y(n2651) );
  OAI21X1 U3887 ( .A(n4659), .B(n9022), .C(n7218), .Y(n2650) );
  OAI21X1 U3889 ( .A(n4659), .B(n9023), .C(n7145), .Y(n2649) );
  OAI21X1 U3891 ( .A(n4659), .B(n9024), .C(n7663), .Y(n2648) );
  OAI21X1 U3893 ( .A(n4659), .B(n9025), .C(n7588), .Y(n2647) );
  OAI21X1 U3895 ( .A(n4659), .B(n9026), .C(n7513), .Y(n2646) );
  OAI21X1 U3897 ( .A(n4659), .B(n9027), .C(n7438), .Y(n2645) );
  OAI21X1 U3899 ( .A(n4659), .B(n9028), .C(n8367), .Y(n2644) );
  OAI21X1 U3901 ( .A(n4659), .B(n9029), .C(n8276), .Y(n2643) );
  OAI21X1 U3903 ( .A(n4659), .B(n9030), .C(n8187), .Y(n2642) );
  OAI21X1 U3905 ( .A(n4659), .B(n9031), .C(n8094), .Y(n2641) );
  OAI21X1 U3907 ( .A(n4659), .B(n9032), .C(n7364), .Y(n2640) );
  OAI21X1 U3909 ( .A(n4659), .B(n9033), .C(n7292), .Y(n2639) );
  OAI21X1 U3911 ( .A(n4659), .B(n9034), .C(n7219), .Y(n2638) );
  OAI21X1 U3913 ( .A(n4659), .B(n9035), .C(n7146), .Y(n2637) );
  OAI21X1 U3915 ( .A(n4659), .B(n9036), .C(n7664), .Y(n2636) );
  OAI21X1 U3917 ( .A(n4659), .B(n9037), .C(n7589), .Y(n2635) );
  OAI21X1 U3919 ( .A(n4659), .B(n9038), .C(n7514), .Y(n2634) );
  OAI21X1 U3921 ( .A(n4659), .B(n9039), .C(n7439), .Y(n2633) );
  OAI21X1 U3923 ( .A(n4659), .B(n9040), .C(n8368), .Y(n2632) );
  OAI21X1 U3925 ( .A(n4659), .B(n9041), .C(n8277), .Y(n2631) );
  OAI21X1 U3927 ( .A(n4659), .B(n9042), .C(n8188), .Y(n2630) );
  OAI21X1 U3929 ( .A(n4659), .B(n9043), .C(n8095), .Y(n2629) );
  OAI21X1 U3931 ( .A(n4659), .B(n9044), .C(n7365), .Y(n2628) );
  OAI21X1 U3933 ( .A(n4659), .B(n9045), .C(n7293), .Y(n2627) );
  OAI21X1 U3935 ( .A(n4659), .B(n9046), .C(n7220), .Y(n2626) );
  OAI21X1 U3937 ( .A(n4659), .B(n9047), .C(n7147), .Y(n2625) );
  OAI21X1 U3939 ( .A(n4659), .B(n9048), .C(n7665), .Y(n2624) );
  OAI21X1 U3941 ( .A(n4659), .B(n9049), .C(n7590), .Y(n2623) );
  OAI21X1 U3943 ( .A(n4659), .B(n9050), .C(n7515), .Y(n2622) );
  OAI21X1 U3945 ( .A(n4659), .B(n9051), .C(n7440), .Y(n2621) );
  OAI21X1 U3947 ( .A(n8243), .B(n8333), .C(n8500), .Y(n4659) );
  OAI21X1 U3948 ( .A(n4701), .B(n9052), .C(n8096), .Y(n2620) );
  OAI21X1 U3950 ( .A(n4701), .B(n9053), .C(n7916), .Y(n2619) );
  OAI21X1 U3952 ( .A(n4701), .B(n9054), .C(n8005), .Y(n2618) );
  OAI21X1 U3954 ( .A(n4701), .B(n9055), .C(n7743), .Y(n2617) );
  OAI21X1 U3956 ( .A(n4701), .B(n9056), .C(n7829), .Y(n2616) );
  OAI21X1 U3958 ( .A(n4701), .B(n9057), .C(n5785), .Y(n2615) );
  OAI21X1 U3960 ( .A(n4701), .B(n9058), .C(n7917), .Y(n2614) );
  OAI21X1 U3962 ( .A(n4701), .B(n9059), .C(n8006), .Y(n2613) );
  OAI21X1 U3964 ( .A(n4701), .B(n9060), .C(n7744), .Y(n2612) );
  OAI21X1 U3966 ( .A(n4701), .B(n9061), .C(n7830), .Y(n2611) );
  OAI21X1 U3968 ( .A(n4701), .B(n9062), .C(n7366), .Y(n2610) );
  OAI21X1 U3970 ( .A(n4701), .B(n9063), .C(n7148), .Y(n2609) );
  OAI21X1 U3972 ( .A(n4701), .B(n9064), .C(n7221), .Y(n2608) );
  OAI21X1 U3974 ( .A(n4701), .B(n9065), .C(n7591), .Y(n2607) );
  OAI21X1 U3976 ( .A(n4701), .B(n9066), .C(n7666), .Y(n2606) );
  OAI21X1 U3978 ( .A(n4701), .B(n9067), .C(n7441), .Y(n2605) );
  OAI21X1 U3980 ( .A(n4701), .B(n9068), .C(n7516), .Y(n2604) );
  OAI21X1 U3982 ( .A(n4701), .B(n9069), .C(n8278), .Y(n2603) );
  OAI21X1 U3984 ( .A(n4701), .B(n9070), .C(n8369), .Y(n2602) );
  OAI21X1 U3986 ( .A(n4701), .B(n9071), .C(n8097), .Y(n2601) );
  OAI21X1 U3988 ( .A(n4701), .B(n9072), .C(n8189), .Y(n2600) );
  OAI21X1 U3990 ( .A(n4701), .B(n9073), .C(n7294), .Y(n2599) );
  OAI21X1 U3992 ( .A(n4701), .B(n9074), .C(n7367), .Y(n2598) );
  OAI21X1 U3994 ( .A(n4701), .B(n9075), .C(n7149), .Y(n2597) );
  OAI21X1 U3996 ( .A(n4701), .B(n9076), .C(n7222), .Y(n2596) );
  OAI21X1 U3998 ( .A(n4701), .B(n9077), .C(n7592), .Y(n2595) );
  OAI21X1 U4000 ( .A(n4701), .B(n9078), .C(n7667), .Y(n2594) );
  OAI21X1 U4002 ( .A(n4701), .B(n9079), .C(n7442), .Y(n2593) );
  OAI21X1 U4004 ( .A(n4701), .B(n9080), .C(n7517), .Y(n2592) );
  OAI21X1 U4006 ( .A(n4701), .B(n9081), .C(n8279), .Y(n2591) );
  OAI21X1 U4008 ( .A(n4701), .B(n9082), .C(n8370), .Y(n2590) );
  OAI21X1 U4010 ( .A(n4701), .B(n9083), .C(n8098), .Y(n2589) );
  OAI21X1 U4012 ( .A(n4701), .B(n9084), .C(n8190), .Y(n2588) );
  OAI21X1 U4014 ( .A(n4701), .B(n9085), .C(n7295), .Y(n2587) );
  OAI21X1 U4016 ( .A(n4701), .B(n9086), .C(n7368), .Y(n2586) );
  OAI21X1 U4018 ( .A(n4701), .B(n9087), .C(n7150), .Y(n2585) );
  OAI21X1 U4020 ( .A(n4701), .B(n9088), .C(n7223), .Y(n2584) );
  OAI21X1 U4022 ( .A(n4701), .B(n9089), .C(n7593), .Y(n2583) );
  OAI21X1 U4024 ( .A(n4701), .B(n9090), .C(n7668), .Y(n2582) );
  OAI21X1 U4026 ( .A(n4701), .B(n9091), .C(n7443), .Y(n2581) );
  OAI21X1 U4028 ( .A(n4701), .B(n9092), .C(n7518), .Y(n2580) );
  OAI21X1 U4030 ( .A(n7970), .B(n8333), .C(n8500), .Y(n4701) );
  OAI21X1 U4031 ( .A(n4743), .B(n9093), .C(n8371), .Y(n2579) );
  OAI21X1 U4033 ( .A(n4743), .B(n9094), .C(n7831), .Y(n2578) );
  OAI21X1 U4035 ( .A(n4743), .B(n9095), .C(n7745), .Y(n2577) );
  OAI21X1 U4037 ( .A(n4743), .B(n9096), .C(n8007), .Y(n2576) );
  OAI21X1 U4039 ( .A(n4743), .B(n9097), .C(n7918), .Y(n2575) );
  OAI21X1 U4041 ( .A(n4743), .B(n9098), .C(n5784), .Y(n2574) );
  OAI21X1 U4043 ( .A(n4743), .B(n9099), .C(n7832), .Y(n2573) );
  OAI21X1 U4045 ( .A(n4743), .B(n9100), .C(n7746), .Y(n2572) );
  OAI21X1 U4047 ( .A(n4743), .B(n9101), .C(n8008), .Y(n2571) );
  OAI21X1 U4049 ( .A(n4743), .B(n9102), .C(n7919), .Y(n2570) );
  OAI21X1 U4051 ( .A(n4743), .B(n9103), .C(n7151), .Y(n2569) );
  OAI21X1 U4053 ( .A(n4743), .B(n9104), .C(n7369), .Y(n2568) );
  OAI21X1 U4055 ( .A(n4743), .B(n9105), .C(n7296), .Y(n2567) );
  OAI21X1 U4057 ( .A(n4743), .B(n9106), .C(n7519), .Y(n2566) );
  OAI21X1 U4059 ( .A(n4743), .B(n9107), .C(n7444), .Y(n2565) );
  OAI21X1 U4061 ( .A(n4743), .B(n9108), .C(n7669), .Y(n2564) );
  OAI21X1 U4063 ( .A(n4743), .B(n9109), .C(n7594), .Y(n2563) );
  OAI21X1 U4065 ( .A(n4743), .B(n9110), .C(n8191), .Y(n2562) );
  OAI21X1 U4067 ( .A(n4743), .B(n9111), .C(n8099), .Y(n2561) );
  OAI21X1 U4069 ( .A(n4743), .B(n9112), .C(n8372), .Y(n2560) );
  OAI21X1 U4071 ( .A(n4743), .B(n9113), .C(n8280), .Y(n2559) );
  OAI21X1 U4073 ( .A(n4743), .B(n9114), .C(n7224), .Y(n2558) );
  OAI21X1 U4075 ( .A(n4743), .B(n9115), .C(n7152), .Y(n2557) );
  OAI21X1 U4077 ( .A(n4743), .B(n9116), .C(n7370), .Y(n2556) );
  OAI21X1 U4079 ( .A(n4743), .B(n9117), .C(n7297), .Y(n2555) );
  OAI21X1 U4081 ( .A(n4743), .B(n9118), .C(n7520), .Y(n2554) );
  OAI21X1 U4083 ( .A(n4743), .B(n9119), .C(n7445), .Y(n2553) );
  OAI21X1 U4085 ( .A(n4743), .B(n9120), .C(n7670), .Y(n2552) );
  OAI21X1 U4087 ( .A(n4743), .B(n9121), .C(n7595), .Y(n2551) );
  OAI21X1 U4089 ( .A(n4743), .B(n9122), .C(n8192), .Y(n2550) );
  OAI21X1 U4091 ( .A(n4743), .B(n9123), .C(n8100), .Y(n2549) );
  OAI21X1 U4093 ( .A(n4743), .B(n9124), .C(n8373), .Y(n2548) );
  OAI21X1 U4095 ( .A(n4743), .B(n9125), .C(n8281), .Y(n2547) );
  OAI21X1 U4097 ( .A(n4743), .B(n9126), .C(n7225), .Y(n2546) );
  OAI21X1 U4099 ( .A(n4743), .B(n9127), .C(n7153), .Y(n2545) );
  OAI21X1 U4101 ( .A(n4743), .B(n9128), .C(n7371), .Y(n2544) );
  OAI21X1 U4103 ( .A(n4743), .B(n9129), .C(n7298), .Y(n2543) );
  OAI21X1 U4105 ( .A(n4743), .B(n9130), .C(n7521), .Y(n2542) );
  OAI21X1 U4107 ( .A(n4743), .B(n9131), .C(n7446), .Y(n2541) );
  OAI21X1 U4109 ( .A(n4743), .B(n9132), .C(n7671), .Y(n2540) );
  OAI21X1 U4111 ( .A(n4743), .B(n9133), .C(n7596), .Y(n2539) );
  OAI21X1 U4113 ( .A(n8061), .B(n8333), .C(n8500), .Y(n4743) );
  OAI21X1 U4114 ( .A(n4785), .B(n9134), .C(n8282), .Y(n2538) );
  OAI21X1 U4116 ( .A(n4785), .B(n9135), .C(n7747), .Y(n2537) );
  OAI21X1 U4118 ( .A(n4785), .B(n9136), .C(n7833), .Y(n2536) );
  OAI21X1 U4120 ( .A(n4785), .B(n9137), .C(n7920), .Y(n2535) );
  OAI21X1 U4122 ( .A(n4785), .B(n9138), .C(n8009), .Y(n2534) );
  OAI21X1 U4124 ( .A(n4785), .B(n9139), .C(n5783), .Y(n2533) );
  OAI21X1 U4126 ( .A(n4785), .B(n9140), .C(n7748), .Y(n2532) );
  OAI21X1 U4128 ( .A(n4785), .B(n9141), .C(n7834), .Y(n2531) );
  OAI21X1 U4130 ( .A(n4785), .B(n9142), .C(n7921), .Y(n2530) );
  OAI21X1 U4132 ( .A(n4785), .B(n9143), .C(n8010), .Y(n2529) );
  OAI21X1 U4134 ( .A(n4785), .B(n9144), .C(n7226), .Y(n2528) );
  OAI21X1 U4136 ( .A(n4785), .B(n9145), .C(n7299), .Y(n2527) );
  OAI21X1 U4138 ( .A(n4785), .B(n9146), .C(n7372), .Y(n2526) );
  OAI21X1 U4140 ( .A(n4785), .B(n9147), .C(n7447), .Y(n2525) );
  OAI21X1 U4142 ( .A(n4785), .B(n9148), .C(n7522), .Y(n2524) );
  OAI21X1 U4144 ( .A(n4785), .B(n9149), .C(n7597), .Y(n2523) );
  OAI21X1 U4146 ( .A(n4785), .B(n9150), .C(n7672), .Y(n2522) );
  OAI21X1 U4148 ( .A(n4785), .B(n9151), .C(n8101), .Y(n2521) );
  OAI21X1 U4150 ( .A(n4785), .B(n9152), .C(n8193), .Y(n2520) );
  OAI21X1 U4152 ( .A(n4785), .B(n9153), .C(n8283), .Y(n2519) );
  OAI21X1 U4154 ( .A(n4785), .B(n9154), .C(n8374), .Y(n2518) );
  OAI21X1 U4156 ( .A(n4785), .B(n9155), .C(n7154), .Y(n2517) );
  OAI21X1 U4158 ( .A(n4785), .B(n9156), .C(n7227), .Y(n2516) );
  OAI21X1 U4160 ( .A(n4785), .B(n9157), .C(n7300), .Y(n2515) );
  OAI21X1 U4162 ( .A(n4785), .B(n9158), .C(n7373), .Y(n2514) );
  OAI21X1 U4164 ( .A(n4785), .B(n9159), .C(n7448), .Y(n2513) );
  OAI21X1 U4166 ( .A(n4785), .B(n9160), .C(n7523), .Y(n2512) );
  OAI21X1 U4168 ( .A(n4785), .B(n9161), .C(n7598), .Y(n2511) );
  OAI21X1 U4170 ( .A(n4785), .B(n9162), .C(n7673), .Y(n2510) );
  OAI21X1 U4172 ( .A(n4785), .B(n9163), .C(n8102), .Y(n2509) );
  OAI21X1 U4174 ( .A(n4785), .B(n9164), .C(n8194), .Y(n2508) );
  OAI21X1 U4176 ( .A(n4785), .B(n9165), .C(n8284), .Y(n2507) );
  OAI21X1 U4178 ( .A(n4785), .B(n9166), .C(n8375), .Y(n2506) );
  OAI21X1 U4180 ( .A(n4785), .B(n9167), .C(n7155), .Y(n2505) );
  OAI21X1 U4182 ( .A(n4785), .B(n9168), .C(n7228), .Y(n2504) );
  OAI21X1 U4184 ( .A(n4785), .B(n9169), .C(n7301), .Y(n2503) );
  OAI21X1 U4186 ( .A(n4785), .B(n9170), .C(n7374), .Y(n2502) );
  OAI21X1 U4188 ( .A(n4785), .B(n9171), .C(n7449), .Y(n2501) );
  OAI21X1 U4190 ( .A(n4785), .B(n9172), .C(n7524), .Y(n2500) );
  OAI21X1 U4192 ( .A(n4785), .B(n9173), .C(n7599), .Y(n2499) );
  OAI21X1 U4194 ( .A(n4785), .B(n9174), .C(n7674), .Y(n2498) );
  OAI21X1 U4196 ( .A(n8152), .B(n8333), .C(n8500), .Y(n4785) );
  NAND3X1 U4197 ( .A(wr_ptr[4]), .B(n8518), .C(put), .Y(n4532) );
  OAI21X1 U4198 ( .A(n4827), .B(n9175), .C(n7229), .Y(n2497) );
  OAI21X1 U4200 ( .A(n4827), .B(n9176), .C(n7675), .Y(n2496) );
  OAI21X1 U4202 ( .A(n4827), .B(n9177), .C(n7600), .Y(n2495) );
  OAI21X1 U4204 ( .A(n4827), .B(n9178), .C(n7525), .Y(n2494) );
  OAI21X1 U4206 ( .A(n4827), .B(n9179), .C(n7450), .Y(n2493) );
  OAI21X1 U4208 ( .A(n4827), .B(n9180), .C(n5782), .Y(n2492) );
  OAI21X1 U4210 ( .A(n4827), .B(n9181), .C(n7676), .Y(n2491) );
  OAI21X1 U4212 ( .A(n4827), .B(n9182), .C(n7601), .Y(n2490) );
  OAI21X1 U4214 ( .A(n4827), .B(n9183), .C(n7526), .Y(n2489) );
  OAI21X1 U4216 ( .A(n4827), .B(n9184), .C(n7451), .Y(n2488) );
  OAI21X1 U4218 ( .A(n4827), .B(n9185), .C(n8285), .Y(n2487) );
  OAI21X1 U4220 ( .A(n4827), .B(n9186), .C(n8195), .Y(n2486) );
  OAI21X1 U4222 ( .A(n4827), .B(n9187), .C(n8103), .Y(n2485) );
  OAI21X1 U4224 ( .A(n4827), .B(n9188), .C(n8011), .Y(n2484) );
  OAI21X1 U4226 ( .A(n4827), .B(n9189), .C(n7922), .Y(n2483) );
  OAI21X1 U4228 ( .A(n4827), .B(n9190), .C(n7835), .Y(n2482) );
  OAI21X1 U4230 ( .A(n4827), .B(n9191), .C(n7749), .Y(n2481) );
  OAI21X1 U4232 ( .A(n4827), .B(n9192), .C(n7375), .Y(n2480) );
  OAI21X1 U4234 ( .A(n4827), .B(n9193), .C(n7302), .Y(n2479) );
  OAI21X1 U4236 ( .A(n4827), .B(n9194), .C(n7230), .Y(n2478) );
  OAI21X1 U4238 ( .A(n4827), .B(n9195), .C(n7156), .Y(n2477) );
  OAI21X1 U4240 ( .A(n4827), .B(n9196), .C(n8376), .Y(n2476) );
  OAI21X1 U4242 ( .A(n4827), .B(n9197), .C(n8286), .Y(n2475) );
  OAI21X1 U4244 ( .A(n4827), .B(n9198), .C(n8196), .Y(n2474) );
  OAI21X1 U4246 ( .A(n4827), .B(n9199), .C(n8104), .Y(n2473) );
  OAI21X1 U4248 ( .A(n4827), .B(n9200), .C(n8012), .Y(n2472) );
  OAI21X1 U4250 ( .A(n4827), .B(n9201), .C(n7923), .Y(n2471) );
  OAI21X1 U4252 ( .A(n4827), .B(n9202), .C(n7836), .Y(n2470) );
  OAI21X1 U4254 ( .A(n4827), .B(n9203), .C(n7750), .Y(n2469) );
  OAI21X1 U4256 ( .A(n4827), .B(n9204), .C(n7376), .Y(n2468) );
  OAI21X1 U4258 ( .A(n4827), .B(n9205), .C(n7303), .Y(n2467) );
  OAI21X1 U4260 ( .A(n4827), .B(n9206), .C(n7231), .Y(n2466) );
  OAI21X1 U4262 ( .A(n4827), .B(n9207), .C(n7157), .Y(n2465) );
  OAI21X1 U4264 ( .A(n4827), .B(n9208), .C(n8377), .Y(n2464) );
  OAI21X1 U4266 ( .A(n4827), .B(n9209), .C(n8287), .Y(n2463) );
  OAI21X1 U4268 ( .A(n4827), .B(n9210), .C(n8197), .Y(n2462) );
  OAI21X1 U4270 ( .A(n4827), .B(n9211), .C(n8105), .Y(n2461) );
  OAI21X1 U4272 ( .A(n4827), .B(n9212), .C(n8013), .Y(n2460) );
  OAI21X1 U4274 ( .A(n4827), .B(n9213), .C(n7924), .Y(n2459) );
  OAI21X1 U4276 ( .A(n4827), .B(n9214), .C(n7837), .Y(n2458) );
  OAI21X1 U4278 ( .A(n4827), .B(n9215), .C(n7751), .Y(n2457) );
  OAI21X1 U4280 ( .A(n8153), .B(n8334), .C(n8500), .Y(n4827) );
  OAI21X1 U4281 ( .A(n4870), .B(n9216), .C(n7158), .Y(n2456) );
  OAI21X1 U4283 ( .A(n4870), .B(n9217), .C(n7602), .Y(n2455) );
  OAI21X1 U4285 ( .A(n4870), .B(n9218), .C(n7677), .Y(n2454) );
  OAI21X1 U4287 ( .A(n4870), .B(n9219), .C(n7452), .Y(n2453) );
  OAI21X1 U4289 ( .A(n4870), .B(n9220), .C(n7527), .Y(n2452) );
  OAI21X1 U4291 ( .A(n4870), .B(n9221), .C(n5781), .Y(n2451) );
  OAI21X1 U4293 ( .A(n4870), .B(n9222), .C(n7603), .Y(n2450) );
  OAI21X1 U4295 ( .A(n4870), .B(n9223), .C(n7678), .Y(n2449) );
  OAI21X1 U4297 ( .A(n4870), .B(n9224), .C(n7453), .Y(n2448) );
  OAI21X1 U4299 ( .A(n4870), .B(n9225), .C(n7528), .Y(n2447) );
  OAI21X1 U4301 ( .A(n4870), .B(n9226), .C(n8378), .Y(n2446) );
  OAI21X1 U4303 ( .A(n4870), .B(n9227), .C(n8106), .Y(n2445) );
  OAI21X1 U4305 ( .A(n4870), .B(n9228), .C(n8198), .Y(n2444) );
  OAI21X1 U4307 ( .A(n4870), .B(n9229), .C(n7925), .Y(n2443) );
  OAI21X1 U4309 ( .A(n4870), .B(n9230), .C(n8014), .Y(n2442) );
  OAI21X1 U4311 ( .A(n4870), .B(n9231), .C(n7752), .Y(n2441) );
  OAI21X1 U4313 ( .A(n4870), .B(n9232), .C(n7838), .Y(n2440) );
  OAI21X1 U4315 ( .A(n4870), .B(n9233), .C(n7304), .Y(n2439) );
  OAI21X1 U4317 ( .A(n4870), .B(n9234), .C(n7377), .Y(n2438) );
  OAI21X1 U4319 ( .A(n4870), .B(n9235), .C(n7159), .Y(n2437) );
  OAI21X1 U4321 ( .A(n4870), .B(n9236), .C(n7232), .Y(n2436) );
  OAI21X1 U4323 ( .A(n4870), .B(n9237), .C(n8288), .Y(n2435) );
  OAI21X1 U4325 ( .A(n4870), .B(n9238), .C(n8379), .Y(n2434) );
  OAI21X1 U4327 ( .A(n4870), .B(n9239), .C(n8107), .Y(n2433) );
  OAI21X1 U4329 ( .A(n4870), .B(n9240), .C(n8199), .Y(n2432) );
  OAI21X1 U4331 ( .A(n4870), .B(n9241), .C(n7926), .Y(n2431) );
  OAI21X1 U4333 ( .A(n4870), .B(n9242), .C(n8015), .Y(n2430) );
  OAI21X1 U4335 ( .A(n4870), .B(n9243), .C(n7753), .Y(n2429) );
  OAI21X1 U4337 ( .A(n4870), .B(n9244), .C(n7839), .Y(n2428) );
  OAI21X1 U4339 ( .A(n4870), .B(n9245), .C(n7305), .Y(n2427) );
  OAI21X1 U4341 ( .A(n4870), .B(n9246), .C(n7378), .Y(n2426) );
  OAI21X1 U4343 ( .A(n4870), .B(n9247), .C(n7160), .Y(n2425) );
  OAI21X1 U4345 ( .A(n4870), .B(n9248), .C(n7233), .Y(n2424) );
  OAI21X1 U4347 ( .A(n4870), .B(n9249), .C(n8289), .Y(n2423) );
  OAI21X1 U4349 ( .A(n4870), .B(n9250), .C(n8380), .Y(n2422) );
  OAI21X1 U4351 ( .A(n4870), .B(n9251), .C(n8108), .Y(n2421) );
  OAI21X1 U4353 ( .A(n4870), .B(n9252), .C(n8200), .Y(n2420) );
  OAI21X1 U4355 ( .A(n4870), .B(n9253), .C(n7927), .Y(n2419) );
  OAI21X1 U4357 ( .A(n4870), .B(n9254), .C(n8016), .Y(n2418) );
  OAI21X1 U4359 ( .A(n4870), .B(n9255), .C(n7754), .Y(n2417) );
  OAI21X1 U4361 ( .A(n4870), .B(n9256), .C(n7840), .Y(n2416) );
  OAI21X1 U4363 ( .A(n8060), .B(n8334), .C(n8500), .Y(n4870) );
  OAI21X1 U4364 ( .A(n4912), .B(n9257), .C(n7379), .Y(n2415) );
  OAI21X1 U4366 ( .A(n4912), .B(n9258), .C(n7529), .Y(n2414) );
  OAI21X1 U4368 ( .A(n4912), .B(n9259), .C(n7454), .Y(n2413) );
  OAI21X1 U4370 ( .A(n4912), .B(n9260), .C(n7679), .Y(n2412) );
  OAI21X1 U4372 ( .A(n4912), .B(n9261), .C(n7604), .Y(n2411) );
  OAI21X1 U4374 ( .A(n4912), .B(n9262), .C(n5780), .Y(n2410) );
  OAI21X1 U4376 ( .A(n4912), .B(n9263), .C(n7530), .Y(n2409) );
  OAI21X1 U4378 ( .A(n4912), .B(n9264), .C(n7455), .Y(n2408) );
  OAI21X1 U4380 ( .A(n4912), .B(n9265), .C(n7680), .Y(n2407) );
  OAI21X1 U4382 ( .A(n4912), .B(n9266), .C(n7605), .Y(n2406) );
  OAI21X1 U4384 ( .A(n4912), .B(n9267), .C(n8109), .Y(n2405) );
  OAI21X1 U4386 ( .A(n4912), .B(n9268), .C(n8381), .Y(n2404) );
  OAI21X1 U4388 ( .A(n4912), .B(n9269), .C(n8290), .Y(n2403) );
  OAI21X1 U4390 ( .A(n4912), .B(n9270), .C(n7841), .Y(n2402) );
  OAI21X1 U4392 ( .A(n4912), .B(n9271), .C(n7755), .Y(n2401) );
  OAI21X1 U4394 ( .A(n4912), .B(n9272), .C(n8017), .Y(n2400) );
  OAI21X1 U4396 ( .A(n4912), .B(n9273), .C(n7928), .Y(n2399) );
  OAI21X1 U4398 ( .A(n4912), .B(n9274), .C(n7234), .Y(n2398) );
  OAI21X1 U4400 ( .A(n4912), .B(n9275), .C(n7161), .Y(n2397) );
  OAI21X1 U4402 ( .A(n4912), .B(n9276), .C(n7380), .Y(n2396) );
  OAI21X1 U4404 ( .A(n4912), .B(n9277), .C(n7306), .Y(n2395) );
  OAI21X1 U4406 ( .A(n4912), .B(n9278), .C(n8201), .Y(n2394) );
  OAI21X1 U4408 ( .A(n4912), .B(n9279), .C(n8110), .Y(n2393) );
  OAI21X1 U4410 ( .A(n4912), .B(n9280), .C(n8382), .Y(n2392) );
  OAI21X1 U4412 ( .A(n4912), .B(n9281), .C(n8291), .Y(n2391) );
  OAI21X1 U4414 ( .A(n4912), .B(n9282), .C(n7842), .Y(n2390) );
  OAI21X1 U4416 ( .A(n4912), .B(n9283), .C(n7756), .Y(n2389) );
  OAI21X1 U4418 ( .A(n4912), .B(n9284), .C(n8018), .Y(n2388) );
  OAI21X1 U4420 ( .A(n4912), .B(n9285), .C(n7929), .Y(n2387) );
  OAI21X1 U4422 ( .A(n4912), .B(n9286), .C(n7235), .Y(n2386) );
  OAI21X1 U4424 ( .A(n4912), .B(n9287), .C(n7162), .Y(n2385) );
  OAI21X1 U4426 ( .A(n4912), .B(n9288), .C(n7381), .Y(n2384) );
  OAI21X1 U4428 ( .A(n4912), .B(n9289), .C(n7307), .Y(n2383) );
  OAI21X1 U4430 ( .A(n4912), .B(n9290), .C(n8202), .Y(n2382) );
  OAI21X1 U4432 ( .A(n4912), .B(n9291), .C(n8111), .Y(n2381) );
  OAI21X1 U4434 ( .A(n4912), .B(n9292), .C(n8383), .Y(n2380) );
  OAI21X1 U4436 ( .A(n4912), .B(n9293), .C(n8292), .Y(n2379) );
  OAI21X1 U4438 ( .A(n4912), .B(n9294), .C(n7843), .Y(n2378) );
  OAI21X1 U4440 ( .A(n4912), .B(n9295), .C(n7757), .Y(n2377) );
  OAI21X1 U4442 ( .A(n4912), .B(n9296), .C(n8019), .Y(n2376) );
  OAI21X1 U4444 ( .A(n4912), .B(n9297), .C(n7930), .Y(n2375) );
  OAI21X1 U4446 ( .A(n7969), .B(n8334), .C(n8500), .Y(n4912) );
  OAI21X1 U4447 ( .A(n4954), .B(n9298), .C(n7308), .Y(n2374) );
  OAI21X1 U4449 ( .A(n4954), .B(n9299), .C(n7456), .Y(n2373) );
  OAI21X1 U4451 ( .A(n4954), .B(n9300), .C(n7531), .Y(n2372) );
  OAI21X1 U4453 ( .A(n4954), .B(n9301), .C(n7606), .Y(n2371) );
  OAI21X1 U4455 ( .A(n4954), .B(n9302), .C(n7681), .Y(n2370) );
  OAI21X1 U4457 ( .A(n4954), .B(n9303), .C(n5779), .Y(n2369) );
  OAI21X1 U4459 ( .A(n4954), .B(n9304), .C(n7457), .Y(n2368) );
  OAI21X1 U4461 ( .A(n4954), .B(n9305), .C(n7532), .Y(n2367) );
  OAI21X1 U4463 ( .A(n4954), .B(n9306), .C(n7607), .Y(n2366) );
  OAI21X1 U4465 ( .A(n4954), .B(n9307), .C(n7682), .Y(n2365) );
  OAI21X1 U4467 ( .A(n4954), .B(n9308), .C(n8203), .Y(n2364) );
  OAI21X1 U4469 ( .A(n4954), .B(n9309), .C(n8293), .Y(n2363) );
  OAI21X1 U4471 ( .A(n4954), .B(n9310), .C(n8384), .Y(n2362) );
  OAI21X1 U4473 ( .A(n4954), .B(n9311), .C(n7758), .Y(n2361) );
  OAI21X1 U4475 ( .A(n4954), .B(n9312), .C(n7844), .Y(n2360) );
  OAI21X1 U4477 ( .A(n4954), .B(n9313), .C(n7931), .Y(n2359) );
  OAI21X1 U4479 ( .A(n4954), .B(n9314), .C(n8020), .Y(n2358) );
  OAI21X1 U4481 ( .A(n4954), .B(n9315), .C(n7163), .Y(n2357) );
  OAI21X1 U4483 ( .A(n4954), .B(n9316), .C(n7236), .Y(n2356) );
  OAI21X1 U4485 ( .A(n4954), .B(n9317), .C(n7309), .Y(n2355) );
  OAI21X1 U4487 ( .A(n4954), .B(n9318), .C(n7382), .Y(n2354) );
  OAI21X1 U4489 ( .A(n4954), .B(n9319), .C(n8112), .Y(n2353) );
  OAI21X1 U4491 ( .A(n4954), .B(n9320), .C(n8204), .Y(n2352) );
  OAI21X1 U4493 ( .A(n4954), .B(n9321), .C(n8294), .Y(n2351) );
  OAI21X1 U4495 ( .A(n4954), .B(n9322), .C(n8385), .Y(n2350) );
  OAI21X1 U4497 ( .A(n4954), .B(n9323), .C(n7759), .Y(n2349) );
  OAI21X1 U4499 ( .A(n4954), .B(n9324), .C(n7845), .Y(n2348) );
  OAI21X1 U4501 ( .A(n4954), .B(n9325), .C(n7932), .Y(n2347) );
  OAI21X1 U4503 ( .A(n4954), .B(n9326), .C(n8021), .Y(n2346) );
  OAI21X1 U4505 ( .A(n4954), .B(n9327), .C(n7164), .Y(n2345) );
  OAI21X1 U4507 ( .A(n4954), .B(n9328), .C(n7237), .Y(n2344) );
  OAI21X1 U4509 ( .A(n4954), .B(n9329), .C(n7310), .Y(n2343) );
  OAI21X1 U4511 ( .A(n4954), .B(n9330), .C(n7383), .Y(n2342) );
  OAI21X1 U4513 ( .A(n4954), .B(n9331), .C(n8113), .Y(n2341) );
  OAI21X1 U4515 ( .A(n4954), .B(n9332), .C(n8205), .Y(n2340) );
  OAI21X1 U4517 ( .A(n4954), .B(n9333), .C(n8295), .Y(n2339) );
  OAI21X1 U4519 ( .A(n4954), .B(n9334), .C(n8386), .Y(n2338) );
  OAI21X1 U4521 ( .A(n4954), .B(n9335), .C(n7760), .Y(n2337) );
  OAI21X1 U4523 ( .A(n4954), .B(n9336), .C(n7846), .Y(n2336) );
  OAI21X1 U4525 ( .A(n4954), .B(n9337), .C(n7933), .Y(n2335) );
  OAI21X1 U4527 ( .A(n4954), .B(n9338), .C(n8022), .Y(n2334) );
  OAI21X1 U4529 ( .A(n8242), .B(n8334), .C(n8500), .Y(n4954) );
  OAI21X1 U4530 ( .A(n4996), .B(n9339), .C(n7533), .Y(n2333) );
  OAI21X1 U4532 ( .A(n4996), .B(n9340), .C(n7384), .Y(n2332) );
  OAI21X1 U4534 ( .A(n4996), .B(n9341), .C(n7311), .Y(n2331) );
  OAI21X1 U4536 ( .A(n4996), .B(n9342), .C(n7238), .Y(n2330) );
  OAI21X1 U4538 ( .A(n4996), .B(n9343), .C(n7165), .Y(n2329) );
  OAI21X1 U4540 ( .A(n4996), .B(n9344), .C(n5778), .Y(n2328) );
  OAI21X1 U4542 ( .A(n4996), .B(n9345), .C(n7385), .Y(n2327) );
  OAI21X1 U4544 ( .A(n4996), .B(n9346), .C(n7312), .Y(n2326) );
  OAI21X1 U4546 ( .A(n4996), .B(n9347), .C(n7239), .Y(n2325) );
  OAI21X1 U4548 ( .A(n4996), .B(n9348), .C(n7166), .Y(n2324) );
  OAI21X1 U4550 ( .A(n4996), .B(n9349), .C(n7934), .Y(n2323) );
  OAI21X1 U4552 ( .A(n4996), .B(n9350), .C(n7847), .Y(n2322) );
  OAI21X1 U4554 ( .A(n4996), .B(n9351), .C(n7761), .Y(n2321) );
  OAI21X1 U4556 ( .A(n4996), .B(n9352), .C(n8387), .Y(n2320) );
  OAI21X1 U4558 ( .A(n4996), .B(n9353), .C(n8296), .Y(n2319) );
  OAI21X1 U4560 ( .A(n4996), .B(n9354), .C(n8206), .Y(n2318) );
  OAI21X1 U4562 ( .A(n4996), .B(n9355), .C(n8114), .Y(n2317) );
  OAI21X1 U4564 ( .A(n4996), .B(n9356), .C(n7683), .Y(n2316) );
  OAI21X1 U4566 ( .A(n4996), .B(n9357), .C(n7608), .Y(n2315) );
  OAI21X1 U4568 ( .A(n4996), .B(n9358), .C(n7534), .Y(n2314) );
  OAI21X1 U4570 ( .A(n4996), .B(n9359), .C(n7458), .Y(n2313) );
  OAI21X1 U4572 ( .A(n4996), .B(n9360), .C(n8023), .Y(n2312) );
  OAI21X1 U4574 ( .A(n4996), .B(n9361), .C(n7935), .Y(n2311) );
  OAI21X1 U4576 ( .A(n4996), .B(n9362), .C(n7848), .Y(n2310) );
  OAI21X1 U4578 ( .A(n4996), .B(n9363), .C(n7762), .Y(n2309) );
  OAI21X1 U4580 ( .A(n4996), .B(n9364), .C(n8388), .Y(n2308) );
  OAI21X1 U4582 ( .A(n4996), .B(n9365), .C(n8297), .Y(n2307) );
  OAI21X1 U4584 ( .A(n4996), .B(n9366), .C(n8207), .Y(n2306) );
  OAI21X1 U4586 ( .A(n4996), .B(n9367), .C(n8115), .Y(n2305) );
  OAI21X1 U4588 ( .A(n4996), .B(n9368), .C(n7684), .Y(n2304) );
  OAI21X1 U4590 ( .A(n4996), .B(n9369), .C(n7609), .Y(n2303) );
  OAI21X1 U4592 ( .A(n4996), .B(n9370), .C(n7535), .Y(n2302) );
  OAI21X1 U4594 ( .A(n4996), .B(n9371), .C(n7459), .Y(n2301) );
  OAI21X1 U4596 ( .A(n4996), .B(n9372), .C(n8024), .Y(n2300) );
  OAI21X1 U4598 ( .A(n4996), .B(n9373), .C(n7936), .Y(n2299) );
  OAI21X1 U4600 ( .A(n4996), .B(n9374), .C(n7849), .Y(n2298) );
  OAI21X1 U4602 ( .A(n4996), .B(n9375), .C(n7763), .Y(n2297) );
  OAI21X1 U4604 ( .A(n4996), .B(n9376), .C(n8389), .Y(n2296) );
  OAI21X1 U4606 ( .A(n4996), .B(n9377), .C(n8298), .Y(n2295) );
  OAI21X1 U4608 ( .A(n4996), .B(n9378), .C(n8208), .Y(n2294) );
  OAI21X1 U4610 ( .A(n4996), .B(n9379), .C(n8116), .Y(n2293) );
  OAI21X1 U4612 ( .A(n8243), .B(n8334), .C(n8500), .Y(n4996) );
  OAI21X1 U4613 ( .A(n5038), .B(n9380), .C(n7460), .Y(n2292) );
  OAI21X1 U4615 ( .A(n5038), .B(n9381), .C(n7313), .Y(n2291) );
  OAI21X1 U4617 ( .A(n5038), .B(n9382), .C(n7386), .Y(n2290) );
  OAI21X1 U4619 ( .A(n5038), .B(n9383), .C(n7167), .Y(n2289) );
  OAI21X1 U4621 ( .A(n5038), .B(n9384), .C(n7240), .Y(n2288) );
  OAI21X1 U4623 ( .A(n5038), .B(n9385), .C(n5777), .Y(n2287) );
  OAI21X1 U4625 ( .A(n5038), .B(n9386), .C(n7314), .Y(n2286) );
  OAI21X1 U4627 ( .A(n5038), .B(n9387), .C(n7387), .Y(n2285) );
  OAI21X1 U4629 ( .A(n5038), .B(n9388), .C(n7168), .Y(n2284) );
  OAI21X1 U4631 ( .A(n5038), .B(n9389), .C(n7241), .Y(n2283) );
  OAI21X1 U4633 ( .A(n5038), .B(n9390), .C(n8025), .Y(n2282) );
  OAI21X1 U4635 ( .A(n5038), .B(n9391), .C(n7764), .Y(n2281) );
  OAI21X1 U4637 ( .A(n5038), .B(n9392), .C(n7850), .Y(n2280) );
  OAI21X1 U4639 ( .A(n5038), .B(n9393), .C(n8299), .Y(n2279) );
  OAI21X1 U4641 ( .A(n5038), .B(n9394), .C(n8390), .Y(n2278) );
  OAI21X1 U4643 ( .A(n5038), .B(n9395), .C(n8117), .Y(n2277) );
  OAI21X1 U4645 ( .A(n5038), .B(n9396), .C(n8209), .Y(n2276) );
  OAI21X1 U4647 ( .A(n5038), .B(n9397), .C(n7610), .Y(n2275) );
  OAI21X1 U4649 ( .A(n5038), .B(n9398), .C(n7685), .Y(n2274) );
  OAI21X1 U4651 ( .A(n5038), .B(n9399), .C(n7461), .Y(n2273) );
  OAI21X1 U4653 ( .A(n5038), .B(n9400), .C(n7536), .Y(n2272) );
  OAI21X1 U4655 ( .A(n5038), .B(n9401), .C(n7937), .Y(n2271) );
  OAI21X1 U4657 ( .A(n5038), .B(n9402), .C(n8026), .Y(n2270) );
  OAI21X1 U4659 ( .A(n5038), .B(n9403), .C(n7765), .Y(n2269) );
  OAI21X1 U4661 ( .A(n5038), .B(n9404), .C(n7851), .Y(n2268) );
  OAI21X1 U4663 ( .A(n5038), .B(n9405), .C(n8300), .Y(n2267) );
  OAI21X1 U4665 ( .A(n5038), .B(n9406), .C(n8391), .Y(n2266) );
  OAI21X1 U4667 ( .A(n5038), .B(n9407), .C(n8118), .Y(n2265) );
  OAI21X1 U4669 ( .A(n5038), .B(n9408), .C(n8210), .Y(n2264) );
  OAI21X1 U4671 ( .A(n5038), .B(n9409), .C(n7611), .Y(n2263) );
  OAI21X1 U4673 ( .A(n5038), .B(n9410), .C(n7686), .Y(n2262) );
  OAI21X1 U4675 ( .A(n5038), .B(n9411), .C(n7462), .Y(n2261) );
  OAI21X1 U4677 ( .A(n5038), .B(n9412), .C(n7537), .Y(n2260) );
  OAI21X1 U4679 ( .A(n5038), .B(n9413), .C(n7938), .Y(n2259) );
  OAI21X1 U4681 ( .A(n5038), .B(n9414), .C(n8027), .Y(n2258) );
  OAI21X1 U4683 ( .A(n5038), .B(n9415), .C(n7766), .Y(n2257) );
  OAI21X1 U4685 ( .A(n5038), .B(n9416), .C(n7852), .Y(n2256) );
  OAI21X1 U4687 ( .A(n5038), .B(n9417), .C(n8301), .Y(n2255) );
  OAI21X1 U4689 ( .A(n5038), .B(n9418), .C(n8392), .Y(n2254) );
  OAI21X1 U4691 ( .A(n5038), .B(n9419), .C(n8119), .Y(n2253) );
  OAI21X1 U4693 ( .A(n5038), .B(n9420), .C(n8211), .Y(n2252) );
  OAI21X1 U4695 ( .A(n7970), .B(n8334), .C(n8500), .Y(n5038) );
  OAI21X1 U4696 ( .A(n5080), .B(n9421), .C(n7687), .Y(n2251) );
  OAI21X1 U4698 ( .A(n5080), .B(n9422), .C(n7242), .Y(n2250) );
  OAI21X1 U4700 ( .A(n5080), .B(n9423), .C(n7169), .Y(n2249) );
  OAI21X1 U4702 ( .A(n5080), .B(n9424), .C(n7388), .Y(n2248) );
  OAI21X1 U4704 ( .A(n5080), .B(n9425), .C(n7315), .Y(n2247) );
  OAI21X1 U4706 ( .A(n5080), .B(n9426), .C(n5776), .Y(n2246) );
  OAI21X1 U4708 ( .A(n5080), .B(n9427), .C(n7243), .Y(n2245) );
  OAI21X1 U4710 ( .A(n5080), .B(n9428), .C(n7170), .Y(n2244) );
  OAI21X1 U4712 ( .A(n5080), .B(n9429), .C(n7389), .Y(n2243) );
  OAI21X1 U4714 ( .A(n5080), .B(n9430), .C(n7316), .Y(n2242) );
  OAI21X1 U4716 ( .A(n5080), .B(n9431), .C(n7767), .Y(n2241) );
  OAI21X1 U4718 ( .A(n5080), .B(n9432), .C(n8028), .Y(n2240) );
  OAI21X1 U4720 ( .A(n5080), .B(n9433), .C(n7939), .Y(n2239) );
  OAI21X1 U4722 ( .A(n5080), .B(n9434), .C(n8212), .Y(n2238) );
  OAI21X1 U4724 ( .A(n5080), .B(n9435), .C(n8120), .Y(n2237) );
  OAI21X1 U4726 ( .A(n5080), .B(n9436), .C(n8393), .Y(n2236) );
  OAI21X1 U4728 ( .A(n5080), .B(n9437), .C(n8302), .Y(n2235) );
  OAI21X1 U4730 ( .A(n5080), .B(n9438), .C(n7538), .Y(n2234) );
  OAI21X1 U4732 ( .A(n5080), .B(n9439), .C(n7463), .Y(n2233) );
  OAI21X1 U4734 ( .A(n5080), .B(n9440), .C(n7688), .Y(n2232) );
  OAI21X1 U4736 ( .A(n5080), .B(n9441), .C(n7612), .Y(n2231) );
  OAI21X1 U4738 ( .A(n5080), .B(n9442), .C(n7853), .Y(n2230) );
  OAI21X1 U4740 ( .A(n5080), .B(n9443), .C(n7768), .Y(n2229) );
  OAI21X1 U4742 ( .A(n5080), .B(n9444), .C(n8029), .Y(n2228) );
  OAI21X1 U4744 ( .A(n5080), .B(n9445), .C(n7940), .Y(n2227) );
  OAI21X1 U4746 ( .A(n5080), .B(n9446), .C(n8213), .Y(n2226) );
  OAI21X1 U4748 ( .A(n5080), .B(n9447), .C(n8121), .Y(n2225) );
  OAI21X1 U4750 ( .A(n5080), .B(n9448), .C(n8394), .Y(n2224) );
  OAI21X1 U4752 ( .A(n5080), .B(n9449), .C(n8303), .Y(n2223) );
  OAI21X1 U4754 ( .A(n5080), .B(n9450), .C(n7539), .Y(n2222) );
  OAI21X1 U4756 ( .A(n5080), .B(n9451), .C(n7464), .Y(n2221) );
  OAI21X1 U4758 ( .A(n5080), .B(n9452), .C(n7689), .Y(n2220) );
  OAI21X1 U4760 ( .A(n5080), .B(n9453), .C(n7613), .Y(n2219) );
  OAI21X1 U4762 ( .A(n5080), .B(n9454), .C(n7854), .Y(n2218) );
  OAI21X1 U4764 ( .A(n5080), .B(n9455), .C(n7769), .Y(n2217) );
  OAI21X1 U4766 ( .A(n5080), .B(n9456), .C(n8030), .Y(n2216) );
  OAI21X1 U4768 ( .A(n5080), .B(n9457), .C(n7941), .Y(n2215) );
  OAI21X1 U4770 ( .A(n5080), .B(n9458), .C(n8214), .Y(n2214) );
  OAI21X1 U4772 ( .A(n5080), .B(n9459), .C(n8122), .Y(n2213) );
  OAI21X1 U4774 ( .A(n5080), .B(n9460), .C(n8395), .Y(n2212) );
  OAI21X1 U4776 ( .A(n5080), .B(n9461), .C(n8304), .Y(n2211) );
  OAI21X1 U4778 ( .A(n8061), .B(n8334), .C(n8500), .Y(n5080) );
  OAI21X1 U4779 ( .A(n5122), .B(n9462), .C(n7614), .Y(n2210) );
  OAI21X1 U4781 ( .A(n5122), .B(n9463), .C(n7171), .Y(n2209) );
  OAI21X1 U4783 ( .A(n5122), .B(n9464), .C(n7244), .Y(n2208) );
  OAI21X1 U4785 ( .A(n5122), .B(n9465), .C(n7317), .Y(n2207) );
  OAI21X1 U4787 ( .A(n5122), .B(n9466), .C(n7390), .Y(n2206) );
  OAI21X1 U4789 ( .A(n5122), .B(n9467), .C(n5775), .Y(n2205) );
  OAI21X1 U4791 ( .A(n5122), .B(n9468), .C(n7172), .Y(n2204) );
  OAI21X1 U4793 ( .A(n5122), .B(n9469), .C(n7245), .Y(n2203) );
  OAI21X1 U4795 ( .A(n5122), .B(n9470), .C(n7318), .Y(n2202) );
  OAI21X1 U4797 ( .A(n5122), .B(n9471), .C(n7391), .Y(n2201) );
  OAI21X1 U4799 ( .A(n5122), .B(n9472), .C(n7855), .Y(n2200) );
  OAI21X1 U4801 ( .A(n5122), .B(n9473), .C(n7942), .Y(n2199) );
  OAI21X1 U4803 ( .A(n5122), .B(n9474), .C(n8031), .Y(n2198) );
  OAI21X1 U4805 ( .A(n5122), .B(n9475), .C(n8123), .Y(n2197) );
  OAI21X1 U4807 ( .A(n5122), .B(n9476), .C(n8215), .Y(n2196) );
  OAI21X1 U4809 ( .A(n5122), .B(n9477), .C(n8305), .Y(n2195) );
  OAI21X1 U4811 ( .A(n5122), .B(n9478), .C(n8396), .Y(n2194) );
  OAI21X1 U4813 ( .A(n5122), .B(n9479), .C(n7465), .Y(n2193) );
  OAI21X1 U4815 ( .A(n5122), .B(n9480), .C(n7540), .Y(n2192) );
  OAI21X1 U4817 ( .A(n5122), .B(n9481), .C(n7615), .Y(n2191) );
  OAI21X1 U4819 ( .A(n5122), .B(n9482), .C(n7690), .Y(n2190) );
  OAI21X1 U4821 ( .A(n5122), .B(n9483), .C(n7770), .Y(n2189) );
  OAI21X1 U4823 ( .A(n5122), .B(n9484), .C(n7856), .Y(n2188) );
  OAI21X1 U4825 ( .A(n5122), .B(n9485), .C(n7943), .Y(n2187) );
  OAI21X1 U4827 ( .A(n5122), .B(n9486), .C(n8032), .Y(n2186) );
  OAI21X1 U4829 ( .A(n5122), .B(n9487), .C(n8124), .Y(n2185) );
  OAI21X1 U4831 ( .A(n5122), .B(n9488), .C(n8216), .Y(n2184) );
  OAI21X1 U4833 ( .A(n5122), .B(n9489), .C(n8306), .Y(n2183) );
  OAI21X1 U4835 ( .A(n5122), .B(n9490), .C(n8397), .Y(n2182) );
  OAI21X1 U4837 ( .A(n5122), .B(n9491), .C(n7466), .Y(n2181) );
  OAI21X1 U4839 ( .A(n5122), .B(n9492), .C(n7541), .Y(n2180) );
  OAI21X1 U4841 ( .A(n5122), .B(n9493), .C(n7616), .Y(n2179) );
  OAI21X1 U4843 ( .A(n5122), .B(n9494), .C(n7691), .Y(n2178) );
  OAI21X1 U4845 ( .A(n5122), .B(n9495), .C(n7771), .Y(n2177) );
  OAI21X1 U4847 ( .A(n5122), .B(n9496), .C(n7857), .Y(n2176) );
  OAI21X1 U4849 ( .A(n5122), .B(n9497), .C(n7944), .Y(n2175) );
  OAI21X1 U4851 ( .A(n5122), .B(n9498), .C(n8033), .Y(n2174) );
  OAI21X1 U4853 ( .A(n5122), .B(n9499), .C(n8125), .Y(n2173) );
  OAI21X1 U4855 ( .A(n5122), .B(n9500), .C(n8217), .Y(n2172) );
  OAI21X1 U4857 ( .A(n5122), .B(n9501), .C(n8307), .Y(n2171) );
  OAI21X1 U4859 ( .A(n5122), .B(n9502), .C(n8398), .Y(n2170) );
  OAI21X1 U4861 ( .A(n8152), .B(n8334), .C(n8500), .Y(n5122) );
  NAND3X1 U4862 ( .A(wr_ptr[3]), .B(n8515), .C(put), .Y(n4869) );
  OAI21X1 U4863 ( .A(n5164), .B(n9503), .C(n7246), .Y(n2169) );
  OAI21X1 U4865 ( .A(n5164), .B(n9504), .C(n7692), .Y(n2168) );
  OAI21X1 U4867 ( .A(n5164), .B(n9505), .C(n7617), .Y(n2167) );
  OAI21X1 U4869 ( .A(n5164), .B(n9506), .C(n7542), .Y(n2166) );
  OAI21X1 U4871 ( .A(n5164), .B(n9507), .C(n7467), .Y(n2165) );
  OAI21X1 U4873 ( .A(n5164), .B(n9508), .C(n5774), .Y(n2164) );
  OAI21X1 U4875 ( .A(n5164), .B(n9509), .C(n7693), .Y(n2163) );
  OAI21X1 U4877 ( .A(n5164), .B(n9510), .C(n7618), .Y(n2162) );
  OAI21X1 U4879 ( .A(n5164), .B(n9511), .C(n7543), .Y(n2161) );
  OAI21X1 U4881 ( .A(n5164), .B(n9512), .C(n7468), .Y(n2160) );
  OAI21X1 U4883 ( .A(n5164), .B(n9513), .C(n8308), .Y(n2159) );
  OAI21X1 U4885 ( .A(n5164), .B(n9514), .C(n8218), .Y(n2158) );
  OAI21X1 U4887 ( .A(n5164), .B(n9515), .C(n8126), .Y(n2157) );
  OAI21X1 U4889 ( .A(n5164), .B(n9516), .C(n8034), .Y(n2156) );
  OAI21X1 U4891 ( .A(n5164), .B(n9517), .C(n7945), .Y(n2155) );
  OAI21X1 U4893 ( .A(n5164), .B(n9518), .C(n7858), .Y(n2154) );
  OAI21X1 U4895 ( .A(n5164), .B(n9519), .C(n7772), .Y(n2153) );
  OAI21X1 U4897 ( .A(n5164), .B(n9520), .C(n7392), .Y(n2152) );
  OAI21X1 U4899 ( .A(n5164), .B(n9521), .C(n7319), .Y(n2151) );
  OAI21X1 U4901 ( .A(n5164), .B(n9522), .C(n7247), .Y(n2150) );
  OAI21X1 U4903 ( .A(n5164), .B(n9523), .C(n7173), .Y(n2149) );
  OAI21X1 U4905 ( .A(n5164), .B(n9524), .C(n8399), .Y(n2148) );
  OAI21X1 U4907 ( .A(n5164), .B(n9525), .C(n8309), .Y(n2147) );
  OAI21X1 U4909 ( .A(n5164), .B(n9526), .C(n8219), .Y(n2146) );
  OAI21X1 U4911 ( .A(n5164), .B(n9527), .C(n8127), .Y(n2145) );
  OAI21X1 U4913 ( .A(n5164), .B(n9528), .C(n8035), .Y(n2144) );
  OAI21X1 U4915 ( .A(n5164), .B(n9529), .C(n7946), .Y(n2143) );
  OAI21X1 U4917 ( .A(n5164), .B(n9530), .C(n7859), .Y(n2142) );
  OAI21X1 U4919 ( .A(n5164), .B(n9531), .C(n7773), .Y(n2141) );
  OAI21X1 U4921 ( .A(n5164), .B(n9532), .C(n7393), .Y(n2140) );
  OAI21X1 U4923 ( .A(n5164), .B(n9533), .C(n7320), .Y(n2139) );
  OAI21X1 U4925 ( .A(n5164), .B(n9534), .C(n7248), .Y(n2138) );
  OAI21X1 U4927 ( .A(n5164), .B(n9535), .C(n7174), .Y(n2137) );
  OAI21X1 U4929 ( .A(n5164), .B(n9536), .C(n8400), .Y(n2136) );
  OAI21X1 U4931 ( .A(n5164), .B(n9537), .C(n8310), .Y(n2135) );
  OAI21X1 U4933 ( .A(n5164), .B(n9538), .C(n8220), .Y(n2134) );
  OAI21X1 U4935 ( .A(n5164), .B(n9539), .C(n8128), .Y(n2133) );
  OAI21X1 U4937 ( .A(n5164), .B(n9540), .C(n8036), .Y(n2132) );
  OAI21X1 U4939 ( .A(n5164), .B(n9541), .C(n7947), .Y(n2131) );
  OAI21X1 U4941 ( .A(n5164), .B(n9542), .C(n7860), .Y(n2130) );
  OAI21X1 U4943 ( .A(n5164), .B(n9543), .C(n7774), .Y(n2129) );
  OAI21X1 U4945 ( .A(n8153), .B(n8426), .C(n8500), .Y(n5164) );
  NAND3X1 U4946 ( .A(wr_ptr[2]), .B(wr_ptr[1]), .C(wr_ptr[0]), .Y(n4105) );
  OAI21X1 U4947 ( .A(n5207), .B(n9544), .C(n7175), .Y(n2128) );
  OAI21X1 U4949 ( .A(n5207), .B(n9545), .C(n7619), .Y(n2127) );
  OAI21X1 U4951 ( .A(n5207), .B(n9546), .C(n7694), .Y(n2126) );
  OAI21X1 U4953 ( .A(n5207), .B(n9547), .C(n7469), .Y(n2125) );
  OAI21X1 U4955 ( .A(n5207), .B(n9548), .C(n7544), .Y(n2124) );
  OAI21X1 U4957 ( .A(n5207), .B(n9549), .C(n5773), .Y(n2123) );
  OAI21X1 U4959 ( .A(n5207), .B(n9550), .C(n7620), .Y(n2122) );
  OAI21X1 U4961 ( .A(n5207), .B(n9551), .C(n7695), .Y(n2121) );
  OAI21X1 U4963 ( .A(n5207), .B(n9552), .C(n7470), .Y(n2120) );
  OAI21X1 U4965 ( .A(n5207), .B(n9553), .C(n7545), .Y(n2119) );
  OAI21X1 U4967 ( .A(n5207), .B(n9554), .C(n8401), .Y(n2118) );
  OAI21X1 U4969 ( .A(n5207), .B(n9555), .C(n8129), .Y(n2117) );
  OAI21X1 U4971 ( .A(n5207), .B(n9556), .C(n8221), .Y(n2116) );
  OAI21X1 U4973 ( .A(n5207), .B(n9557), .C(n7948), .Y(n2115) );
  OAI21X1 U4975 ( .A(n5207), .B(n9558), .C(n8037), .Y(n2114) );
  OAI21X1 U4977 ( .A(n5207), .B(n9559), .C(n7775), .Y(n2113) );
  OAI21X1 U4979 ( .A(n5207), .B(n9560), .C(n7861), .Y(n2112) );
  OAI21X1 U4981 ( .A(n5207), .B(n9561), .C(n7321), .Y(n2111) );
  OAI21X1 U4983 ( .A(n5207), .B(n9562), .C(n7394), .Y(n2110) );
  OAI21X1 U4985 ( .A(n5207), .B(n9563), .C(n7176), .Y(n2109) );
  OAI21X1 U4987 ( .A(n5207), .B(n9564), .C(n7249), .Y(n2108) );
  OAI21X1 U4989 ( .A(n5207), .B(n9565), .C(n8311), .Y(n2107) );
  OAI21X1 U4991 ( .A(n5207), .B(n9566), .C(n8402), .Y(n2106) );
  OAI21X1 U4993 ( .A(n5207), .B(n9567), .C(n8130), .Y(n2105) );
  OAI21X1 U4995 ( .A(n5207), .B(n9568), .C(n8222), .Y(n2104) );
  OAI21X1 U4997 ( .A(n5207), .B(n9569), .C(n7949), .Y(n2103) );
  OAI21X1 U4999 ( .A(n5207), .B(n9570), .C(n8038), .Y(n2102) );
  OAI21X1 U5001 ( .A(n5207), .B(n9571), .C(n7776), .Y(n2101) );
  OAI21X1 U5003 ( .A(n5207), .B(n9572), .C(n7862), .Y(n2100) );
  OAI21X1 U5005 ( .A(n5207), .B(n9573), .C(n7322), .Y(n2099) );
  OAI21X1 U5007 ( .A(n5207), .B(n9574), .C(n7395), .Y(n2098) );
  OAI21X1 U5009 ( .A(n5207), .B(n9575), .C(n7177), .Y(n2097) );
  OAI21X1 U5011 ( .A(n5207), .B(n9576), .C(n7250), .Y(n2096) );
  OAI21X1 U5013 ( .A(n5207), .B(n9577), .C(n8312), .Y(n2095) );
  OAI21X1 U5015 ( .A(n5207), .B(n9578), .C(n8403), .Y(n2094) );
  OAI21X1 U5017 ( .A(n5207), .B(n9579), .C(n8131), .Y(n2093) );
  OAI21X1 U5019 ( .A(n5207), .B(n9580), .C(n8223), .Y(n2092) );
  OAI21X1 U5021 ( .A(n5207), .B(n9581), .C(n7950), .Y(n2091) );
  OAI21X1 U5023 ( .A(n5207), .B(n9582), .C(n8039), .Y(n2090) );
  OAI21X1 U5025 ( .A(n5207), .B(n9583), .C(n7777), .Y(n2089) );
  OAI21X1 U5027 ( .A(n5207), .B(n9584), .C(n7863), .Y(n2088) );
  OAI21X1 U5029 ( .A(n8060), .B(n8426), .C(n8500), .Y(n5207) );
  NAND3X1 U5030 ( .A(wr_ptr[1]), .B(n8506), .C(wr_ptr[2]), .Y(n4232) );
  OAI21X1 U5031 ( .A(n5249), .B(n9585), .C(n7396), .Y(n2087) );
  OAI21X1 U5033 ( .A(n5249), .B(n9586), .C(n7546), .Y(n2086) );
  OAI21X1 U5035 ( .A(n5249), .B(n9587), .C(n7471), .Y(n2085) );
  OAI21X1 U5037 ( .A(n5249), .B(n9588), .C(n7696), .Y(n2084) );
  OAI21X1 U5039 ( .A(n5249), .B(n9589), .C(n7621), .Y(n2083) );
  OAI21X1 U5041 ( .A(n5249), .B(n9590), .C(n5772), .Y(n2082) );
  OAI21X1 U5043 ( .A(n5249), .B(n9591), .C(n7547), .Y(n2081) );
  OAI21X1 U5045 ( .A(n5249), .B(n9592), .C(n7472), .Y(n2080) );
  OAI21X1 U5047 ( .A(n5249), .B(n9593), .C(n7697), .Y(n2079) );
  OAI21X1 U5049 ( .A(n5249), .B(n9594), .C(n7622), .Y(n2078) );
  OAI21X1 U5051 ( .A(n5249), .B(n9595), .C(n8132), .Y(n2077) );
  OAI21X1 U5053 ( .A(n5249), .B(n9596), .C(n8404), .Y(n2076) );
  OAI21X1 U5055 ( .A(n5249), .B(n9597), .C(n8313), .Y(n2075) );
  OAI21X1 U5057 ( .A(n5249), .B(n9598), .C(n7864), .Y(n2074) );
  OAI21X1 U5059 ( .A(n5249), .B(n9599), .C(n7778), .Y(n2073) );
  OAI21X1 U5061 ( .A(n5249), .B(n9600), .C(n8040), .Y(n2072) );
  OAI21X1 U5063 ( .A(n5249), .B(n9601), .C(n7951), .Y(n2071) );
  OAI21X1 U5065 ( .A(n5249), .B(n9602), .C(n7251), .Y(n2070) );
  OAI21X1 U5067 ( .A(n5249), .B(n9603), .C(n7178), .Y(n2069) );
  OAI21X1 U5069 ( .A(n5249), .B(n9604), .C(n7397), .Y(n2068) );
  OAI21X1 U5071 ( .A(n5249), .B(n9605), .C(n7323), .Y(n2067) );
  OAI21X1 U5073 ( .A(n5249), .B(n9606), .C(n8224), .Y(n2066) );
  OAI21X1 U5075 ( .A(n5249), .B(n9607), .C(n8133), .Y(n2065) );
  OAI21X1 U5077 ( .A(n5249), .B(n9608), .C(n8405), .Y(n2064) );
  OAI21X1 U5079 ( .A(n5249), .B(n9609), .C(n8314), .Y(n2063) );
  OAI21X1 U5081 ( .A(n5249), .B(n9610), .C(n7865), .Y(n2062) );
  OAI21X1 U5083 ( .A(n5249), .B(n9611), .C(n7779), .Y(n2061) );
  OAI21X1 U5085 ( .A(n5249), .B(n9612), .C(n8041), .Y(n2060) );
  OAI21X1 U5087 ( .A(n5249), .B(n9613), .C(n7952), .Y(n2059) );
  OAI21X1 U5089 ( .A(n5249), .B(n9614), .C(n7252), .Y(n2058) );
  OAI21X1 U5091 ( .A(n5249), .B(n9615), .C(n7179), .Y(n2057) );
  OAI21X1 U5093 ( .A(n5249), .B(n9616), .C(n7398), .Y(n2056) );
  OAI21X1 U5095 ( .A(n5249), .B(n9617), .C(n7324), .Y(n2055) );
  OAI21X1 U5097 ( .A(n5249), .B(n9618), .C(n8225), .Y(n2054) );
  OAI21X1 U5099 ( .A(n5249), .B(n9619), .C(n8134), .Y(n2053) );
  OAI21X1 U5101 ( .A(n5249), .B(n9620), .C(n8406), .Y(n2052) );
  OAI21X1 U5103 ( .A(n5249), .B(n9621), .C(n8315), .Y(n2051) );
  OAI21X1 U5105 ( .A(n5249), .B(n9622), .C(n7866), .Y(n2050) );
  OAI21X1 U5107 ( .A(n5249), .B(n9623), .C(n7780), .Y(n2049) );
  OAI21X1 U5109 ( .A(n5249), .B(n9624), .C(n8042), .Y(n2048) );
  OAI21X1 U5111 ( .A(n5249), .B(n9625), .C(n7953), .Y(n2047) );
  OAI21X1 U5113 ( .A(n7969), .B(n8426), .C(n8500), .Y(n5249) );
  NAND3X1 U5114 ( .A(wr_ptr[2]), .B(n8516), .C(wr_ptr[0]), .Y(n4275) );
  OAI21X1 U5115 ( .A(n5291), .B(n9626), .C(n7325), .Y(n2046) );
  OAI21X1 U5117 ( .A(n5291), .B(n9627), .C(n7473), .Y(n2045) );
  OAI21X1 U5119 ( .A(n5291), .B(n9628), .C(n7548), .Y(n2044) );
  OAI21X1 U5121 ( .A(n5291), .B(n9629), .C(n7623), .Y(n2043) );
  OAI21X1 U5123 ( .A(n5291), .B(n9630), .C(n7698), .Y(n2042) );
  OAI21X1 U5125 ( .A(n5291), .B(n9631), .C(n5771), .Y(n2041) );
  OAI21X1 U5127 ( .A(n5291), .B(n9632), .C(n7474), .Y(n2040) );
  OAI21X1 U5129 ( .A(n5291), .B(n9633), .C(n7549), .Y(n2039) );
  OAI21X1 U5131 ( .A(n5291), .B(n9634), .C(n7624), .Y(n2038) );
  OAI21X1 U5133 ( .A(n5291), .B(n9635), .C(n7699), .Y(n2037) );
  OAI21X1 U5135 ( .A(n5291), .B(n9636), .C(n8226), .Y(n2036) );
  OAI21X1 U5137 ( .A(n5291), .B(n9637), .C(n8316), .Y(n2035) );
  OAI21X1 U5139 ( .A(n5291), .B(n9638), .C(n8407), .Y(n2034) );
  OAI21X1 U5141 ( .A(n5291), .B(n9639), .C(n7781), .Y(n2033) );
  OAI21X1 U5143 ( .A(n5291), .B(n9640), .C(n7867), .Y(n2032) );
  OAI21X1 U5145 ( .A(n5291), .B(n9641), .C(n7954), .Y(n2031) );
  OAI21X1 U5147 ( .A(n5291), .B(n9642), .C(n8043), .Y(n2030) );
  OAI21X1 U5149 ( .A(n5291), .B(n9643), .C(n7180), .Y(n2029) );
  OAI21X1 U5151 ( .A(n5291), .B(n9644), .C(n7253), .Y(n2028) );
  OAI21X1 U5153 ( .A(n5291), .B(n9645), .C(n7326), .Y(n2027) );
  OAI21X1 U5155 ( .A(n5291), .B(n9646), .C(n7399), .Y(n2026) );
  OAI21X1 U5157 ( .A(n5291), .B(n9647), .C(n8135), .Y(n2025) );
  OAI21X1 U5159 ( .A(n5291), .B(n9648), .C(n8227), .Y(n2024) );
  OAI21X1 U5161 ( .A(n5291), .B(n9649), .C(n8317), .Y(n2023) );
  OAI21X1 U5163 ( .A(n5291), .B(n9650), .C(n8408), .Y(n2022) );
  OAI21X1 U5165 ( .A(n5291), .B(n9651), .C(n7782), .Y(n2021) );
  OAI21X1 U5167 ( .A(n5291), .B(n9652), .C(n7868), .Y(n2020) );
  OAI21X1 U5169 ( .A(n5291), .B(n9653), .C(n7955), .Y(n2019) );
  OAI21X1 U5171 ( .A(n5291), .B(n9654), .C(n8044), .Y(n2018) );
  OAI21X1 U5173 ( .A(n5291), .B(n9655), .C(n7181), .Y(n2017) );
  OAI21X1 U5175 ( .A(n5291), .B(n9656), .C(n7254), .Y(n2016) );
  OAI21X1 U5177 ( .A(n5291), .B(n9657), .C(n7327), .Y(n2015) );
  OAI21X1 U5179 ( .A(n5291), .B(n9658), .C(n7400), .Y(n2014) );
  OAI21X1 U5181 ( .A(n5291), .B(n9659), .C(n8136), .Y(n2013) );
  OAI21X1 U5183 ( .A(n5291), .B(n9660), .C(n8228), .Y(n2012) );
  OAI21X1 U5185 ( .A(n5291), .B(n9661), .C(n8318), .Y(n2011) );
  OAI21X1 U5187 ( .A(n5291), .B(n9662), .C(n8409), .Y(n2010) );
  OAI21X1 U5189 ( .A(n5291), .B(n9663), .C(n7783), .Y(n2009) );
  OAI21X1 U5191 ( .A(n5291), .B(n9664), .C(n7869), .Y(n2008) );
  OAI21X1 U5193 ( .A(n5291), .B(n9665), .C(n7956), .Y(n2007) );
  OAI21X1 U5195 ( .A(n5291), .B(n9666), .C(n8045), .Y(n2006) );
  OAI21X1 U5197 ( .A(n8242), .B(n8426), .C(n8500), .Y(n5291) );
  NAND3X1 U5198 ( .A(n8506), .B(n8516), .C(wr_ptr[2]), .Y(n4318) );
  OAI21X1 U5199 ( .A(n5333), .B(n9667), .C(n7550), .Y(n2005) );
  OAI21X1 U5201 ( .A(n5333), .B(n9668), .C(n7401), .Y(n2004) );
  OAI21X1 U5203 ( .A(n5333), .B(n9669), .C(n7328), .Y(n2003) );
  OAI21X1 U5205 ( .A(n5333), .B(n9670), .C(n7255), .Y(n2002) );
  OAI21X1 U5207 ( .A(n5333), .B(n9671), .C(n7182), .Y(n2001) );
  OAI21X1 U5209 ( .A(n5333), .B(n9672), .C(n5770), .Y(n2000) );
  OAI21X1 U5211 ( .A(n5333), .B(n9673), .C(n7402), .Y(n1999) );
  OAI21X1 U5213 ( .A(n5333), .B(n9674), .C(n7329), .Y(n1998) );
  OAI21X1 U5215 ( .A(n5333), .B(n9675), .C(n7256), .Y(n1997) );
  OAI21X1 U5217 ( .A(n5333), .B(n9676), .C(n7183), .Y(n1996) );
  OAI21X1 U5219 ( .A(n5333), .B(n9677), .C(n7957), .Y(n1995) );
  OAI21X1 U5221 ( .A(n5333), .B(n9678), .C(n7870), .Y(n1994) );
  OAI21X1 U5223 ( .A(n5333), .B(n9679), .C(n7784), .Y(n1993) );
  OAI21X1 U5225 ( .A(n5333), .B(n9680), .C(n8410), .Y(n1992) );
  OAI21X1 U5227 ( .A(n5333), .B(n9681), .C(n8319), .Y(n1991) );
  OAI21X1 U5229 ( .A(n5333), .B(n9682), .C(n8229), .Y(n1990) );
  OAI21X1 U5231 ( .A(n5333), .B(n9683), .C(n8137), .Y(n1989) );
  OAI21X1 U5233 ( .A(n5333), .B(n9684), .C(n7700), .Y(n1988) );
  OAI21X1 U5235 ( .A(n5333), .B(n9685), .C(n7625), .Y(n1987) );
  OAI21X1 U5237 ( .A(n5333), .B(n9686), .C(n7551), .Y(n1986) );
  OAI21X1 U5239 ( .A(n5333), .B(n9687), .C(n7475), .Y(n1985) );
  OAI21X1 U5241 ( .A(n5333), .B(n9688), .C(n8046), .Y(n1984) );
  OAI21X1 U5243 ( .A(n5333), .B(n9689), .C(n7958), .Y(n1983) );
  OAI21X1 U5245 ( .A(n5333), .B(n9690), .C(n7871), .Y(n1982) );
  OAI21X1 U5247 ( .A(n5333), .B(n9691), .C(n7785), .Y(n1981) );
  OAI21X1 U5249 ( .A(n5333), .B(n9692), .C(n8411), .Y(n1980) );
  OAI21X1 U5251 ( .A(n5333), .B(n9693), .C(n8320), .Y(n1979) );
  OAI21X1 U5253 ( .A(n5333), .B(n9694), .C(n8230), .Y(n1978) );
  OAI21X1 U5255 ( .A(n5333), .B(n9695), .C(n8138), .Y(n1977) );
  OAI21X1 U5257 ( .A(n5333), .B(n9696), .C(n7701), .Y(n1976) );
  OAI21X1 U5259 ( .A(n5333), .B(n9697), .C(n7626), .Y(n1975) );
  OAI21X1 U5261 ( .A(n5333), .B(n9698), .C(n7552), .Y(n1974) );
  OAI21X1 U5263 ( .A(n5333), .B(n9699), .C(n7476), .Y(n1973) );
  OAI21X1 U5265 ( .A(n5333), .B(n9700), .C(n8047), .Y(n1972) );
  OAI21X1 U5267 ( .A(n5333), .B(n9701), .C(n7959), .Y(n1971) );
  OAI21X1 U5269 ( .A(n5333), .B(n9702), .C(n7872), .Y(n1970) );
  OAI21X1 U5271 ( .A(n5333), .B(n9703), .C(n7786), .Y(n1969) );
  OAI21X1 U5273 ( .A(n5333), .B(n9704), .C(n8412), .Y(n1968) );
  OAI21X1 U5275 ( .A(n5333), .B(n9705), .C(n8321), .Y(n1967) );
  OAI21X1 U5277 ( .A(n5333), .B(n9706), .C(n8231), .Y(n1966) );
  OAI21X1 U5279 ( .A(n5333), .B(n9707), .C(n8139), .Y(n1965) );
  OAI21X1 U5281 ( .A(n8243), .B(n8426), .C(n8500), .Y(n5333) );
  NAND3X1 U5282 ( .A(wr_ptr[1]), .B(n8517), .C(wr_ptr[0]), .Y(n4103) );
  OAI21X1 U5283 ( .A(n5375), .B(n9708), .C(n7477), .Y(n1964) );
  OAI21X1 U5285 ( .A(n5375), .B(n9709), .C(n7330), .Y(n1963) );
  OAI21X1 U5287 ( .A(n5375), .B(n9710), .C(n7403), .Y(n1962) );
  OAI21X1 U5289 ( .A(n5375), .B(n9711), .C(n7184), .Y(n1961) );
  OAI21X1 U5291 ( .A(n5375), .B(n9712), .C(n7257), .Y(n1960) );
  OAI21X1 U5293 ( .A(n5375), .B(n9713), .C(n5769), .Y(n1959) );
  OAI21X1 U5295 ( .A(n5375), .B(n9714), .C(n7331), .Y(n1958) );
  OAI21X1 U5297 ( .A(n5375), .B(n9715), .C(n7404), .Y(n1957) );
  OAI21X1 U5299 ( .A(n5375), .B(n9716), .C(n7185), .Y(n1956) );
  OAI21X1 U5301 ( .A(n5375), .B(n9717), .C(n7258), .Y(n1955) );
  OAI21X1 U5303 ( .A(n5375), .B(n9718), .C(n8048), .Y(n1954) );
  OAI21X1 U5305 ( .A(n5375), .B(n9719), .C(n7787), .Y(n1953) );
  OAI21X1 U5307 ( .A(n5375), .B(n9720), .C(n7873), .Y(n1952) );
  OAI21X1 U5309 ( .A(n5375), .B(n9721), .C(n8322), .Y(n1951) );
  OAI21X1 U5311 ( .A(n5375), .B(n9722), .C(n8413), .Y(n1950) );
  OAI21X1 U5313 ( .A(n5375), .B(n9723), .C(n8140), .Y(n1949) );
  OAI21X1 U5315 ( .A(n5375), .B(n9724), .C(n8232), .Y(n1948) );
  OAI21X1 U5317 ( .A(n5375), .B(n9725), .C(n7627), .Y(n1947) );
  OAI21X1 U5319 ( .A(n5375), .B(n9726), .C(n7702), .Y(n1946) );
  OAI21X1 U5321 ( .A(n5375), .B(n9727), .C(n7478), .Y(n1945) );
  OAI21X1 U5323 ( .A(n5375), .B(n9728), .C(n7553), .Y(n1944) );
  OAI21X1 U5325 ( .A(n5375), .B(n9729), .C(n7960), .Y(n1943) );
  OAI21X1 U5327 ( .A(n5375), .B(n9730), .C(n8049), .Y(n1942) );
  OAI21X1 U5329 ( .A(n5375), .B(n9731), .C(n7788), .Y(n1941) );
  OAI21X1 U5331 ( .A(n5375), .B(n9732), .C(n7874), .Y(n1940) );
  OAI21X1 U5333 ( .A(n5375), .B(n9733), .C(n8323), .Y(n1939) );
  OAI21X1 U5335 ( .A(n5375), .B(n9734), .C(n8414), .Y(n1938) );
  OAI21X1 U5337 ( .A(n5375), .B(n9735), .C(n8141), .Y(n1937) );
  OAI21X1 U5339 ( .A(n5375), .B(n9736), .C(n8233), .Y(n1936) );
  OAI21X1 U5341 ( .A(n5375), .B(n9737), .C(n7628), .Y(n1935) );
  OAI21X1 U5343 ( .A(n5375), .B(n9738), .C(n7703), .Y(n1934) );
  OAI21X1 U5345 ( .A(n5375), .B(n9739), .C(n7479), .Y(n1933) );
  OAI21X1 U5347 ( .A(n5375), .B(n9740), .C(n7554), .Y(n1932) );
  OAI21X1 U5349 ( .A(n5375), .B(n9741), .C(n7961), .Y(n1931) );
  OAI21X1 U5351 ( .A(n5375), .B(n9742), .C(n8050), .Y(n1930) );
  OAI21X1 U5353 ( .A(n5375), .B(n9743), .C(n7789), .Y(n1929) );
  OAI21X1 U5355 ( .A(n5375), .B(n9744), .C(n7875), .Y(n1928) );
  OAI21X1 U5357 ( .A(n5375), .B(n9745), .C(n8324), .Y(n1927) );
  OAI21X1 U5359 ( .A(n5375), .B(n9746), .C(n8415), .Y(n1926) );
  OAI21X1 U5361 ( .A(n5375), .B(n9747), .C(n8142), .Y(n1925) );
  OAI21X1 U5363 ( .A(n5375), .B(n9748), .C(n8234), .Y(n1924) );
  OAI21X1 U5365 ( .A(n7970), .B(n8426), .C(n8500), .Y(n5375) );
  NAND3X1 U5366 ( .A(n8506), .B(n8517), .C(wr_ptr[1]), .Y(n4403) );
  OAI21X1 U5367 ( .A(n5417), .B(n9749), .C(n7704), .Y(n1923) );
  OAI21X1 U5369 ( .A(n5417), .B(n9750), .C(n7259), .Y(n1922) );
  OAI21X1 U5371 ( .A(n5417), .B(n9751), .C(n7186), .Y(n1921) );
  OAI21X1 U5373 ( .A(n5417), .B(n9752), .C(n7405), .Y(n1920) );
  OAI21X1 U5375 ( .A(n5417), .B(n9753), .C(n7332), .Y(n1919) );
  OAI21X1 U5377 ( .A(n5417), .B(n9754), .C(n5768), .Y(n1918) );
  OAI21X1 U5379 ( .A(n5417), .B(n9755), .C(n7260), .Y(n1917) );
  OAI21X1 U5381 ( .A(n5417), .B(n9756), .C(n7187), .Y(n1916) );
  OAI21X1 U5383 ( .A(n5417), .B(n9757), .C(n7406), .Y(n1915) );
  OAI21X1 U5385 ( .A(n5417), .B(n9758), .C(n7333), .Y(n1914) );
  OAI21X1 U5387 ( .A(n5417), .B(n9759), .C(n7790), .Y(n1913) );
  OAI21X1 U5389 ( .A(n5417), .B(n9760), .C(n8051), .Y(n1912) );
  OAI21X1 U5391 ( .A(n5417), .B(n9761), .C(n7962), .Y(n1911) );
  OAI21X1 U5393 ( .A(n5417), .B(n9762), .C(n8235), .Y(n1910) );
  OAI21X1 U5395 ( .A(n5417), .B(n9763), .C(n8143), .Y(n1909) );
  OAI21X1 U5397 ( .A(n5417), .B(n9764), .C(n8416), .Y(n1908) );
  OAI21X1 U5399 ( .A(n5417), .B(n9765), .C(n8325), .Y(n1907) );
  OAI21X1 U5401 ( .A(n5417), .B(n9766), .C(n7555), .Y(n1906) );
  OAI21X1 U5403 ( .A(n5417), .B(n9767), .C(n7480), .Y(n1905) );
  OAI21X1 U5405 ( .A(n5417), .B(n9768), .C(n7705), .Y(n1904) );
  OAI21X1 U5407 ( .A(n5417), .B(n9769), .C(n7629), .Y(n1903) );
  OAI21X1 U5409 ( .A(n5417), .B(n9770), .C(n7876), .Y(n1902) );
  OAI21X1 U5411 ( .A(n5417), .B(n9771), .C(n7791), .Y(n1901) );
  OAI21X1 U5413 ( .A(n5417), .B(n9772), .C(n8052), .Y(n1900) );
  OAI21X1 U5415 ( .A(n5417), .B(n9773), .C(n7963), .Y(n1899) );
  OAI21X1 U5417 ( .A(n5417), .B(n9774), .C(n8236), .Y(n1898) );
  OAI21X1 U5419 ( .A(n5417), .B(n9775), .C(n8144), .Y(n1897) );
  OAI21X1 U5421 ( .A(n5417), .B(n9776), .C(n8417), .Y(n1896) );
  OAI21X1 U5423 ( .A(n5417), .B(n9777), .C(n8326), .Y(n1895) );
  OAI21X1 U5425 ( .A(n5417), .B(n9778), .C(n7556), .Y(n1894) );
  OAI21X1 U5427 ( .A(n5417), .B(n9779), .C(n7481), .Y(n1893) );
  OAI21X1 U5429 ( .A(n5417), .B(n9780), .C(n7706), .Y(n1892) );
  OAI21X1 U5431 ( .A(n5417), .B(n9781), .C(n7630), .Y(n1891) );
  OAI21X1 U5433 ( .A(n5417), .B(n9782), .C(n7877), .Y(n1890) );
  OAI21X1 U5435 ( .A(n5417), .B(n9783), .C(n7792), .Y(n1889) );
  OAI21X1 U5437 ( .A(n5417), .B(n9784), .C(n8053), .Y(n1888) );
  OAI21X1 U5439 ( .A(n5417), .B(n9785), .C(n7964), .Y(n1887) );
  OAI21X1 U5441 ( .A(n5417), .B(n9786), .C(n8237), .Y(n1886) );
  OAI21X1 U5443 ( .A(n5417), .B(n9787), .C(n8145), .Y(n1885) );
  OAI21X1 U5445 ( .A(n5417), .B(n9788), .C(n8418), .Y(n1884) );
  OAI21X1 U5447 ( .A(n5417), .B(n9789), .C(n8327), .Y(n1883) );
  OAI21X1 U5449 ( .A(n8061), .B(n8426), .C(n8500), .Y(n5417) );
  NAND3X1 U5450 ( .A(n8516), .B(n8517), .C(wr_ptr[0]), .Y(n4446) );
  OAI21X1 U5451 ( .A(n5459), .B(n9790), .C(n7631), .Y(n1882) );
  OAI21X1 U5453 ( .A(n5459), .B(n9791), .C(n7188), .Y(n1881) );
  OAI21X1 U5455 ( .A(n5459), .B(n9792), .C(n7261), .Y(n1880) );
  OAI21X1 U5457 ( .A(n5459), .B(n9793), .C(n7334), .Y(n1879) );
  OAI21X1 U5459 ( .A(n5459), .B(n9794), .C(n7407), .Y(n1878) );
  OAI21X1 U5461 ( .A(n5459), .B(n9795), .C(n5767), .Y(n1877) );
  OAI21X1 U5463 ( .A(n5459), .B(n9796), .C(n7189), .Y(n1876) );
  OAI21X1 U5465 ( .A(n5459), .B(n9797), .C(n7262), .Y(n1875) );
  OAI21X1 U5467 ( .A(n5459), .B(n9798), .C(n7335), .Y(n1874) );
  OAI21X1 U5469 ( .A(n5459), .B(n9799), .C(n7408), .Y(n1873) );
  OAI21X1 U5471 ( .A(n5459), .B(n9800), .C(n7878), .Y(n1872) );
  OAI21X1 U5473 ( .A(n5459), .B(n9801), .C(n7965), .Y(n1871) );
  OAI21X1 U5475 ( .A(n5459), .B(n9802), .C(n8054), .Y(n1870) );
  OAI21X1 U5477 ( .A(n5459), .B(n9803), .C(n8146), .Y(n1869) );
  OAI21X1 U5479 ( .A(n5459), .B(n9804), .C(n8238), .Y(n1868) );
  OAI21X1 U5481 ( .A(n5459), .B(n9805), .C(n8328), .Y(n1867) );
  OAI21X1 U5483 ( .A(n5459), .B(n9806), .C(n8419), .Y(n1866) );
  OAI21X1 U5485 ( .A(n5459), .B(n9807), .C(n7482), .Y(n1865) );
  OAI21X1 U5487 ( .A(n5459), .B(n9808), .C(n7557), .Y(n1864) );
  OAI21X1 U5489 ( .A(n5459), .B(n9809), .C(n7632), .Y(n1863) );
  OAI21X1 U5491 ( .A(n5459), .B(n9810), .C(n7707), .Y(n1862) );
  OAI21X1 U5493 ( .A(n5459), .B(n9811), .C(n7793), .Y(n1861) );
  OAI21X1 U5495 ( .A(n5459), .B(n9812), .C(n7879), .Y(n1860) );
  OAI21X1 U5497 ( .A(n5459), .B(n9813), .C(n7966), .Y(n1859) );
  OAI21X1 U5499 ( .A(n5459), .B(n9814), .C(n8055), .Y(n1858) );
  OAI21X1 U5501 ( .A(n5459), .B(n9815), .C(n8147), .Y(n1857) );
  OAI21X1 U5503 ( .A(n5459), .B(n9816), .C(n8239), .Y(n1856) );
  OAI21X1 U5505 ( .A(n5459), .B(n9817), .C(n8329), .Y(n1855) );
  OAI21X1 U5507 ( .A(n5459), .B(n9818), .C(n8420), .Y(n1854) );
  OAI21X1 U5509 ( .A(n5459), .B(n9819), .C(n7483), .Y(n1853) );
  OAI21X1 U5511 ( .A(n5459), .B(n9820), .C(n7558), .Y(n1852) );
  OAI21X1 U5513 ( .A(n5459), .B(n9821), .C(n7633), .Y(n1851) );
  OAI21X1 U5515 ( .A(n5459), .B(n9822), .C(n7708), .Y(n1850) );
  OAI21X1 U5517 ( .A(n5459), .B(n9823), .C(n7794), .Y(n1849) );
  OAI21X1 U5519 ( .A(n5459), .B(n9824), .C(n7880), .Y(n1848) );
  OAI21X1 U5521 ( .A(n5459), .B(n9825), .C(n7967), .Y(n1847) );
  OAI21X1 U5523 ( .A(n5459), .B(n9826), .C(n8056), .Y(n1846) );
  OAI21X1 U5525 ( .A(n5459), .B(n9827), .C(n8148), .Y(n1845) );
  OAI21X1 U5527 ( .A(n5459), .B(n9828), .C(n8240), .Y(n1844) );
  OAI21X1 U5529 ( .A(n5459), .B(n9829), .C(n8330), .Y(n1843) );
  OAI21X1 U5531 ( .A(n5459), .B(n9830), .C(n8421), .Y(n1842) );
  OAI21X1 U5533 ( .A(n8152), .B(n8426), .C(n8500), .Y(n5459) );
  NAND3X1 U5534 ( .A(n8518), .B(n8515), .C(put), .Y(n5206) );
  NAND3X1 U5535 ( .A(n8516), .B(n8517), .C(n8506), .Y(n4489) );
  XNOR2X1 U5536 ( .A(n8503), .B(n4094), .Y(fillcount[4]) );
  XNOR2X1 U5537 ( .A(n16), .B(n8515), .Y(n4094) );
  AOI21X1 U5538 ( .A(n8514), .B(n5501), .C(n6127), .Y(n1343) );
  AOI21X1 U5539 ( .A(n8504), .B(n15), .C(n8518), .Y(n5502) );
  XOR2X1 U5540 ( .A(n5501), .B(n4091), .Y(fillcount[3]) );
  XNOR2X1 U5541 ( .A(n15), .B(wr_ptr[3]), .Y(n4091) );
  OAI21X1 U5542 ( .A(n14), .B(n7881), .C(n5504), .Y(n5501) );
  OAI21X1 U5543 ( .A(n8505), .B(n8513), .C(wr_ptr[2]), .Y(n5504) );
  XOR2X1 U5544 ( .A(n8505), .B(n4090), .Y(fillcount[2]) );
  XNOR2X1 U5545 ( .A(n14), .B(wr_ptr[2]), .Y(n4090) );
  AOI21X1 U5546 ( .A(n8512), .B(n8423), .C(n7882), .Y(n5503) );
  AOI21X1 U5547 ( .A(n5505), .B(n13), .C(n8516), .Y(n5506) );
  XNOR2X1 U5548 ( .A(n8423), .B(n4093), .Y(fillcount[1]) );
  XNOR2X1 U5549 ( .A(n13), .B(n8516), .Y(n4093) );
  OAI21X1 U5550 ( .A(n12), .B(n8506), .C(n8423), .Y(fillcount[0]) );
  OR2X1 U3 ( .A(n5857), .B(n6021), .Y(n3564) );
  OR2X1 U4 ( .A(n5858), .B(n6022), .Y(n3565) );
  OR2X1 U5 ( .A(n5856), .B(n6020), .Y(n3563) );
  OR2X1 U6 ( .A(n5941), .B(n6105), .Y(n1528) );
  OR2X1 U7 ( .A(n5942), .B(n6106), .Y(n1529) );
  OR2X1 U8 ( .A(n5940), .B(n6104), .Y(n1527) );
  OR2X1 U9 ( .A(n5861), .B(n6025), .Y(n3530) );
  OR2X1 U10 ( .A(n5862), .B(n6026), .Y(n3531) );
  OR2X1 U11 ( .A(n5860), .B(n6024), .Y(n3529) );
  OR2X1 U12 ( .A(n5945), .B(n6109), .Y(n1494) );
  OR2X1 U13 ( .A(n5946), .B(n6110), .Y(n1495) );
  OR2X1 U14 ( .A(n5944), .B(n6108), .Y(n1493) );
  OR2X1 U15 ( .A(n5865), .B(n6029), .Y(n3496) );
  OR2X1 U16 ( .A(n5866), .B(n6030), .Y(n3497) );
  OR2X1 U17 ( .A(n5864), .B(n6028), .Y(n3495) );
  OR2X1 U18 ( .A(n5949), .B(n6113), .Y(n1460) );
  OR2X1 U19 ( .A(n5950), .B(n6114), .Y(n1461) );
  OR2X1 U20 ( .A(n5948), .B(n6112), .Y(n1459) );
  OR2X1 U21 ( .A(n5869), .B(n6033), .Y(n3462) );
  OR2X1 U22 ( .A(n5870), .B(n6034), .Y(n3463) );
  OR2X1 U23 ( .A(n5868), .B(n6032), .Y(n3461) );
  OR2X1 U24 ( .A(n5953), .B(n6117), .Y(n1426) );
  OR2X1 U25 ( .A(n5954), .B(n6118), .Y(n1427) );
  OR2X1 U26 ( .A(n5952), .B(n6116), .Y(n1425) );
  OR2X1 U27 ( .A(n5873), .B(n6037), .Y(n3428) );
  OR2X1 U28 ( .A(n5874), .B(n6038), .Y(n3429) );
  OR2X1 U29 ( .A(n5872), .B(n6036), .Y(n3427) );
  OR2X1 U30 ( .A(n5957), .B(n6121), .Y(n1392) );
  OR2X1 U31 ( .A(n5958), .B(n6122), .Y(n1393) );
  OR2X1 U32 ( .A(n5956), .B(n6120), .Y(n1391) );
  OR2X1 U33 ( .A(n5877), .B(n6041), .Y(n3394) );
  OR2X1 U34 ( .A(n5878), .B(n6042), .Y(n3395) );
  OR2X1 U35 ( .A(n5876), .B(n6040), .Y(n3393) );
  OR2X1 U36 ( .A(n5961), .B(n6125), .Y(n1348) );
  OR2X1 U37 ( .A(n5962), .B(n6126), .Y(n1349) );
  OR2X1 U38 ( .A(n5960), .B(n6124), .Y(n1347) );
  OR2X1 U39 ( .A(n5800), .B(n5964), .Y(n4039) );
  OR2X1 U40 ( .A(n5801), .B(n5965), .Y(n4040) );
  OR2X1 U41 ( .A(n5802), .B(n5966), .Y(n4041) );
  OR2X1 U42 ( .A(n5804), .B(n5968), .Y(n4005) );
  OR2X1 U43 ( .A(n5805), .B(n5969), .Y(n4006) );
  OR2X1 U44 ( .A(n5806), .B(n5970), .Y(n4007) );
  OR2X1 U45 ( .A(n5808), .B(n5972), .Y(n3971) );
  OR2X1 U46 ( .A(n5809), .B(n5973), .Y(n3972) );
  OR2X1 U47 ( .A(n5810), .B(n5974), .Y(n3973) );
  OR2X1 U48 ( .A(n5812), .B(n5976), .Y(n3937) );
  OR2X1 U49 ( .A(n5813), .B(n5977), .Y(n3938) );
  OR2X1 U50 ( .A(n5814), .B(n5978), .Y(n3939) );
  OR2X1 U51 ( .A(n5816), .B(n5980), .Y(n3903) );
  OR2X1 U52 ( .A(n5817), .B(n5981), .Y(n3904) );
  OR2X1 U53 ( .A(n5818), .B(n5982), .Y(n3905) );
  OR2X1 U54 ( .A(n5820), .B(n5984), .Y(n3869) );
  OR2X1 U55 ( .A(n5821), .B(n5985), .Y(n3870) );
  OR2X1 U56 ( .A(n5822), .B(n5986), .Y(n3871) );
  OR2X1 U57 ( .A(n5824), .B(n5988), .Y(n3835) );
  OR2X1 U58 ( .A(n5825), .B(n5989), .Y(n3836) );
  OR2X1 U59 ( .A(n5826), .B(n5990), .Y(n3837) );
  OR2X1 U60 ( .A(n5828), .B(n5992), .Y(n3801) );
  OR2X1 U61 ( .A(n5829), .B(n5993), .Y(n3802) );
  OR2X1 U62 ( .A(n5830), .B(n5994), .Y(n3803) );
  OR2X1 U63 ( .A(n5832), .B(n5996), .Y(n3767) );
  OR2X1 U64 ( .A(n5833), .B(n5997), .Y(n3768) );
  OR2X1 U65 ( .A(n5834), .B(n5998), .Y(n3769) );
  OR2X1 U66 ( .A(n5836), .B(n6000), .Y(n3733) );
  OR2X1 U67 ( .A(n5837), .B(n6001), .Y(n3734) );
  OR2X1 U68 ( .A(n5838), .B(n6002), .Y(n3735) );
  OR2X1 U69 ( .A(n5840), .B(n6004), .Y(n3699) );
  OR2X1 U70 ( .A(n5841), .B(n6005), .Y(n3700) );
  OR2X1 U71 ( .A(n5842), .B(n6006), .Y(n3701) );
  OR2X1 U72 ( .A(n5844), .B(n6008), .Y(n3665) );
  OR2X1 U73 ( .A(n5845), .B(n6009), .Y(n3666) );
  OR2X1 U74 ( .A(n5846), .B(n6010), .Y(n3667) );
  OR2X1 U75 ( .A(n5885), .B(n6049), .Y(n3326) );
  OR2X1 U76 ( .A(n5886), .B(n6050), .Y(n3327) );
  OR2X1 U77 ( .A(n5884), .B(n6048), .Y(n3325) );
  OR2X1 U78 ( .A(n5889), .B(n6053), .Y(n3292) );
  OR2X1 U79 ( .A(n5890), .B(n6054), .Y(n3293) );
  OR2X1 U80 ( .A(n5888), .B(n6052), .Y(n3291) );
  OR2X1 U81 ( .A(n5893), .B(n6057), .Y(n3258) );
  OR2X1 U82 ( .A(n5894), .B(n6058), .Y(n3259) );
  OR2X1 U83 ( .A(n5892), .B(n6056), .Y(n3257) );
  OR2X1 U84 ( .A(n5897), .B(n6061), .Y(n3224) );
  OR2X1 U85 ( .A(n5898), .B(n6062), .Y(n3225) );
  OR2X1 U86 ( .A(n5896), .B(n6060), .Y(n3223) );
  OR2X1 U87 ( .A(n5901), .B(n6065), .Y(n3190) );
  OR2X1 U88 ( .A(n5902), .B(n6066), .Y(n3191) );
  OR2X1 U89 ( .A(n5900), .B(n6064), .Y(n3189) );
  OR2X1 U90 ( .A(n5905), .B(n6069), .Y(n1834) );
  OR2X1 U91 ( .A(n5906), .B(n6070), .Y(n1835) );
  OR2X1 U92 ( .A(n5904), .B(n6068), .Y(n1833) );
  OR2X1 U93 ( .A(n5909), .B(n6073), .Y(n1800) );
  OR2X1 U94 ( .A(n5910), .B(n6074), .Y(n1801) );
  OR2X1 U95 ( .A(n5908), .B(n6072), .Y(n1799) );
  OR2X1 U96 ( .A(n5913), .B(n6077), .Y(n1766) );
  OR2X1 U97 ( .A(n5914), .B(n6078), .Y(n1767) );
  OR2X1 U98 ( .A(n5912), .B(n6076), .Y(n1765) );
  OR2X1 U99 ( .A(n5917), .B(n6081), .Y(n1732) );
  OR2X1 U100 ( .A(n5918), .B(n6082), .Y(n1733) );
  OR2X1 U101 ( .A(n5916), .B(n6080), .Y(n1731) );
  OR2X1 U102 ( .A(n5921), .B(n6085), .Y(n1698) );
  OR2X1 U103 ( .A(n5922), .B(n6086), .Y(n1699) );
  OR2X1 U104 ( .A(n5920), .B(n6084), .Y(n1697) );
  OR2X1 U105 ( .A(n5925), .B(n6089), .Y(n1664) );
  OR2X1 U106 ( .A(n5926), .B(n6090), .Y(n1665) );
  OR2X1 U107 ( .A(n5924), .B(n6088), .Y(n1663) );
  OR2X1 U108 ( .A(n5929), .B(n6093), .Y(n1630) );
  OR2X1 U109 ( .A(n5930), .B(n6094), .Y(n1631) );
  OR2X1 U110 ( .A(n5928), .B(n6092), .Y(n1629) );
  OR2X1 U111 ( .A(n5933), .B(n6097), .Y(n1596) );
  OR2X1 U112 ( .A(n5934), .B(n6098), .Y(n1597) );
  OR2X1 U113 ( .A(n5932), .B(n6096), .Y(n1595) );
  OR2X1 U114 ( .A(n5849), .B(n6013), .Y(n3632) );
  OR2X1 U115 ( .A(n5850), .B(n6014), .Y(n3633) );
  OR2X1 U116 ( .A(n5848), .B(n6012), .Y(n3631) );
  OR2X1 U117 ( .A(n5881), .B(n6045), .Y(n3360) );
  OR2X1 U118 ( .A(n5882), .B(n6046), .Y(n3361) );
  OR2X1 U119 ( .A(n5880), .B(n6044), .Y(n3359) );
  OR2X1 U120 ( .A(n5937), .B(n6101), .Y(n1562) );
  OR2X1 U121 ( .A(n5938), .B(n6102), .Y(n1563) );
  OR2X1 U122 ( .A(n5936), .B(n6100), .Y(n1561) );
  OR2X1 U123 ( .A(n5853), .B(n6017), .Y(n3598) );
  OR2X1 U124 ( .A(n5854), .B(n6018), .Y(n3599) );
  OR2X1 U125 ( .A(n5852), .B(n6016), .Y(n3597) );
  AND2X1 U126 ( .A(get), .B(empty_bar), .Y(n4089) );
  OR2X1 U127 ( .A(n5855), .B(n6019), .Y(n3561) );
  OR2X1 U128 ( .A(n5939), .B(n6103), .Y(n1525) );
  OR2X1 U129 ( .A(n5859), .B(n6023), .Y(n3527) );
  OR2X1 U130 ( .A(n5943), .B(n6107), .Y(n1491) );
  OR2X1 U131 ( .A(n5863), .B(n6027), .Y(n3493) );
  OR2X1 U132 ( .A(n5947), .B(n6111), .Y(n1457) );
  OR2X1 U133 ( .A(n5867), .B(n6031), .Y(n3459) );
  OR2X1 U134 ( .A(n5951), .B(n6115), .Y(n1423) );
  OR2X1 U135 ( .A(n5871), .B(n6035), .Y(n3425) );
  OR2X1 U136 ( .A(n5955), .B(n6119), .Y(n1389) );
  OR2X1 U137 ( .A(n5875), .B(n6039), .Y(n3391) );
  OR2X1 U138 ( .A(n5959), .B(n6123), .Y(n1345) );
  OR2X1 U139 ( .A(n5799), .B(n5963), .Y(n4037) );
  OR2X1 U140 ( .A(n5803), .B(n5967), .Y(n4003) );
  OR2X1 U141 ( .A(n5807), .B(n5971), .Y(n3969) );
  OR2X1 U142 ( .A(n5811), .B(n5975), .Y(n3935) );
  OR2X1 U143 ( .A(n5815), .B(n5979), .Y(n3901) );
  OR2X1 U144 ( .A(n5819), .B(n5983), .Y(n3867) );
  OR2X1 U145 ( .A(n5823), .B(n5987), .Y(n3833) );
  OR2X1 U146 ( .A(n5827), .B(n5991), .Y(n3799) );
  OR2X1 U147 ( .A(n5831), .B(n5995), .Y(n3765) );
  OR2X1 U148 ( .A(n5835), .B(n5999), .Y(n3731) );
  OR2X1 U149 ( .A(n5839), .B(n6003), .Y(n3697) );
  OR2X1 U150 ( .A(n5843), .B(n6007), .Y(n3663) );
  OR2X1 U151 ( .A(n5883), .B(n6047), .Y(n3323) );
  OR2X1 U152 ( .A(n5887), .B(n6051), .Y(n3289) );
  OR2X1 U153 ( .A(n5891), .B(n6055), .Y(n3255) );
  OR2X1 U154 ( .A(n5895), .B(n6059), .Y(n3221) );
  OR2X1 U155 ( .A(n5899), .B(n6063), .Y(n3187) );
  OR2X1 U156 ( .A(n5903), .B(n6067), .Y(n1831) );
  OR2X1 U157 ( .A(n5907), .B(n6071), .Y(n1797) );
  OR2X1 U158 ( .A(n5911), .B(n6075), .Y(n1763) );
  OR2X1 U159 ( .A(n5915), .B(n6079), .Y(n1729) );
  OR2X1 U160 ( .A(n5919), .B(n6083), .Y(n1695) );
  OR2X1 U161 ( .A(n5923), .B(n6087), .Y(n1661) );
  OR2X1 U162 ( .A(n5927), .B(n6091), .Y(n1627) );
  OR2X1 U163 ( .A(n5931), .B(n6095), .Y(n1593) );
  OR2X1 U164 ( .A(n5847), .B(n6011), .Y(n3629) );
  OR2X1 U165 ( .A(n5879), .B(n6043), .Y(n3357) );
  OR2X1 U166 ( .A(n5935), .B(n6099), .Y(n1559) );
  OR2X1 U167 ( .A(n5851), .B(n6015), .Y(n3595) );
  OR2X1 U168 ( .A(n8243), .B(n8424), .Y(n4102) );
  OR2X1 U169 ( .A(n8332), .B(n8506), .Y(n4077) );
  AND2X1 U170 ( .A(reset), .B(n8150), .Y(n4082) );
  AND2X1 U171 ( .A(n8500), .B(n8149), .Y(n4062) );
  AND2X1 U172 ( .A(n8500), .B(n8332), .Y(n4076) );
  BUFX2 U173 ( .A(n3162), .Y(n5723) );
  BUFX2 U174 ( .A(n5547), .Y(n5724) );
  BUFX2 U175 ( .A(n5546), .Y(n5725) );
  BUFX2 U176 ( .A(n5545), .Y(n5726) );
  BUFX2 U177 ( .A(n5544), .Y(n5727) );
  BUFX2 U178 ( .A(n5543), .Y(n5728) );
  BUFX2 U179 ( .A(n5542), .Y(n5729) );
  BUFX2 U180 ( .A(n5541), .Y(n5730) );
  BUFX2 U181 ( .A(n5540), .Y(n5731) );
  BUFX2 U182 ( .A(n5539), .Y(n5732) );
  BUFX2 U183 ( .A(n5538), .Y(n5733) );
  BUFX2 U184 ( .A(n5537), .Y(n5734) );
  BUFX2 U185 ( .A(n5536), .Y(n5735) );
  BUFX2 U186 ( .A(n5535), .Y(n5736) );
  BUFX2 U187 ( .A(n5534), .Y(n5737) );
  BUFX2 U188 ( .A(n5533), .Y(n5738) );
  BUFX2 U189 ( .A(n5532), .Y(n5739) );
  BUFX2 U190 ( .A(n5531), .Y(n5740) );
  BUFX2 U191 ( .A(n5530), .Y(n5741) );
  BUFX2 U192 ( .A(n5529), .Y(n5742) );
  BUFX2 U193 ( .A(n5528), .Y(n5743) );
  BUFX2 U194 ( .A(n5527), .Y(n5744) );
  BUFX2 U195 ( .A(n5526), .Y(n5745) );
  BUFX2 U196 ( .A(n5525), .Y(n5746) );
  BUFX2 U197 ( .A(n5524), .Y(n5747) );
  BUFX2 U198 ( .A(n5523), .Y(n5748) );
  BUFX2 U199 ( .A(n5522), .Y(n5749) );
  BUFX2 U200 ( .A(n5521), .Y(n5750) );
  BUFX2 U201 ( .A(n5520), .Y(n5751) );
  BUFX2 U202 ( .A(n5519), .Y(n5752) );
  BUFX2 U203 ( .A(n5518), .Y(n5753) );
  BUFX2 U204 ( .A(n5517), .Y(n5754) );
  BUFX2 U205 ( .A(n5516), .Y(n5755) );
  BUFX2 U206 ( .A(n5515), .Y(n5756) );
  BUFX2 U207 ( .A(n5514), .Y(n5757) );
  BUFX2 U208 ( .A(n5513), .Y(n5758) );
  BUFX2 U209 ( .A(n5512), .Y(n5759) );
  BUFX2 U210 ( .A(n5511), .Y(n5760) );
  BUFX2 U211 ( .A(n5510), .Y(n5761) );
  BUFX2 U212 ( .A(n5509), .Y(n5762) );
  BUFX2 U213 ( .A(n5508), .Y(n5763) );
  BUFX2 U214 ( .A(n5507), .Y(n5764) );
  BUFX2 U215 ( .A(n4088), .Y(n5765) );
  BUFX2 U216 ( .A(n4085), .Y(n5766) );
  AND2X1 U217 ( .A(n4118), .B(n5459), .Y(n5465) );
  INVX1 U218 ( .A(n5465), .Y(n5767) );
  AND2X1 U219 ( .A(n4118), .B(n5417), .Y(n5423) );
  INVX1 U220 ( .A(n5423), .Y(n5768) );
  AND2X1 U221 ( .A(n4118), .B(n5375), .Y(n5381) );
  INVX1 U222 ( .A(n5381), .Y(n5769) );
  AND2X1 U223 ( .A(n4118), .B(n5333), .Y(n5339) );
  INVX1 U224 ( .A(n5339), .Y(n5770) );
  AND2X1 U225 ( .A(n4118), .B(n5291), .Y(n5297) );
  INVX1 U226 ( .A(n5297), .Y(n5771) );
  AND2X1 U227 ( .A(n4118), .B(n5249), .Y(n5255) );
  INVX1 U228 ( .A(n5255), .Y(n5772) );
  AND2X1 U229 ( .A(n4118), .B(n5207), .Y(n5213) );
  INVX1 U230 ( .A(n5213), .Y(n5773) );
  AND2X1 U231 ( .A(n4118), .B(n5164), .Y(n5170) );
  INVX1 U232 ( .A(n5170), .Y(n5774) );
  AND2X1 U233 ( .A(n4118), .B(n5122), .Y(n5128) );
  INVX1 U234 ( .A(n5128), .Y(n5775) );
  AND2X1 U235 ( .A(n4118), .B(n5080), .Y(n5086) );
  INVX1 U236 ( .A(n5086), .Y(n5776) );
  AND2X1 U237 ( .A(n4118), .B(n5038), .Y(n5044) );
  INVX1 U238 ( .A(n5044), .Y(n5777) );
  AND2X1 U239 ( .A(n4118), .B(n4996), .Y(n5002) );
  INVX1 U240 ( .A(n5002), .Y(n5778) );
  AND2X1 U241 ( .A(n4118), .B(n4954), .Y(n4960) );
  INVX1 U242 ( .A(n4960), .Y(n5779) );
  AND2X1 U243 ( .A(n4118), .B(n4912), .Y(n4918) );
  INVX1 U244 ( .A(n4918), .Y(n5780) );
  AND2X1 U245 ( .A(n4118), .B(n4870), .Y(n4876) );
  INVX1 U246 ( .A(n4876), .Y(n5781) );
  AND2X1 U247 ( .A(n4118), .B(n4827), .Y(n4833) );
  INVX1 U248 ( .A(n4833), .Y(n5782) );
  AND2X1 U249 ( .A(n4118), .B(n4785), .Y(n4791) );
  INVX1 U250 ( .A(n4791), .Y(n5783) );
  AND2X1 U251 ( .A(n4118), .B(n4743), .Y(n4749) );
  INVX1 U252 ( .A(n4749), .Y(n5784) );
  AND2X1 U253 ( .A(n4118), .B(n4701), .Y(n4707) );
  INVX1 U254 ( .A(n4707), .Y(n5785) );
  AND2X1 U255 ( .A(n4118), .B(n4659), .Y(n4665) );
  INVX1 U256 ( .A(n4665), .Y(n5786) );
  AND2X1 U257 ( .A(n4118), .B(n4617), .Y(n4623) );
  INVX1 U258 ( .A(n4623), .Y(n5787) );
  AND2X1 U259 ( .A(n4118), .B(n4575), .Y(n4581) );
  INVX1 U260 ( .A(n4581), .Y(n5788) );
  AND2X1 U261 ( .A(n4118), .B(n4533), .Y(n4539) );
  INVX1 U262 ( .A(n4539), .Y(n5789) );
  AND2X1 U263 ( .A(n4118), .B(n4490), .Y(n4496) );
  INVX1 U264 ( .A(n4496), .Y(n5790) );
  AND2X1 U265 ( .A(n4118), .B(n4447), .Y(n4453) );
  INVX1 U266 ( .A(n4453), .Y(n5791) );
  AND2X1 U267 ( .A(n4118), .B(n4404), .Y(n4410) );
  INVX1 U268 ( .A(n4410), .Y(n5792) );
  AND2X1 U269 ( .A(n4118), .B(n4361), .Y(n4367) );
  INVX1 U270 ( .A(n4367), .Y(n5793) );
  AND2X1 U271 ( .A(n4118), .B(n4319), .Y(n4325) );
  INVX1 U272 ( .A(n4325), .Y(n5794) );
  AND2X1 U273 ( .A(n4118), .B(n4276), .Y(n4282) );
  INVX1 U274 ( .A(n4282), .Y(n5795) );
  AND2X1 U275 ( .A(n4118), .B(n4233), .Y(n4239) );
  INVX1 U276 ( .A(n4239), .Y(n5796) );
  AND2X1 U277 ( .A(n4118), .B(n4190), .Y(n4196) );
  INVX1 U278 ( .A(n4196), .Y(n5797) );
  AND2X1 U279 ( .A(n4118), .B(n4106), .Y(n4117) );
  INVX1 U280 ( .A(n4117), .Y(n5798) );
  BUFX2 U281 ( .A(n4066), .Y(n5799) );
  BUFX2 U282 ( .A(n4058), .Y(n5800) );
  BUFX2 U283 ( .A(n4050), .Y(n5801) );
  BUFX2 U284 ( .A(n4042), .Y(n5802) );
  BUFX2 U285 ( .A(n4029), .Y(n5803) );
  BUFX2 U286 ( .A(n4022), .Y(n5804) );
  BUFX2 U287 ( .A(n4015), .Y(n5805) );
  BUFX2 U288 ( .A(n4008), .Y(n5806) );
  BUFX2 U289 ( .A(n3995), .Y(n5807) );
  BUFX2 U290 ( .A(n3988), .Y(n5808) );
  BUFX2 U291 ( .A(n3981), .Y(n5809) );
  BUFX2 U292 ( .A(n3974), .Y(n5810) );
  BUFX2 U293 ( .A(n3961), .Y(n5811) );
  BUFX2 U294 ( .A(n3954), .Y(n5812) );
  BUFX2 U295 ( .A(n3947), .Y(n5813) );
  BUFX2 U296 ( .A(n3940), .Y(n5814) );
  BUFX2 U297 ( .A(n3927), .Y(n5815) );
  BUFX2 U298 ( .A(n3920), .Y(n5816) );
  BUFX2 U299 ( .A(n3913), .Y(n5817) );
  BUFX2 U300 ( .A(n3906), .Y(n5818) );
  BUFX2 U301 ( .A(n3893), .Y(n5819) );
  BUFX2 U302 ( .A(n3886), .Y(n5820) );
  BUFX2 U303 ( .A(n3879), .Y(n5821) );
  BUFX2 U304 ( .A(n3872), .Y(n5822) );
  BUFX2 U305 ( .A(n3859), .Y(n5823) );
  BUFX2 U306 ( .A(n3852), .Y(n5824) );
  BUFX2 U307 ( .A(n3845), .Y(n5825) );
  BUFX2 U308 ( .A(n3838), .Y(n5826) );
  BUFX2 U309 ( .A(n3825), .Y(n5827) );
  BUFX2 U310 ( .A(n3818), .Y(n5828) );
  BUFX2 U311 ( .A(n3811), .Y(n5829) );
  BUFX2 U312 ( .A(n3804), .Y(n5830) );
  BUFX2 U313 ( .A(n3791), .Y(n5831) );
  BUFX2 U314 ( .A(n3784), .Y(n5832) );
  BUFX2 U315 ( .A(n3777), .Y(n5833) );
  BUFX2 U316 ( .A(n3770), .Y(n5834) );
  BUFX2 U317 ( .A(n3757), .Y(n5835) );
  BUFX2 U318 ( .A(n3750), .Y(n5836) );
  BUFX2 U319 ( .A(n3743), .Y(n5837) );
  BUFX2 U320 ( .A(n3736), .Y(n5838) );
  BUFX2 U321 ( .A(n3723), .Y(n5839) );
  BUFX2 U322 ( .A(n3716), .Y(n5840) );
  BUFX2 U323 ( .A(n3709), .Y(n5841) );
  BUFX2 U324 ( .A(n3702), .Y(n5842) );
  BUFX2 U325 ( .A(n3689), .Y(n5843) );
  BUFX2 U326 ( .A(n3682), .Y(n5844) );
  BUFX2 U327 ( .A(n3675), .Y(n5845) );
  BUFX2 U328 ( .A(n3668), .Y(n5846) );
  BUFX2 U329 ( .A(n3655), .Y(n5847) );
  BUFX2 U330 ( .A(n3648), .Y(n5848) );
  BUFX2 U331 ( .A(n3641), .Y(n5849) );
  BUFX2 U332 ( .A(n3634), .Y(n5850) );
  BUFX2 U333 ( .A(n3621), .Y(n5851) );
  BUFX2 U334 ( .A(n3614), .Y(n5852) );
  BUFX2 U335 ( .A(n3607), .Y(n5853) );
  BUFX2 U336 ( .A(n3600), .Y(n5854) );
  BUFX2 U337 ( .A(n3587), .Y(n5855) );
  BUFX2 U338 ( .A(n3580), .Y(n5856) );
  BUFX2 U339 ( .A(n3573), .Y(n5857) );
  BUFX2 U340 ( .A(n3566), .Y(n5858) );
  BUFX2 U341 ( .A(n3553), .Y(n5859) );
  BUFX2 U342 ( .A(n3546), .Y(n5860) );
  BUFX2 U343 ( .A(n3539), .Y(n5861) );
  BUFX2 U344 ( .A(n3532), .Y(n5862) );
  BUFX2 U345 ( .A(n3519), .Y(n5863) );
  BUFX2 U346 ( .A(n3512), .Y(n5864) );
  BUFX2 U347 ( .A(n3505), .Y(n5865) );
  BUFX2 U348 ( .A(n3498), .Y(n5866) );
  BUFX2 U349 ( .A(n3485), .Y(n5867) );
  BUFX2 U350 ( .A(n3478), .Y(n5868) );
  BUFX2 U351 ( .A(n3471), .Y(n5869) );
  BUFX2 U352 ( .A(n3464), .Y(n5870) );
  BUFX2 U353 ( .A(n3451), .Y(n5871) );
  BUFX2 U354 ( .A(n3444), .Y(n5872) );
  BUFX2 U355 ( .A(n3437), .Y(n5873) );
  BUFX2 U356 ( .A(n3430), .Y(n5874) );
  BUFX2 U357 ( .A(n3417), .Y(n5875) );
  BUFX2 U358 ( .A(n3410), .Y(n5876) );
  BUFX2 U359 ( .A(n3403), .Y(n5877) );
  BUFX2 U360 ( .A(n3396), .Y(n5878) );
  BUFX2 U361 ( .A(n3383), .Y(n5879) );
  BUFX2 U362 ( .A(n3376), .Y(n5880) );
  BUFX2 U363 ( .A(n3369), .Y(n5881) );
  BUFX2 U364 ( .A(n3362), .Y(n5882) );
  BUFX2 U365 ( .A(n3349), .Y(n5883) );
  BUFX2 U366 ( .A(n3342), .Y(n5884) );
  BUFX2 U367 ( .A(n3335), .Y(n5885) );
  BUFX2 U368 ( .A(n3328), .Y(n5886) );
  BUFX2 U369 ( .A(n3315), .Y(n5887) );
  BUFX2 U370 ( .A(n3308), .Y(n5888) );
  BUFX2 U371 ( .A(n3301), .Y(n5889) );
  BUFX2 U372 ( .A(n3294), .Y(n5890) );
  BUFX2 U373 ( .A(n3281), .Y(n5891) );
  BUFX2 U374 ( .A(n3274), .Y(n5892) );
  BUFX2 U375 ( .A(n3267), .Y(n5893) );
  BUFX2 U376 ( .A(n3260), .Y(n5894) );
  BUFX2 U377 ( .A(n3247), .Y(n5895) );
  BUFX2 U378 ( .A(n3240), .Y(n5896) );
  BUFX2 U379 ( .A(n3233), .Y(n5897) );
  BUFX2 U380 ( .A(n3226), .Y(n5898) );
  BUFX2 U381 ( .A(n3213), .Y(n5899) );
  BUFX2 U382 ( .A(n3206), .Y(n5900) );
  BUFX2 U383 ( .A(n3199), .Y(n5901) );
  BUFX2 U384 ( .A(n3192), .Y(n5902) );
  BUFX2 U385 ( .A(n3179), .Y(n5903) );
  BUFX2 U386 ( .A(n3172), .Y(n5904) );
  BUFX2 U387 ( .A(n3165), .Y(n5905) );
  BUFX2 U388 ( .A(n1836), .Y(n5906) );
  BUFX2 U389 ( .A(n1823), .Y(n5907) );
  BUFX2 U390 ( .A(n1816), .Y(n5908) );
  BUFX2 U391 ( .A(n1809), .Y(n5909) );
  BUFX2 U392 ( .A(n1802), .Y(n5910) );
  BUFX2 U393 ( .A(n1789), .Y(n5911) );
  BUFX2 U394 ( .A(n1782), .Y(n5912) );
  BUFX2 U395 ( .A(n1775), .Y(n5913) );
  BUFX2 U396 ( .A(n1768), .Y(n5914) );
  BUFX2 U397 ( .A(n1755), .Y(n5915) );
  BUFX2 U398 ( .A(n1748), .Y(n5916) );
  BUFX2 U399 ( .A(n1741), .Y(n5917) );
  BUFX2 U400 ( .A(n1734), .Y(n5918) );
  BUFX2 U401 ( .A(n1721), .Y(n5919) );
  BUFX2 U402 ( .A(n1714), .Y(n5920) );
  BUFX2 U403 ( .A(n1707), .Y(n5921) );
  BUFX2 U404 ( .A(n1700), .Y(n5922) );
  BUFX2 U405 ( .A(n1687), .Y(n5923) );
  BUFX2 U406 ( .A(n1680), .Y(n5924) );
  BUFX2 U407 ( .A(n1673), .Y(n5925) );
  BUFX2 U408 ( .A(n1666), .Y(n5926) );
  BUFX2 U409 ( .A(n1653), .Y(n5927) );
  BUFX2 U410 ( .A(n1646), .Y(n5928) );
  BUFX2 U411 ( .A(n1639), .Y(n5929) );
  BUFX2 U412 ( .A(n1632), .Y(n5930) );
  BUFX2 U413 ( .A(n1619), .Y(n5931) );
  BUFX2 U414 ( .A(n1612), .Y(n5932) );
  BUFX2 U415 ( .A(n1605), .Y(n5933) );
  BUFX2 U416 ( .A(n1598), .Y(n5934) );
  BUFX2 U417 ( .A(n1585), .Y(n5935) );
  BUFX2 U418 ( .A(n1578), .Y(n5936) );
  BUFX2 U419 ( .A(n1571), .Y(n5937) );
  BUFX2 U420 ( .A(n1564), .Y(n5938) );
  BUFX2 U421 ( .A(n1551), .Y(n5939) );
  BUFX2 U422 ( .A(n1544), .Y(n5940) );
  BUFX2 U423 ( .A(n1537), .Y(n5941) );
  BUFX2 U424 ( .A(n1530), .Y(n5942) );
  BUFX2 U425 ( .A(n1517), .Y(n5943) );
  BUFX2 U426 ( .A(n1510), .Y(n5944) );
  BUFX2 U427 ( .A(n1503), .Y(n5945) );
  BUFX2 U428 ( .A(n1496), .Y(n5946) );
  BUFX2 U429 ( .A(n1483), .Y(n5947) );
  BUFX2 U430 ( .A(n1476), .Y(n5948) );
  BUFX2 U431 ( .A(n1469), .Y(n5949) );
  BUFX2 U432 ( .A(n1462), .Y(n5950) );
  BUFX2 U433 ( .A(n1449), .Y(n5951) );
  BUFX2 U434 ( .A(n1442), .Y(n5952) );
  BUFX2 U435 ( .A(n1435), .Y(n5953) );
  BUFX2 U436 ( .A(n1428), .Y(n5954) );
  BUFX2 U437 ( .A(n1415), .Y(n5955) );
  BUFX2 U438 ( .A(n1408), .Y(n5956) );
  BUFX2 U439 ( .A(n1401), .Y(n5957) );
  BUFX2 U440 ( .A(n1394), .Y(n5958) );
  BUFX2 U441 ( .A(n1380), .Y(n5959) );
  BUFX2 U442 ( .A(n1372), .Y(n5960) );
  BUFX2 U443 ( .A(n1364), .Y(n5961) );
  BUFX2 U444 ( .A(n1350), .Y(n5962) );
  BUFX2 U445 ( .A(n4067), .Y(n5963) );
  BUFX2 U446 ( .A(n4059), .Y(n5964) );
  BUFX2 U447 ( .A(n4051), .Y(n5965) );
  BUFX2 U448 ( .A(n4043), .Y(n5966) );
  BUFX2 U449 ( .A(n4030), .Y(n5967) );
  BUFX2 U450 ( .A(n4023), .Y(n5968) );
  BUFX2 U451 ( .A(n4016), .Y(n5969) );
  BUFX2 U452 ( .A(n4009), .Y(n5970) );
  BUFX2 U453 ( .A(n3996), .Y(n5971) );
  BUFX2 U454 ( .A(n3989), .Y(n5972) );
  BUFX2 U455 ( .A(n3982), .Y(n5973) );
  BUFX2 U456 ( .A(n3975), .Y(n5974) );
  BUFX2 U457 ( .A(n3962), .Y(n5975) );
  BUFX2 U458 ( .A(n3955), .Y(n5976) );
  BUFX2 U459 ( .A(n3948), .Y(n5977) );
  BUFX2 U460 ( .A(n3941), .Y(n5978) );
  BUFX2 U461 ( .A(n3928), .Y(n5979) );
  BUFX2 U462 ( .A(n3921), .Y(n5980) );
  BUFX2 U463 ( .A(n3914), .Y(n5981) );
  BUFX2 U464 ( .A(n3907), .Y(n5982) );
  BUFX2 U465 ( .A(n3894), .Y(n5983) );
  BUFX2 U466 ( .A(n3887), .Y(n5984) );
  BUFX2 U467 ( .A(n3880), .Y(n5985) );
  BUFX2 U468 ( .A(n3873), .Y(n5986) );
  BUFX2 U469 ( .A(n3860), .Y(n5987) );
  BUFX2 U470 ( .A(n3853), .Y(n5988) );
  BUFX2 U471 ( .A(n3846), .Y(n5989) );
  BUFX2 U472 ( .A(n3839), .Y(n5990) );
  BUFX2 U473 ( .A(n3826), .Y(n5991) );
  BUFX2 U474 ( .A(n3819), .Y(n5992) );
  BUFX2 U475 ( .A(n3812), .Y(n5993) );
  BUFX2 U476 ( .A(n3805), .Y(n5994) );
  BUFX2 U477 ( .A(n3792), .Y(n5995) );
  BUFX2 U478 ( .A(n3785), .Y(n5996) );
  BUFX2 U479 ( .A(n3778), .Y(n5997) );
  BUFX2 U480 ( .A(n3771), .Y(n5998) );
  BUFX2 U481 ( .A(n3758), .Y(n5999) );
  BUFX2 U482 ( .A(n3751), .Y(n6000) );
  BUFX2 U483 ( .A(n3744), .Y(n6001) );
  BUFX2 U484 ( .A(n3737), .Y(n6002) );
  BUFX2 U485 ( .A(n3724), .Y(n6003) );
  BUFX2 U486 ( .A(n3717), .Y(n6004) );
  BUFX2 U487 ( .A(n3710), .Y(n6005) );
  BUFX2 U488 ( .A(n3703), .Y(n6006) );
  BUFX2 U489 ( .A(n3690), .Y(n6007) );
  BUFX2 U490 ( .A(n3683), .Y(n6008) );
  BUFX2 U491 ( .A(n3676), .Y(n6009) );
  BUFX2 U492 ( .A(n3669), .Y(n6010) );
  BUFX2 U493 ( .A(n3656), .Y(n6011) );
  BUFX2 U494 ( .A(n3649), .Y(n6012) );
  BUFX2 U495 ( .A(n3642), .Y(n6013) );
  BUFX2 U496 ( .A(n3635), .Y(n6014) );
  BUFX2 U497 ( .A(n3622), .Y(n6015) );
  BUFX2 U498 ( .A(n3615), .Y(n6016) );
  BUFX2 U499 ( .A(n3608), .Y(n6017) );
  BUFX2 U500 ( .A(n3601), .Y(n6018) );
  BUFX2 U501 ( .A(n3588), .Y(n6019) );
  BUFX2 U502 ( .A(n3581), .Y(n6020) );
  BUFX2 U503 ( .A(n3574), .Y(n6021) );
  BUFX2 U504 ( .A(n3567), .Y(n6022) );
  BUFX2 U505 ( .A(n3554), .Y(n6023) );
  BUFX2 U506 ( .A(n3547), .Y(n6024) );
  BUFX2 U507 ( .A(n3540), .Y(n6025) );
  BUFX2 U508 ( .A(n3533), .Y(n6026) );
  BUFX2 U509 ( .A(n3520), .Y(n6027) );
  BUFX2 U510 ( .A(n3513), .Y(n6028) );
  BUFX2 U511 ( .A(n3506), .Y(n6029) );
  BUFX2 U512 ( .A(n3499), .Y(n6030) );
  BUFX2 U513 ( .A(n3486), .Y(n6031) );
  BUFX2 U514 ( .A(n3479), .Y(n6032) );
  BUFX2 U515 ( .A(n3472), .Y(n6033) );
  BUFX2 U516 ( .A(n3465), .Y(n6034) );
  BUFX2 U517 ( .A(n3452), .Y(n6035) );
  BUFX2 U518 ( .A(n3445), .Y(n6036) );
  BUFX2 U519 ( .A(n3438), .Y(n6037) );
  BUFX2 U520 ( .A(n3431), .Y(n6038) );
  BUFX2 U521 ( .A(n3418), .Y(n6039) );
  BUFX2 U522 ( .A(n3411), .Y(n6040) );
  BUFX2 U523 ( .A(n3404), .Y(n6041) );
  BUFX2 U524 ( .A(n3397), .Y(n6042) );
  BUFX2 U525 ( .A(n3384), .Y(n6043) );
  BUFX2 U526 ( .A(n3377), .Y(n6044) );
  BUFX2 U527 ( .A(n3370), .Y(n6045) );
  BUFX2 U528 ( .A(n3363), .Y(n6046) );
  BUFX2 U529 ( .A(n3350), .Y(n6047) );
  BUFX2 U530 ( .A(n3343), .Y(n6048) );
  BUFX2 U531 ( .A(n3336), .Y(n6049) );
  BUFX2 U532 ( .A(n3329), .Y(n6050) );
  BUFX2 U533 ( .A(n3316), .Y(n6051) );
  BUFX2 U534 ( .A(n3309), .Y(n6052) );
  BUFX2 U535 ( .A(n3302), .Y(n6053) );
  BUFX2 U536 ( .A(n3295), .Y(n6054) );
  BUFX2 U537 ( .A(n3282), .Y(n6055) );
  BUFX2 U538 ( .A(n3275), .Y(n6056) );
  BUFX2 U539 ( .A(n3268), .Y(n6057) );
  BUFX2 U540 ( .A(n3261), .Y(n6058) );
  BUFX2 U541 ( .A(n3248), .Y(n6059) );
  BUFX2 U542 ( .A(n3241), .Y(n6060) );
  BUFX2 U543 ( .A(n3234), .Y(n6061) );
  BUFX2 U544 ( .A(n3227), .Y(n6062) );
  BUFX2 U545 ( .A(n3214), .Y(n6063) );
  BUFX2 U546 ( .A(n3207), .Y(n6064) );
  BUFX2 U547 ( .A(n3200), .Y(n6065) );
  BUFX2 U548 ( .A(n3193), .Y(n6066) );
  BUFX2 U549 ( .A(n3180), .Y(n6067) );
  BUFX2 U550 ( .A(n3173), .Y(n6068) );
  BUFX2 U551 ( .A(n3166), .Y(n6069) );
  BUFX2 U552 ( .A(n1837), .Y(n6070) );
  BUFX2 U553 ( .A(n1824), .Y(n6071) );
  BUFX2 U554 ( .A(n1817), .Y(n6072) );
  BUFX2 U555 ( .A(n1810), .Y(n6073) );
  BUFX2 U556 ( .A(n1803), .Y(n6074) );
  BUFX2 U557 ( .A(n1790), .Y(n6075) );
  BUFX2 U558 ( .A(n1783), .Y(n6076) );
  BUFX2 U559 ( .A(n1776), .Y(n6077) );
  BUFX2 U560 ( .A(n1769), .Y(n6078) );
  BUFX2 U561 ( .A(n1756), .Y(n6079) );
  BUFX2 U562 ( .A(n1749), .Y(n6080) );
  BUFX2 U563 ( .A(n1742), .Y(n6081) );
  BUFX2 U564 ( .A(n1735), .Y(n6082) );
  BUFX2 U565 ( .A(n1722), .Y(n6083) );
  BUFX2 U566 ( .A(n1715), .Y(n6084) );
  BUFX2 U567 ( .A(n1708), .Y(n6085) );
  BUFX2 U568 ( .A(n1701), .Y(n6086) );
  BUFX2 U569 ( .A(n1688), .Y(n6087) );
  BUFX2 U570 ( .A(n1681), .Y(n6088) );
  BUFX2 U571 ( .A(n1674), .Y(n6089) );
  BUFX2 U572 ( .A(n1667), .Y(n6090) );
  BUFX2 U573 ( .A(n1654), .Y(n6091) );
  BUFX2 U574 ( .A(n1647), .Y(n6092) );
  BUFX2 U575 ( .A(n1640), .Y(n6093) );
  BUFX2 U576 ( .A(n1633), .Y(n6094) );
  BUFX2 U577 ( .A(n1620), .Y(n6095) );
  BUFX2 U578 ( .A(n1613), .Y(n6096) );
  BUFX2 U579 ( .A(n1606), .Y(n6097) );
  BUFX2 U580 ( .A(n1599), .Y(n6098) );
  BUFX2 U581 ( .A(n1586), .Y(n6099) );
  BUFX2 U582 ( .A(n1579), .Y(n6100) );
  BUFX2 U583 ( .A(n1572), .Y(n6101) );
  BUFX2 U584 ( .A(n1565), .Y(n6102) );
  BUFX2 U585 ( .A(n1552), .Y(n6103) );
  BUFX2 U586 ( .A(n1545), .Y(n6104) );
  BUFX2 U587 ( .A(n1538), .Y(n6105) );
  BUFX2 U588 ( .A(n1531), .Y(n6106) );
  BUFX2 U589 ( .A(n1518), .Y(n6107) );
  BUFX2 U590 ( .A(n1511), .Y(n6108) );
  BUFX2 U591 ( .A(n1504), .Y(n6109) );
  BUFX2 U592 ( .A(n1497), .Y(n6110) );
  BUFX2 U593 ( .A(n1484), .Y(n6111) );
  BUFX2 U594 ( .A(n1477), .Y(n6112) );
  BUFX2 U595 ( .A(n1470), .Y(n6113) );
  BUFX2 U596 ( .A(n1463), .Y(n6114) );
  BUFX2 U597 ( .A(n1450), .Y(n6115) );
  BUFX2 U598 ( .A(n1443), .Y(n6116) );
  BUFX2 U599 ( .A(n1436), .Y(n6117) );
  BUFX2 U600 ( .A(n1429), .Y(n6118) );
  BUFX2 U601 ( .A(n1416), .Y(n6119) );
  BUFX2 U602 ( .A(n1409), .Y(n6120) );
  BUFX2 U603 ( .A(n1402), .Y(n6121) );
  BUFX2 U604 ( .A(n1395), .Y(n6122) );
  BUFX2 U605 ( .A(n1381), .Y(n6123) );
  BUFX2 U606 ( .A(n1373), .Y(n6124) );
  BUFX2 U607 ( .A(n1365), .Y(n6125) );
  BUFX2 U608 ( .A(n1351), .Y(n6126) );
  BUFX2 U609 ( .A(n5502), .Y(n6127) );
  BUFX2 U610 ( .A(n4070), .Y(n6128) );
  BUFX2 U611 ( .A(n4063), .Y(n6129) );
  BUFX2 U612 ( .A(n4055), .Y(n6130) );
  BUFX2 U613 ( .A(n4047), .Y(n6131) );
  BUFX2 U614 ( .A(n4033), .Y(n6132) );
  BUFX2 U615 ( .A(n4026), .Y(n6133) );
  BUFX2 U616 ( .A(n4019), .Y(n6134) );
  BUFX2 U617 ( .A(n4012), .Y(n6135) );
  BUFX2 U618 ( .A(n3999), .Y(n6136) );
  BUFX2 U619 ( .A(n3992), .Y(n6137) );
  BUFX2 U620 ( .A(n3985), .Y(n6138) );
  BUFX2 U621 ( .A(n3978), .Y(n6139) );
  BUFX2 U622 ( .A(n3965), .Y(n6140) );
  BUFX2 U623 ( .A(n3958), .Y(n6141) );
  BUFX2 U624 ( .A(n3951), .Y(n6142) );
  BUFX2 U625 ( .A(n3944), .Y(n6143) );
  BUFX2 U626 ( .A(n3931), .Y(n6144) );
  BUFX2 U627 ( .A(n3924), .Y(n6145) );
  BUFX2 U628 ( .A(n3917), .Y(n6146) );
  BUFX2 U629 ( .A(n3910), .Y(n6147) );
  BUFX2 U630 ( .A(n3897), .Y(n6148) );
  BUFX2 U631 ( .A(n3890), .Y(n6149) );
  BUFX2 U632 ( .A(n3883), .Y(n6150) );
  BUFX2 U633 ( .A(n3876), .Y(n6151) );
  BUFX2 U634 ( .A(n3863), .Y(n6152) );
  BUFX2 U635 ( .A(n3856), .Y(n6153) );
  BUFX2 U636 ( .A(n3849), .Y(n6154) );
  BUFX2 U637 ( .A(n3842), .Y(n6155) );
  BUFX2 U638 ( .A(n3829), .Y(n6156) );
  BUFX2 U639 ( .A(n3822), .Y(n6157) );
  BUFX2 U640 ( .A(n3815), .Y(n6158) );
  BUFX2 U641 ( .A(n3808), .Y(n6159) );
  BUFX2 U642 ( .A(n3795), .Y(n6160) );
  BUFX2 U643 ( .A(n3788), .Y(n6161) );
  BUFX2 U644 ( .A(n3781), .Y(n6162) );
  BUFX2 U645 ( .A(n3774), .Y(n6163) );
  BUFX2 U646 ( .A(n3761), .Y(n6164) );
  BUFX2 U647 ( .A(n3754), .Y(n6165) );
  BUFX2 U648 ( .A(n3747), .Y(n6166) );
  BUFX2 U649 ( .A(n3740), .Y(n6167) );
  BUFX2 U650 ( .A(n3727), .Y(n6168) );
  BUFX2 U651 ( .A(n3720), .Y(n6169) );
  BUFX2 U652 ( .A(n3713), .Y(n6170) );
  BUFX2 U653 ( .A(n3706), .Y(n6171) );
  BUFX2 U654 ( .A(n3693), .Y(n6172) );
  BUFX2 U655 ( .A(n3686), .Y(n6173) );
  BUFX2 U656 ( .A(n3679), .Y(n6174) );
  BUFX2 U657 ( .A(n3672), .Y(n6175) );
  BUFX2 U658 ( .A(n3659), .Y(n6176) );
  BUFX2 U659 ( .A(n3652), .Y(n6177) );
  BUFX2 U660 ( .A(n3645), .Y(n6178) );
  BUFX2 U661 ( .A(n3638), .Y(n6179) );
  BUFX2 U662 ( .A(n3625), .Y(n6180) );
  BUFX2 U663 ( .A(n3618), .Y(n6181) );
  BUFX2 U664 ( .A(n3611), .Y(n6182) );
  BUFX2 U665 ( .A(n3604), .Y(n6183) );
  BUFX2 U666 ( .A(n3591), .Y(n6184) );
  BUFX2 U667 ( .A(n3584), .Y(n6185) );
  BUFX2 U668 ( .A(n3577), .Y(n6186) );
  BUFX2 U669 ( .A(n3570), .Y(n6187) );
  BUFX2 U670 ( .A(n3557), .Y(n6188) );
  BUFX2 U671 ( .A(n3550), .Y(n6189) );
  BUFX2 U672 ( .A(n3543), .Y(n6190) );
  BUFX2 U673 ( .A(n3536), .Y(n6191) );
  BUFX2 U674 ( .A(n3523), .Y(n6192) );
  BUFX2 U675 ( .A(n3516), .Y(n6193) );
  BUFX2 U676 ( .A(n3509), .Y(n6194) );
  BUFX2 U677 ( .A(n3502), .Y(n6195) );
  BUFX2 U678 ( .A(n3489), .Y(n6196) );
  BUFX2 U679 ( .A(n3482), .Y(n6197) );
  BUFX2 U680 ( .A(n3475), .Y(n6198) );
  BUFX2 U681 ( .A(n3468), .Y(n6199) );
  BUFX2 U682 ( .A(n3455), .Y(n6200) );
  BUFX2 U683 ( .A(n3448), .Y(n6201) );
  BUFX2 U684 ( .A(n3441), .Y(n6202) );
  BUFX2 U685 ( .A(n3434), .Y(n6203) );
  BUFX2 U686 ( .A(n3421), .Y(n6204) );
  BUFX2 U687 ( .A(n3414), .Y(n6205) );
  BUFX2 U688 ( .A(n3407), .Y(n6206) );
  BUFX2 U689 ( .A(n3400), .Y(n6207) );
  BUFX2 U690 ( .A(n3387), .Y(n6208) );
  BUFX2 U691 ( .A(n3380), .Y(n6209) );
  BUFX2 U692 ( .A(n3373), .Y(n6210) );
  BUFX2 U693 ( .A(n3366), .Y(n6211) );
  BUFX2 U694 ( .A(n3353), .Y(n6212) );
  BUFX2 U695 ( .A(n3346), .Y(n6213) );
  BUFX2 U696 ( .A(n3339), .Y(n6214) );
  BUFX2 U697 ( .A(n3332), .Y(n6215) );
  BUFX2 U698 ( .A(n3319), .Y(n6216) );
  BUFX2 U699 ( .A(n3312), .Y(n6217) );
  BUFX2 U700 ( .A(n3305), .Y(n6218) );
  BUFX2 U701 ( .A(n3298), .Y(n6219) );
  BUFX2 U702 ( .A(n3285), .Y(n6220) );
  BUFX2 U703 ( .A(n3278), .Y(n6221) );
  BUFX2 U704 ( .A(n3271), .Y(n6222) );
  BUFX2 U705 ( .A(n3264), .Y(n6223) );
  BUFX2 U706 ( .A(n3251), .Y(n6224) );
  BUFX2 U707 ( .A(n3244), .Y(n6225) );
  BUFX2 U708 ( .A(n3237), .Y(n6226) );
  BUFX2 U709 ( .A(n3230), .Y(n6227) );
  BUFX2 U710 ( .A(n3217), .Y(n6228) );
  BUFX2 U711 ( .A(n3210), .Y(n6229) );
  BUFX2 U712 ( .A(n3203), .Y(n6230) );
  BUFX2 U713 ( .A(n3196), .Y(n6231) );
  BUFX2 U714 ( .A(n3183), .Y(n6232) );
  BUFX2 U715 ( .A(n3176), .Y(n6233) );
  BUFX2 U716 ( .A(n3169), .Y(n6234) );
  BUFX2 U717 ( .A(n1840), .Y(n6235) );
  BUFX2 U718 ( .A(n1827), .Y(n6236) );
  BUFX2 U719 ( .A(n1820), .Y(n6237) );
  BUFX2 U720 ( .A(n1813), .Y(n6238) );
  BUFX2 U721 ( .A(n1806), .Y(n6239) );
  BUFX2 U722 ( .A(n1793), .Y(n6240) );
  BUFX2 U723 ( .A(n1786), .Y(n6241) );
  BUFX2 U724 ( .A(n1779), .Y(n6242) );
  BUFX2 U725 ( .A(n1772), .Y(n6243) );
  BUFX2 U726 ( .A(n1759), .Y(n6244) );
  BUFX2 U727 ( .A(n1752), .Y(n6245) );
  BUFX2 U728 ( .A(n1745), .Y(n6246) );
  BUFX2 U729 ( .A(n1738), .Y(n6247) );
  BUFX2 U730 ( .A(n1725), .Y(n6248) );
  BUFX2 U731 ( .A(n1718), .Y(n6249) );
  BUFX2 U732 ( .A(n1711), .Y(n6250) );
  BUFX2 U733 ( .A(n1704), .Y(n6251) );
  BUFX2 U734 ( .A(n1691), .Y(n6252) );
  BUFX2 U735 ( .A(n1684), .Y(n6253) );
  BUFX2 U736 ( .A(n1677), .Y(n6254) );
  BUFX2 U737 ( .A(n1670), .Y(n6255) );
  BUFX2 U738 ( .A(n1657), .Y(n6256) );
  BUFX2 U739 ( .A(n1650), .Y(n6257) );
  BUFX2 U740 ( .A(n1643), .Y(n6258) );
  BUFX2 U741 ( .A(n1636), .Y(n6259) );
  BUFX2 U742 ( .A(n1623), .Y(n6260) );
  BUFX2 U743 ( .A(n1616), .Y(n6261) );
  BUFX2 U744 ( .A(n1609), .Y(n6262) );
  BUFX2 U745 ( .A(n1602), .Y(n6263) );
  BUFX2 U746 ( .A(n1589), .Y(n6264) );
  BUFX2 U747 ( .A(n1582), .Y(n6265) );
  BUFX2 U748 ( .A(n1575), .Y(n6266) );
  BUFX2 U749 ( .A(n1568), .Y(n6267) );
  BUFX2 U750 ( .A(n1555), .Y(n6268) );
  BUFX2 U751 ( .A(n1548), .Y(n6269) );
  BUFX2 U752 ( .A(n1541), .Y(n6270) );
  BUFX2 U753 ( .A(n1534), .Y(n6271) );
  BUFX2 U754 ( .A(n1521), .Y(n6272) );
  BUFX2 U755 ( .A(n1514), .Y(n6273) );
  BUFX2 U756 ( .A(n1507), .Y(n6274) );
  BUFX2 U757 ( .A(n1500), .Y(n6275) );
  BUFX2 U758 ( .A(n1487), .Y(n6276) );
  BUFX2 U759 ( .A(n1480), .Y(n6277) );
  BUFX2 U760 ( .A(n1473), .Y(n6278) );
  BUFX2 U761 ( .A(n1466), .Y(n6279) );
  BUFX2 U762 ( .A(n1453), .Y(n6280) );
  BUFX2 U763 ( .A(n1446), .Y(n6281) );
  BUFX2 U764 ( .A(n1439), .Y(n6282) );
  BUFX2 U765 ( .A(n1432), .Y(n6283) );
  BUFX2 U766 ( .A(n1419), .Y(n6284) );
  BUFX2 U767 ( .A(n1412), .Y(n6285) );
  BUFX2 U768 ( .A(n1405), .Y(n6286) );
  BUFX2 U769 ( .A(n1398), .Y(n6287) );
  BUFX2 U770 ( .A(n1385), .Y(n6288) );
  BUFX2 U771 ( .A(n1377), .Y(n6289) );
  BUFX2 U772 ( .A(n1369), .Y(n6290) );
  BUFX2 U773 ( .A(n1356), .Y(n6291) );
  AND2X1 U774 ( .A(n1382), .B(n8428), .Y(n4079) );
  INVX1 U775 ( .A(n4079), .Y(n6292) );
  AND2X1 U776 ( .A(data_out[12]), .B(n4082), .Y(n4036) );
  INVX1 U777 ( .A(n4036), .Y(n6293) );
  AND2X1 U778 ( .A(data_out[13]), .B(n4082), .Y(n4002) );
  INVX1 U779 ( .A(n4002), .Y(n6294) );
  AND2X1 U780 ( .A(data_out[14]), .B(n4082), .Y(n3968) );
  INVX1 U781 ( .A(n3968), .Y(n6295) );
  AND2X1 U782 ( .A(data_out[15]), .B(n4082), .Y(n3934) );
  INVX1 U783 ( .A(n3934), .Y(n6296) );
  AND2X1 U784 ( .A(data_out[16]), .B(n4082), .Y(n3900) );
  INVX1 U785 ( .A(n3900), .Y(n6297) );
  AND2X1 U786 ( .A(data_out[17]), .B(n4082), .Y(n3866) );
  INVX1 U787 ( .A(n3866), .Y(n6298) );
  AND2X1 U788 ( .A(data_out[18]), .B(n4082), .Y(n3832) );
  INVX1 U789 ( .A(n3832), .Y(n6299) );
  AND2X1 U790 ( .A(data_out[19]), .B(n4082), .Y(n3798) );
  INVX1 U791 ( .A(n3798), .Y(n6300) );
  AND2X1 U792 ( .A(data_out[20]), .B(n4082), .Y(n3764) );
  INVX1 U793 ( .A(n3764), .Y(n6301) );
  AND2X1 U794 ( .A(data_out[21]), .B(n4082), .Y(n3730) );
  INVX1 U795 ( .A(n3730), .Y(n6302) );
  AND2X1 U796 ( .A(data_out[22]), .B(n4082), .Y(n3696) );
  INVX1 U797 ( .A(n3696), .Y(n6303) );
  AND2X1 U798 ( .A(data_out[23]), .B(n4082), .Y(n3662) );
  INVX1 U799 ( .A(n3662), .Y(n6304) );
  AND2X1 U800 ( .A(data_out[37]), .B(n4082), .Y(n3628) );
  INVX1 U801 ( .A(n3628), .Y(n6305) );
  AND2X1 U802 ( .A(data_out[40]), .B(n4082), .Y(n3594) );
  INVX1 U803 ( .A(n3594), .Y(n6306) );
  AND2X1 U804 ( .A(data_out[0]), .B(n4082), .Y(n3560) );
  INVX1 U805 ( .A(n3560), .Y(n6307) );
  AND2X1 U806 ( .A(data_out[2]), .B(n4082), .Y(n3526) );
  INVX1 U807 ( .A(n3526), .Y(n6308) );
  AND2X1 U808 ( .A(data_out[4]), .B(n4082), .Y(n3492) );
  INVX1 U809 ( .A(n3492), .Y(n6309) );
  AND2X1 U810 ( .A(data_out[6]), .B(n4082), .Y(n3458) );
  INVX1 U811 ( .A(n3458), .Y(n6310) );
  AND2X1 U812 ( .A(data_out[8]), .B(n4082), .Y(n3424) );
  INVX1 U813 ( .A(n3424), .Y(n6311) );
  AND2X1 U814 ( .A(data_out[10]), .B(n4082), .Y(n3390) );
  INVX1 U815 ( .A(n3390), .Y(n6312) );
  AND2X1 U816 ( .A(data_out[38]), .B(n4082), .Y(n3356) );
  INVX1 U817 ( .A(n3356), .Y(n6313) );
  AND2X1 U818 ( .A(data_out[24]), .B(n4082), .Y(n3322) );
  INVX1 U819 ( .A(n3322), .Y(n6314) );
  AND2X1 U820 ( .A(data_out[25]), .B(n4082), .Y(n3288) );
  INVX1 U821 ( .A(n3288), .Y(n6315) );
  AND2X1 U822 ( .A(data_out[26]), .B(n4082), .Y(n3254) );
  INVX1 U823 ( .A(n3254), .Y(n6316) );
  AND2X1 U824 ( .A(data_out[27]), .B(n4082), .Y(n3220) );
  INVX1 U825 ( .A(n3220), .Y(n6317) );
  AND2X1 U826 ( .A(data_out[28]), .B(n4082), .Y(n3186) );
  INVX1 U827 ( .A(n3186), .Y(n6318) );
  AND2X1 U828 ( .A(data_out[29]), .B(n4082), .Y(n1830) );
  INVX1 U829 ( .A(n1830), .Y(n6319) );
  AND2X1 U830 ( .A(data_out[30]), .B(n4082), .Y(n1796) );
  INVX1 U831 ( .A(n1796), .Y(n6320) );
  AND2X1 U832 ( .A(data_out[31]), .B(n4082), .Y(n1762) );
  INVX1 U833 ( .A(n1762), .Y(n6321) );
  AND2X1 U834 ( .A(data_out[32]), .B(n4082), .Y(n1728) );
  INVX1 U835 ( .A(n1728), .Y(n6322) );
  AND2X1 U836 ( .A(data_out[33]), .B(n4082), .Y(n1694) );
  INVX1 U837 ( .A(n1694), .Y(n6323) );
  AND2X1 U838 ( .A(data_out[34]), .B(n4082), .Y(n1660) );
  INVX1 U839 ( .A(n1660), .Y(n6324) );
  AND2X1 U840 ( .A(data_out[35]), .B(n4082), .Y(n1626) );
  INVX1 U841 ( .A(n1626), .Y(n6325) );
  AND2X1 U842 ( .A(data_out[36]), .B(n4082), .Y(n1592) );
  INVX1 U843 ( .A(n1592), .Y(n6326) );
  AND2X1 U844 ( .A(data_out[39]), .B(n4082), .Y(n1558) );
  INVX1 U845 ( .A(n1558), .Y(n6327) );
  AND2X1 U846 ( .A(data_out[1]), .B(n4082), .Y(n1524) );
  INVX1 U847 ( .A(n1524), .Y(n6328) );
  AND2X1 U848 ( .A(data_out[3]), .B(n4082), .Y(n1490) );
  INVX1 U849 ( .A(n1490), .Y(n6329) );
  AND2X1 U850 ( .A(data_out[5]), .B(n4082), .Y(n1456) );
  INVX1 U851 ( .A(n1456), .Y(n6330) );
  AND2X1 U852 ( .A(data_out[7]), .B(n4082), .Y(n1422) );
  INVX1 U853 ( .A(n1422), .Y(n6331) );
  AND2X1 U854 ( .A(data_out[9]), .B(n4082), .Y(n1388) );
  INVX1 U855 ( .A(n1388), .Y(n6332) );
  AND2X1 U856 ( .A(data_out[11]), .B(n4082), .Y(n1344) );
  INVX1 U857 ( .A(n1344), .Y(n6333) );
  BUFX2 U858 ( .A(n4087), .Y(n6334) );
  AND2X1 U859 ( .A(n1361), .B(n9326), .Y(n4071) );
  INVX1 U860 ( .A(n4071), .Y(n6335) );
  AND2X1 U861 ( .A(n8430), .B(n9203), .Y(n4068) );
  INVX1 U862 ( .A(n4068), .Y(n6336) );
  AND2X1 U863 ( .A(n1361), .B(n9654), .Y(n4064) );
  INVX1 U864 ( .A(n4064), .Y(n6337) );
  AND2X1 U865 ( .A(n8429), .B(n9531), .Y(n4060) );
  INVX1 U866 ( .A(n4060), .Y(n6338) );
  AND2X1 U867 ( .A(n1361), .B(n8670), .Y(n4056) );
  INVX1 U868 ( .A(n4056), .Y(n6339) );
  AND2X1 U869 ( .A(n8429), .B(n8547), .Y(n4052) );
  INVX1 U870 ( .A(n4052), .Y(n6340) );
  AND2X1 U871 ( .A(n1361), .B(n8998), .Y(n4048) );
  INVX1 U872 ( .A(n4048), .Y(n6341) );
  AND2X1 U873 ( .A(n8429), .B(n8875), .Y(n4044) );
  INVX1 U874 ( .A(n4044), .Y(n6342) );
  AND2X1 U875 ( .A(n1361), .B(n9325), .Y(n4034) );
  INVX1 U876 ( .A(n4034), .Y(n6343) );
  AND2X1 U877 ( .A(n8428), .B(n9202), .Y(n4031) );
  INVX1 U878 ( .A(n4031), .Y(n6344) );
  AND2X1 U879 ( .A(n1361), .B(n9653), .Y(n4027) );
  INVX1 U880 ( .A(n4027), .Y(n6345) );
  AND2X1 U881 ( .A(n8430), .B(n9530), .Y(n4024) );
  INVX1 U882 ( .A(n4024), .Y(n6346) );
  AND2X1 U883 ( .A(n1361), .B(n8669), .Y(n4020) );
  INVX1 U884 ( .A(n4020), .Y(n6347) );
  AND2X1 U885 ( .A(n8430), .B(n8546), .Y(n4017) );
  INVX1 U886 ( .A(n4017), .Y(n6348) );
  AND2X1 U887 ( .A(n1361), .B(n8997), .Y(n4013) );
  INVX1 U888 ( .A(n4013), .Y(n6349) );
  AND2X1 U889 ( .A(n8428), .B(n8874), .Y(n4010) );
  INVX1 U890 ( .A(n4010), .Y(n6350) );
  AND2X1 U891 ( .A(n8462), .B(n9324), .Y(n4000) );
  INVX1 U892 ( .A(n4000), .Y(n6351) );
  AND2X1 U893 ( .A(n8428), .B(n9201), .Y(n3997) );
  INVX1 U894 ( .A(n3997), .Y(n6352) );
  AND2X1 U895 ( .A(n8462), .B(n9652), .Y(n3993) );
  INVX1 U896 ( .A(n3993), .Y(n6353) );
  AND2X1 U897 ( .A(n8427), .B(n9529), .Y(n3990) );
  INVX1 U898 ( .A(n3990), .Y(n6354) );
  AND2X1 U899 ( .A(n8462), .B(n8668), .Y(n3986) );
  INVX1 U900 ( .A(n3986), .Y(n6355) );
  AND2X1 U901 ( .A(n8428), .B(n8545), .Y(n3983) );
  INVX1 U902 ( .A(n3983), .Y(n6356) );
  AND2X1 U903 ( .A(n8462), .B(n8996), .Y(n3979) );
  INVX1 U904 ( .A(n3979), .Y(n6357) );
  AND2X1 U905 ( .A(n8427), .B(n8873), .Y(n3976) );
  INVX1 U906 ( .A(n3976), .Y(n6358) );
  AND2X1 U907 ( .A(n8462), .B(n9323), .Y(n3966) );
  INVX1 U908 ( .A(n3966), .Y(n6359) );
  AND2X1 U909 ( .A(n8430), .B(n9200), .Y(n3963) );
  INVX1 U910 ( .A(n3963), .Y(n6360) );
  AND2X1 U911 ( .A(n8462), .B(n9651), .Y(n3959) );
  INVX1 U912 ( .A(n3959), .Y(n6361) );
  AND2X1 U913 ( .A(n8430), .B(n9528), .Y(n3956) );
  INVX1 U914 ( .A(n3956), .Y(n6362) );
  AND2X1 U915 ( .A(n8462), .B(n8667), .Y(n3952) );
  INVX1 U916 ( .A(n3952), .Y(n6363) );
  AND2X1 U917 ( .A(n8430), .B(n8544), .Y(n3949) );
  INVX1 U918 ( .A(n3949), .Y(n6364) );
  AND2X1 U919 ( .A(n8462), .B(n8995), .Y(n3945) );
  INVX1 U920 ( .A(n3945), .Y(n6365) );
  AND2X1 U921 ( .A(n8430), .B(n8872), .Y(n3942) );
  INVX1 U922 ( .A(n3942), .Y(n6366) );
  AND2X1 U923 ( .A(n8462), .B(n9322), .Y(n3932) );
  INVX1 U924 ( .A(n3932), .Y(n6367) );
  AND2X1 U925 ( .A(n8430), .B(n9199), .Y(n3929) );
  INVX1 U926 ( .A(n3929), .Y(n6368) );
  AND2X1 U927 ( .A(n8462), .B(n9650), .Y(n3925) );
  INVX1 U928 ( .A(n3925), .Y(n6369) );
  AND2X1 U929 ( .A(n8430), .B(n9527), .Y(n3922) );
  INVX1 U930 ( .A(n3922), .Y(n6370) );
  AND2X1 U931 ( .A(n8462), .B(n8666), .Y(n3918) );
  INVX1 U932 ( .A(n3918), .Y(n6371) );
  AND2X1 U933 ( .A(n8430), .B(n8543), .Y(n3915) );
  INVX1 U934 ( .A(n3915), .Y(n6372) );
  AND2X1 U935 ( .A(n8462), .B(n8994), .Y(n3911) );
  INVX1 U936 ( .A(n3911), .Y(n6373) );
  AND2X1 U937 ( .A(n8430), .B(n8871), .Y(n3908) );
  INVX1 U938 ( .A(n3908), .Y(n6374) );
  AND2X1 U939 ( .A(n8461), .B(n9321), .Y(n3898) );
  INVX1 U940 ( .A(n3898), .Y(n6375) );
  AND2X1 U941 ( .A(n8430), .B(n9198), .Y(n3895) );
  INVX1 U942 ( .A(n3895), .Y(n6376) );
  AND2X1 U943 ( .A(n8461), .B(n9649), .Y(n3891) );
  INVX1 U944 ( .A(n3891), .Y(n6377) );
  AND2X1 U945 ( .A(n8430), .B(n9526), .Y(n3888) );
  INVX1 U946 ( .A(n3888), .Y(n6378) );
  AND2X1 U947 ( .A(n8461), .B(n8665), .Y(n3884) );
  INVX1 U948 ( .A(n3884), .Y(n6379) );
  AND2X1 U949 ( .A(n8430), .B(n8542), .Y(n3881) );
  INVX1 U950 ( .A(n3881), .Y(n6380) );
  AND2X1 U951 ( .A(n8461), .B(n8993), .Y(n3877) );
  INVX1 U952 ( .A(n3877), .Y(n6381) );
  AND2X1 U953 ( .A(n8430), .B(n8870), .Y(n3874) );
  INVX1 U954 ( .A(n3874), .Y(n6382) );
  AND2X1 U955 ( .A(n8461), .B(n9320), .Y(n3864) );
  INVX1 U956 ( .A(n3864), .Y(n6383) );
  AND2X1 U957 ( .A(n8430), .B(n9197), .Y(n3861) );
  INVX1 U958 ( .A(n3861), .Y(n6384) );
  AND2X1 U959 ( .A(n8461), .B(n9648), .Y(n3857) );
  INVX1 U960 ( .A(n3857), .Y(n6385) );
  AND2X1 U961 ( .A(n8430), .B(n9525), .Y(n3854) );
  INVX1 U962 ( .A(n3854), .Y(n6386) );
  AND2X1 U963 ( .A(n8461), .B(n8664), .Y(n3850) );
  INVX1 U964 ( .A(n3850), .Y(n6387) );
  AND2X1 U965 ( .A(n8430), .B(n8541), .Y(n3847) );
  INVX1 U966 ( .A(n3847), .Y(n6388) );
  AND2X1 U967 ( .A(n8461), .B(n8992), .Y(n3843) );
  INVX1 U968 ( .A(n3843), .Y(n6389) );
  AND2X1 U969 ( .A(n8430), .B(n8869), .Y(n3840) );
  INVX1 U970 ( .A(n3840), .Y(n6390) );
  AND2X1 U971 ( .A(n8461), .B(n9319), .Y(n3830) );
  INVX1 U972 ( .A(n3830), .Y(n6391) );
  AND2X1 U973 ( .A(n8430), .B(n9196), .Y(n3827) );
  INVX1 U974 ( .A(n3827), .Y(n6392) );
  AND2X1 U975 ( .A(n8461), .B(n9647), .Y(n3823) );
  INVX1 U976 ( .A(n3823), .Y(n6393) );
  AND2X1 U977 ( .A(n8429), .B(n9524), .Y(n3820) );
  INVX1 U978 ( .A(n3820), .Y(n6394) );
  AND2X1 U979 ( .A(n8461), .B(n8663), .Y(n3816) );
  INVX1 U980 ( .A(n3816), .Y(n6395) );
  AND2X1 U981 ( .A(n8429), .B(n8540), .Y(n3813) );
  INVX1 U982 ( .A(n3813), .Y(n6396) );
  AND2X1 U983 ( .A(n8461), .B(n8991), .Y(n3809) );
  INVX1 U984 ( .A(n3809), .Y(n6397) );
  AND2X1 U985 ( .A(n8429), .B(n8868), .Y(n3806) );
  INVX1 U986 ( .A(n3806), .Y(n6398) );
  AND2X1 U987 ( .A(n8460), .B(n9318), .Y(n3796) );
  INVX1 U988 ( .A(n3796), .Y(n6399) );
  AND2X1 U989 ( .A(n8429), .B(n9195), .Y(n3793) );
  INVX1 U990 ( .A(n3793), .Y(n6400) );
  AND2X1 U991 ( .A(n8460), .B(n9646), .Y(n3789) );
  INVX1 U992 ( .A(n3789), .Y(n6401) );
  AND2X1 U993 ( .A(n8429), .B(n9523), .Y(n3786) );
  INVX1 U994 ( .A(n3786), .Y(n6402) );
  AND2X1 U995 ( .A(n8460), .B(n8662), .Y(n3782) );
  INVX1 U996 ( .A(n3782), .Y(n6403) );
  AND2X1 U997 ( .A(n8429), .B(n8539), .Y(n3779) );
  INVX1 U998 ( .A(n3779), .Y(n6404) );
  AND2X1 U999 ( .A(n8460), .B(n8990), .Y(n3775) );
  INVX1 U1000 ( .A(n3775), .Y(n6405) );
  AND2X1 U1001 ( .A(n8429), .B(n8867), .Y(n3772) );
  INVX1 U1002 ( .A(n3772), .Y(n6406) );
  AND2X1 U1003 ( .A(n8460), .B(n9317), .Y(n3762) );
  INVX1 U1004 ( .A(n3762), .Y(n6407) );
  AND2X1 U1005 ( .A(n8429), .B(n9194), .Y(n3759) );
  INVX1 U1006 ( .A(n3759), .Y(n6408) );
  AND2X1 U1007 ( .A(n8460), .B(n9645), .Y(n3755) );
  INVX1 U1008 ( .A(n3755), .Y(n6409) );
  AND2X1 U1009 ( .A(n8429), .B(n9522), .Y(n3752) );
  INVX1 U1010 ( .A(n3752), .Y(n6410) );
  AND2X1 U1011 ( .A(n8460), .B(n8661), .Y(n3748) );
  INVX1 U1012 ( .A(n3748), .Y(n6411) );
  AND2X1 U1013 ( .A(n8429), .B(n8538), .Y(n3745) );
  INVX1 U1014 ( .A(n3745), .Y(n6412) );
  AND2X1 U1015 ( .A(n8460), .B(n8989), .Y(n3741) );
  INVX1 U1016 ( .A(n3741), .Y(n6413) );
  AND2X1 U1017 ( .A(n8429), .B(n8866), .Y(n3738) );
  INVX1 U1018 ( .A(n3738), .Y(n6414) );
  AND2X1 U1019 ( .A(n8460), .B(n9316), .Y(n3728) );
  INVX1 U1020 ( .A(n3728), .Y(n6415) );
  AND2X1 U1021 ( .A(n8429), .B(n9193), .Y(n3725) );
  INVX1 U1022 ( .A(n3725), .Y(n6416) );
  AND2X1 U1023 ( .A(n8460), .B(n9644), .Y(n3721) );
  INVX1 U1024 ( .A(n3721), .Y(n6417) );
  AND2X1 U1025 ( .A(n8429), .B(n9521), .Y(n3718) );
  INVX1 U1026 ( .A(n3718), .Y(n6418) );
  AND2X1 U1027 ( .A(n8460), .B(n8660), .Y(n3714) );
  INVX1 U1028 ( .A(n3714), .Y(n6419) );
  AND2X1 U1029 ( .A(n8429), .B(n8537), .Y(n3711) );
  INVX1 U1030 ( .A(n3711), .Y(n6420) );
  AND2X1 U1031 ( .A(n8460), .B(n8988), .Y(n3707) );
  INVX1 U1032 ( .A(n3707), .Y(n6421) );
  AND2X1 U1033 ( .A(n8429), .B(n8865), .Y(n3704) );
  INVX1 U1034 ( .A(n3704), .Y(n6422) );
  AND2X1 U1035 ( .A(n8459), .B(n9315), .Y(n3694) );
  INVX1 U1036 ( .A(n3694), .Y(n6423) );
  AND2X1 U1037 ( .A(n8429), .B(n9192), .Y(n3691) );
  INVX1 U1038 ( .A(n3691), .Y(n6424) );
  AND2X1 U1039 ( .A(n8459), .B(n9643), .Y(n3687) );
  INVX1 U1040 ( .A(n3687), .Y(n6425) );
  AND2X1 U1041 ( .A(n8429), .B(n9520), .Y(n3684) );
  INVX1 U1042 ( .A(n3684), .Y(n6426) );
  AND2X1 U1043 ( .A(n8459), .B(n8659), .Y(n3680) );
  INVX1 U1044 ( .A(n3680), .Y(n6427) );
  AND2X1 U1045 ( .A(n8427), .B(n8536), .Y(n3677) );
  INVX1 U1046 ( .A(n3677), .Y(n6428) );
  AND2X1 U1047 ( .A(n8459), .B(n8987), .Y(n3673) );
  INVX1 U1048 ( .A(n3673), .Y(n6429) );
  AND2X1 U1049 ( .A(n8428), .B(n8864), .Y(n3670) );
  INVX1 U1050 ( .A(n3670), .Y(n6430) );
  AND2X1 U1051 ( .A(n8459), .B(n9301), .Y(n3660) );
  INVX1 U1052 ( .A(n3660), .Y(n6431) );
  AND2X1 U1053 ( .A(n8428), .B(n9178), .Y(n3657) );
  INVX1 U1054 ( .A(n3657), .Y(n6432) );
  AND2X1 U1055 ( .A(n8459), .B(n9629), .Y(n3653) );
  INVX1 U1056 ( .A(n3653), .Y(n6433) );
  AND2X1 U1057 ( .A(n8427), .B(n9506), .Y(n3650) );
  INVX1 U1058 ( .A(n3650), .Y(n6434) );
  AND2X1 U1059 ( .A(n8459), .B(n8645), .Y(n3646) );
  INVX1 U1060 ( .A(n3646), .Y(n6435) );
  AND2X1 U1061 ( .A(n8428), .B(n8522), .Y(n3643) );
  INVX1 U1062 ( .A(n3643), .Y(n6436) );
  AND2X1 U1063 ( .A(n8459), .B(n8973), .Y(n3639) );
  INVX1 U1064 ( .A(n3639), .Y(n6437) );
  AND2X1 U1065 ( .A(n8429), .B(n8850), .Y(n3636) );
  INVX1 U1066 ( .A(n3636), .Y(n6438) );
  AND2X1 U1067 ( .A(n8459), .B(n9298), .Y(n3626) );
  INVX1 U1068 ( .A(n3626), .Y(n6439) );
  AND2X1 U1069 ( .A(n8430), .B(n9175), .Y(n3623) );
  INVX1 U1070 ( .A(n3623), .Y(n6440) );
  AND2X1 U1071 ( .A(n8459), .B(n9626), .Y(n3619) );
  INVX1 U1072 ( .A(n3619), .Y(n6441) );
  AND2X1 U1073 ( .A(n8429), .B(n9503), .Y(n3616) );
  INVX1 U1074 ( .A(n3616), .Y(n6442) );
  AND2X1 U1075 ( .A(n8459), .B(n8642), .Y(n3612) );
  INVX1 U1076 ( .A(n3612), .Y(n6443) );
  AND2X1 U1077 ( .A(n8428), .B(n8519), .Y(n3609) );
  INVX1 U1078 ( .A(n3609), .Y(n6444) );
  AND2X1 U1079 ( .A(n8459), .B(n8970), .Y(n3605) );
  INVX1 U1080 ( .A(n3605), .Y(n6445) );
  AND2X1 U1081 ( .A(n8430), .B(n8847), .Y(n3602) );
  INVX1 U1082 ( .A(n3602), .Y(n6446) );
  AND2X1 U1083 ( .A(n8458), .B(n9338), .Y(n3592) );
  INVX1 U1084 ( .A(n3592), .Y(n6447) );
  AND2X1 U1085 ( .A(n8429), .B(n9215), .Y(n3589) );
  INVX1 U1086 ( .A(n3589), .Y(n6448) );
  AND2X1 U1087 ( .A(n8458), .B(n9666), .Y(n3585) );
  INVX1 U1088 ( .A(n3585), .Y(n6449) );
  AND2X1 U1089 ( .A(n8430), .B(n9543), .Y(n3582) );
  INVX1 U1090 ( .A(n3582), .Y(n6450) );
  AND2X1 U1091 ( .A(n8458), .B(n8682), .Y(n3578) );
  INVX1 U1092 ( .A(n3578), .Y(n6451) );
  AND2X1 U1093 ( .A(n8429), .B(n8559), .Y(n3575) );
  INVX1 U1094 ( .A(n3575), .Y(n6452) );
  AND2X1 U1095 ( .A(n8458), .B(n9010), .Y(n3571) );
  INVX1 U1096 ( .A(n3571), .Y(n6453) );
  AND2X1 U1097 ( .A(n8429), .B(n8887), .Y(n3568) );
  INVX1 U1098 ( .A(n3568), .Y(n6454) );
  AND2X1 U1099 ( .A(n8458), .B(n9336), .Y(n3558) );
  INVX1 U1100 ( .A(n3558), .Y(n6455) );
  AND2X1 U1101 ( .A(n8430), .B(n9213), .Y(n3555) );
  INVX1 U1102 ( .A(n3555), .Y(n6456) );
  AND2X1 U1103 ( .A(n8458), .B(n9664), .Y(n3551) );
  INVX1 U1104 ( .A(n3551), .Y(n6457) );
  AND2X1 U1105 ( .A(n8427), .B(n9541), .Y(n3548) );
  INVX1 U1106 ( .A(n3548), .Y(n6458) );
  AND2X1 U1107 ( .A(n8458), .B(n8680), .Y(n3544) );
  INVX1 U1108 ( .A(n3544), .Y(n6459) );
  AND2X1 U1109 ( .A(n8430), .B(n8557), .Y(n3541) );
  INVX1 U1110 ( .A(n3541), .Y(n6460) );
  AND2X1 U1111 ( .A(n8458), .B(n9008), .Y(n3537) );
  INVX1 U1112 ( .A(n3537), .Y(n6461) );
  AND2X1 U1113 ( .A(n8428), .B(n8885), .Y(n3534) );
  INVX1 U1114 ( .A(n3534), .Y(n6462) );
  AND2X1 U1115 ( .A(n8458), .B(n9334), .Y(n3524) );
  INVX1 U1116 ( .A(n3524), .Y(n6463) );
  AND2X1 U1117 ( .A(n8427), .B(n9211), .Y(n3521) );
  INVX1 U1118 ( .A(n3521), .Y(n6464) );
  AND2X1 U1119 ( .A(n8458), .B(n9662), .Y(n3517) );
  INVX1 U1120 ( .A(n3517), .Y(n6465) );
  AND2X1 U1121 ( .A(n8429), .B(n9539), .Y(n3514) );
  INVX1 U1122 ( .A(n3514), .Y(n6466) );
  AND2X1 U1123 ( .A(n8458), .B(n8678), .Y(n3510) );
  INVX1 U1124 ( .A(n3510), .Y(n6467) );
  AND2X1 U1125 ( .A(n8430), .B(n8555), .Y(n3507) );
  INVX1 U1126 ( .A(n3507), .Y(n6468) );
  AND2X1 U1127 ( .A(n8458), .B(n9006), .Y(n3503) );
  INVX1 U1128 ( .A(n3503), .Y(n6469) );
  AND2X1 U1129 ( .A(n8430), .B(n8883), .Y(n3500) );
  INVX1 U1130 ( .A(n3500), .Y(n6470) );
  AND2X1 U1131 ( .A(n8457), .B(n9332), .Y(n3490) );
  INVX1 U1132 ( .A(n3490), .Y(n6471) );
  AND2X1 U1133 ( .A(n8430), .B(n9209), .Y(n3487) );
  INVX1 U1134 ( .A(n3487), .Y(n6472) );
  AND2X1 U1135 ( .A(n8457), .B(n9660), .Y(n3483) );
  INVX1 U1136 ( .A(n3483), .Y(n6473) );
  AND2X1 U1137 ( .A(n8430), .B(n9537), .Y(n3480) );
  INVX1 U1138 ( .A(n3480), .Y(n6474) );
  AND2X1 U1139 ( .A(n8457), .B(n8676), .Y(n3476) );
  INVX1 U1140 ( .A(n3476), .Y(n6475) );
  AND2X1 U1141 ( .A(n8429), .B(n8553), .Y(n3473) );
  INVX1 U1142 ( .A(n3473), .Y(n6476) );
  AND2X1 U1143 ( .A(n8457), .B(n9004), .Y(n3469) );
  INVX1 U1144 ( .A(n3469), .Y(n6477) );
  AND2X1 U1145 ( .A(n8429), .B(n8881), .Y(n3466) );
  INVX1 U1146 ( .A(n3466), .Y(n6478) );
  AND2X1 U1147 ( .A(n8457), .B(n9330), .Y(n3456) );
  INVX1 U1148 ( .A(n3456), .Y(n6479) );
  AND2X1 U1149 ( .A(n8429), .B(n9207), .Y(n3453) );
  INVX1 U1150 ( .A(n3453), .Y(n6480) );
  AND2X1 U1151 ( .A(n8457), .B(n9658), .Y(n3449) );
  INVX1 U1152 ( .A(n3449), .Y(n6481) );
  AND2X1 U1153 ( .A(n8427), .B(n9535), .Y(n3446) );
  INVX1 U1154 ( .A(n3446), .Y(n6482) );
  AND2X1 U1155 ( .A(n8457), .B(n8674), .Y(n3442) );
  INVX1 U1156 ( .A(n3442), .Y(n6483) );
  AND2X1 U1157 ( .A(n8430), .B(n8551), .Y(n3439) );
  INVX1 U1158 ( .A(n3439), .Y(n6484) );
  AND2X1 U1159 ( .A(n8457), .B(n9002), .Y(n3435) );
  INVX1 U1160 ( .A(n3435), .Y(n6485) );
  AND2X1 U1161 ( .A(n8430), .B(n8879), .Y(n3432) );
  INVX1 U1162 ( .A(n3432), .Y(n6486) );
  AND2X1 U1163 ( .A(n8457), .B(n9328), .Y(n3422) );
  INVX1 U1164 ( .A(n3422), .Y(n6487) );
  AND2X1 U1165 ( .A(n8430), .B(n9205), .Y(n3419) );
  INVX1 U1166 ( .A(n3419), .Y(n6488) );
  AND2X1 U1167 ( .A(n8457), .B(n9656), .Y(n3415) );
  INVX1 U1168 ( .A(n3415), .Y(n6489) );
  AND2X1 U1169 ( .A(n8428), .B(n9533), .Y(n3412) );
  INVX1 U1170 ( .A(n3412), .Y(n6490) );
  AND2X1 U1171 ( .A(n8457), .B(n8672), .Y(n3408) );
  INVX1 U1172 ( .A(n3408), .Y(n6491) );
  AND2X1 U1173 ( .A(n8427), .B(n8549), .Y(n3405) );
  INVX1 U1174 ( .A(n3405), .Y(n6492) );
  AND2X1 U1175 ( .A(n8457), .B(n9000), .Y(n3401) );
  INVX1 U1176 ( .A(n3401), .Y(n6493) );
  AND2X1 U1177 ( .A(n8427), .B(n8877), .Y(n3398) );
  INVX1 U1178 ( .A(n3398), .Y(n6494) );
  AND2X1 U1179 ( .A(n8456), .B(n9300), .Y(n3388) );
  INVX1 U1180 ( .A(n3388), .Y(n6495) );
  AND2X1 U1181 ( .A(n8428), .B(n9177), .Y(n3385) );
  INVX1 U1182 ( .A(n3385), .Y(n6496) );
  AND2X1 U1183 ( .A(n8456), .B(n9628), .Y(n3381) );
  INVX1 U1184 ( .A(n3381), .Y(n6497) );
  AND2X1 U1185 ( .A(n8429), .B(n9505), .Y(n3378) );
  INVX1 U1186 ( .A(n3378), .Y(n6498) );
  AND2X1 U1187 ( .A(n8456), .B(n8644), .Y(n3374) );
  INVX1 U1188 ( .A(n3374), .Y(n6499) );
  AND2X1 U1189 ( .A(n8429), .B(n8521), .Y(n3371) );
  INVX1 U1190 ( .A(n3371), .Y(n6500) );
  AND2X1 U1191 ( .A(n8456), .B(n8972), .Y(n3367) );
  INVX1 U1192 ( .A(n3367), .Y(n6501) );
  AND2X1 U1193 ( .A(n8427), .B(n8849), .Y(n3364) );
  INVX1 U1194 ( .A(n3364), .Y(n6502) );
  AND2X1 U1195 ( .A(n8456), .B(n9314), .Y(n3354) );
  INVX1 U1196 ( .A(n3354), .Y(n6503) );
  AND2X1 U1197 ( .A(n8427), .B(n9191), .Y(n3351) );
  INVX1 U1198 ( .A(n3351), .Y(n6504) );
  AND2X1 U1199 ( .A(n8456), .B(n9642), .Y(n3347) );
  INVX1 U1200 ( .A(n3347), .Y(n6505) );
  AND2X1 U1201 ( .A(n8430), .B(n9519), .Y(n3344) );
  INVX1 U1202 ( .A(n3344), .Y(n6506) );
  AND2X1 U1203 ( .A(n8456), .B(n8658), .Y(n3340) );
  INVX1 U1204 ( .A(n3340), .Y(n6507) );
  AND2X1 U1205 ( .A(n8430), .B(n8535), .Y(n3337) );
  INVX1 U1206 ( .A(n3337), .Y(n6508) );
  AND2X1 U1207 ( .A(n8456), .B(n8986), .Y(n3333) );
  INVX1 U1208 ( .A(n3333), .Y(n6509) );
  AND2X1 U1209 ( .A(n8427), .B(n8863), .Y(n3330) );
  INVX1 U1210 ( .A(n3330), .Y(n6510) );
  AND2X1 U1211 ( .A(n8456), .B(n9313), .Y(n3320) );
  INVX1 U1212 ( .A(n3320), .Y(n6511) );
  AND2X1 U1213 ( .A(n8428), .B(n9190), .Y(n3317) );
  INVX1 U1214 ( .A(n3317), .Y(n6512) );
  AND2X1 U1215 ( .A(n8456), .B(n9641), .Y(n3313) );
  INVX1 U1216 ( .A(n3313), .Y(n6513) );
  AND2X1 U1217 ( .A(n8428), .B(n9518), .Y(n3310) );
  INVX1 U1218 ( .A(n3310), .Y(n6514) );
  AND2X1 U1219 ( .A(n8456), .B(n8657), .Y(n3306) );
  INVX1 U1220 ( .A(n3306), .Y(n6515) );
  AND2X1 U1221 ( .A(n8428), .B(n8534), .Y(n3303) );
  INVX1 U1222 ( .A(n3303), .Y(n6516) );
  AND2X1 U1223 ( .A(n8456), .B(n8985), .Y(n3299) );
  INVX1 U1224 ( .A(n3299), .Y(n6517) );
  AND2X1 U1225 ( .A(n8427), .B(n8862), .Y(n3296) );
  INVX1 U1226 ( .A(n3296), .Y(n6518) );
  AND2X1 U1227 ( .A(n8455), .B(n9312), .Y(n3286) );
  INVX1 U1228 ( .A(n3286), .Y(n6519) );
  AND2X1 U1229 ( .A(n8427), .B(n9189), .Y(n3283) );
  INVX1 U1230 ( .A(n3283), .Y(n6520) );
  AND2X1 U1231 ( .A(n8455), .B(n9640), .Y(n3279) );
  INVX1 U1232 ( .A(n3279), .Y(n6521) );
  AND2X1 U1233 ( .A(n8428), .B(n9517), .Y(n3276) );
  INVX1 U1234 ( .A(n3276), .Y(n6522) );
  AND2X1 U1235 ( .A(n8455), .B(n8656), .Y(n3272) );
  INVX1 U1236 ( .A(n3272), .Y(n6523) );
  AND2X1 U1237 ( .A(n8427), .B(n8533), .Y(n3269) );
  INVX1 U1238 ( .A(n3269), .Y(n6524) );
  AND2X1 U1239 ( .A(n8455), .B(n8984), .Y(n3265) );
  INVX1 U1240 ( .A(n3265), .Y(n6525) );
  AND2X1 U1241 ( .A(n8429), .B(n8861), .Y(n3262) );
  INVX1 U1242 ( .A(n3262), .Y(n6526) );
  AND2X1 U1243 ( .A(n8455), .B(n9311), .Y(n3252) );
  INVX1 U1244 ( .A(n3252), .Y(n6527) );
  AND2X1 U1245 ( .A(n8429), .B(n9188), .Y(n3249) );
  INVX1 U1246 ( .A(n3249), .Y(n6528) );
  AND2X1 U1247 ( .A(n8455), .B(n9639), .Y(n3245) );
  INVX1 U1248 ( .A(n3245), .Y(n6529) );
  AND2X1 U1249 ( .A(n8430), .B(n9516), .Y(n3242) );
  INVX1 U1250 ( .A(n3242), .Y(n6530) );
  AND2X1 U1251 ( .A(n8455), .B(n8655), .Y(n3238) );
  INVX1 U1252 ( .A(n3238), .Y(n6531) );
  AND2X1 U1253 ( .A(n8429), .B(n8532), .Y(n3235) );
  INVX1 U1254 ( .A(n3235), .Y(n6532) );
  AND2X1 U1255 ( .A(n8455), .B(n8983), .Y(n3231) );
  INVX1 U1256 ( .A(n3231), .Y(n6533) );
  AND2X1 U1257 ( .A(n8430), .B(n8860), .Y(n3228) );
  INVX1 U1258 ( .A(n3228), .Y(n6534) );
  AND2X1 U1259 ( .A(n8455), .B(n9310), .Y(n3218) );
  INVX1 U1260 ( .A(n3218), .Y(n6535) );
  AND2X1 U1261 ( .A(n8430), .B(n9187), .Y(n3215) );
  INVX1 U1262 ( .A(n3215), .Y(n6536) );
  AND2X1 U1263 ( .A(n8455), .B(n9638), .Y(n3211) );
  INVX1 U1264 ( .A(n3211), .Y(n6537) );
  AND2X1 U1265 ( .A(n8428), .B(n9515), .Y(n3208) );
  INVX1 U1266 ( .A(n3208), .Y(n6538) );
  AND2X1 U1267 ( .A(n8455), .B(n8654), .Y(n3204) );
  INVX1 U1268 ( .A(n3204), .Y(n6539) );
  AND2X1 U1269 ( .A(n8430), .B(n8531), .Y(n3201) );
  INVX1 U1270 ( .A(n3201), .Y(n6540) );
  AND2X1 U1271 ( .A(n8455), .B(n8982), .Y(n3197) );
  INVX1 U1272 ( .A(n3197), .Y(n6541) );
  AND2X1 U1273 ( .A(n8428), .B(n8859), .Y(n3194) );
  INVX1 U1274 ( .A(n3194), .Y(n6542) );
  AND2X1 U1275 ( .A(n8454), .B(n9309), .Y(n3184) );
  INVX1 U1276 ( .A(n3184), .Y(n6543) );
  AND2X1 U1277 ( .A(n8428), .B(n9186), .Y(n3181) );
  INVX1 U1278 ( .A(n3181), .Y(n6544) );
  AND2X1 U1279 ( .A(n8454), .B(n9637), .Y(n3177) );
  INVX1 U1280 ( .A(n3177), .Y(n6545) );
  AND2X1 U1281 ( .A(n8427), .B(n9514), .Y(n3174) );
  INVX1 U1282 ( .A(n3174), .Y(n6546) );
  AND2X1 U1283 ( .A(n8454), .B(n8653), .Y(n3170) );
  INVX1 U1284 ( .A(n3170), .Y(n6547) );
  AND2X1 U1285 ( .A(n8428), .B(n8530), .Y(n3167) );
  INVX1 U1286 ( .A(n3167), .Y(n6548) );
  AND2X1 U1287 ( .A(n8454), .B(n8981), .Y(n1841) );
  INVX1 U1288 ( .A(n1841), .Y(n6549) );
  AND2X1 U1289 ( .A(n8427), .B(n8858), .Y(n1838) );
  INVX1 U1290 ( .A(n1838), .Y(n6550) );
  AND2X1 U1291 ( .A(n8454), .B(n9308), .Y(n1828) );
  INVX1 U1292 ( .A(n1828), .Y(n6551) );
  AND2X1 U1293 ( .A(n8427), .B(n9185), .Y(n1825) );
  INVX1 U1294 ( .A(n1825), .Y(n6552) );
  AND2X1 U1295 ( .A(n8454), .B(n9636), .Y(n1821) );
  INVX1 U1296 ( .A(n1821), .Y(n6553) );
  AND2X1 U1297 ( .A(n8429), .B(n9513), .Y(n1818) );
  INVX1 U1298 ( .A(n1818), .Y(n6554) );
  AND2X1 U1299 ( .A(n8454), .B(n8652), .Y(n1814) );
  INVX1 U1300 ( .A(n1814), .Y(n6555) );
  AND2X1 U1301 ( .A(n8427), .B(n8529), .Y(n1811) );
  INVX1 U1302 ( .A(n1811), .Y(n6556) );
  AND2X1 U1303 ( .A(n8454), .B(n8980), .Y(n1807) );
  INVX1 U1304 ( .A(n1807), .Y(n6557) );
  AND2X1 U1305 ( .A(n8429), .B(n8857), .Y(n1804) );
  INVX1 U1306 ( .A(n1804), .Y(n6558) );
  AND2X1 U1307 ( .A(n8454), .B(n9307), .Y(n1794) );
  INVX1 U1308 ( .A(n1794), .Y(n6559) );
  AND2X1 U1309 ( .A(n8429), .B(n9184), .Y(n1791) );
  INVX1 U1310 ( .A(n1791), .Y(n6560) );
  AND2X1 U1311 ( .A(n8454), .B(n9635), .Y(n1787) );
  INVX1 U1312 ( .A(n1787), .Y(n6561) );
  AND2X1 U1313 ( .A(n8428), .B(n9512), .Y(n1784) );
  INVX1 U1314 ( .A(n1784), .Y(n6562) );
  AND2X1 U1315 ( .A(n8454), .B(n8651), .Y(n1780) );
  INVX1 U1316 ( .A(n1780), .Y(n6563) );
  AND2X1 U1317 ( .A(n8428), .B(n8528), .Y(n1777) );
  INVX1 U1318 ( .A(n1777), .Y(n6564) );
  AND2X1 U1319 ( .A(n8454), .B(n8979), .Y(n1773) );
  INVX1 U1320 ( .A(n1773), .Y(n6565) );
  AND2X1 U1321 ( .A(n8428), .B(n8856), .Y(n1770) );
  INVX1 U1322 ( .A(n1770), .Y(n6566) );
  AND2X1 U1323 ( .A(n1361), .B(n9306), .Y(n1760) );
  INVX1 U1324 ( .A(n1760), .Y(n6567) );
  AND2X1 U1325 ( .A(n8428), .B(n9183), .Y(n1757) );
  INVX1 U1326 ( .A(n1757), .Y(n6568) );
  AND2X1 U1327 ( .A(n1361), .B(n9634), .Y(n1753) );
  INVX1 U1328 ( .A(n1753), .Y(n6569) );
  AND2X1 U1329 ( .A(n8428), .B(n9511), .Y(n1750) );
  INVX1 U1330 ( .A(n1750), .Y(n6570) );
  AND2X1 U1331 ( .A(n1361), .B(n8650), .Y(n1746) );
  INVX1 U1332 ( .A(n1746), .Y(n6571) );
  AND2X1 U1333 ( .A(n8428), .B(n8527), .Y(n1743) );
  INVX1 U1334 ( .A(n1743), .Y(n6572) );
  AND2X1 U1335 ( .A(n1361), .B(n8978), .Y(n1739) );
  INVX1 U1336 ( .A(n1739), .Y(n6573) );
  AND2X1 U1337 ( .A(n8428), .B(n8855), .Y(n1736) );
  INVX1 U1338 ( .A(n1736), .Y(n6574) );
  AND2X1 U1339 ( .A(n1361), .B(n9305), .Y(n1726) );
  INVX1 U1340 ( .A(n1726), .Y(n6575) );
  AND2X1 U1341 ( .A(n8428), .B(n9182), .Y(n1723) );
  INVX1 U1342 ( .A(n1723), .Y(n6576) );
  AND2X1 U1343 ( .A(n1361), .B(n9633), .Y(n1719) );
  INVX1 U1344 ( .A(n1719), .Y(n6577) );
  AND2X1 U1345 ( .A(n8428), .B(n9510), .Y(n1716) );
  INVX1 U1346 ( .A(n1716), .Y(n6578) );
  AND2X1 U1347 ( .A(n1361), .B(n8649), .Y(n1712) );
  INVX1 U1348 ( .A(n1712), .Y(n6579) );
  AND2X1 U1349 ( .A(n8428), .B(n8526), .Y(n1709) );
  INVX1 U1350 ( .A(n1709), .Y(n6580) );
  AND2X1 U1351 ( .A(n1361), .B(n8977), .Y(n1705) );
  INVX1 U1352 ( .A(n1705), .Y(n6581) );
  AND2X1 U1353 ( .A(n8428), .B(n8854), .Y(n1702) );
  INVX1 U1354 ( .A(n1702), .Y(n6582) );
  AND2X1 U1355 ( .A(n1361), .B(n9304), .Y(n1692) );
  INVX1 U1356 ( .A(n1692), .Y(n6583) );
  AND2X1 U1357 ( .A(n8428), .B(n9181), .Y(n1689) );
  INVX1 U1358 ( .A(n1689), .Y(n6584) );
  AND2X1 U1359 ( .A(n1361), .B(n9632), .Y(n1685) );
  INVX1 U1360 ( .A(n1685), .Y(n6585) );
  AND2X1 U1361 ( .A(n8428), .B(n9509), .Y(n1682) );
  INVX1 U1362 ( .A(n1682), .Y(n6586) );
  AND2X1 U1363 ( .A(n1361), .B(n8648), .Y(n1678) );
  INVX1 U1364 ( .A(n1678), .Y(n6587) );
  AND2X1 U1365 ( .A(n8428), .B(n8525), .Y(n1675) );
  INVX1 U1366 ( .A(n1675), .Y(n6588) );
  AND2X1 U1367 ( .A(n1361), .B(n8976), .Y(n1671) );
  INVX1 U1368 ( .A(n1671), .Y(n6589) );
  AND2X1 U1369 ( .A(n8428), .B(n8853), .Y(n1668) );
  INVX1 U1370 ( .A(n1668), .Y(n6590) );
  AND2X1 U1371 ( .A(n1361), .B(n9303), .Y(n1658) );
  INVX1 U1372 ( .A(n1658), .Y(n6591) );
  AND2X1 U1373 ( .A(n8428), .B(n9180), .Y(n1655) );
  INVX1 U1374 ( .A(n1655), .Y(n6592) );
  AND2X1 U1375 ( .A(n1361), .B(n9631), .Y(n1651) );
  INVX1 U1376 ( .A(n1651), .Y(n6593) );
  AND2X1 U1377 ( .A(n8428), .B(n9508), .Y(n1648) );
  INVX1 U1378 ( .A(n1648), .Y(n6594) );
  AND2X1 U1379 ( .A(n1361), .B(n8647), .Y(n1644) );
  INVX1 U1380 ( .A(n1644), .Y(n6595) );
  AND2X1 U1381 ( .A(n8427), .B(n8524), .Y(n1641) );
  INVX1 U1382 ( .A(n1641), .Y(n6596) );
  AND2X1 U1383 ( .A(n1361), .B(n8975), .Y(n1637) );
  INVX1 U1384 ( .A(n1637), .Y(n6597) );
  AND2X1 U1385 ( .A(n8427), .B(n8852), .Y(n1634) );
  INVX1 U1386 ( .A(n1634), .Y(n6598) );
  AND2X1 U1387 ( .A(n1361), .B(n9302), .Y(n1624) );
  INVX1 U1388 ( .A(n1624), .Y(n6599) );
  AND2X1 U1389 ( .A(n8427), .B(n9179), .Y(n1621) );
  INVX1 U1390 ( .A(n1621), .Y(n6600) );
  AND2X1 U1391 ( .A(n1361), .B(n9630), .Y(n1617) );
  INVX1 U1392 ( .A(n1617), .Y(n6601) );
  AND2X1 U1393 ( .A(n8427), .B(n9507), .Y(n1614) );
  INVX1 U1394 ( .A(n1614), .Y(n6602) );
  AND2X1 U1395 ( .A(n1361), .B(n8646), .Y(n1610) );
  INVX1 U1396 ( .A(n1610), .Y(n6603) );
  AND2X1 U1397 ( .A(n8427), .B(n8523), .Y(n1607) );
  INVX1 U1398 ( .A(n1607), .Y(n6604) );
  AND2X1 U1399 ( .A(n1361), .B(n8974), .Y(n1603) );
  INVX1 U1400 ( .A(n1603), .Y(n6605) );
  AND2X1 U1401 ( .A(n8427), .B(n8851), .Y(n1600) );
  INVX1 U1402 ( .A(n1600), .Y(n6606) );
  AND2X1 U1403 ( .A(n1361), .B(n9299), .Y(n1590) );
  INVX1 U1404 ( .A(n1590), .Y(n6607) );
  AND2X1 U1405 ( .A(n8427), .B(n9176), .Y(n1587) );
  INVX1 U1406 ( .A(n1587), .Y(n6608) );
  AND2X1 U1407 ( .A(n1361), .B(n9627), .Y(n1583) );
  INVX1 U1408 ( .A(n1583), .Y(n6609) );
  AND2X1 U1409 ( .A(n8427), .B(n9504), .Y(n1580) );
  INVX1 U1410 ( .A(n1580), .Y(n6610) );
  AND2X1 U1411 ( .A(n1361), .B(n8643), .Y(n1576) );
  INVX1 U1412 ( .A(n1576), .Y(n6611) );
  AND2X1 U1413 ( .A(n8427), .B(n8520), .Y(n1573) );
  INVX1 U1414 ( .A(n1573), .Y(n6612) );
  AND2X1 U1415 ( .A(n1361), .B(n8971), .Y(n1569) );
  INVX1 U1416 ( .A(n1569), .Y(n6613) );
  AND2X1 U1417 ( .A(n8427), .B(n8848), .Y(n1566) );
  INVX1 U1418 ( .A(n1566), .Y(n6614) );
  AND2X1 U1419 ( .A(n1361), .B(n9337), .Y(n1556) );
  INVX1 U1420 ( .A(n1556), .Y(n6615) );
  AND2X1 U1421 ( .A(n8427), .B(n9214), .Y(n1553) );
  INVX1 U1422 ( .A(n1553), .Y(n6616) );
  AND2X1 U1423 ( .A(n1361), .B(n9665), .Y(n1549) );
  INVX1 U1424 ( .A(n1549), .Y(n6617) );
  AND2X1 U1425 ( .A(n8427), .B(n9542), .Y(n1546) );
  INVX1 U1426 ( .A(n1546), .Y(n6618) );
  AND2X1 U1427 ( .A(n1361), .B(n8681), .Y(n1542) );
  INVX1 U1428 ( .A(n1542), .Y(n6619) );
  AND2X1 U1429 ( .A(n8427), .B(n8558), .Y(n1539) );
  INVX1 U1430 ( .A(n1539), .Y(n6620) );
  AND2X1 U1431 ( .A(n1361), .B(n9009), .Y(n1535) );
  INVX1 U1432 ( .A(n1535), .Y(n6621) );
  AND2X1 U1437 ( .A(n8427), .B(n8886), .Y(n1532) );
  INVX1 U1440 ( .A(n1532), .Y(n6622) );
  AND2X1 U1443 ( .A(n1361), .B(n9335), .Y(n1522) );
  INVX1 U1445 ( .A(n1522), .Y(n6623) );
  AND2X1 U1448 ( .A(n8427), .B(n9212), .Y(n1519) );
  INVX1 U1451 ( .A(n1519), .Y(n6624) );
  AND2X1 U1453 ( .A(n1361), .B(n9663), .Y(n1515) );
  INVX1 U1456 ( .A(n1515), .Y(n6625) );
  AND2X1 U1459 ( .A(n8427), .B(n9540), .Y(n1512) );
  INVX1 U1463 ( .A(n1512), .Y(n6626) );
  AND2X1 U1466 ( .A(n1361), .B(n8679), .Y(n1508) );
  INVX1 U1468 ( .A(n1508), .Y(n6627) );
  AND2X1 U1471 ( .A(n8427), .B(n8556), .Y(n1505) );
  INVX1 U1474 ( .A(n1505), .Y(n6628) );
  AND2X1 U1477 ( .A(n1361), .B(n9007), .Y(n1501) );
  INVX1 U1479 ( .A(n1501), .Y(n6629) );
  AND2X1 U1482 ( .A(n8427), .B(n8884), .Y(n1498) );
  INVX1 U1485 ( .A(n1498), .Y(n6630) );
  AND2X1 U1487 ( .A(n1361), .B(n9333), .Y(n1488) );
  INVX1 U1490 ( .A(n1488), .Y(n6631) );
  AND2X1 U1493 ( .A(n8430), .B(n9210), .Y(n1485) );
  INVX1 U1497 ( .A(n1485), .Y(n6632) );
  AND2X1 U1500 ( .A(n1361), .B(n9661), .Y(n1481) );
  INVX1 U1502 ( .A(n1481), .Y(n6633) );
  AND2X1 U1505 ( .A(n8427), .B(n9538), .Y(n1478) );
  INVX1 U1508 ( .A(n1478), .Y(n6634) );
  AND2X1 U1511 ( .A(n1361), .B(n8677), .Y(n1474) );
  INVX1 U1513 ( .A(n1474), .Y(n6635) );
  AND2X1 U1516 ( .A(n8428), .B(n8554), .Y(n1471) );
  INVX1 U1519 ( .A(n1471), .Y(n6636) );
  AND2X1 U1521 ( .A(n1361), .B(n9005), .Y(n1467) );
  INVX1 U1524 ( .A(n1467), .Y(n6637) );
  AND2X1 U1527 ( .A(n8429), .B(n8882), .Y(n1464) );
  INVX1 U1531 ( .A(n1464), .Y(n6638) );
  AND2X1 U1534 ( .A(n1361), .B(n9331), .Y(n1454) );
  INVX1 U1536 ( .A(n1454), .Y(n6639) );
  AND2X1 U1539 ( .A(n8429), .B(n9208), .Y(n1451) );
  INVX1 U1542 ( .A(n1451), .Y(n6640) );
  AND2X1 U1545 ( .A(n1361), .B(n9659), .Y(n1447) );
  INVX1 U1547 ( .A(n1447), .Y(n6641) );
  AND2X1 U1550 ( .A(n8427), .B(n9536), .Y(n1444) );
  INVX1 U1553 ( .A(n1444), .Y(n6642) );
  AND2X1 U1555 ( .A(n1361), .B(n8675), .Y(n1440) );
  INVX1 U1558 ( .A(n1440), .Y(n6643) );
  AND2X1 U1561 ( .A(n8429), .B(n8552), .Y(n1437) );
  INVX1 U1565 ( .A(n1437), .Y(n6644) );
  AND2X1 U1568 ( .A(n1361), .B(n9003), .Y(n1433) );
  INVX1 U1570 ( .A(n1433), .Y(n6645) );
  AND2X1 U1573 ( .A(n8428), .B(n8880), .Y(n1430) );
  INVX1 U1576 ( .A(n1430), .Y(n6646) );
  AND2X1 U1579 ( .A(n1361), .B(n9329), .Y(n1420) );
  INVX1 U1581 ( .A(n1420), .Y(n6647) );
  AND2X1 U1584 ( .A(n8428), .B(n9206), .Y(n1417) );
  INVX1 U1587 ( .A(n1417), .Y(n6648) );
  AND2X1 U1589 ( .A(n1361), .B(n9657), .Y(n1413) );
  INVX1 U1592 ( .A(n1413), .Y(n6649) );
  AND2X1 U1595 ( .A(n8428), .B(n9534), .Y(n1410) );
  INVX1 U1599 ( .A(n1410), .Y(n6650) );
  AND2X1 U1602 ( .A(n1361), .B(n8673), .Y(n1406) );
  INVX1 U1604 ( .A(n1406), .Y(n6651) );
  AND2X1 U1607 ( .A(n8427), .B(n8550), .Y(n1403) );
  INVX1 U1610 ( .A(n1403), .Y(n6652) );
  AND2X1 U1613 ( .A(n1361), .B(n9001), .Y(n1399) );
  INVX1 U1615 ( .A(n1399), .Y(n6653) );
  AND2X1 U1618 ( .A(n8430), .B(n8878), .Y(n1396) );
  INVX1 U1621 ( .A(n1396), .Y(n6654) );
  AND2X1 U1623 ( .A(n1361), .B(n9327), .Y(n1386) );
  INVX1 U1626 ( .A(n1386), .Y(n6655) );
  AND2X1 U1629 ( .A(n8429), .B(n9204), .Y(n1383) );
  INVX1 U1633 ( .A(n1383), .Y(n6656) );
  AND2X1 U1636 ( .A(n1361), .B(n9655), .Y(n1378) );
  INVX1 U1638 ( .A(n1378), .Y(n6657) );
  AND2X1 U1641 ( .A(n8429), .B(n9532), .Y(n1375) );
  INVX1 U1644 ( .A(n1375), .Y(n6658) );
  AND2X1 U1647 ( .A(n1361), .B(n8671), .Y(n1370) );
  INVX1 U1649 ( .A(n1370), .Y(n6659) );
  AND2X1 U1652 ( .A(n8430), .B(n8548), .Y(n1367) );
  INVX1 U1655 ( .A(n1367), .Y(n6660) );
  AND2X1 U1657 ( .A(n1361), .B(n8999), .Y(n1357) );
  INVX1 U1660 ( .A(n1357), .Y(n6661) );
  AND2X1 U1663 ( .A(n8430), .B(n8876), .Y(n1352) );
  INVX1 U1667 ( .A(n1352), .Y(n6662) );
  BUFX2 U1670 ( .A(n4080), .Y(n6663) );
  BUFX2 U1672 ( .A(n4072), .Y(n6664) );
  BUFX2 U1675 ( .A(n4069), .Y(n6665) );
  BUFX2 U1678 ( .A(n4065), .Y(n6666) );
  BUFX2 U1681 ( .A(n4061), .Y(n6667) );
  BUFX2 U1683 ( .A(n4057), .Y(n6668) );
  BUFX2 U1686 ( .A(n4053), .Y(n6669) );
  BUFX2 U1689 ( .A(n4049), .Y(n6670) );
  BUFX2 U1691 ( .A(n4045), .Y(n6671) );
  BUFX2 U1694 ( .A(n4035), .Y(n6672) );
  BUFX2 U1697 ( .A(n4032), .Y(n6673) );
  BUFX2 U1701 ( .A(n4028), .Y(n6674) );
  BUFX2 U1704 ( .A(n4025), .Y(n6675) );
  BUFX2 U1706 ( .A(n4021), .Y(n6676) );
  BUFX2 U1709 ( .A(n4018), .Y(n6677) );
  BUFX2 U1712 ( .A(n4014), .Y(n6678) );
  BUFX2 U1715 ( .A(n4011), .Y(n6679) );
  BUFX2 U1717 ( .A(n4001), .Y(n6680) );
  BUFX2 U1720 ( .A(n3998), .Y(n6681) );
  BUFX2 U1723 ( .A(n3994), .Y(n6682) );
  BUFX2 U1725 ( .A(n3991), .Y(n6683) );
  BUFX2 U1728 ( .A(n3987), .Y(n6684) );
  BUFX2 U1731 ( .A(n3984), .Y(n6685) );
  BUFX2 U1735 ( .A(n3980), .Y(n6686) );
  BUFX2 U1738 ( .A(n3977), .Y(n6687) );
  BUFX2 U1740 ( .A(n3967), .Y(n6688) );
  BUFX2 U1743 ( .A(n3964), .Y(n6689) );
  BUFX2 U1746 ( .A(n3960), .Y(n6690) );
  BUFX2 U1749 ( .A(n3957), .Y(n6691) );
  BUFX2 U1751 ( .A(n3953), .Y(n6692) );
  BUFX2 U1754 ( .A(n3950), .Y(n6693) );
  BUFX2 U1757 ( .A(n3946), .Y(n6694) );
  BUFX2 U1759 ( .A(n3943), .Y(n6695) );
  BUFX2 U1762 ( .A(n3933), .Y(n6696) );
  BUFX2 U1765 ( .A(n3930), .Y(n6697) );
  BUFX2 U1769 ( .A(n3926), .Y(n6698) );
  BUFX2 U1772 ( .A(n3923), .Y(n6699) );
  BUFX2 U1774 ( .A(n3919), .Y(n6700) );
  BUFX2 U1777 ( .A(n3916), .Y(n6701) );
  BUFX2 U1780 ( .A(n3912), .Y(n6702) );
  BUFX2 U1783 ( .A(n3909), .Y(n6703) );
  BUFX2 U1785 ( .A(n3899), .Y(n6704) );
  BUFX2 U1788 ( .A(n3896), .Y(n6705) );
  BUFX2 U1791 ( .A(n3892), .Y(n6706) );
  BUFX2 U1793 ( .A(n3889), .Y(n6707) );
  BUFX2 U1796 ( .A(n3885), .Y(n6708) );
  BUFX2 U1799 ( .A(n3882), .Y(n6709) );
  BUFX2 U1803 ( .A(n3878), .Y(n6710) );
  BUFX2 U1806 ( .A(n3875), .Y(n6711) );
  BUFX2 U1808 ( .A(n3865), .Y(n6712) );
  BUFX2 U1811 ( .A(n3862), .Y(n6713) );
  BUFX2 U1814 ( .A(n3858), .Y(n6714) );
  BUFX2 U1817 ( .A(n3855), .Y(n6715) );
  BUFX2 U1819 ( .A(n3851), .Y(n6716) );
  BUFX2 U1822 ( .A(n3848), .Y(n6717) );
  BUFX2 U1825 ( .A(n3844), .Y(n6718) );
  BUFX2 U1827 ( .A(n3841), .Y(n6719) );
  BUFX2 U1830 ( .A(n3831), .Y(n6720) );
  BUFX2 U1833 ( .A(n3828), .Y(n6721) );
  BUFX2 U1837 ( .A(n3824), .Y(n6722) );
  BUFX2 U1840 ( .A(n3821), .Y(n6723) );
  BUFX2 U1842 ( .A(n3817), .Y(n6724) );
  BUFX2 U1845 ( .A(n3814), .Y(n6725) );
  BUFX2 U1848 ( .A(n3810), .Y(n6726) );
  BUFX2 U1851 ( .A(n3807), .Y(n6727) );
  BUFX2 U1853 ( .A(n3797), .Y(n6728) );
  BUFX2 U1856 ( .A(n3794), .Y(n6729) );
  BUFX2 U1859 ( .A(n3790), .Y(n6730) );
  BUFX2 U1861 ( .A(n3787), .Y(n6731) );
  BUFX2 U1864 ( .A(n3783), .Y(n6732) );
  BUFX2 U1867 ( .A(n3780), .Y(n6733) );
  BUFX2 U1871 ( .A(n3776), .Y(n6734) );
  BUFX2 U1874 ( .A(n3773), .Y(n6735) );
  BUFX2 U1876 ( .A(n3763), .Y(n6736) );
  BUFX2 U1879 ( .A(n3760), .Y(n6737) );
  BUFX2 U1882 ( .A(n3756), .Y(n6738) );
  BUFX2 U1885 ( .A(n3753), .Y(n6739) );
  BUFX2 U1887 ( .A(n3749), .Y(n6740) );
  BUFX2 U1890 ( .A(n3746), .Y(n6741) );
  BUFX2 U1893 ( .A(n3742), .Y(n6742) );
  BUFX2 U1895 ( .A(n3739), .Y(n6743) );
  BUFX2 U1898 ( .A(n3729), .Y(n6744) );
  BUFX2 U1901 ( .A(n3726), .Y(n6745) );
  BUFX2 U1905 ( .A(n3722), .Y(n6746) );
  BUFX2 U1908 ( .A(n3719), .Y(n6747) );
  BUFX2 U1910 ( .A(n3715), .Y(n6748) );
  BUFX2 U1913 ( .A(n3712), .Y(n6749) );
  BUFX2 U1916 ( .A(n3708), .Y(n6750) );
  BUFX2 U1919 ( .A(n3705), .Y(n6751) );
  BUFX2 U1921 ( .A(n3695), .Y(n6752) );
  BUFX2 U1924 ( .A(n3692), .Y(n6753) );
  BUFX2 U1927 ( .A(n3688), .Y(n6754) );
  BUFX2 U1929 ( .A(n3685), .Y(n6755) );
  BUFX2 U1932 ( .A(n3681), .Y(n6756) );
  BUFX2 U1935 ( .A(n3678), .Y(n6757) );
  BUFX2 U1939 ( .A(n3674), .Y(n6758) );
  BUFX2 U1942 ( .A(n3671), .Y(n6759) );
  BUFX2 U1944 ( .A(n3661), .Y(n6760) );
  BUFX2 U1947 ( .A(n3658), .Y(n6761) );
  BUFX2 U1950 ( .A(n3654), .Y(n6762) );
  BUFX2 U1953 ( .A(n3651), .Y(n6763) );
  BUFX2 U1955 ( .A(n3647), .Y(n6764) );
  BUFX2 U1958 ( .A(n3644), .Y(n6765) );
  BUFX2 U1961 ( .A(n3640), .Y(n6766) );
  BUFX2 U1963 ( .A(n3637), .Y(n6767) );
  BUFX2 U1966 ( .A(n3627), .Y(n6768) );
  BUFX2 U1969 ( .A(n3624), .Y(n6769) );
  BUFX2 U1973 ( .A(n3620), .Y(n6770) );
  BUFX2 U1976 ( .A(n3617), .Y(n6771) );
  BUFX2 U1978 ( .A(n3613), .Y(n6772) );
  BUFX2 U1981 ( .A(n3610), .Y(n6773) );
  BUFX2 U1984 ( .A(n3606), .Y(n6774) );
  BUFX2 U1987 ( .A(n3603), .Y(n6775) );
  BUFX2 U1989 ( .A(n3593), .Y(n6776) );
  BUFX2 U1992 ( .A(n3590), .Y(n6777) );
  BUFX2 U1995 ( .A(n3586), .Y(n6778) );
  BUFX2 U1997 ( .A(n3583), .Y(n6779) );
  BUFX2 U2000 ( .A(n3579), .Y(n6780) );
  BUFX2 U2003 ( .A(n3576), .Y(n6781) );
  BUFX2 U2007 ( .A(n3572), .Y(n6782) );
  BUFX2 U2010 ( .A(n3569), .Y(n6783) );
  BUFX2 U2012 ( .A(n3559), .Y(n6784) );
  BUFX2 U2015 ( .A(n3556), .Y(n6785) );
  BUFX2 U2018 ( .A(n3552), .Y(n6786) );
  BUFX2 U2021 ( .A(n3549), .Y(n6787) );
  BUFX2 U2023 ( .A(n3545), .Y(n6788) );
  BUFX2 U2026 ( .A(n3542), .Y(n6789) );
  BUFX2 U2029 ( .A(n3538), .Y(n6790) );
  BUFX2 U2031 ( .A(n3535), .Y(n6791) );
  BUFX2 U2034 ( .A(n3525), .Y(n6792) );
  BUFX2 U2037 ( .A(n3522), .Y(n6793) );
  BUFX2 U2041 ( .A(n3518), .Y(n6794) );
  BUFX2 U2044 ( .A(n3515), .Y(n6795) );
  BUFX2 U2046 ( .A(n3511), .Y(n6796) );
  BUFX2 U2049 ( .A(n3508), .Y(n6797) );
  BUFX2 U2052 ( .A(n3504), .Y(n6798) );
  BUFX2 U2055 ( .A(n3501), .Y(n6799) );
  BUFX2 U2057 ( .A(n3491), .Y(n6800) );
  BUFX2 U2060 ( .A(n3488), .Y(n6801) );
  BUFX2 U2063 ( .A(n3484), .Y(n6802) );
  BUFX2 U2065 ( .A(n3481), .Y(n6803) );
  BUFX2 U2068 ( .A(n3477), .Y(n6804) );
  BUFX2 U2071 ( .A(n3474), .Y(n6805) );
  BUFX2 U2075 ( .A(n3470), .Y(n6806) );
  BUFX2 U2078 ( .A(n3467), .Y(n6807) );
  BUFX2 U2080 ( .A(n3457), .Y(n6808) );
  BUFX2 U2083 ( .A(n3454), .Y(n6809) );
  BUFX2 U2086 ( .A(n3450), .Y(n6810) );
  BUFX2 U2089 ( .A(n3447), .Y(n6811) );
  BUFX2 U2091 ( .A(n3443), .Y(n6812) );
  BUFX2 U2094 ( .A(n3440), .Y(n6813) );
  BUFX2 U2097 ( .A(n3436), .Y(n6814) );
  BUFX2 U2099 ( .A(n3433), .Y(n6815) );
  BUFX2 U2102 ( .A(n3423), .Y(n6816) );
  BUFX2 U2105 ( .A(n3420), .Y(n6817) );
  BUFX2 U2109 ( .A(n3416), .Y(n6818) );
  BUFX2 U2112 ( .A(n3413), .Y(n6819) );
  BUFX2 U2114 ( .A(n3409), .Y(n6820) );
  BUFX2 U2117 ( .A(n3406), .Y(n6821) );
  BUFX2 U2120 ( .A(n3402), .Y(n6822) );
  BUFX2 U2123 ( .A(n3399), .Y(n6823) );
  BUFX2 U2125 ( .A(n3389), .Y(n6824) );
  BUFX2 U2128 ( .A(n3386), .Y(n6825) );
  BUFX2 U2131 ( .A(n3382), .Y(n6826) );
  BUFX2 U2133 ( .A(n3379), .Y(n6827) );
  BUFX2 U2136 ( .A(n3375), .Y(n6828) );
  BUFX2 U2139 ( .A(n3372), .Y(n6829) );
  BUFX2 U2143 ( .A(n3368), .Y(n6830) );
  BUFX2 U2146 ( .A(n3365), .Y(n6831) );
  BUFX2 U2148 ( .A(n3355), .Y(n6832) );
  BUFX2 U2151 ( .A(n3352), .Y(n6833) );
  BUFX2 U2154 ( .A(n3348), .Y(n6834) );
  BUFX2 U2157 ( .A(n3345), .Y(n6835) );
  BUFX2 U2159 ( .A(n3341), .Y(n6836) );
  BUFX2 U2162 ( .A(n3338), .Y(n6837) );
  BUFX2 U2165 ( .A(n3334), .Y(n6838) );
  BUFX2 U2167 ( .A(n3331), .Y(n6839) );
  BUFX2 U2170 ( .A(n3321), .Y(n6840) );
  BUFX2 U2173 ( .A(n3318), .Y(n6841) );
  BUFX2 U2177 ( .A(n3314), .Y(n6842) );
  BUFX2 U2180 ( .A(n3311), .Y(n6843) );
  BUFX2 U2182 ( .A(n3307), .Y(n6844) );
  BUFX2 U2185 ( .A(n3304), .Y(n6845) );
  BUFX2 U2188 ( .A(n3300), .Y(n6846) );
  BUFX2 U2191 ( .A(n3297), .Y(n6847) );
  BUFX2 U2193 ( .A(n3287), .Y(n6848) );
  BUFX2 U2196 ( .A(n3284), .Y(n6849) );
  BUFX2 U2199 ( .A(n3280), .Y(n6850) );
  BUFX2 U2201 ( .A(n3277), .Y(n6851) );
  BUFX2 U2204 ( .A(n3273), .Y(n6852) );
  BUFX2 U2207 ( .A(n3270), .Y(n6853) );
  BUFX2 U2211 ( .A(n3266), .Y(n6854) );
  BUFX2 U2214 ( .A(n3263), .Y(n6855) );
  BUFX2 U2216 ( .A(n3253), .Y(n6856) );
  BUFX2 U2219 ( .A(n3250), .Y(n6857) );
  BUFX2 U2222 ( .A(n3246), .Y(n6858) );
  BUFX2 U2225 ( .A(n3243), .Y(n6859) );
  BUFX2 U2227 ( .A(n3239), .Y(n6860) );
  BUFX2 U2230 ( .A(n3236), .Y(n6861) );
  BUFX2 U2233 ( .A(n3232), .Y(n6862) );
  BUFX2 U2235 ( .A(n3229), .Y(n6863) );
  BUFX2 U2238 ( .A(n3219), .Y(n6864) );
  BUFX2 U2241 ( .A(n3216), .Y(n6865) );
  BUFX2 U2245 ( .A(n3212), .Y(n6866) );
  BUFX2 U2248 ( .A(n3209), .Y(n6867) );
  BUFX2 U2250 ( .A(n3205), .Y(n6868) );
  BUFX2 U2253 ( .A(n3202), .Y(n6869) );
  BUFX2 U2256 ( .A(n3198), .Y(n6870) );
  BUFX2 U2259 ( .A(n3195), .Y(n6871) );
  BUFX2 U2261 ( .A(n3185), .Y(n6872) );
  BUFX2 U2264 ( .A(n3182), .Y(n6873) );
  BUFX2 U2267 ( .A(n3178), .Y(n6874) );
  BUFX2 U2269 ( .A(n3175), .Y(n6875) );
  BUFX2 U2272 ( .A(n3171), .Y(n6876) );
  BUFX2 U2275 ( .A(n3168), .Y(n6877) );
  BUFX2 U2279 ( .A(n3164), .Y(n6878) );
  BUFX2 U2282 ( .A(n1839), .Y(n6879) );
  BUFX2 U2284 ( .A(n1829), .Y(n6880) );
  BUFX2 U2287 ( .A(n1826), .Y(n6881) );
  BUFX2 U2290 ( .A(n1822), .Y(n6882) );
  BUFX2 U2293 ( .A(n1819), .Y(n6883) );
  BUFX2 U2295 ( .A(n1815), .Y(n6884) );
  BUFX2 U2298 ( .A(n1812), .Y(n6885) );
  BUFX2 U2301 ( .A(n1808), .Y(n6886) );
  BUFX2 U2303 ( .A(n1805), .Y(n6887) );
  BUFX2 U2306 ( .A(n1795), .Y(n6888) );
  BUFX2 U2309 ( .A(n1792), .Y(n6889) );
  BUFX2 U2313 ( .A(n1788), .Y(n6890) );
  BUFX2 U2316 ( .A(n1785), .Y(n6891) );
  BUFX2 U2318 ( .A(n1781), .Y(n6892) );
  BUFX2 U2321 ( .A(n1778), .Y(n6893) );
  BUFX2 U2324 ( .A(n1774), .Y(n6894) );
  BUFX2 U2327 ( .A(n1771), .Y(n6895) );
  BUFX2 U2329 ( .A(n1761), .Y(n6896) );
  BUFX2 U2332 ( .A(n1758), .Y(n6897) );
  BUFX2 U2335 ( .A(n1754), .Y(n6898) );
  BUFX2 U2337 ( .A(n1751), .Y(n6899) );
  BUFX2 U2340 ( .A(n1747), .Y(n6900) );
  BUFX2 U2343 ( .A(n1744), .Y(n6901) );
  BUFX2 U2347 ( .A(n1740), .Y(n6902) );
  BUFX2 U2350 ( .A(n1737), .Y(n6903) );
  BUFX2 U2352 ( .A(n1727), .Y(n6904) );
  BUFX2 U2355 ( .A(n1724), .Y(n6905) );
  BUFX2 U2358 ( .A(n1720), .Y(n6906) );
  BUFX2 U2361 ( .A(n1717), .Y(n6907) );
  BUFX2 U2363 ( .A(n1713), .Y(n6908) );
  BUFX2 U2366 ( .A(n1710), .Y(n6909) );
  BUFX2 U2369 ( .A(n1706), .Y(n6910) );
  BUFX2 U2371 ( .A(n1703), .Y(n6911) );
  BUFX2 U2374 ( .A(n1693), .Y(n6912) );
  BUFX2 U2377 ( .A(n1690), .Y(n6913) );
  BUFX2 U2381 ( .A(n1686), .Y(n6914) );
  BUFX2 U2384 ( .A(n1683), .Y(n6915) );
  BUFX2 U2386 ( .A(n1679), .Y(n6916) );
  BUFX2 U2389 ( .A(n1676), .Y(n6917) );
  BUFX2 U2392 ( .A(n1672), .Y(n6918) );
  BUFX2 U2395 ( .A(n1669), .Y(n6919) );
  BUFX2 U2397 ( .A(n1659), .Y(n6920) );
  BUFX2 U2400 ( .A(n1656), .Y(n6921) );
  BUFX2 U2403 ( .A(n1652), .Y(n6922) );
  BUFX2 U2405 ( .A(n1649), .Y(n6923) );
  BUFX2 U2408 ( .A(n1645), .Y(n6924) );
  BUFX2 U2411 ( .A(n1642), .Y(n6925) );
  BUFX2 U2415 ( .A(n1638), .Y(n6926) );
  BUFX2 U2418 ( .A(n1635), .Y(n6927) );
  BUFX2 U2420 ( .A(n1625), .Y(n6928) );
  BUFX2 U2423 ( .A(n1622), .Y(n6929) );
  BUFX2 U2426 ( .A(n1618), .Y(n6930) );
  BUFX2 U2429 ( .A(n1615), .Y(n6931) );
  BUFX2 U2431 ( .A(n1611), .Y(n6932) );
  BUFX2 U2434 ( .A(n1608), .Y(n6933) );
  BUFX2 U2437 ( .A(n1604), .Y(n6934) );
  BUFX2 U2439 ( .A(n1601), .Y(n6935) );
  BUFX2 U2442 ( .A(n1591), .Y(n6936) );
  BUFX2 U2445 ( .A(n1588), .Y(n6937) );
  BUFX2 U2449 ( .A(n1584), .Y(n6938) );
  BUFX2 U2452 ( .A(n1581), .Y(n6939) );
  BUFX2 U2454 ( .A(n1577), .Y(n6940) );
  BUFX2 U2457 ( .A(n1574), .Y(n6941) );
  BUFX2 U2460 ( .A(n1570), .Y(n6942) );
  BUFX2 U2463 ( .A(n1567), .Y(n6943) );
  BUFX2 U2465 ( .A(n1557), .Y(n6944) );
  BUFX2 U2468 ( .A(n1554), .Y(n6945) );
  BUFX2 U2471 ( .A(n1550), .Y(n6946) );
  BUFX2 U2473 ( .A(n1547), .Y(n6947) );
  BUFX2 U2476 ( .A(n1543), .Y(n6948) );
  BUFX2 U2479 ( .A(n1540), .Y(n6949) );
  BUFX2 U2483 ( .A(n1536), .Y(n6950) );
  BUFX2 U2486 ( .A(n1533), .Y(n6951) );
  BUFX2 U2488 ( .A(n1523), .Y(n6952) );
  BUFX2 U2491 ( .A(n1520), .Y(n6953) );
  BUFX2 U2494 ( .A(n1516), .Y(n6954) );
  BUFX2 U2497 ( .A(n1513), .Y(n6955) );
  BUFX2 U2499 ( .A(n1509), .Y(n6956) );
  BUFX2 U2502 ( .A(n1506), .Y(n6957) );
  BUFX2 U2505 ( .A(n1502), .Y(n6958) );
  BUFX2 U2507 ( .A(n1499), .Y(n6959) );
  BUFX2 U2510 ( .A(n1489), .Y(n6960) );
  BUFX2 U2513 ( .A(n1486), .Y(n6961) );
  BUFX2 U2517 ( .A(n1482), .Y(n6962) );
  BUFX2 U2520 ( .A(n1479), .Y(n6963) );
  BUFX2 U2522 ( .A(n1475), .Y(n6964) );
  BUFX2 U2525 ( .A(n1472), .Y(n6965) );
  BUFX2 U2528 ( .A(n1468), .Y(n6966) );
  BUFX2 U2531 ( .A(n1465), .Y(n6967) );
  BUFX2 U2533 ( .A(n1455), .Y(n6968) );
  BUFX2 U2536 ( .A(n1452), .Y(n6969) );
  BUFX2 U2539 ( .A(n1448), .Y(n6970) );
  BUFX2 U2541 ( .A(n1445), .Y(n6971) );
  BUFX2 U2544 ( .A(n1441), .Y(n6972) );
  BUFX2 U2547 ( .A(n1438), .Y(n6973) );
  BUFX2 U2551 ( .A(n1434), .Y(n6974) );
  BUFX2 U2554 ( .A(n1431), .Y(n6975) );
  BUFX2 U2556 ( .A(n1421), .Y(n6976) );
  BUFX2 U2559 ( .A(n1418), .Y(n6977) );
  BUFX2 U2562 ( .A(n1414), .Y(n6978) );
  BUFX2 U2565 ( .A(n1411), .Y(n6979) );
  BUFX2 U2567 ( .A(n1407), .Y(n6980) );
  BUFX2 U2570 ( .A(n1404), .Y(n6981) );
  BUFX2 U2573 ( .A(n1400), .Y(n6982) );
  BUFX2 U2575 ( .A(n1397), .Y(n6983) );
  BUFX2 U2578 ( .A(n1387), .Y(n6984) );
  BUFX2 U2581 ( .A(n1384), .Y(n6985) );
  BUFX2 U2585 ( .A(n1379), .Y(n6986) );
  BUFX2 U2588 ( .A(n1376), .Y(n6987) );
  BUFX2 U2590 ( .A(n1371), .Y(n6988) );
  BUFX2 U2593 ( .A(n1368), .Y(n6989) );
  BUFX2 U2596 ( .A(n1358), .Y(n6990) );
  BUFX2 U2599 ( .A(n1353), .Y(n6991) );
  INVX1 U2601 ( .A(n4039), .Y(n6992) );
  INVX1 U2604 ( .A(n4005), .Y(n6993) );
  INVX1 U2607 ( .A(n3971), .Y(n6994) );
  INVX1 U2609 ( .A(n3937), .Y(n6995) );
  INVX1 U2612 ( .A(n3903), .Y(n6996) );
  INVX1 U2615 ( .A(n3869), .Y(n6997) );
  INVX1 U2619 ( .A(n3835), .Y(n6998) );
  INVX1 U2622 ( .A(n3801), .Y(n6999) );
  INVX1 U2624 ( .A(n3767), .Y(n7000) );
  INVX1 U2627 ( .A(n3733), .Y(n7001) );
  INVX1 U2630 ( .A(n3699), .Y(n7002) );
  INVX1 U2633 ( .A(n3665), .Y(n7003) );
  INVX1 U2635 ( .A(n3631), .Y(n7004) );
  INVX1 U2638 ( .A(n3597), .Y(n7005) );
  INVX1 U2641 ( .A(n3563), .Y(n7006) );
  INVX1 U2643 ( .A(n3529), .Y(n7007) );
  INVX1 U2646 ( .A(n3495), .Y(n7008) );
  INVX1 U2649 ( .A(n3461), .Y(n7009) );
  INVX1 U2653 ( .A(n3427), .Y(n7010) );
  INVX1 U2656 ( .A(n3393), .Y(n7011) );
  INVX1 U2658 ( .A(n3359), .Y(n7012) );
  INVX1 U2661 ( .A(n3325), .Y(n7013) );
  INVX1 U2664 ( .A(n3291), .Y(n7014) );
  INVX1 U2667 ( .A(n3257), .Y(n7015) );
  INVX1 U2669 ( .A(n3223), .Y(n7016) );
  INVX1 U2672 ( .A(n3189), .Y(n7017) );
  INVX1 U2675 ( .A(n1833), .Y(n7018) );
  INVX1 U2677 ( .A(n1799), .Y(n7019) );
  INVX1 U2680 ( .A(n1765), .Y(n7020) );
  INVX1 U2683 ( .A(n1731), .Y(n7021) );
  INVX1 U2687 ( .A(n1697), .Y(n7022) );
  INVX1 U2690 ( .A(n1663), .Y(n7023) );
  INVX1 U2692 ( .A(n1629), .Y(n7024) );
  INVX1 U2695 ( .A(n1595), .Y(n7025) );
  INVX1 U2698 ( .A(n1561), .Y(n7026) );
  INVX1 U2701 ( .A(n1527), .Y(n7027) );
  INVX1 U2703 ( .A(n1493), .Y(n7028) );
  INVX1 U2706 ( .A(n1459), .Y(n7029) );
  INVX1 U2709 ( .A(n1425), .Y(n7030) );
  INVX1 U2711 ( .A(n1391), .Y(n7031) );
  INVX1 U2714 ( .A(n1347), .Y(n7032) );
  INVX1 U2717 ( .A(n4040), .Y(n7033) );
  INVX1 U2721 ( .A(n4006), .Y(n7034) );
  INVX1 U2724 ( .A(n3972), .Y(n7035) );
  INVX1 U2726 ( .A(n3938), .Y(n7036) );
  INVX1 U2729 ( .A(n3904), .Y(n7037) );
  INVX1 U2732 ( .A(n3870), .Y(n7038) );
  INVX1 U2735 ( .A(n3836), .Y(n7039) );
  INVX1 U2737 ( .A(n3802), .Y(n7040) );
  INVX1 U2740 ( .A(n3768), .Y(n7041) );
  INVX1 U2743 ( .A(n3734), .Y(n7042) );
  INVX1 U2745 ( .A(n3700), .Y(n7043) );
  INVX1 U2748 ( .A(n3666), .Y(n7044) );
  INVX1 U2751 ( .A(n3632), .Y(n7045) );
  INVX1 U2755 ( .A(n3598), .Y(n7046) );
  INVX1 U2758 ( .A(n3564), .Y(n7047) );
  INVX1 U2760 ( .A(n3530), .Y(n7048) );
  INVX1 U2763 ( .A(n3496), .Y(n7049) );
  INVX1 U2766 ( .A(n3462), .Y(n7050) );
  INVX1 U2769 ( .A(n3428), .Y(n7051) );
  INVX1 U2771 ( .A(n3394), .Y(n7052) );
  INVX1 U2774 ( .A(n3360), .Y(n7053) );
  INVX1 U2777 ( .A(n3326), .Y(n7054) );
  INVX1 U2779 ( .A(n3292), .Y(n7055) );
  INVX1 U2782 ( .A(n3258), .Y(n7056) );
  INVX1 U2785 ( .A(n3224), .Y(n7057) );
  INVX1 U2789 ( .A(n3190), .Y(n7058) );
  INVX1 U2792 ( .A(n1834), .Y(n7059) );
  INVX1 U2794 ( .A(n1800), .Y(n7060) );
  INVX1 U2797 ( .A(n1766), .Y(n7061) );
  INVX1 U2800 ( .A(n1732), .Y(n7062) );
  INVX1 U2803 ( .A(n1698), .Y(n7063) );
  INVX1 U2805 ( .A(n1664), .Y(n7064) );
  INVX1 U2808 ( .A(n1630), .Y(n7065) );
  INVX1 U2811 ( .A(n1596), .Y(n7066) );
  INVX1 U2813 ( .A(n1562), .Y(n7067) );
  INVX1 U2816 ( .A(n1528), .Y(n7068) );
  INVX1 U2820 ( .A(n1494), .Y(n7069) );
  INVX1 U2825 ( .A(n1460), .Y(n7070) );
  INVX1 U2828 ( .A(n1426), .Y(n7071) );
  INVX1 U2830 ( .A(n1392), .Y(n7072) );
  INVX1 U2835 ( .A(n1348), .Y(n7073) );
  INVX1 U2836 ( .A(n4041), .Y(n7074) );
  INVX1 U2839 ( .A(n4007), .Y(n7075) );
  INVX1 U2849 ( .A(n3973), .Y(n7076) );
  INVX1 U2850 ( .A(n3939), .Y(n7077) );
  INVX1 U2851 ( .A(n3905), .Y(n7078) );
  INVX1 U2856 ( .A(n3871), .Y(n7079) );
  INVX1 U2866 ( .A(n3837), .Y(n7080) );
  INVX1 U2867 ( .A(n3803), .Y(n7081) );
  INVX1 U2869 ( .A(n3769), .Y(n7082) );
  INVX1 U2871 ( .A(n3735), .Y(n7083) );
  INVX1 U2873 ( .A(n3701), .Y(n7084) );
  INVX1 U2875 ( .A(n3667), .Y(n7085) );
  INVX1 U2877 ( .A(n3633), .Y(n7086) );
  INVX1 U2879 ( .A(n3599), .Y(n7087) );
  INVX1 U2881 ( .A(n3565), .Y(n7088) );
  INVX1 U2883 ( .A(n3531), .Y(n7089) );
  INVX1 U2885 ( .A(n3497), .Y(n7090) );
  INVX1 U2887 ( .A(n3463), .Y(n7091) );
  INVX1 U2889 ( .A(n3429), .Y(n7092) );
  INVX1 U2891 ( .A(n3395), .Y(n7093) );
  INVX1 U2893 ( .A(n3361), .Y(n7094) );
  INVX1 U2895 ( .A(n3327), .Y(n7095) );
  INVX1 U2897 ( .A(n3293), .Y(n7096) );
  INVX1 U2899 ( .A(n3259), .Y(n7097) );
  INVX1 U2901 ( .A(n3225), .Y(n7098) );
  INVX1 U2903 ( .A(n3191), .Y(n7099) );
  INVX1 U2905 ( .A(n1835), .Y(n7100) );
  INVX1 U2907 ( .A(n1801), .Y(n7101) );
  INVX1 U2909 ( .A(n1767), .Y(n7102) );
  INVX1 U2911 ( .A(n1733), .Y(n7103) );
  INVX1 U2913 ( .A(n1699), .Y(n7104) );
  INVX1 U2915 ( .A(n1665), .Y(n7105) );
  INVX1 U2917 ( .A(n1631), .Y(n7106) );
  INVX1 U2919 ( .A(n1597), .Y(n7107) );
  INVX1 U2921 ( .A(n1563), .Y(n7108) );
  INVX1 U2923 ( .A(n1529), .Y(n7109) );
  INVX1 U2925 ( .A(n1495), .Y(n7110) );
  INVX1 U2927 ( .A(n1461), .Y(n7111) );
  INVX1 U2929 ( .A(n1427), .Y(n7112) );
  INVX1 U2931 ( .A(n1393), .Y(n7113) );
  INVX1 U2933 ( .A(n1349), .Y(n7114) );
  BUFX2 U2935 ( .A(n1343), .Y(n7115) );
  BUFX2 U2937 ( .A(n4084), .Y(n7116) );
  AND2X1 U2939 ( .A(n4132), .B(n4106), .Y(n4131) );
  INVX1 U2941 ( .A(n4131), .Y(n7117) );
  AND2X1 U2943 ( .A(n4156), .B(n4106), .Y(n4155) );
  INVX1 U2945 ( .A(n4155), .Y(n7118) );
  AND2X1 U2947 ( .A(n4180), .B(n4106), .Y(n4179) );
  INVX1 U2949 ( .A(n4179), .Y(n7119) );
  AND2X1 U2952 ( .A(n4130), .B(n4190), .Y(n4202) );
  INVX1 U2954 ( .A(n4202), .Y(n7120) );
  AND2X1 U2956 ( .A(n4154), .B(n4190), .Y(n4214) );
  INVX1 U2958 ( .A(n4214), .Y(n7121) );
  AND2X1 U2960 ( .A(n4178), .B(n4190), .Y(n4226) );
  INVX1 U2962 ( .A(n4226), .Y(n7122) );
  AND2X1 U2964 ( .A(n4128), .B(n4233), .Y(n4244) );
  INVX1 U2966 ( .A(n4244), .Y(n7123) );
  AND2X1 U2968 ( .A(n4152), .B(n4233), .Y(n4256) );
  INVX1 U2970 ( .A(n4256), .Y(n7124) );
  AND2X1 U2972 ( .A(n4176), .B(n4233), .Y(n4268) );
  INVX1 U2974 ( .A(n4268), .Y(n7125) );
  AND2X1 U2976 ( .A(n4150), .B(n4276), .Y(n4298) );
  INVX1 U2978 ( .A(n4298), .Y(n7126) );
  AND2X1 U2980 ( .A(n4174), .B(n4276), .Y(n4310) );
  INVX1 U2982 ( .A(n4310), .Y(n7127) );
  AND2X1 U2984 ( .A(n4148), .B(n4319), .Y(n4340) );
  INVX1 U2986 ( .A(n4340), .Y(n7128) );
  AND2X1 U2988 ( .A(n4172), .B(n4319), .Y(n4352) );
  INVX1 U2990 ( .A(n4352), .Y(n7129) );
  AND2X1 U2992 ( .A(n4108), .B(n4361), .Y(n4362) );
  INVX1 U2994 ( .A(n4362), .Y(n7130) );
  AND2X1 U2996 ( .A(n4146), .B(n4361), .Y(n4381) );
  INVX1 U2998 ( .A(n4381), .Y(n7131) );
  AND2X1 U3000 ( .A(n4170), .B(n4361), .Y(n4393) );
  INVX1 U3002 ( .A(n4393), .Y(n7132) );
  AND2X1 U3004 ( .A(n4144), .B(n4404), .Y(n4423) );
  INVX1 U3006 ( .A(n4423), .Y(n7133) );
  AND2X1 U3008 ( .A(n4168), .B(n4404), .Y(n4435) );
  INVX1 U3010 ( .A(n4435), .Y(n7134) );
  AND2X1 U3012 ( .A(n4142), .B(n4447), .Y(n4465) );
  INVX1 U3014 ( .A(n4465), .Y(n7135) );
  AND2X1 U3016 ( .A(n4166), .B(n4447), .Y(n4477) );
  INVX1 U3018 ( .A(n4477), .Y(n7136) );
  AND2X1 U3020 ( .A(n4116), .B(n4490), .Y(n4495) );
  INVX1 U3022 ( .A(n4495), .Y(n7137) );
  AND2X1 U3024 ( .A(n4126), .B(n4490), .Y(n4500) );
  INVX1 U3026 ( .A(n4500), .Y(n7138) );
  AND2X1 U3028 ( .A(n4114), .B(n4533), .Y(n4537) );
  INVX1 U3030 ( .A(n4537), .Y(n7139) );
  AND2X1 U3032 ( .A(n4124), .B(n4533), .Y(n4542) );
  INVX1 U3035 ( .A(n4542), .Y(n7140) );
  AND2X1 U3037 ( .A(n4112), .B(n4575), .Y(n4578) );
  INVX1 U3039 ( .A(n4578), .Y(n7141) );
  AND2X1 U3041 ( .A(n4122), .B(n4575), .Y(n4583) );
  INVX1 U3043 ( .A(n4583), .Y(n7142) );
  AND2X1 U3045 ( .A(n4110), .B(n4617), .Y(n4619) );
  INVX1 U3047 ( .A(n4619), .Y(n7143) );
  AND2X1 U3049 ( .A(n4120), .B(n4617), .Y(n4624) );
  INVX1 U3051 ( .A(n4624), .Y(n7144) );
  AND2X1 U3053 ( .A(n4132), .B(n4659), .Y(n4672) );
  INVX1 U3055 ( .A(n4672), .Y(n7145) );
  AND2X1 U3057 ( .A(n4156), .B(n4659), .Y(n4684) );
  INVX1 U3059 ( .A(n4684), .Y(n7146) );
  AND2X1 U3061 ( .A(n4180), .B(n4659), .Y(n4696) );
  INVX1 U3063 ( .A(n4696), .Y(n7147) );
  AND2X1 U3065 ( .A(n4130), .B(n4701), .Y(n4713) );
  INVX1 U3067 ( .A(n4713), .Y(n7148) );
  AND2X1 U3069 ( .A(n4154), .B(n4701), .Y(n4725) );
  INVX1 U3071 ( .A(n4725), .Y(n7149) );
  AND2X1 U3073 ( .A(n4178), .B(n4701), .Y(n4737) );
  INVX1 U3075 ( .A(n4737), .Y(n7150) );
  AND2X1 U3077 ( .A(n4128), .B(n4743), .Y(n4754) );
  INVX1 U3079 ( .A(n4754), .Y(n7151) );
  AND2X1 U3081 ( .A(n4152), .B(n4743), .Y(n4766) );
  INVX1 U3083 ( .A(n4766), .Y(n7152) );
  AND2X1 U3085 ( .A(n4176), .B(n4743), .Y(n4778) );
  INVX1 U3087 ( .A(n4778), .Y(n7153) );
  AND2X1 U3089 ( .A(n4150), .B(n4785), .Y(n4807) );
  INVX1 U3091 ( .A(n4807), .Y(n7154) );
  AND2X1 U3093 ( .A(n4174), .B(n4785), .Y(n4819) );
  INVX1 U3095 ( .A(n4819), .Y(n7155) );
  AND2X1 U3097 ( .A(n4148), .B(n4827), .Y(n4848) );
  INVX1 U3099 ( .A(n4848), .Y(n7156) );
  AND2X1 U3101 ( .A(n4172), .B(n4827), .Y(n4860) );
  INVX1 U3103 ( .A(n4860), .Y(n7157) );
  AND2X1 U3105 ( .A(n4108), .B(n4870), .Y(n4871) );
  INVX1 U3107 ( .A(n4871), .Y(n7158) );
  AND2X1 U3109 ( .A(n4146), .B(n4870), .Y(n4890) );
  INVX1 U3111 ( .A(n4890), .Y(n7159) );
  AND2X1 U3113 ( .A(n4170), .B(n4870), .Y(n4902) );
  INVX1 U3115 ( .A(n4902), .Y(n7160) );
  AND2X1 U3118 ( .A(n4144), .B(n4912), .Y(n4931) );
  INVX1 U3120 ( .A(n4931), .Y(n7161) );
  AND2X1 U3122 ( .A(n4168), .B(n4912), .Y(n4943) );
  INVX1 U3124 ( .A(n4943), .Y(n7162) );
  AND2X1 U3126 ( .A(n4142), .B(n4954), .Y(n4972) );
  INVX1 U3128 ( .A(n4972), .Y(n7163) );
  AND2X1 U3130 ( .A(n4166), .B(n4954), .Y(n4984) );
  INVX1 U3132 ( .A(n4984), .Y(n7164) );
  AND2X1 U3134 ( .A(n4116), .B(n4996), .Y(n5001) );
  INVX1 U3136 ( .A(n5001), .Y(n7165) );
  AND2X1 U3138 ( .A(n4126), .B(n4996), .Y(n5006) );
  INVX1 U3140 ( .A(n5006), .Y(n7166) );
  AND2X1 U3142 ( .A(n4114), .B(n5038), .Y(n5042) );
  INVX1 U3144 ( .A(n5042), .Y(n7167) );
  AND2X1 U3146 ( .A(n4124), .B(n5038), .Y(n5047) );
  INVX1 U3148 ( .A(n5047), .Y(n7168) );
  AND2X1 U3150 ( .A(n4112), .B(n5080), .Y(n5083) );
  INVX1 U3152 ( .A(n5083), .Y(n7169) );
  AND2X1 U3154 ( .A(n4122), .B(n5080), .Y(n5088) );
  INVX1 U3156 ( .A(n5088), .Y(n7170) );
  AND2X1 U3158 ( .A(n4110), .B(n5122), .Y(n5124) );
  INVX1 U3160 ( .A(n5124), .Y(n7171) );
  AND2X1 U3162 ( .A(n4120), .B(n5122), .Y(n5129) );
  INVX1 U3164 ( .A(n5129), .Y(n7172) );
  AND2X1 U3166 ( .A(n4148), .B(n5164), .Y(n5185) );
  INVX1 U3168 ( .A(n5185), .Y(n7173) );
  AND2X1 U3170 ( .A(n4172), .B(n5164), .Y(n5197) );
  INVX1 U3172 ( .A(n5197), .Y(n7174) );
  AND2X1 U3174 ( .A(n4108), .B(n5207), .Y(n5208) );
  INVX1 U3176 ( .A(n5208), .Y(n7175) );
  AND2X1 U3178 ( .A(n4146), .B(n5207), .Y(n5227) );
  INVX1 U3180 ( .A(n5227), .Y(n7176) );
  AND2X1 U3182 ( .A(n4170), .B(n5207), .Y(n5239) );
  INVX1 U3184 ( .A(n5239), .Y(n7177) );
  AND2X1 U3186 ( .A(n4144), .B(n5249), .Y(n5268) );
  INVX1 U3188 ( .A(n5268), .Y(n7178) );
  AND2X1 U3190 ( .A(n4168), .B(n5249), .Y(n5280) );
  INVX1 U3192 ( .A(n5280), .Y(n7179) );
  AND2X1 U3194 ( .A(n4142), .B(n5291), .Y(n5309) );
  INVX1 U3196 ( .A(n5309), .Y(n7180) );
  AND2X1 U3198 ( .A(n4166), .B(n5291), .Y(n5321) );
  INVX1 U3201 ( .A(n5321), .Y(n7181) );
  AND2X1 U3203 ( .A(n4116), .B(n5333), .Y(n5338) );
  INVX1 U3205 ( .A(n5338), .Y(n7182) );
  AND2X1 U3207 ( .A(n4126), .B(n5333), .Y(n5343) );
  INVX1 U3209 ( .A(n5343), .Y(n7183) );
  AND2X1 U3211 ( .A(n4114), .B(n5375), .Y(n5379) );
  INVX1 U3213 ( .A(n5379), .Y(n7184) );
  AND2X1 U3215 ( .A(n4124), .B(n5375), .Y(n5384) );
  INVX1 U3217 ( .A(n5384), .Y(n7185) );
  AND2X1 U3219 ( .A(n4112), .B(n5417), .Y(n5420) );
  INVX1 U3221 ( .A(n5420), .Y(n7186) );
  AND2X1 U3223 ( .A(n4122), .B(n5417), .Y(n5425) );
  INVX1 U3225 ( .A(n5425), .Y(n7187) );
  AND2X1 U3227 ( .A(n4110), .B(n5459), .Y(n5461) );
  INVX1 U3229 ( .A(n5461), .Y(n7188) );
  AND2X1 U3231 ( .A(n4120), .B(n5459), .Y(n5466) );
  INVX1 U3233 ( .A(n5466), .Y(n7189) );
  AND2X1 U3235 ( .A(n4130), .B(n4106), .Y(n4129) );
  INVX1 U3237 ( .A(n4129), .Y(n7190) );
  AND2X1 U3239 ( .A(n4154), .B(n4106), .Y(n4153) );
  INVX1 U3241 ( .A(n4153), .Y(n7191) );
  AND2X1 U3243 ( .A(n4178), .B(n4106), .Y(n4177) );
  INVX1 U3245 ( .A(n4177), .Y(n7192) );
  AND2X1 U3247 ( .A(n4132), .B(n4190), .Y(n4203) );
  INVX1 U3249 ( .A(n4203), .Y(n7193) );
  AND2X1 U3251 ( .A(n4156), .B(n4190), .Y(n4215) );
  INVX1 U3253 ( .A(n4215), .Y(n7194) );
  AND2X1 U3255 ( .A(n4180), .B(n4190), .Y(n4227) );
  INVX1 U3257 ( .A(n4227), .Y(n7195) );
  AND2X1 U3259 ( .A(n4150), .B(n4233), .Y(n4255) );
  INVX1 U3261 ( .A(n4255), .Y(n7196) );
  AND2X1 U3263 ( .A(n4174), .B(n4233), .Y(n4267) );
  INVX1 U3265 ( .A(n4267), .Y(n7197) );
  AND2X1 U3267 ( .A(n4128), .B(n4276), .Y(n4287) );
  INVX1 U3269 ( .A(n4287), .Y(n7198) );
  AND2X1 U3271 ( .A(n4152), .B(n4276), .Y(n4299) );
  INVX1 U3273 ( .A(n4299), .Y(n7199) );
  AND2X1 U3275 ( .A(n4176), .B(n4276), .Y(n4311) );
  INVX1 U3277 ( .A(n4311), .Y(n7200) );
  AND2X1 U3279 ( .A(n4108), .B(n4319), .Y(n4320) );
  INVX1 U3281 ( .A(n4320), .Y(n7201) );
  AND2X1 U3284 ( .A(n4146), .B(n4319), .Y(n4339) );
  INVX1 U3286 ( .A(n4339), .Y(n7202) );
  AND2X1 U3288 ( .A(n4170), .B(n4319), .Y(n4351) );
  INVX1 U3290 ( .A(n4351), .Y(n7203) );
  AND2X1 U3292 ( .A(n4148), .B(n4361), .Y(n4382) );
  INVX1 U3294 ( .A(n4382), .Y(n7204) );
  AND2X1 U3296 ( .A(n4172), .B(n4361), .Y(n4394) );
  INVX1 U3298 ( .A(n4394), .Y(n7205) );
  AND2X1 U3300 ( .A(n4142), .B(n4404), .Y(n4422) );
  INVX1 U3302 ( .A(n4422), .Y(n7206) );
  AND2X1 U3304 ( .A(n4166), .B(n4404), .Y(n4434) );
  INVX1 U3306 ( .A(n4434), .Y(n7207) );
  AND2X1 U3308 ( .A(n4144), .B(n4447), .Y(n4466) );
  INVX1 U3310 ( .A(n4466), .Y(n7208) );
  AND2X1 U3312 ( .A(n4168), .B(n4447), .Y(n4478) );
  INVX1 U3314 ( .A(n4478), .Y(n7209) );
  AND2X1 U3316 ( .A(n4114), .B(n4490), .Y(n4494) );
  INVX1 U3318 ( .A(n4494), .Y(n7210) );
  AND2X1 U3320 ( .A(n4124), .B(n4490), .Y(n4499) );
  INVX1 U3322 ( .A(n4499), .Y(n7211) );
  AND2X1 U3324 ( .A(n4116), .B(n4533), .Y(n4538) );
  INVX1 U3326 ( .A(n4538), .Y(n7212) );
  AND2X1 U3328 ( .A(n4126), .B(n4533), .Y(n4543) );
  INVX1 U3330 ( .A(n4543), .Y(n7213) );
  AND2X1 U3332 ( .A(n4110), .B(n4575), .Y(n4577) );
  INVX1 U3334 ( .A(n4577), .Y(n7214) );
  AND2X1 U3336 ( .A(n4120), .B(n4575), .Y(n4582) );
  INVX1 U3338 ( .A(n4582), .Y(n7215) );
  AND2X1 U3340 ( .A(n4112), .B(n4617), .Y(n4620) );
  INVX1 U3342 ( .A(n4620), .Y(n7216) );
  AND2X1 U3344 ( .A(n4122), .B(n4617), .Y(n4625) );
  INVX1 U3346 ( .A(n4625), .Y(n7217) );
  AND2X1 U3348 ( .A(n4130), .B(n4659), .Y(n4671) );
  INVX1 U3350 ( .A(n4671), .Y(n7218) );
  AND2X1 U3352 ( .A(n4154), .B(n4659), .Y(n4683) );
  INVX1 U3354 ( .A(n4683), .Y(n7219) );
  AND2X1 U3356 ( .A(n4178), .B(n4659), .Y(n4695) );
  INVX1 U3358 ( .A(n4695), .Y(n7220) );
  AND2X1 U3360 ( .A(n4132), .B(n4701), .Y(n4714) );
  INVX1 U3362 ( .A(n4714), .Y(n7221) );
  AND2X1 U3364 ( .A(n4156), .B(n4701), .Y(n4726) );
  INVX1 U3367 ( .A(n4726), .Y(n7222) );
  AND2X1 U3369 ( .A(n4180), .B(n4701), .Y(n4738) );
  INVX1 U3371 ( .A(n4738), .Y(n7223) );
  AND2X1 U3373 ( .A(n4150), .B(n4743), .Y(n4765) );
  INVX1 U3375 ( .A(n4765), .Y(n7224) );
  AND2X1 U3377 ( .A(n4174), .B(n4743), .Y(n4777) );
  INVX1 U3379 ( .A(n4777), .Y(n7225) );
  AND2X1 U3381 ( .A(n4128), .B(n4785), .Y(n4796) );
  INVX1 U3383 ( .A(n4796), .Y(n7226) );
  AND2X1 U3385 ( .A(n4152), .B(n4785), .Y(n4808) );
  INVX1 U3387 ( .A(n4808), .Y(n7227) );
  AND2X1 U3389 ( .A(n4176), .B(n4785), .Y(n4820) );
  INVX1 U3391 ( .A(n4820), .Y(n7228) );
  AND2X1 U3393 ( .A(n4108), .B(n4827), .Y(n4828) );
  INVX1 U3395 ( .A(n4828), .Y(n7229) );
  AND2X1 U3397 ( .A(n4146), .B(n4827), .Y(n4847) );
  INVX1 U3399 ( .A(n4847), .Y(n7230) );
  AND2X1 U3401 ( .A(n4170), .B(n4827), .Y(n4859) );
  INVX1 U3403 ( .A(n4859), .Y(n7231) );
  AND2X1 U3405 ( .A(n4148), .B(n4870), .Y(n4891) );
  INVX1 U3407 ( .A(n4891), .Y(n7232) );
  AND2X1 U3409 ( .A(n4172), .B(n4870), .Y(n4903) );
  INVX1 U3411 ( .A(n4903), .Y(n7233) );
  AND2X1 U3413 ( .A(n4142), .B(n4912), .Y(n4930) );
  INVX1 U3415 ( .A(n4930), .Y(n7234) );
  AND2X1 U3417 ( .A(n4166), .B(n4912), .Y(n4942) );
  INVX1 U3419 ( .A(n4942), .Y(n7235) );
  AND2X1 U3421 ( .A(n4144), .B(n4954), .Y(n4973) );
  INVX1 U3423 ( .A(n4973), .Y(n7236) );
  AND2X1 U3425 ( .A(n4168), .B(n4954), .Y(n4985) );
  INVX1 U3427 ( .A(n4985), .Y(n7237) );
  AND2X1 U3429 ( .A(n4114), .B(n4996), .Y(n5000) );
  INVX1 U3431 ( .A(n5000), .Y(n7238) );
  AND2X1 U3433 ( .A(n4124), .B(n4996), .Y(n5005) );
  INVX1 U3435 ( .A(n5005), .Y(n7239) );
  AND2X1 U3437 ( .A(n4116), .B(n5038), .Y(n5043) );
  INVX1 U3439 ( .A(n5043), .Y(n7240) );
  AND2X1 U3441 ( .A(n4126), .B(n5038), .Y(n5048) );
  INVX1 U3443 ( .A(n5048), .Y(n7241) );
  AND2X1 U3445 ( .A(n4110), .B(n5080), .Y(n5082) );
  INVX1 U3447 ( .A(n5082), .Y(n7242) );
  AND2X1 U3450 ( .A(n4120), .B(n5080), .Y(n5087) );
  INVX1 U3452 ( .A(n5087), .Y(n7243) );
  AND2X1 U3454 ( .A(n4112), .B(n5122), .Y(n5125) );
  INVX1 U3456 ( .A(n5125), .Y(n7244) );
  AND2X1 U3458 ( .A(n4122), .B(n5122), .Y(n5130) );
  INVX1 U3460 ( .A(n5130), .Y(n7245) );
  AND2X1 U3462 ( .A(n4108), .B(n5164), .Y(n5165) );
  INVX1 U3464 ( .A(n5165), .Y(n7246) );
  AND2X1 U3466 ( .A(n4146), .B(n5164), .Y(n5184) );
  INVX1 U3468 ( .A(n5184), .Y(n7247) );
  AND2X1 U3470 ( .A(n4170), .B(n5164), .Y(n5196) );
  INVX1 U3472 ( .A(n5196), .Y(n7248) );
  AND2X1 U3474 ( .A(n4148), .B(n5207), .Y(n5228) );
  INVX1 U3476 ( .A(n5228), .Y(n7249) );
  AND2X1 U3478 ( .A(n4172), .B(n5207), .Y(n5240) );
  INVX1 U3480 ( .A(n5240), .Y(n7250) );
  AND2X1 U3482 ( .A(n4142), .B(n5249), .Y(n5267) );
  INVX1 U3484 ( .A(n5267), .Y(n7251) );
  AND2X1 U3486 ( .A(n4166), .B(n5249), .Y(n5279) );
  INVX1 U3488 ( .A(n5279), .Y(n7252) );
  AND2X1 U3490 ( .A(n4144), .B(n5291), .Y(n5310) );
  INVX1 U3492 ( .A(n5310), .Y(n7253) );
  AND2X1 U3494 ( .A(n4168), .B(n5291), .Y(n5322) );
  INVX1 U3496 ( .A(n5322), .Y(n7254) );
  AND2X1 U3498 ( .A(n4114), .B(n5333), .Y(n5337) );
  INVX1 U3500 ( .A(n5337), .Y(n7255) );
  AND2X1 U3502 ( .A(n4124), .B(n5333), .Y(n5342) );
  INVX1 U3504 ( .A(n5342), .Y(n7256) );
  AND2X1 U3506 ( .A(n4116), .B(n5375), .Y(n5380) );
  INVX1 U3508 ( .A(n5380), .Y(n7257) );
  AND2X1 U3510 ( .A(n4126), .B(n5375), .Y(n5385) );
  INVX1 U3512 ( .A(n5385), .Y(n7258) );
  AND2X1 U3514 ( .A(n4110), .B(n5417), .Y(n5419) );
  INVX1 U3516 ( .A(n5419), .Y(n7259) );
  AND2X1 U3518 ( .A(n4120), .B(n5417), .Y(n5424) );
  INVX1 U3520 ( .A(n5424), .Y(n7260) );
  AND2X1 U3522 ( .A(n4112), .B(n5459), .Y(n5462) );
  INVX1 U3524 ( .A(n5462), .Y(n7261) );
  AND2X1 U3526 ( .A(n4122), .B(n5459), .Y(n5467) );
  INVX1 U3528 ( .A(n5467), .Y(n7262) );
  AND2X1 U3530 ( .A(n4128), .B(n4106), .Y(n4127) );
  INVX1 U3534 ( .A(n4127), .Y(n7263) );
  AND2X1 U3536 ( .A(n4152), .B(n4106), .Y(n4151) );
  INVX1 U3538 ( .A(n4151), .Y(n7264) );
  AND2X1 U3540 ( .A(n4176), .B(n4106), .Y(n4175) );
  INVX1 U3542 ( .A(n4175), .Y(n7265) );
  AND2X1 U3544 ( .A(n4150), .B(n4190), .Y(n4212) );
  INVX1 U3546 ( .A(n4212), .Y(n7266) );
  AND2X1 U3548 ( .A(n4174), .B(n4190), .Y(n4224) );
  INVX1 U3550 ( .A(n4224), .Y(n7267) );
  AND2X1 U3552 ( .A(n4132), .B(n4233), .Y(n4246) );
  INVX1 U3554 ( .A(n4246), .Y(n7268) );
  AND2X1 U3556 ( .A(n4156), .B(n4233), .Y(n4258) );
  INVX1 U3558 ( .A(n4258), .Y(n7269) );
  AND2X1 U3560 ( .A(n4180), .B(n4233), .Y(n4270) );
  INVX1 U3562 ( .A(n4270), .Y(n7270) );
  AND2X1 U3564 ( .A(n4130), .B(n4276), .Y(n4288) );
  INVX1 U3566 ( .A(n4288), .Y(n7271) );
  AND2X1 U3568 ( .A(n4154), .B(n4276), .Y(n4300) );
  INVX1 U3570 ( .A(n4300), .Y(n7272) );
  AND2X1 U3572 ( .A(n4178), .B(n4276), .Y(n4312) );
  INVX1 U3574 ( .A(n4312), .Y(n7273) );
  AND2X1 U3576 ( .A(n4144), .B(n4319), .Y(n4338) );
  INVX1 U3578 ( .A(n4338), .Y(n7274) );
  AND2X1 U3580 ( .A(n4168), .B(n4319), .Y(n4350) );
  INVX1 U3582 ( .A(n4350), .Y(n7275) );
  AND2X1 U3584 ( .A(n4142), .B(n4361), .Y(n4379) );
  INVX1 U3586 ( .A(n4379), .Y(n7276) );
  AND2X1 U3588 ( .A(n4166), .B(n4361), .Y(n4391) );
  INVX1 U3590 ( .A(n4391), .Y(n7277) );
  AND2X1 U3592 ( .A(n4148), .B(n4404), .Y(n4425) );
  INVX1 U3594 ( .A(n4425), .Y(n7278) );
  AND2X1 U3596 ( .A(n4172), .B(n4404), .Y(n4437) );
  INVX1 U3598 ( .A(n4437), .Y(n7279) );
  AND2X1 U3600 ( .A(n4108), .B(n4447), .Y(n4448) );
  INVX1 U3602 ( .A(n4448), .Y(n7280) );
  AND2X1 U3604 ( .A(n4146), .B(n4447), .Y(n4467) );
  INVX1 U3606 ( .A(n4467), .Y(n7281) );
  AND2X1 U3608 ( .A(n4170), .B(n4447), .Y(n4479) );
  INVX1 U3610 ( .A(n4479), .Y(n7282) );
  AND2X1 U3612 ( .A(n4112), .B(n4490), .Y(n4493) );
  INVX1 U3614 ( .A(n4493), .Y(n7283) );
  AND2X1 U3617 ( .A(n4122), .B(n4490), .Y(n4498) );
  INVX1 U3619 ( .A(n4498), .Y(n7284) );
  AND2X1 U3621 ( .A(n4110), .B(n4533), .Y(n4535) );
  INVX1 U3623 ( .A(n4535), .Y(n7285) );
  AND2X1 U3625 ( .A(n4120), .B(n4533), .Y(n4540) );
  INVX1 U3627 ( .A(n4540), .Y(n7286) );
  AND2X1 U3629 ( .A(n4116), .B(n4575), .Y(n4580) );
  INVX1 U3631 ( .A(n4580), .Y(n7287) );
  AND2X1 U3633 ( .A(n4126), .B(n4575), .Y(n4585) );
  INVX1 U3635 ( .A(n4585), .Y(n7288) );
  AND2X1 U3637 ( .A(n4114), .B(n4617), .Y(n4621) );
  INVX1 U3639 ( .A(n4621), .Y(n7289) );
  AND2X1 U3641 ( .A(n4124), .B(n4617), .Y(n4626) );
  INVX1 U3643 ( .A(n4626), .Y(n7290) );
  AND2X1 U3645 ( .A(n4128), .B(n4659), .Y(n4670) );
  INVX1 U3647 ( .A(n4670), .Y(n7291) );
  AND2X1 U3649 ( .A(n4152), .B(n4659), .Y(n4682) );
  INVX1 U3651 ( .A(n4682), .Y(n7292) );
  AND2X1 U3653 ( .A(n4176), .B(n4659), .Y(n4694) );
  INVX1 U3655 ( .A(n4694), .Y(n7293) );
  AND2X1 U3657 ( .A(n4150), .B(n4701), .Y(n4723) );
  INVX1 U3659 ( .A(n4723), .Y(n7294) );
  AND2X1 U3661 ( .A(n4174), .B(n4701), .Y(n4735) );
  INVX1 U3663 ( .A(n4735), .Y(n7295) );
  AND2X1 U3665 ( .A(n4132), .B(n4743), .Y(n4756) );
  INVX1 U3667 ( .A(n4756), .Y(n7296) );
  AND2X1 U3669 ( .A(n4156), .B(n4743), .Y(n4768) );
  INVX1 U3671 ( .A(n4768), .Y(n7297) );
  AND2X1 U3673 ( .A(n4180), .B(n4743), .Y(n4780) );
  INVX1 U3675 ( .A(n4780), .Y(n7298) );
  AND2X1 U3677 ( .A(n4130), .B(n4785), .Y(n4797) );
  INVX1 U3679 ( .A(n4797), .Y(n7299) );
  AND2X1 U3681 ( .A(n4154), .B(n4785), .Y(n4809) );
  INVX1 U3683 ( .A(n4809), .Y(n7300) );
  AND2X1 U3685 ( .A(n4178), .B(n4785), .Y(n4821) );
  INVX1 U3687 ( .A(n4821), .Y(n7301) );
  AND2X1 U3689 ( .A(n4144), .B(n4827), .Y(n4846) );
  INVX1 U3691 ( .A(n4846), .Y(n7302) );
  AND2X1 U3693 ( .A(n4168), .B(n4827), .Y(n4858) );
  INVX1 U3695 ( .A(n4858), .Y(n7303) );
  AND2X1 U3697 ( .A(n4142), .B(n4870), .Y(n4888) );
  INVX1 U3700 ( .A(n4888), .Y(n7304) );
  AND2X1 U3702 ( .A(n4166), .B(n4870), .Y(n4900) );
  INVX1 U3704 ( .A(n4900), .Y(n7305) );
  AND2X1 U3706 ( .A(n4148), .B(n4912), .Y(n4933) );
  INVX1 U3708 ( .A(n4933), .Y(n7306) );
  AND2X1 U3710 ( .A(n4172), .B(n4912), .Y(n4945) );
  INVX1 U3712 ( .A(n4945), .Y(n7307) );
  AND2X1 U3714 ( .A(n4108), .B(n4954), .Y(n4955) );
  INVX1 U3716 ( .A(n4955), .Y(n7308) );
  AND2X1 U3718 ( .A(n4146), .B(n4954), .Y(n4974) );
  INVX1 U3720 ( .A(n4974), .Y(n7309) );
  AND2X1 U3722 ( .A(n4170), .B(n4954), .Y(n4986) );
  INVX1 U3724 ( .A(n4986), .Y(n7310) );
  AND2X1 U3726 ( .A(n4112), .B(n4996), .Y(n4999) );
  INVX1 U3728 ( .A(n4999), .Y(n7311) );
  AND2X1 U3730 ( .A(n4122), .B(n4996), .Y(n5004) );
  INVX1 U3732 ( .A(n5004), .Y(n7312) );
  AND2X1 U3734 ( .A(n4110), .B(n5038), .Y(n5040) );
  INVX1 U3736 ( .A(n5040), .Y(n7313) );
  AND2X1 U3738 ( .A(n4120), .B(n5038), .Y(n5045) );
  INVX1 U3740 ( .A(n5045), .Y(n7314) );
  AND2X1 U3742 ( .A(n4116), .B(n5080), .Y(n5085) );
  INVX1 U3744 ( .A(n5085), .Y(n7315) );
  AND2X1 U3746 ( .A(n4126), .B(n5080), .Y(n5090) );
  INVX1 U3748 ( .A(n5090), .Y(n7316) );
  AND2X1 U3750 ( .A(n4114), .B(n5122), .Y(n5126) );
  INVX1 U3752 ( .A(n5126), .Y(n7317) );
  AND2X1 U3754 ( .A(n4124), .B(n5122), .Y(n5131) );
  INVX1 U3756 ( .A(n5131), .Y(n7318) );
  AND2X1 U3758 ( .A(n4144), .B(n5164), .Y(n5183) );
  INVX1 U3760 ( .A(n5183), .Y(n7319) );
  AND2X1 U3762 ( .A(n4168), .B(n5164), .Y(n5195) );
  INVX1 U3764 ( .A(n5195), .Y(n7320) );
  AND2X1 U3766 ( .A(n4142), .B(n5207), .Y(n5225) );
  INVX1 U3768 ( .A(n5225), .Y(n7321) );
  AND2X1 U3770 ( .A(n4166), .B(n5207), .Y(n5237) );
  INVX1 U3772 ( .A(n5237), .Y(n7322) );
  AND2X1 U3774 ( .A(n4148), .B(n5249), .Y(n5270) );
  INVX1 U3776 ( .A(n5270), .Y(n7323) );
  AND2X1 U3778 ( .A(n4172), .B(n5249), .Y(n5282) );
  INVX1 U3780 ( .A(n5282), .Y(n7324) );
  AND2X1 U3783 ( .A(n4108), .B(n5291), .Y(n5292) );
  INVX1 U3785 ( .A(n5292), .Y(n7325) );
  AND2X1 U3787 ( .A(n4146), .B(n5291), .Y(n5311) );
  INVX1 U3789 ( .A(n5311), .Y(n7326) );
  AND2X1 U3791 ( .A(n4170), .B(n5291), .Y(n5323) );
  INVX1 U3793 ( .A(n5323), .Y(n7327) );
  AND2X1 U3795 ( .A(n4112), .B(n5333), .Y(n5336) );
  INVX1 U3797 ( .A(n5336), .Y(n7328) );
  AND2X1 U3799 ( .A(n4122), .B(n5333), .Y(n5341) );
  INVX1 U3801 ( .A(n5341), .Y(n7329) );
  AND2X1 U3803 ( .A(n4110), .B(n5375), .Y(n5377) );
  INVX1 U3805 ( .A(n5377), .Y(n7330) );
  AND2X1 U3807 ( .A(n4120), .B(n5375), .Y(n5382) );
  INVX1 U3809 ( .A(n5382), .Y(n7331) );
  AND2X1 U3811 ( .A(n4116), .B(n5417), .Y(n5422) );
  INVX1 U3813 ( .A(n5422), .Y(n7332) );
  AND2X1 U3815 ( .A(n4126), .B(n5417), .Y(n5427) );
  INVX1 U3817 ( .A(n5427), .Y(n7333) );
  AND2X1 U3819 ( .A(n4114), .B(n5459), .Y(n5463) );
  INVX1 U3821 ( .A(n5463), .Y(n7334) );
  AND2X1 U3823 ( .A(n4124), .B(n5459), .Y(n5468) );
  INVX1 U3825 ( .A(n5468), .Y(n7335) );
  AND2X1 U3827 ( .A(n4150), .B(n4106), .Y(n4149) );
  INVX1 U3829 ( .A(n4149), .Y(n7336) );
  AND2X1 U3831 ( .A(n4174), .B(n4106), .Y(n4173) );
  INVX1 U3833 ( .A(n4173), .Y(n7337) );
  AND2X1 U3835 ( .A(n4128), .B(n4190), .Y(n4201) );
  INVX1 U3837 ( .A(n4201), .Y(n7338) );
  AND2X1 U3839 ( .A(n4152), .B(n4190), .Y(n4213) );
  INVX1 U3841 ( .A(n4213), .Y(n7339) );
  AND2X1 U3843 ( .A(n4176), .B(n4190), .Y(n4225) );
  INVX1 U3845 ( .A(n4225), .Y(n7340) );
  AND2X1 U3847 ( .A(n4130), .B(n4233), .Y(n4245) );
  INVX1 U3849 ( .A(n4245), .Y(n7341) );
  AND2X1 U3851 ( .A(n4154), .B(n4233), .Y(n4257) );
  INVX1 U3853 ( .A(n4257), .Y(n7342) );
  AND2X1 U3855 ( .A(n4178), .B(n4233), .Y(n4269) );
  INVX1 U3857 ( .A(n4269), .Y(n7343) );
  AND2X1 U3859 ( .A(n4132), .B(n4276), .Y(n4289) );
  INVX1 U3861 ( .A(n4289), .Y(n7344) );
  AND2X1 U3863 ( .A(n4156), .B(n4276), .Y(n4301) );
  INVX1 U3866 ( .A(n4301), .Y(n7345) );
  AND2X1 U3868 ( .A(n4180), .B(n4276), .Y(n4313) );
  INVX1 U3870 ( .A(n4313), .Y(n7346) );
  AND2X1 U3872 ( .A(n4142), .B(n4319), .Y(n4337) );
  INVX1 U3874 ( .A(n4337), .Y(n7347) );
  AND2X1 U3876 ( .A(n4166), .B(n4319), .Y(n4349) );
  INVX1 U3878 ( .A(n4349), .Y(n7348) );
  AND2X1 U3880 ( .A(n4144), .B(n4361), .Y(n4380) );
  INVX1 U3882 ( .A(n4380), .Y(n7349) );
  AND2X1 U3884 ( .A(n4168), .B(n4361), .Y(n4392) );
  INVX1 U3886 ( .A(n4392), .Y(n7350) );
  AND2X1 U3888 ( .A(n4108), .B(n4404), .Y(n4405) );
  INVX1 U3890 ( .A(n4405), .Y(n7351) );
  AND2X1 U3892 ( .A(n4146), .B(n4404), .Y(n4424) );
  INVX1 U3894 ( .A(n4424), .Y(n7352) );
  AND2X1 U3896 ( .A(n4170), .B(n4404), .Y(n4436) );
  INVX1 U3898 ( .A(n4436), .Y(n7353) );
  AND2X1 U3900 ( .A(n4148), .B(n4447), .Y(n4468) );
  INVX1 U3902 ( .A(n4468), .Y(n7354) );
  AND2X1 U3904 ( .A(n4172), .B(n4447), .Y(n4480) );
  INVX1 U3906 ( .A(n4480), .Y(n7355) );
  AND2X1 U3908 ( .A(n4110), .B(n4490), .Y(n4492) );
  INVX1 U3910 ( .A(n4492), .Y(n7356) );
  AND2X1 U3912 ( .A(n4120), .B(n4490), .Y(n4497) );
  INVX1 U3914 ( .A(n4497), .Y(n7357) );
  AND2X1 U3916 ( .A(n4112), .B(n4533), .Y(n4536) );
  INVX1 U3918 ( .A(n4536), .Y(n7358) );
  AND2X1 U3920 ( .A(n4122), .B(n4533), .Y(n4541) );
  INVX1 U3922 ( .A(n4541), .Y(n7359) );
  AND2X1 U3924 ( .A(n4114), .B(n4575), .Y(n4579) );
  INVX1 U3926 ( .A(n4579), .Y(n7360) );
  AND2X1 U3928 ( .A(n4124), .B(n4575), .Y(n4584) );
  INVX1 U3930 ( .A(n4584), .Y(n7361) );
  AND2X1 U3932 ( .A(n4116), .B(n4617), .Y(n4622) );
  INVX1 U3934 ( .A(n4622), .Y(n7362) );
  AND2X1 U3936 ( .A(n4126), .B(n4617), .Y(n4627) );
  INVX1 U3938 ( .A(n4627), .Y(n7363) );
  AND2X1 U3940 ( .A(n4150), .B(n4659), .Y(n4681) );
  INVX1 U3942 ( .A(n4681), .Y(n7364) );
  AND2X1 U3944 ( .A(n4174), .B(n4659), .Y(n4693) );
  INVX1 U3946 ( .A(n4693), .Y(n7365) );
  AND2X1 U3949 ( .A(n4128), .B(n4701), .Y(n4712) );
  INVX1 U3951 ( .A(n4712), .Y(n7366) );
  AND2X1 U3953 ( .A(n4152), .B(n4701), .Y(n4724) );
  INVX1 U3955 ( .A(n4724), .Y(n7367) );
  AND2X1 U3957 ( .A(n4176), .B(n4701), .Y(n4736) );
  INVX1 U3959 ( .A(n4736), .Y(n7368) );
  AND2X1 U3961 ( .A(n4130), .B(n4743), .Y(n4755) );
  INVX1 U3963 ( .A(n4755), .Y(n7369) );
  AND2X1 U3965 ( .A(n4154), .B(n4743), .Y(n4767) );
  INVX1 U3967 ( .A(n4767), .Y(n7370) );
  AND2X1 U3969 ( .A(n4178), .B(n4743), .Y(n4779) );
  INVX1 U3971 ( .A(n4779), .Y(n7371) );
  AND2X1 U3973 ( .A(n4132), .B(n4785), .Y(n4798) );
  INVX1 U3975 ( .A(n4798), .Y(n7372) );
  AND2X1 U3977 ( .A(n4156), .B(n4785), .Y(n4810) );
  INVX1 U3979 ( .A(n4810), .Y(n7373) );
  AND2X1 U3981 ( .A(n4180), .B(n4785), .Y(n4822) );
  INVX1 U3983 ( .A(n4822), .Y(n7374) );
  AND2X1 U3985 ( .A(n4142), .B(n4827), .Y(n4845) );
  INVX1 U3987 ( .A(n4845), .Y(n7375) );
  AND2X1 U3989 ( .A(n4166), .B(n4827), .Y(n4857) );
  INVX1 U3991 ( .A(n4857), .Y(n7376) );
  AND2X1 U3993 ( .A(n4144), .B(n4870), .Y(n4889) );
  INVX1 U3995 ( .A(n4889), .Y(n7377) );
  AND2X1 U3997 ( .A(n4168), .B(n4870), .Y(n4901) );
  INVX1 U3999 ( .A(n4901), .Y(n7378) );
  AND2X1 U4001 ( .A(n4108), .B(n4912), .Y(n4913) );
  INVX1 U4003 ( .A(n4913), .Y(n7379) );
  AND2X1 U4005 ( .A(n4146), .B(n4912), .Y(n4932) );
  INVX1 U4007 ( .A(n4932), .Y(n7380) );
  AND2X1 U4009 ( .A(n4170), .B(n4912), .Y(n4944) );
  INVX1 U4011 ( .A(n4944), .Y(n7381) );
  AND2X1 U4013 ( .A(n4148), .B(n4954), .Y(n4975) );
  INVX1 U4015 ( .A(n4975), .Y(n7382) );
  AND2X1 U4017 ( .A(n4172), .B(n4954), .Y(n4987) );
  INVX1 U4019 ( .A(n4987), .Y(n7383) );
  AND2X1 U4021 ( .A(n4110), .B(n4996), .Y(n4998) );
  INVX1 U4023 ( .A(n4998), .Y(n7384) );
  AND2X1 U4025 ( .A(n4120), .B(n4996), .Y(n5003) );
  INVX1 U4027 ( .A(n5003), .Y(n7385) );
  AND2X1 U4029 ( .A(n4112), .B(n5038), .Y(n5041) );
  INVX1 U4032 ( .A(n5041), .Y(n7386) );
  AND2X1 U4034 ( .A(n4122), .B(n5038), .Y(n5046) );
  INVX1 U4036 ( .A(n5046), .Y(n7387) );
  AND2X1 U4038 ( .A(n4114), .B(n5080), .Y(n5084) );
  INVX1 U4040 ( .A(n5084), .Y(n7388) );
  AND2X1 U4042 ( .A(n4124), .B(n5080), .Y(n5089) );
  INVX1 U4044 ( .A(n5089), .Y(n7389) );
  AND2X1 U4046 ( .A(n4116), .B(n5122), .Y(n5127) );
  INVX1 U4048 ( .A(n5127), .Y(n7390) );
  AND2X1 U4050 ( .A(n4126), .B(n5122), .Y(n5132) );
  INVX1 U4052 ( .A(n5132), .Y(n7391) );
  AND2X1 U4054 ( .A(n4142), .B(n5164), .Y(n5182) );
  INVX1 U4056 ( .A(n5182), .Y(n7392) );
  AND2X1 U4058 ( .A(n4166), .B(n5164), .Y(n5194) );
  INVX1 U4060 ( .A(n5194), .Y(n7393) );
  AND2X1 U4062 ( .A(n4144), .B(n5207), .Y(n5226) );
  INVX1 U4064 ( .A(n5226), .Y(n7394) );
  AND2X1 U4066 ( .A(n4168), .B(n5207), .Y(n5238) );
  INVX1 U4068 ( .A(n5238), .Y(n7395) );
  AND2X1 U4070 ( .A(n4108), .B(n5249), .Y(n5250) );
  INVX1 U4072 ( .A(n5250), .Y(n7396) );
  AND2X1 U4074 ( .A(n4146), .B(n5249), .Y(n5269) );
  INVX1 U4076 ( .A(n5269), .Y(n7397) );
  AND2X1 U4078 ( .A(n4170), .B(n5249), .Y(n5281) );
  INVX1 U4080 ( .A(n5281), .Y(n7398) );
  AND2X1 U4082 ( .A(n4148), .B(n5291), .Y(n5312) );
  INVX1 U4084 ( .A(n5312), .Y(n7399) );
  AND2X1 U4086 ( .A(n4172), .B(n5291), .Y(n5324) );
  INVX1 U4088 ( .A(n5324), .Y(n7400) );
  AND2X1 U4090 ( .A(n4110), .B(n5333), .Y(n5335) );
  INVX1 U4092 ( .A(n5335), .Y(n7401) );
  AND2X1 U4094 ( .A(n4120), .B(n5333), .Y(n5340) );
  INVX1 U4096 ( .A(n5340), .Y(n7402) );
  AND2X1 U4098 ( .A(n4112), .B(n5375), .Y(n5378) );
  INVX1 U4100 ( .A(n5378), .Y(n7403) );
  AND2X1 U4102 ( .A(n4122), .B(n5375), .Y(n5383) );
  INVX1 U4104 ( .A(n5383), .Y(n7404) );
  AND2X1 U4106 ( .A(n4114), .B(n5417), .Y(n5421) );
  INVX1 U4108 ( .A(n5421), .Y(n7405) );
  AND2X1 U4110 ( .A(n4124), .B(n5417), .Y(n5426) );
  INVX1 U4112 ( .A(n5426), .Y(n7406) );
  AND2X1 U4115 ( .A(n4116), .B(n5459), .Y(n5464) );
  INVX1 U4117 ( .A(n5464), .Y(n7407) );
  AND2X1 U4119 ( .A(n4126), .B(n5459), .Y(n5469) );
  INVX1 U4121 ( .A(n5469), .Y(n7408) );
  AND2X1 U4123 ( .A(n4140), .B(n4106), .Y(n4139) );
  INVX1 U4125 ( .A(n4139), .Y(n7409) );
  AND2X1 U4127 ( .A(n4164), .B(n4106), .Y(n4163) );
  INVX1 U4129 ( .A(n4163), .Y(n7410) );
  AND2X1 U4131 ( .A(n4188), .B(n4106), .Y(n4187) );
  INVX1 U4133 ( .A(n4187), .Y(n7411) );
  AND2X1 U4135 ( .A(n4138), .B(n4190), .Y(n4206) );
  INVX1 U4137 ( .A(n4206), .Y(n7412) );
  AND2X1 U4139 ( .A(n4162), .B(n4190), .Y(n4218) );
  INVX1 U4141 ( .A(n4218), .Y(n7413) );
  AND2X1 U4143 ( .A(n4186), .B(n4190), .Y(n4230) );
  INVX1 U4145 ( .A(n4230), .Y(n7414) );
  AND2X1 U4147 ( .A(n4136), .B(n4233), .Y(n4248) );
  INVX1 U4149 ( .A(n4248), .Y(n7415) );
  AND2X1 U4151 ( .A(n4160), .B(n4233), .Y(n4260) );
  INVX1 U4153 ( .A(n4260), .Y(n7416) );
  AND2X1 U4155 ( .A(n4184), .B(n4233), .Y(n4272) );
  INVX1 U4157 ( .A(n4272), .Y(n7417) );
  AND2X1 U4159 ( .A(n4134), .B(n4276), .Y(n4290) );
  INVX1 U4161 ( .A(n4290), .Y(n7418) );
  AND2X1 U4163 ( .A(n4158), .B(n4276), .Y(n4302) );
  INVX1 U4165 ( .A(n4302), .Y(n7419) );
  AND2X1 U4167 ( .A(n4182), .B(n4276), .Y(n4314) );
  INVX1 U4169 ( .A(n4314), .Y(n7420) );
  AND2X1 U4171 ( .A(n4116), .B(n4319), .Y(n4324) );
  INVX1 U4173 ( .A(n4324), .Y(n7421) );
  AND2X1 U4175 ( .A(n4126), .B(n4319), .Y(n4329) );
  INVX1 U4177 ( .A(n4329), .Y(n7422) );
  AND2X1 U4179 ( .A(n4114), .B(n4361), .Y(n4365) );
  INVX1 U4181 ( .A(n4365), .Y(n7423) );
  AND2X1 U4183 ( .A(n4124), .B(n4361), .Y(n4370) );
  INVX1 U4185 ( .A(n4370), .Y(n7424) );
  AND2X1 U4187 ( .A(n4112), .B(n4404), .Y(n4407) );
  INVX1 U4189 ( .A(n4407), .Y(n7425) );
  AND2X1 U4191 ( .A(n4122), .B(n4404), .Y(n4412) );
  INVX1 U4193 ( .A(n4412), .Y(n7426) );
  AND2X1 U4195 ( .A(n4110), .B(n4447), .Y(n4449) );
  INVX1 U4199 ( .A(n4449), .Y(n7427) );
  AND2X1 U4201 ( .A(n4120), .B(n4447), .Y(n4454) );
  INVX1 U4203 ( .A(n4454), .Y(n7428) );
  AND2X1 U4205 ( .A(n4148), .B(n4490), .Y(n4511) );
  INVX1 U4207 ( .A(n4511), .Y(n7429) );
  AND2X1 U4209 ( .A(n4172), .B(n4490), .Y(n4523) );
  INVX1 U4211 ( .A(n4523), .Y(n7430) );
  AND2X1 U4213 ( .A(n4108), .B(n4533), .Y(n4534) );
  INVX1 U4215 ( .A(n4534), .Y(n7431) );
  AND2X1 U4217 ( .A(n4146), .B(n4533), .Y(n4553) );
  INVX1 U4219 ( .A(n4553), .Y(n7432) );
  AND2X1 U4221 ( .A(n4170), .B(n4533), .Y(n4565) );
  INVX1 U4223 ( .A(n4565), .Y(n7433) );
  AND2X1 U4225 ( .A(n4144), .B(n4575), .Y(n4594) );
  INVX1 U4227 ( .A(n4594), .Y(n7434) );
  AND2X1 U4229 ( .A(n4168), .B(n4575), .Y(n4606) );
  INVX1 U4231 ( .A(n4606), .Y(n7435) );
  AND2X1 U4233 ( .A(n4142), .B(n4617), .Y(n4635) );
  INVX1 U4235 ( .A(n4635), .Y(n7436) );
  AND2X1 U4237 ( .A(n4166), .B(n4617), .Y(n4647) );
  INVX1 U4239 ( .A(n4647), .Y(n7437) );
  AND2X1 U4241 ( .A(n4140), .B(n4659), .Y(n4676) );
  INVX1 U4243 ( .A(n4676), .Y(n7438) );
  AND2X1 U4245 ( .A(n4164), .B(n4659), .Y(n4688) );
  INVX1 U4247 ( .A(n4688), .Y(n7439) );
  AND2X1 U4249 ( .A(n4188), .B(n4659), .Y(n4700) );
  INVX1 U4251 ( .A(n4700), .Y(n7440) );
  AND2X1 U4253 ( .A(n4138), .B(n4701), .Y(n4717) );
  INVX1 U4255 ( .A(n4717), .Y(n7441) );
  AND2X1 U4257 ( .A(n4162), .B(n4701), .Y(n4729) );
  INVX1 U4259 ( .A(n4729), .Y(n7442) );
  AND2X1 U4261 ( .A(n4186), .B(n4701), .Y(n4741) );
  INVX1 U4263 ( .A(n4741), .Y(n7443) );
  AND2X1 U4265 ( .A(n4136), .B(n4743), .Y(n4758) );
  INVX1 U4267 ( .A(n4758), .Y(n7444) );
  AND2X1 U4269 ( .A(n4160), .B(n4743), .Y(n4770) );
  INVX1 U4271 ( .A(n4770), .Y(n7445) );
  AND2X1 U4273 ( .A(n4184), .B(n4743), .Y(n4782) );
  INVX1 U4275 ( .A(n4782), .Y(n7446) );
  AND2X1 U4277 ( .A(n4134), .B(n4785), .Y(n4799) );
  INVX1 U4279 ( .A(n4799), .Y(n7447) );
  AND2X1 U4282 ( .A(n4158), .B(n4785), .Y(n4811) );
  INVX1 U4284 ( .A(n4811), .Y(n7448) );
  AND2X1 U4286 ( .A(n4182), .B(n4785), .Y(n4823) );
  INVX1 U4288 ( .A(n4823), .Y(n7449) );
  AND2X1 U4290 ( .A(n4116), .B(n4827), .Y(n4832) );
  INVX1 U4292 ( .A(n4832), .Y(n7450) );
  AND2X1 U4294 ( .A(n4126), .B(n4827), .Y(n4837) );
  INVX1 U4296 ( .A(n4837), .Y(n7451) );
  AND2X1 U4298 ( .A(n4114), .B(n4870), .Y(n4874) );
  INVX1 U4300 ( .A(n4874), .Y(n7452) );
  AND2X1 U4302 ( .A(n4124), .B(n4870), .Y(n4879) );
  INVX1 U4304 ( .A(n4879), .Y(n7453) );
  AND2X1 U4306 ( .A(n4112), .B(n4912), .Y(n4915) );
  INVX1 U4308 ( .A(n4915), .Y(n7454) );
  AND2X1 U4310 ( .A(n4122), .B(n4912), .Y(n4920) );
  INVX1 U4312 ( .A(n4920), .Y(n7455) );
  AND2X1 U4314 ( .A(n4110), .B(n4954), .Y(n4956) );
  INVX1 U4316 ( .A(n4956), .Y(n7456) );
  AND2X1 U4318 ( .A(n4120), .B(n4954), .Y(n4961) );
  INVX1 U4320 ( .A(n4961), .Y(n7457) );
  AND2X1 U4322 ( .A(n4148), .B(n4996), .Y(n5017) );
  INVX1 U4324 ( .A(n5017), .Y(n7458) );
  AND2X1 U4326 ( .A(n4172), .B(n4996), .Y(n5029) );
  INVX1 U4328 ( .A(n5029), .Y(n7459) );
  AND2X1 U4330 ( .A(n4108), .B(n5038), .Y(n5039) );
  INVX1 U4332 ( .A(n5039), .Y(n7460) );
  AND2X1 U4334 ( .A(n4146), .B(n5038), .Y(n5058) );
  INVX1 U4336 ( .A(n5058), .Y(n7461) );
  AND2X1 U4338 ( .A(n4170), .B(n5038), .Y(n5070) );
  INVX1 U4340 ( .A(n5070), .Y(n7462) );
  AND2X1 U4342 ( .A(n4144), .B(n5080), .Y(n5099) );
  INVX1 U4344 ( .A(n5099), .Y(n7463) );
  AND2X1 U4346 ( .A(n4168), .B(n5080), .Y(n5111) );
  INVX1 U4348 ( .A(n5111), .Y(n7464) );
  AND2X1 U4350 ( .A(n4142), .B(n5122), .Y(n5140) );
  INVX1 U4352 ( .A(n5140), .Y(n7465) );
  AND2X1 U4354 ( .A(n4166), .B(n5122), .Y(n5152) );
  INVX1 U4356 ( .A(n5152), .Y(n7466) );
  AND2X1 U4358 ( .A(n4116), .B(n5164), .Y(n5169) );
  INVX1 U4360 ( .A(n5169), .Y(n7467) );
  AND2X1 U4362 ( .A(n4126), .B(n5164), .Y(n5174) );
  INVX1 U4365 ( .A(n5174), .Y(n7468) );
  AND2X1 U4367 ( .A(n4114), .B(n5207), .Y(n5211) );
  INVX1 U4369 ( .A(n5211), .Y(n7469) );
  AND2X1 U4371 ( .A(n4124), .B(n5207), .Y(n5216) );
  INVX1 U4373 ( .A(n5216), .Y(n7470) );
  AND2X1 U4375 ( .A(n4112), .B(n5249), .Y(n5252) );
  INVX1 U4377 ( .A(n5252), .Y(n7471) );
  AND2X1 U4379 ( .A(n4122), .B(n5249), .Y(n5257) );
  INVX1 U4381 ( .A(n5257), .Y(n7472) );
  AND2X1 U4383 ( .A(n4110), .B(n5291), .Y(n5293) );
  INVX1 U4385 ( .A(n5293), .Y(n7473) );
  AND2X1 U4387 ( .A(n4120), .B(n5291), .Y(n5298) );
  INVX1 U4389 ( .A(n5298), .Y(n7474) );
  AND2X1 U4391 ( .A(n4148), .B(n5333), .Y(n5354) );
  INVX1 U4393 ( .A(n5354), .Y(n7475) );
  AND2X1 U4395 ( .A(n4172), .B(n5333), .Y(n5366) );
  INVX1 U4397 ( .A(n5366), .Y(n7476) );
  AND2X1 U4399 ( .A(n4108), .B(n5375), .Y(n5376) );
  INVX1 U4401 ( .A(n5376), .Y(n7477) );
  AND2X1 U4403 ( .A(n4146), .B(n5375), .Y(n5395) );
  INVX1 U4405 ( .A(n5395), .Y(n7478) );
  AND2X1 U4407 ( .A(n4170), .B(n5375), .Y(n5407) );
  INVX1 U4409 ( .A(n5407), .Y(n7479) );
  AND2X1 U4411 ( .A(n4144), .B(n5417), .Y(n5436) );
  INVX1 U4413 ( .A(n5436), .Y(n7480) );
  AND2X1 U4415 ( .A(n4168), .B(n5417), .Y(n5448) );
  INVX1 U4417 ( .A(n5448), .Y(n7481) );
  AND2X1 U4419 ( .A(n4142), .B(n5459), .Y(n5477) );
  INVX1 U4421 ( .A(n5477), .Y(n7482) );
  AND2X1 U4423 ( .A(n4166), .B(n5459), .Y(n5489) );
  INVX1 U4425 ( .A(n5489), .Y(n7483) );
  AND2X1 U4427 ( .A(n4138), .B(n4106), .Y(n4137) );
  INVX1 U4429 ( .A(n4137), .Y(n7484) );
  AND2X1 U4431 ( .A(n4162), .B(n4106), .Y(n4161) );
  INVX1 U4433 ( .A(n4161), .Y(n7485) );
  AND2X1 U4435 ( .A(n4186), .B(n4106), .Y(n4185) );
  INVX1 U4437 ( .A(n4185), .Y(n7486) );
  AND2X1 U4439 ( .A(n4140), .B(n4190), .Y(n4207) );
  INVX1 U4441 ( .A(n4207), .Y(n7487) );
  AND2X1 U4443 ( .A(n4164), .B(n4190), .Y(n4219) );
  INVX1 U4445 ( .A(n4219), .Y(n7488) );
  AND2X1 U4448 ( .A(n4188), .B(n4190), .Y(n4231) );
  INVX1 U4450 ( .A(n4231), .Y(n7489) );
  AND2X1 U4452 ( .A(n4134), .B(n4233), .Y(n4247) );
  INVX1 U4454 ( .A(n4247), .Y(n7490) );
  AND2X1 U4456 ( .A(n4158), .B(n4233), .Y(n4259) );
  INVX1 U4458 ( .A(n4259), .Y(n7491) );
  AND2X1 U4460 ( .A(n4182), .B(n4233), .Y(n4271) );
  INVX1 U4462 ( .A(n4271), .Y(n7492) );
  AND2X1 U4464 ( .A(n4136), .B(n4276), .Y(n4291) );
  INVX1 U4466 ( .A(n4291), .Y(n7493) );
  AND2X1 U4468 ( .A(n4160), .B(n4276), .Y(n4303) );
  INVX1 U4470 ( .A(n4303), .Y(n7494) );
  AND2X1 U4472 ( .A(n4184), .B(n4276), .Y(n4315) );
  INVX1 U4474 ( .A(n4315), .Y(n7495) );
  AND2X1 U4476 ( .A(n4114), .B(n4319), .Y(n4323) );
  INVX1 U4478 ( .A(n4323), .Y(n7496) );
  AND2X1 U4480 ( .A(n4124), .B(n4319), .Y(n4328) );
  INVX1 U4482 ( .A(n4328), .Y(n7497) );
  AND2X1 U4484 ( .A(n4116), .B(n4361), .Y(n4366) );
  INVX1 U4486 ( .A(n4366), .Y(n7498) );
  AND2X1 U4488 ( .A(n4126), .B(n4361), .Y(n4371) );
  INVX1 U4490 ( .A(n4371), .Y(n7499) );
  AND2X1 U4492 ( .A(n4110), .B(n4404), .Y(n4406) );
  INVX1 U4494 ( .A(n4406), .Y(n7500) );
  AND2X1 U4496 ( .A(n4120), .B(n4404), .Y(n4411) );
  INVX1 U4498 ( .A(n4411), .Y(n7501) );
  AND2X1 U4500 ( .A(n4112), .B(n4447), .Y(n4450) );
  INVX1 U4502 ( .A(n4450), .Y(n7502) );
  AND2X1 U4504 ( .A(n4122), .B(n4447), .Y(n4455) );
  INVX1 U4506 ( .A(n4455), .Y(n7503) );
  AND2X1 U4508 ( .A(n4108), .B(n4490), .Y(n4491) );
  INVX1 U4510 ( .A(n4491), .Y(n7504) );
  AND2X1 U4512 ( .A(n4146), .B(n4490), .Y(n4510) );
  INVX1 U4514 ( .A(n4510), .Y(n7505) );
  AND2X1 U4516 ( .A(n4170), .B(n4490), .Y(n4522) );
  INVX1 U4518 ( .A(n4522), .Y(n7506) );
  AND2X1 U4520 ( .A(n4148), .B(n4533), .Y(n4554) );
  INVX1 U4522 ( .A(n4554), .Y(n7507) );
  AND2X1 U4524 ( .A(n4172), .B(n4533), .Y(n4566) );
  INVX1 U4526 ( .A(n4566), .Y(n7508) );
  AND2X1 U4528 ( .A(n4142), .B(n4575), .Y(n4593) );
  INVX1 U4531 ( .A(n4593), .Y(n7509) );
  AND2X1 U4533 ( .A(n4166), .B(n4575), .Y(n4605) );
  INVX1 U4535 ( .A(n4605), .Y(n7510) );
  AND2X1 U4537 ( .A(n4144), .B(n4617), .Y(n4636) );
  INVX1 U4539 ( .A(n4636), .Y(n7511) );
  AND2X1 U4541 ( .A(n4168), .B(n4617), .Y(n4648) );
  INVX1 U4543 ( .A(n4648), .Y(n7512) );
  AND2X1 U4545 ( .A(n4138), .B(n4659), .Y(n4675) );
  INVX1 U4547 ( .A(n4675), .Y(n7513) );
  AND2X1 U4549 ( .A(n4162), .B(n4659), .Y(n4687) );
  INVX1 U4551 ( .A(n4687), .Y(n7514) );
  AND2X1 U4553 ( .A(n4186), .B(n4659), .Y(n4699) );
  INVX1 U4555 ( .A(n4699), .Y(n7515) );
  AND2X1 U4557 ( .A(n4140), .B(n4701), .Y(n4718) );
  INVX1 U4559 ( .A(n4718), .Y(n7516) );
  AND2X1 U4561 ( .A(n4164), .B(n4701), .Y(n4730) );
  INVX1 U4563 ( .A(n4730), .Y(n7517) );
  AND2X1 U4565 ( .A(n4188), .B(n4701), .Y(n4742) );
  INVX1 U4567 ( .A(n4742), .Y(n7518) );
  AND2X1 U4569 ( .A(n4134), .B(n4743), .Y(n4757) );
  INVX1 U4571 ( .A(n4757), .Y(n7519) );
  AND2X1 U4573 ( .A(n4158), .B(n4743), .Y(n4769) );
  INVX1 U4575 ( .A(n4769), .Y(n7520) );
  AND2X1 U4577 ( .A(n4182), .B(n4743), .Y(n4781) );
  INVX1 U4579 ( .A(n4781), .Y(n7521) );
  AND2X1 U4581 ( .A(n4136), .B(n4785), .Y(n4800) );
  INVX1 U4583 ( .A(n4800), .Y(n7522) );
  AND2X1 U4585 ( .A(n4160), .B(n4785), .Y(n4812) );
  INVX1 U4587 ( .A(n4812), .Y(n7523) );
  AND2X1 U4589 ( .A(n4184), .B(n4785), .Y(n4824) );
  INVX1 U4591 ( .A(n4824), .Y(n7524) );
  AND2X1 U4593 ( .A(n4114), .B(n4827), .Y(n4831) );
  INVX1 U4595 ( .A(n4831), .Y(n7525) );
  AND2X1 U4597 ( .A(n4124), .B(n4827), .Y(n4836) );
  INVX1 U4599 ( .A(n4836), .Y(n7526) );
  AND2X1 U4601 ( .A(n4116), .B(n4870), .Y(n4875) );
  INVX1 U4603 ( .A(n4875), .Y(n7527) );
  AND2X1 U4605 ( .A(n4126), .B(n4870), .Y(n4880) );
  INVX1 U4607 ( .A(n4880), .Y(n7528) );
  AND2X1 U4609 ( .A(n4110), .B(n4912), .Y(n4914) );
  INVX1 U4611 ( .A(n4914), .Y(n7529) );
  AND2X1 U4614 ( .A(n4120), .B(n4912), .Y(n4919) );
  INVX1 U4616 ( .A(n4919), .Y(n7530) );
  AND2X1 U4618 ( .A(n4112), .B(n4954), .Y(n4957) );
  INVX1 U4620 ( .A(n4957), .Y(n7531) );
  AND2X1 U4622 ( .A(n4122), .B(n4954), .Y(n4962) );
  INVX1 U4624 ( .A(n4962), .Y(n7532) );
  AND2X1 U4626 ( .A(n4108), .B(n4996), .Y(n4997) );
  INVX1 U4628 ( .A(n4997), .Y(n7533) );
  AND2X1 U4630 ( .A(n4146), .B(n4996), .Y(n5016) );
  INVX1 U4632 ( .A(n5016), .Y(n7534) );
  AND2X1 U4634 ( .A(n4170), .B(n4996), .Y(n5028) );
  INVX1 U4636 ( .A(n5028), .Y(n7535) );
  AND2X1 U4638 ( .A(n4148), .B(n5038), .Y(n5059) );
  INVX1 U4640 ( .A(n5059), .Y(n7536) );
  AND2X1 U4642 ( .A(n4172), .B(n5038), .Y(n5071) );
  INVX1 U4644 ( .A(n5071), .Y(n7537) );
  AND2X1 U4646 ( .A(n4142), .B(n5080), .Y(n5098) );
  INVX1 U4648 ( .A(n5098), .Y(n7538) );
  AND2X1 U4650 ( .A(n4166), .B(n5080), .Y(n5110) );
  INVX1 U4652 ( .A(n5110), .Y(n7539) );
  AND2X1 U4654 ( .A(n4144), .B(n5122), .Y(n5141) );
  INVX1 U4656 ( .A(n5141), .Y(n7540) );
  AND2X1 U4658 ( .A(n4168), .B(n5122), .Y(n5153) );
  INVX1 U4660 ( .A(n5153), .Y(n7541) );
  AND2X1 U4662 ( .A(n4114), .B(n5164), .Y(n5168) );
  INVX1 U4664 ( .A(n5168), .Y(n7542) );
  AND2X1 U4666 ( .A(n4124), .B(n5164), .Y(n5173) );
  INVX1 U4668 ( .A(n5173), .Y(n7543) );
  AND2X1 U4670 ( .A(n4116), .B(n5207), .Y(n5212) );
  INVX1 U4672 ( .A(n5212), .Y(n7544) );
  AND2X1 U4674 ( .A(n4126), .B(n5207), .Y(n5217) );
  INVX1 U4676 ( .A(n5217), .Y(n7545) );
  AND2X1 U4678 ( .A(n4110), .B(n5249), .Y(n5251) );
  INVX1 U4680 ( .A(n5251), .Y(n7546) );
  AND2X1 U4682 ( .A(n4120), .B(n5249), .Y(n5256) );
  INVX1 U4684 ( .A(n5256), .Y(n7547) );
  AND2X1 U4686 ( .A(n4112), .B(n5291), .Y(n5294) );
  INVX1 U4688 ( .A(n5294), .Y(n7548) );
  AND2X1 U4690 ( .A(n4122), .B(n5291), .Y(n5299) );
  INVX1 U4692 ( .A(n5299), .Y(n7549) );
  AND2X1 U4694 ( .A(n4108), .B(n5333), .Y(n5334) );
  INVX1 U4697 ( .A(n5334), .Y(n7550) );
  AND2X1 U4699 ( .A(n4146), .B(n5333), .Y(n5353) );
  INVX1 U4701 ( .A(n5353), .Y(n7551) );
  AND2X1 U4703 ( .A(n4170), .B(n5333), .Y(n5365) );
  INVX1 U4705 ( .A(n5365), .Y(n7552) );
  AND2X1 U4707 ( .A(n4148), .B(n5375), .Y(n5396) );
  INVX1 U4709 ( .A(n5396), .Y(n7553) );
  AND2X1 U4711 ( .A(n4172), .B(n5375), .Y(n5408) );
  INVX1 U4713 ( .A(n5408), .Y(n7554) );
  AND2X1 U4715 ( .A(n4142), .B(n5417), .Y(n5435) );
  INVX1 U4717 ( .A(n5435), .Y(n7555) );
  AND2X1 U4719 ( .A(n4166), .B(n5417), .Y(n5447) );
  INVX1 U4721 ( .A(n5447), .Y(n7556) );
  AND2X1 U4723 ( .A(n4144), .B(n5459), .Y(n5478) );
  INVX1 U4725 ( .A(n5478), .Y(n7557) );
  AND2X1 U4727 ( .A(n4168), .B(n5459), .Y(n5490) );
  INVX1 U4729 ( .A(n5490), .Y(n7558) );
  AND2X1 U4731 ( .A(n4136), .B(n4106), .Y(n4135) );
  INVX1 U4733 ( .A(n4135), .Y(n7559) );
  AND2X1 U4735 ( .A(n4160), .B(n4106), .Y(n4159) );
  INVX1 U4737 ( .A(n4159), .Y(n7560) );
  AND2X1 U4739 ( .A(n4184), .B(n4106), .Y(n4183) );
  INVX1 U4741 ( .A(n4183), .Y(n7561) );
  AND2X1 U4743 ( .A(n4134), .B(n4190), .Y(n4204) );
  INVX1 U4745 ( .A(n4204), .Y(n7562) );
  AND2X1 U4747 ( .A(n4158), .B(n4190), .Y(n4216) );
  INVX1 U4749 ( .A(n4216), .Y(n7563) );
  AND2X1 U4751 ( .A(n4182), .B(n4190), .Y(n4228) );
  INVX1 U4753 ( .A(n4228), .Y(n7564) );
  AND2X1 U4755 ( .A(n4140), .B(n4233), .Y(n4250) );
  INVX1 U4757 ( .A(n4250), .Y(n7565) );
  AND2X1 U4759 ( .A(n4164), .B(n4233), .Y(n4262) );
  INVX1 U4761 ( .A(n4262), .Y(n7566) );
  AND2X1 U4763 ( .A(n4188), .B(n4233), .Y(n4274) );
  INVX1 U4765 ( .A(n4274), .Y(n7567) );
  AND2X1 U4767 ( .A(n4138), .B(n4276), .Y(n4292) );
  INVX1 U4769 ( .A(n4292), .Y(n7568) );
  AND2X1 U4771 ( .A(n4162), .B(n4276), .Y(n4304) );
  INVX1 U4773 ( .A(n4304), .Y(n7569) );
  AND2X1 U4775 ( .A(n4186), .B(n4276), .Y(n4316) );
  INVX1 U4777 ( .A(n4316), .Y(n7570) );
  AND2X1 U4780 ( .A(n4112), .B(n4319), .Y(n4322) );
  INVX1 U4782 ( .A(n4322), .Y(n7571) );
  AND2X1 U4784 ( .A(n4122), .B(n4319), .Y(n4327) );
  INVX1 U4786 ( .A(n4327), .Y(n7572) );
  AND2X1 U4788 ( .A(n4110), .B(n4361), .Y(n4363) );
  INVX1 U4790 ( .A(n4363), .Y(n7573) );
  AND2X1 U4792 ( .A(n4120), .B(n4361), .Y(n4368) );
  INVX1 U4794 ( .A(n4368), .Y(n7574) );
  AND2X1 U4796 ( .A(n4116), .B(n4404), .Y(n4409) );
  INVX1 U4798 ( .A(n4409), .Y(n7575) );
  AND2X1 U4800 ( .A(n4126), .B(n4404), .Y(n4414) );
  INVX1 U4802 ( .A(n4414), .Y(n7576) );
  AND2X1 U4804 ( .A(n4114), .B(n4447), .Y(n4451) );
  INVX1 U4806 ( .A(n4451), .Y(n7577) );
  AND2X1 U4808 ( .A(n4124), .B(n4447), .Y(n4456) );
  INVX1 U4810 ( .A(n4456), .Y(n7578) );
  AND2X1 U4812 ( .A(n4144), .B(n4490), .Y(n4509) );
  INVX1 U4814 ( .A(n4509), .Y(n7579) );
  AND2X1 U4816 ( .A(n4168), .B(n4490), .Y(n4521) );
  INVX1 U4818 ( .A(n4521), .Y(n7580) );
  AND2X1 U4820 ( .A(n4142), .B(n4533), .Y(n4551) );
  INVX1 U4822 ( .A(n4551), .Y(n7581) );
  AND2X1 U4824 ( .A(n4166), .B(n4533), .Y(n4563) );
  INVX1 U4826 ( .A(n4563), .Y(n7582) );
  AND2X1 U4828 ( .A(n4148), .B(n4575), .Y(n4596) );
  INVX1 U4830 ( .A(n4596), .Y(n7583) );
  AND2X1 U4832 ( .A(n4172), .B(n4575), .Y(n4608) );
  INVX1 U4834 ( .A(n4608), .Y(n7584) );
  AND2X1 U4836 ( .A(n4108), .B(n4617), .Y(n4618) );
  INVX1 U4838 ( .A(n4618), .Y(n7585) );
  AND2X1 U4840 ( .A(n4146), .B(n4617), .Y(n4637) );
  INVX1 U4842 ( .A(n4637), .Y(n7586) );
  AND2X1 U4844 ( .A(n4170), .B(n4617), .Y(n4649) );
  INVX1 U4846 ( .A(n4649), .Y(n7587) );
  AND2X1 U4848 ( .A(n4136), .B(n4659), .Y(n4674) );
  INVX1 U4850 ( .A(n4674), .Y(n7588) );
  AND2X1 U4852 ( .A(n4160), .B(n4659), .Y(n4686) );
  INVX1 U4854 ( .A(n4686), .Y(n7589) );
  AND2X1 U4856 ( .A(n4184), .B(n4659), .Y(n4698) );
  INVX1 U4858 ( .A(n4698), .Y(n7590) );
  AND2X1 U4860 ( .A(n4134), .B(n4701), .Y(n4715) );
  INVX1 U4864 ( .A(n4715), .Y(n7591) );
  AND2X1 U4866 ( .A(n4158), .B(n4701), .Y(n4727) );
  INVX1 U4868 ( .A(n4727), .Y(n7592) );
  AND2X1 U4870 ( .A(n4182), .B(n4701), .Y(n4739) );
  INVX1 U4872 ( .A(n4739), .Y(n7593) );
  AND2X1 U4874 ( .A(n4140), .B(n4743), .Y(n4760) );
  INVX1 U4876 ( .A(n4760), .Y(n7594) );
  AND2X1 U4878 ( .A(n4164), .B(n4743), .Y(n4772) );
  INVX1 U4880 ( .A(n4772), .Y(n7595) );
  AND2X1 U4882 ( .A(n4188), .B(n4743), .Y(n4784) );
  INVX1 U4884 ( .A(n4784), .Y(n7596) );
  AND2X1 U4886 ( .A(n4138), .B(n4785), .Y(n4801) );
  INVX1 U4888 ( .A(n4801), .Y(n7597) );
  AND2X1 U4890 ( .A(n4162), .B(n4785), .Y(n4813) );
  INVX1 U4892 ( .A(n4813), .Y(n7598) );
  AND2X1 U4894 ( .A(n4186), .B(n4785), .Y(n4825) );
  INVX1 U4896 ( .A(n4825), .Y(n7599) );
  AND2X1 U4898 ( .A(n4112), .B(n4827), .Y(n4830) );
  INVX1 U4900 ( .A(n4830), .Y(n7600) );
  AND2X1 U4902 ( .A(n4122), .B(n4827), .Y(n4835) );
  INVX1 U4904 ( .A(n4835), .Y(n7601) );
  AND2X1 U4906 ( .A(n4110), .B(n4870), .Y(n4872) );
  INVX1 U4908 ( .A(n4872), .Y(n7602) );
  AND2X1 U4910 ( .A(n4120), .B(n4870), .Y(n4877) );
  INVX1 U4912 ( .A(n4877), .Y(n7603) );
  AND2X1 U4914 ( .A(n4116), .B(n4912), .Y(n4917) );
  INVX1 U4916 ( .A(n4917), .Y(n7604) );
  AND2X1 U4918 ( .A(n4126), .B(n4912), .Y(n4922) );
  INVX1 U4920 ( .A(n4922), .Y(n7605) );
  AND2X1 U4922 ( .A(n4114), .B(n4954), .Y(n4958) );
  INVX1 U4924 ( .A(n4958), .Y(n7606) );
  AND2X1 U4926 ( .A(n4124), .B(n4954), .Y(n4963) );
  INVX1 U4928 ( .A(n4963), .Y(n7607) );
  AND2X1 U4930 ( .A(n4144), .B(n4996), .Y(n5015) );
  INVX1 U4932 ( .A(n5015), .Y(n7608) );
  AND2X1 U4934 ( .A(n4168), .B(n4996), .Y(n5027) );
  INVX1 U4936 ( .A(n5027), .Y(n7609) );
  AND2X1 U4938 ( .A(n4142), .B(n5038), .Y(n5056) );
  INVX1 U4940 ( .A(n5056), .Y(n7610) );
  AND2X1 U4942 ( .A(n4166), .B(n5038), .Y(n5068) );
  INVX1 U4944 ( .A(n5068), .Y(n7611) );
  AND2X1 U4948 ( .A(n4148), .B(n5080), .Y(n5101) );
  INVX1 U4950 ( .A(n5101), .Y(n7612) );
  AND2X1 U4952 ( .A(n4172), .B(n5080), .Y(n5113) );
  INVX1 U4954 ( .A(n5113), .Y(n7613) );
  AND2X1 U4956 ( .A(n4108), .B(n5122), .Y(n5123) );
  INVX1 U4958 ( .A(n5123), .Y(n7614) );
  AND2X1 U4960 ( .A(n4146), .B(n5122), .Y(n5142) );
  INVX1 U4962 ( .A(n5142), .Y(n7615) );
  AND2X1 U4964 ( .A(n4170), .B(n5122), .Y(n5154) );
  INVX1 U4966 ( .A(n5154), .Y(n7616) );
  AND2X1 U4968 ( .A(n4112), .B(n5164), .Y(n5167) );
  INVX1 U4970 ( .A(n5167), .Y(n7617) );
  AND2X1 U4972 ( .A(n4122), .B(n5164), .Y(n5172) );
  INVX1 U4974 ( .A(n5172), .Y(n7618) );
  AND2X1 U4976 ( .A(n4110), .B(n5207), .Y(n5209) );
  INVX1 U4978 ( .A(n5209), .Y(n7619) );
  AND2X1 U4980 ( .A(n4120), .B(n5207), .Y(n5214) );
  INVX1 U4982 ( .A(n5214), .Y(n7620) );
  AND2X1 U4984 ( .A(n4116), .B(n5249), .Y(n5254) );
  INVX1 U4986 ( .A(n5254), .Y(n7621) );
  AND2X1 U4988 ( .A(n4126), .B(n5249), .Y(n5259) );
  INVX1 U4990 ( .A(n5259), .Y(n7622) );
  AND2X1 U4992 ( .A(n4114), .B(n5291), .Y(n5295) );
  INVX1 U4994 ( .A(n5295), .Y(n7623) );
  AND2X1 U4996 ( .A(n4124), .B(n5291), .Y(n5300) );
  INVX1 U4998 ( .A(n5300), .Y(n7624) );
  AND2X1 U5000 ( .A(n4144), .B(n5333), .Y(n5352) );
  INVX1 U5002 ( .A(n5352), .Y(n7625) );
  AND2X1 U5004 ( .A(n4168), .B(n5333), .Y(n5364) );
  INVX1 U5006 ( .A(n5364), .Y(n7626) );
  AND2X1 U5008 ( .A(n4142), .B(n5375), .Y(n5393) );
  INVX1 U5010 ( .A(n5393), .Y(n7627) );
  AND2X1 U5012 ( .A(n4166), .B(n5375), .Y(n5405) );
  INVX1 U5014 ( .A(n5405), .Y(n7628) );
  AND2X1 U5016 ( .A(n4148), .B(n5417), .Y(n5438) );
  INVX1 U5018 ( .A(n5438), .Y(n7629) );
  AND2X1 U5020 ( .A(n4172), .B(n5417), .Y(n5450) );
  INVX1 U5022 ( .A(n5450), .Y(n7630) );
  AND2X1 U5024 ( .A(n4108), .B(n5459), .Y(n5460) );
  INVX1 U5026 ( .A(n5460), .Y(n7631) );
  AND2X1 U5028 ( .A(n4146), .B(n5459), .Y(n5479) );
  INVX1 U5032 ( .A(n5479), .Y(n7632) );
  AND2X1 U5034 ( .A(n4170), .B(n5459), .Y(n5491) );
  INVX1 U5036 ( .A(n5491), .Y(n7633) );
  AND2X1 U5038 ( .A(n4134), .B(n4106), .Y(n4133) );
  INVX1 U5040 ( .A(n4133), .Y(n7634) );
  AND2X1 U5042 ( .A(n4158), .B(n4106), .Y(n4157) );
  INVX1 U5044 ( .A(n4157), .Y(n7635) );
  AND2X1 U5046 ( .A(n4182), .B(n4106), .Y(n4181) );
  INVX1 U5048 ( .A(n4181), .Y(n7636) );
  AND2X1 U5050 ( .A(n4136), .B(n4190), .Y(n4205) );
  INVX1 U5052 ( .A(n4205), .Y(n7637) );
  AND2X1 U5054 ( .A(n4160), .B(n4190), .Y(n4217) );
  INVX1 U5056 ( .A(n4217), .Y(n7638) );
  AND2X1 U5058 ( .A(n4184), .B(n4190), .Y(n4229) );
  INVX1 U5060 ( .A(n4229), .Y(n7639) );
  AND2X1 U5062 ( .A(n4138), .B(n4233), .Y(n4249) );
  INVX1 U5064 ( .A(n4249), .Y(n7640) );
  AND2X1 U5066 ( .A(n4162), .B(n4233), .Y(n4261) );
  INVX1 U5068 ( .A(n4261), .Y(n7641) );
  AND2X1 U5070 ( .A(n4186), .B(n4233), .Y(n4273) );
  INVX1 U5072 ( .A(n4273), .Y(n7642) );
  AND2X1 U5074 ( .A(n4140), .B(n4276), .Y(n4293) );
  INVX1 U5076 ( .A(n4293), .Y(n7643) );
  AND2X1 U5078 ( .A(n4164), .B(n4276), .Y(n4305) );
  INVX1 U5080 ( .A(n4305), .Y(n7644) );
  AND2X1 U5082 ( .A(n4188), .B(n4276), .Y(n4317) );
  INVX1 U5084 ( .A(n4317), .Y(n7645) );
  AND2X1 U5086 ( .A(n4110), .B(n4319), .Y(n4321) );
  INVX1 U5088 ( .A(n4321), .Y(n7646) );
  AND2X1 U5090 ( .A(n4120), .B(n4319), .Y(n4326) );
  INVX1 U5092 ( .A(n4326), .Y(n7647) );
  AND2X1 U5094 ( .A(n4112), .B(n4361), .Y(n4364) );
  INVX1 U5096 ( .A(n4364), .Y(n7648) );
  AND2X1 U5098 ( .A(n4122), .B(n4361), .Y(n4369) );
  INVX1 U5100 ( .A(n4369), .Y(n7649) );
  AND2X1 U5102 ( .A(n4114), .B(n4404), .Y(n4408) );
  INVX1 U5104 ( .A(n4408), .Y(n7650) );
  AND2X1 U5106 ( .A(n4124), .B(n4404), .Y(n4413) );
  INVX1 U5108 ( .A(n4413), .Y(n7651) );
  AND2X1 U5110 ( .A(n4116), .B(n4447), .Y(n4452) );
  INVX1 U5112 ( .A(n4452), .Y(n7652) );
  AND2X1 U5116 ( .A(n4126), .B(n4447), .Y(n4457) );
  INVX1 U5118 ( .A(n4457), .Y(n7653) );
  AND2X1 U5120 ( .A(n4142), .B(n4490), .Y(n4508) );
  INVX1 U5122 ( .A(n4508), .Y(n7654) );
  AND2X1 U5124 ( .A(n4166), .B(n4490), .Y(n4520) );
  INVX1 U5126 ( .A(n4520), .Y(n7655) );
  AND2X1 U5128 ( .A(n4144), .B(n4533), .Y(n4552) );
  INVX1 U5130 ( .A(n4552), .Y(n7656) );
  AND2X1 U5132 ( .A(n4168), .B(n4533), .Y(n4564) );
  INVX1 U5134 ( .A(n4564), .Y(n7657) );
  AND2X1 U5136 ( .A(n4108), .B(n4575), .Y(n4576) );
  INVX1 U5138 ( .A(n4576), .Y(n7658) );
  AND2X1 U5140 ( .A(n4146), .B(n4575), .Y(n4595) );
  INVX1 U5142 ( .A(n4595), .Y(n7659) );
  AND2X1 U5144 ( .A(n4170), .B(n4575), .Y(n4607) );
  INVX1 U5146 ( .A(n4607), .Y(n7660) );
  AND2X1 U5148 ( .A(n4148), .B(n4617), .Y(n4638) );
  INVX1 U5150 ( .A(n4638), .Y(n7661) );
  AND2X1 U5152 ( .A(n4172), .B(n4617), .Y(n4650) );
  INVX1 U5154 ( .A(n4650), .Y(n7662) );
  AND2X1 U5156 ( .A(n4134), .B(n4659), .Y(n4673) );
  INVX1 U5158 ( .A(n4673), .Y(n7663) );
  AND2X1 U5160 ( .A(n4158), .B(n4659), .Y(n4685) );
  INVX1 U5162 ( .A(n4685), .Y(n7664) );
  AND2X1 U5164 ( .A(n4182), .B(n4659), .Y(n4697) );
  INVX1 U5166 ( .A(n4697), .Y(n7665) );
  AND2X1 U5168 ( .A(n4136), .B(n4701), .Y(n4716) );
  INVX1 U5170 ( .A(n4716), .Y(n7666) );
  AND2X1 U5172 ( .A(n4160), .B(n4701), .Y(n4728) );
  INVX1 U5174 ( .A(n4728), .Y(n7667) );
  AND2X1 U5176 ( .A(n4184), .B(n4701), .Y(n4740) );
  INVX1 U5178 ( .A(n4740), .Y(n7668) );
  AND2X1 U5180 ( .A(n4138), .B(n4743), .Y(n4759) );
  INVX1 U5182 ( .A(n4759), .Y(n7669) );
  AND2X1 U5184 ( .A(n4162), .B(n4743), .Y(n4771) );
  INVX1 U5186 ( .A(n4771), .Y(n7670) );
  AND2X1 U5188 ( .A(n4186), .B(n4743), .Y(n4783) );
  INVX1 U5190 ( .A(n4783), .Y(n7671) );
  AND2X1 U5192 ( .A(n4140), .B(n4785), .Y(n4802) );
  INVX1 U5194 ( .A(n4802), .Y(n7672) );
  AND2X1 U5196 ( .A(n4164), .B(n4785), .Y(n4814) );
  INVX1 U5200 ( .A(n4814), .Y(n7673) );
  AND2X1 U5202 ( .A(n4188), .B(n4785), .Y(n4826) );
  INVX1 U5204 ( .A(n4826), .Y(n7674) );
  AND2X1 U5206 ( .A(n4110), .B(n4827), .Y(n4829) );
  INVX1 U5208 ( .A(n4829), .Y(n7675) );
  AND2X1 U5210 ( .A(n4120), .B(n4827), .Y(n4834) );
  INVX1 U5212 ( .A(n4834), .Y(n7676) );
  AND2X1 U5214 ( .A(n4112), .B(n4870), .Y(n4873) );
  INVX1 U5216 ( .A(n4873), .Y(n7677) );
  AND2X1 U5218 ( .A(n4122), .B(n4870), .Y(n4878) );
  INVX1 U5220 ( .A(n4878), .Y(n7678) );
  AND2X1 U5222 ( .A(n4114), .B(n4912), .Y(n4916) );
  INVX1 U5224 ( .A(n4916), .Y(n7679) );
  AND2X1 U5226 ( .A(n4124), .B(n4912), .Y(n4921) );
  INVX1 U5228 ( .A(n4921), .Y(n7680) );
  AND2X1 U5230 ( .A(n4116), .B(n4954), .Y(n4959) );
  INVX1 U5232 ( .A(n4959), .Y(n7681) );
  AND2X1 U5234 ( .A(n4126), .B(n4954), .Y(n4964) );
  INVX1 U5236 ( .A(n4964), .Y(n7682) );
  AND2X1 U5238 ( .A(n4142), .B(n4996), .Y(n5014) );
  INVX1 U5240 ( .A(n5014), .Y(n7683) );
  AND2X1 U5242 ( .A(n4166), .B(n4996), .Y(n5026) );
  INVX1 U5244 ( .A(n5026), .Y(n7684) );
  AND2X1 U5246 ( .A(n4144), .B(n5038), .Y(n5057) );
  INVX1 U5248 ( .A(n5057), .Y(n7685) );
  AND2X1 U5250 ( .A(n4168), .B(n5038), .Y(n5069) );
  INVX1 U5252 ( .A(n5069), .Y(n7686) );
  AND2X1 U5254 ( .A(n4108), .B(n5080), .Y(n5081) );
  INVX1 U5256 ( .A(n5081), .Y(n7687) );
  AND2X1 U5258 ( .A(n4146), .B(n5080), .Y(n5100) );
  INVX1 U5260 ( .A(n5100), .Y(n7688) );
  AND2X1 U5262 ( .A(n4170), .B(n5080), .Y(n5112) );
  INVX1 U5264 ( .A(n5112), .Y(n7689) );
  AND2X1 U5266 ( .A(n4148), .B(n5122), .Y(n5143) );
  INVX1 U5268 ( .A(n5143), .Y(n7690) );
  AND2X1 U5270 ( .A(n4172), .B(n5122), .Y(n5155) );
  INVX1 U5272 ( .A(n5155), .Y(n7691) );
  AND2X1 U5274 ( .A(n4110), .B(n5164), .Y(n5166) );
  INVX1 U5276 ( .A(n5166), .Y(n7692) );
  AND2X1 U5278 ( .A(n4120), .B(n5164), .Y(n5171) );
  INVX1 U5280 ( .A(n5171), .Y(n7693) );
  AND2X1 U5284 ( .A(n4112), .B(n5207), .Y(n5210) );
  INVX1 U5286 ( .A(n5210), .Y(n7694) );
  AND2X1 U5288 ( .A(n4122), .B(n5207), .Y(n5215) );
  INVX1 U5290 ( .A(n5215), .Y(n7695) );
  AND2X1 U5292 ( .A(n4114), .B(n5249), .Y(n5253) );
  INVX1 U5294 ( .A(n5253), .Y(n7696) );
  AND2X1 U5296 ( .A(n4124), .B(n5249), .Y(n5258) );
  INVX1 U5298 ( .A(n5258), .Y(n7697) );
  AND2X1 U5300 ( .A(n4116), .B(n5291), .Y(n5296) );
  INVX1 U5302 ( .A(n5296), .Y(n7698) );
  AND2X1 U5304 ( .A(n4126), .B(n5291), .Y(n5301) );
  INVX1 U5306 ( .A(n5301), .Y(n7699) );
  AND2X1 U5308 ( .A(n4142), .B(n5333), .Y(n5351) );
  INVX1 U5310 ( .A(n5351), .Y(n7700) );
  AND2X1 U5312 ( .A(n4166), .B(n5333), .Y(n5363) );
  INVX1 U5314 ( .A(n5363), .Y(n7701) );
  AND2X1 U5316 ( .A(n4144), .B(n5375), .Y(n5394) );
  INVX1 U5318 ( .A(n5394), .Y(n7702) );
  AND2X1 U5320 ( .A(n4168), .B(n5375), .Y(n5406) );
  INVX1 U5322 ( .A(n5406), .Y(n7703) );
  AND2X1 U5324 ( .A(n4108), .B(n5417), .Y(n5418) );
  INVX1 U5326 ( .A(n5418), .Y(n7704) );
  AND2X1 U5328 ( .A(n4146), .B(n5417), .Y(n5437) );
  INVX1 U5330 ( .A(n5437), .Y(n7705) );
  AND2X1 U5332 ( .A(n4170), .B(n5417), .Y(n5449) );
  INVX1 U5334 ( .A(n5449), .Y(n7706) );
  AND2X1 U5336 ( .A(n4148), .B(n5459), .Y(n5480) );
  INVX1 U5338 ( .A(n5480), .Y(n7707) );
  AND2X1 U5340 ( .A(n4172), .B(n5459), .Y(n5492) );
  INVX1 U5342 ( .A(n5492), .Y(n7708) );
  BUFX2 U5344 ( .A(n4099), .Y(n7709) );
  AND2X1 U5346 ( .A(n4116), .B(n4106), .Y(n4115) );
  INVX1 U5348 ( .A(n4115), .Y(n7710) );
  AND2X1 U5350 ( .A(n4126), .B(n4106), .Y(n4125) );
  INVX1 U5352 ( .A(n4125), .Y(n7711) );
  AND2X1 U5354 ( .A(n4114), .B(n4190), .Y(n4194) );
  INVX1 U5356 ( .A(n4194), .Y(n7712) );
  AND2X1 U5358 ( .A(n4124), .B(n4190), .Y(n4199) );
  INVX1 U5360 ( .A(n4199), .Y(n7713) );
  AND2X1 U5362 ( .A(n4112), .B(n4233), .Y(n4236) );
  INVX1 U5364 ( .A(n4236), .Y(n7714) );
  AND2X1 U5368 ( .A(n4122), .B(n4233), .Y(n4241) );
  INVX1 U5370 ( .A(n4241), .Y(n7715) );
  AND2X1 U5372 ( .A(n4110), .B(n4276), .Y(n4278) );
  INVX1 U5374 ( .A(n4278), .Y(n7716) );
  AND2X1 U5376 ( .A(n4120), .B(n4276), .Y(n4283) );
  INVX1 U5378 ( .A(n4283), .Y(n7717) );
  AND2X1 U5380 ( .A(n4140), .B(n4319), .Y(n4336) );
  INVX1 U5382 ( .A(n4336), .Y(n7718) );
  AND2X1 U5384 ( .A(n4164), .B(n4319), .Y(n4348) );
  INVX1 U5386 ( .A(n4348), .Y(n7719) );
  AND2X1 U5388 ( .A(n4188), .B(n4319), .Y(n4360) );
  INVX1 U5390 ( .A(n4360), .Y(n7720) );
  AND2X1 U5392 ( .A(n4138), .B(n4361), .Y(n4377) );
  INVX1 U5394 ( .A(n4377), .Y(n7721) );
  AND2X1 U5396 ( .A(n4162), .B(n4361), .Y(n4389) );
  INVX1 U5398 ( .A(n4389), .Y(n7722) );
  AND2X1 U5400 ( .A(n4186), .B(n4361), .Y(n4401) );
  INVX1 U5402 ( .A(n4401), .Y(n7723) );
  AND2X1 U5404 ( .A(n4136), .B(n4404), .Y(n4419) );
  INVX1 U5406 ( .A(n4419), .Y(n7724) );
  AND2X1 U5408 ( .A(n4160), .B(n4404), .Y(n4431) );
  INVX1 U5410 ( .A(n4431), .Y(n7725) );
  AND2X1 U5412 ( .A(n4184), .B(n4404), .Y(n4443) );
  INVX1 U5414 ( .A(n4443), .Y(n7726) );
  AND2X1 U5416 ( .A(n4134), .B(n4447), .Y(n4461) );
  INVX1 U5418 ( .A(n4461), .Y(n7727) );
  AND2X1 U5420 ( .A(n4158), .B(n4447), .Y(n4473) );
  INVX1 U5422 ( .A(n4473), .Y(n7728) );
  AND2X1 U5424 ( .A(n4182), .B(n4447), .Y(n4485) );
  INVX1 U5426 ( .A(n4485), .Y(n7729) );
  AND2X1 U5428 ( .A(n4132), .B(n4490), .Y(n4503) );
  INVX1 U5430 ( .A(n4503), .Y(n7730) );
  AND2X1 U5432 ( .A(n4156), .B(n4490), .Y(n4515) );
  INVX1 U5434 ( .A(n4515), .Y(n7731) );
  AND2X1 U5436 ( .A(n4180), .B(n4490), .Y(n4527) );
  INVX1 U5438 ( .A(n4527), .Y(n7732) );
  AND2X1 U5440 ( .A(n4130), .B(n4533), .Y(n4545) );
  INVX1 U5442 ( .A(n4545), .Y(n7733) );
  AND2X1 U5444 ( .A(n4154), .B(n4533), .Y(n4557) );
  INVX1 U5446 ( .A(n4557), .Y(n7734) );
  AND2X1 U5448 ( .A(n4178), .B(n4533), .Y(n4569) );
  INVX1 U5452 ( .A(n4569), .Y(n7735) );
  AND2X1 U5454 ( .A(n4128), .B(n4575), .Y(n4586) );
  INVX1 U5456 ( .A(n4586), .Y(n7736) );
  AND2X1 U5458 ( .A(n4152), .B(n4575), .Y(n4598) );
  INVX1 U5460 ( .A(n4598), .Y(n7737) );
  AND2X1 U5462 ( .A(n4176), .B(n4575), .Y(n4610) );
  INVX1 U5464 ( .A(n4610), .Y(n7738) );
  AND2X1 U5466 ( .A(n4150), .B(n4617), .Y(n4639) );
  INVX1 U5468 ( .A(n4639), .Y(n7739) );
  AND2X1 U5470 ( .A(n4174), .B(n4617), .Y(n4651) );
  INVX1 U5472 ( .A(n4651), .Y(n7740) );
  AND2X1 U5474 ( .A(n4116), .B(n4659), .Y(n4664) );
  INVX1 U5476 ( .A(n4664), .Y(n7741) );
  AND2X1 U5478 ( .A(n4126), .B(n4659), .Y(n4669) );
  INVX1 U5480 ( .A(n4669), .Y(n7742) );
  AND2X1 U5482 ( .A(n4114), .B(n4701), .Y(n4705) );
  INVX1 U5484 ( .A(n4705), .Y(n7743) );
  AND2X1 U5486 ( .A(n4124), .B(n4701), .Y(n4710) );
  INVX1 U5488 ( .A(n4710), .Y(n7744) );
  AND2X1 U5490 ( .A(n4112), .B(n4743), .Y(n4746) );
  INVX1 U5492 ( .A(n4746), .Y(n7745) );
  AND2X1 U5494 ( .A(n4122), .B(n4743), .Y(n4751) );
  INVX1 U5496 ( .A(n4751), .Y(n7746) );
  AND2X1 U5498 ( .A(n4110), .B(n4785), .Y(n4787) );
  INVX1 U5500 ( .A(n4787), .Y(n7747) );
  AND2X1 U5502 ( .A(n4120), .B(n4785), .Y(n4792) );
  INVX1 U5504 ( .A(n4792), .Y(n7748) );
  AND2X1 U5506 ( .A(n4140), .B(n4827), .Y(n4844) );
  INVX1 U5508 ( .A(n4844), .Y(n7749) );
  AND2X1 U5510 ( .A(n4164), .B(n4827), .Y(n4856) );
  INVX1 U5512 ( .A(n4856), .Y(n7750) );
  AND2X1 U5514 ( .A(n4188), .B(n4827), .Y(n4868) );
  INVX1 U5516 ( .A(n4868), .Y(n7751) );
  AND2X1 U5518 ( .A(n4138), .B(n4870), .Y(n4886) );
  INVX1 U5520 ( .A(n4886), .Y(n7752) );
  AND2X1 U5522 ( .A(n4162), .B(n4870), .Y(n4898) );
  INVX1 U5524 ( .A(n4898), .Y(n7753) );
  AND2X1 U5526 ( .A(n4186), .B(n4870), .Y(n4910) );
  INVX1 U5528 ( .A(n4910), .Y(n7754) );
  AND2X1 U5530 ( .A(n4136), .B(n4912), .Y(n4927) );
  INVX1 U5532 ( .A(n4927), .Y(n7755) );
  AND2X1 U5551 ( .A(n4160), .B(n4912), .Y(n4939) );
  INVX1 U5552 ( .A(n4939), .Y(n7756) );
  AND2X1 U5553 ( .A(n4184), .B(n4912), .Y(n4951) );
  INVX1 U5554 ( .A(n4951), .Y(n7757) );
  AND2X1 U5555 ( .A(n4134), .B(n4954), .Y(n4968) );
  INVX1 U5556 ( .A(n4968), .Y(n7758) );
  AND2X1 U5557 ( .A(n4158), .B(n4954), .Y(n4980) );
  INVX1 U5558 ( .A(n4980), .Y(n7759) );
  AND2X1 U5559 ( .A(n4182), .B(n4954), .Y(n4992) );
  INVX1 U5560 ( .A(n4992), .Y(n7760) );
  AND2X1 U5561 ( .A(n4132), .B(n4996), .Y(n5009) );
  INVX1 U5562 ( .A(n5009), .Y(n7761) );
  AND2X1 U5563 ( .A(n4156), .B(n4996), .Y(n5021) );
  INVX1 U5564 ( .A(n5021), .Y(n7762) );
  AND2X1 U5565 ( .A(n4180), .B(n4996), .Y(n5033) );
  INVX1 U5566 ( .A(n5033), .Y(n7763) );
  AND2X1 U5567 ( .A(n4130), .B(n5038), .Y(n5050) );
  INVX1 U5568 ( .A(n5050), .Y(n7764) );
  AND2X1 U5569 ( .A(n4154), .B(n5038), .Y(n5062) );
  INVX1 U5570 ( .A(n5062), .Y(n7765) );
  AND2X1 U5571 ( .A(n4178), .B(n5038), .Y(n5074) );
  INVX1 U5572 ( .A(n5074), .Y(n7766) );
  AND2X1 U5573 ( .A(n4128), .B(n5080), .Y(n5091) );
  INVX1 U5574 ( .A(n5091), .Y(n7767) );
  AND2X1 U5575 ( .A(n4152), .B(n5080), .Y(n5103) );
  INVX1 U5576 ( .A(n5103), .Y(n7768) );
  AND2X1 U5577 ( .A(n4176), .B(n5080), .Y(n5115) );
  INVX1 U5578 ( .A(n5115), .Y(n7769) );
  AND2X1 U5579 ( .A(n4150), .B(n5122), .Y(n5144) );
  INVX1 U5580 ( .A(n5144), .Y(n7770) );
  AND2X1 U5581 ( .A(n4174), .B(n5122), .Y(n5156) );
  INVX1 U5582 ( .A(n5156), .Y(n7771) );
  AND2X1 U5583 ( .A(n4140), .B(n5164), .Y(n5181) );
  INVX1 U5584 ( .A(n5181), .Y(n7772) );
  AND2X1 U5585 ( .A(n4164), .B(n5164), .Y(n5193) );
  INVX1 U5586 ( .A(n5193), .Y(n7773) );
  AND2X1 U5587 ( .A(n4188), .B(n5164), .Y(n5205) );
  INVX1 U5588 ( .A(n5205), .Y(n7774) );
  AND2X1 U5589 ( .A(n4138), .B(n5207), .Y(n5223) );
  INVX1 U5590 ( .A(n5223), .Y(n7775) );
  AND2X1 U5591 ( .A(n4162), .B(n5207), .Y(n5235) );
  INVX1 U5592 ( .A(n5235), .Y(n7776) );
  AND2X1 U5593 ( .A(n4186), .B(n5207), .Y(n5247) );
  INVX1 U5594 ( .A(n5247), .Y(n7777) );
  AND2X1 U5595 ( .A(n4136), .B(n5249), .Y(n5264) );
  INVX1 U5596 ( .A(n5264), .Y(n7778) );
  AND2X1 U5597 ( .A(n4160), .B(n5249), .Y(n5276) );
  INVX1 U5598 ( .A(n5276), .Y(n7779) );
  AND2X1 U5599 ( .A(n4184), .B(n5249), .Y(n5288) );
  INVX1 U5600 ( .A(n5288), .Y(n7780) );
  AND2X1 U5601 ( .A(n4134), .B(n5291), .Y(n5305) );
  INVX1 U5602 ( .A(n5305), .Y(n7781) );
  AND2X1 U5603 ( .A(n4158), .B(n5291), .Y(n5317) );
  INVX1 U5604 ( .A(n5317), .Y(n7782) );
  AND2X1 U5605 ( .A(n4182), .B(n5291), .Y(n5329) );
  INVX1 U5606 ( .A(n5329), .Y(n7783) );
  AND2X1 U5607 ( .A(n4132), .B(n5333), .Y(n5346) );
  INVX1 U5608 ( .A(n5346), .Y(n7784) );
  AND2X1 U5609 ( .A(n4156), .B(n5333), .Y(n5358) );
  INVX1 U5610 ( .A(n5358), .Y(n7785) );
  AND2X1 U5611 ( .A(n4180), .B(n5333), .Y(n5370) );
  INVX1 U5612 ( .A(n5370), .Y(n7786) );
  AND2X1 U5613 ( .A(n4130), .B(n5375), .Y(n5387) );
  INVX1 U5614 ( .A(n5387), .Y(n7787) );
  AND2X1 U5615 ( .A(n4154), .B(n5375), .Y(n5399) );
  INVX1 U5616 ( .A(n5399), .Y(n7788) );
  AND2X1 U5617 ( .A(n4178), .B(n5375), .Y(n5411) );
  INVX1 U5618 ( .A(n5411), .Y(n7789) );
  AND2X1 U5619 ( .A(n4128), .B(n5417), .Y(n5428) );
  INVX1 U5620 ( .A(n5428), .Y(n7790) );
  AND2X1 U5621 ( .A(n4152), .B(n5417), .Y(n5440) );
  INVX1 U5622 ( .A(n5440), .Y(n7791) );
  AND2X1 U5623 ( .A(n4176), .B(n5417), .Y(n5452) );
  INVX1 U5624 ( .A(n5452), .Y(n7792) );
  AND2X1 U5625 ( .A(n4150), .B(n5459), .Y(n5481) );
  INVX1 U5626 ( .A(n5481), .Y(n7793) );
  AND2X1 U5627 ( .A(n4174), .B(n5459), .Y(n5493) );
  INVX1 U5628 ( .A(n5493), .Y(n7794) );
  BUFX2 U5629 ( .A(n4101), .Y(n7795) );
  AND2X1 U5630 ( .A(n4114), .B(n4106), .Y(n4113) );
  INVX1 U5631 ( .A(n4113), .Y(n7796) );
  AND2X1 U5632 ( .A(n4124), .B(n4106), .Y(n4123) );
  INVX1 U5633 ( .A(n4123), .Y(n7797) );
  AND2X1 U5634 ( .A(n4116), .B(n4190), .Y(n4195) );
  INVX1 U5635 ( .A(n4195), .Y(n7798) );
  AND2X1 U5636 ( .A(n4126), .B(n4190), .Y(n4200) );
  INVX1 U5637 ( .A(n4200), .Y(n7799) );
  AND2X1 U5638 ( .A(n4110), .B(n4233), .Y(n4235) );
  INVX1 U5639 ( .A(n4235), .Y(n7800) );
  AND2X1 U5640 ( .A(n4120), .B(n4233), .Y(n4240) );
  INVX1 U5641 ( .A(n4240), .Y(n7801) );
  AND2X1 U5642 ( .A(n4112), .B(n4276), .Y(n4279) );
  INVX1 U5643 ( .A(n4279), .Y(n7802) );
  AND2X1 U5644 ( .A(n4122), .B(n4276), .Y(n4284) );
  INVX1 U5645 ( .A(n4284), .Y(n7803) );
  AND2X1 U5646 ( .A(n4138), .B(n4319), .Y(n4335) );
  INVX1 U5647 ( .A(n4335), .Y(n7804) );
  AND2X1 U5648 ( .A(n4162), .B(n4319), .Y(n4347) );
  INVX1 U5649 ( .A(n4347), .Y(n7805) );
  AND2X1 U5650 ( .A(n4186), .B(n4319), .Y(n4359) );
  INVX1 U5651 ( .A(n4359), .Y(n7806) );
  AND2X1 U5652 ( .A(n4140), .B(n4361), .Y(n4378) );
  INVX1 U5653 ( .A(n4378), .Y(n7807) );
  AND2X1 U5654 ( .A(n4164), .B(n4361), .Y(n4390) );
  INVX1 U5655 ( .A(n4390), .Y(n7808) );
  AND2X1 U5656 ( .A(n4188), .B(n4361), .Y(n4402) );
  INVX1 U5657 ( .A(n4402), .Y(n7809) );
  AND2X1 U5658 ( .A(n4134), .B(n4404), .Y(n4418) );
  INVX1 U5659 ( .A(n4418), .Y(n7810) );
  AND2X1 U5660 ( .A(n4158), .B(n4404), .Y(n4430) );
  INVX1 U5661 ( .A(n4430), .Y(n7811) );
  AND2X1 U5662 ( .A(n4182), .B(n4404), .Y(n4442) );
  INVX1 U5663 ( .A(n4442), .Y(n7812) );
  AND2X1 U5664 ( .A(n4136), .B(n4447), .Y(n4462) );
  INVX1 U5665 ( .A(n4462), .Y(n7813) );
  AND2X1 U5666 ( .A(n4160), .B(n4447), .Y(n4474) );
  INVX1 U5667 ( .A(n4474), .Y(n7814) );
  AND2X1 U5668 ( .A(n4184), .B(n4447), .Y(n4486) );
  INVX1 U5669 ( .A(n4486), .Y(n7815) );
  AND2X1 U5670 ( .A(n4130), .B(n4490), .Y(n4502) );
  INVX1 U5671 ( .A(n4502), .Y(n7816) );
  AND2X1 U5672 ( .A(n4154), .B(n4490), .Y(n4514) );
  INVX1 U5673 ( .A(n4514), .Y(n7817) );
  AND2X1 U5674 ( .A(n4178), .B(n4490), .Y(n4526) );
  INVX1 U5675 ( .A(n4526), .Y(n7818) );
  AND2X1 U5676 ( .A(n4132), .B(n4533), .Y(n4546) );
  INVX1 U5677 ( .A(n4546), .Y(n7819) );
  AND2X1 U5678 ( .A(n4156), .B(n4533), .Y(n4558) );
  INVX1 U5679 ( .A(n4558), .Y(n7820) );
  AND2X1 U5680 ( .A(n4180), .B(n4533), .Y(n4570) );
  INVX1 U5681 ( .A(n4570), .Y(n7821) );
  AND2X1 U5682 ( .A(n4150), .B(n4575), .Y(n4597) );
  INVX1 U5683 ( .A(n4597), .Y(n7822) );
  AND2X1 U5684 ( .A(n4174), .B(n4575), .Y(n4609) );
  INVX1 U5685 ( .A(n4609), .Y(n7823) );
  AND2X1 U5686 ( .A(n4128), .B(n4617), .Y(n4628) );
  INVX1 U5687 ( .A(n4628), .Y(n7824) );
  AND2X1 U5688 ( .A(n4152), .B(n4617), .Y(n4640) );
  INVX1 U5689 ( .A(n4640), .Y(n7825) );
  AND2X1 U5690 ( .A(n4176), .B(n4617), .Y(n4652) );
  INVX1 U5691 ( .A(n4652), .Y(n7826) );
  AND2X1 U5692 ( .A(n4114), .B(n4659), .Y(n4663) );
  INVX1 U5693 ( .A(n4663), .Y(n7827) );
  AND2X1 U5694 ( .A(n4124), .B(n4659), .Y(n4668) );
  INVX1 U5695 ( .A(n4668), .Y(n7828) );
  AND2X1 U5696 ( .A(n4116), .B(n4701), .Y(n4706) );
  INVX1 U5697 ( .A(n4706), .Y(n7829) );
  AND2X1 U5698 ( .A(n4126), .B(n4701), .Y(n4711) );
  INVX1 U5699 ( .A(n4711), .Y(n7830) );
  AND2X1 U5700 ( .A(n4110), .B(n4743), .Y(n4745) );
  INVX1 U5701 ( .A(n4745), .Y(n7831) );
  AND2X1 U5702 ( .A(n4120), .B(n4743), .Y(n4750) );
  INVX1 U5703 ( .A(n4750), .Y(n7832) );
  AND2X1 U5704 ( .A(n4112), .B(n4785), .Y(n4788) );
  INVX1 U5705 ( .A(n4788), .Y(n7833) );
  AND2X1 U5706 ( .A(n4122), .B(n4785), .Y(n4793) );
  INVX1 U5707 ( .A(n4793), .Y(n7834) );
  AND2X1 U5708 ( .A(n4138), .B(n4827), .Y(n4843) );
  INVX1 U5709 ( .A(n4843), .Y(n7835) );
  AND2X1 U5710 ( .A(n4162), .B(n4827), .Y(n4855) );
  INVX1 U5711 ( .A(n4855), .Y(n7836) );
  AND2X1 U5712 ( .A(n4186), .B(n4827), .Y(n4867) );
  INVX1 U5713 ( .A(n4867), .Y(n7837) );
  AND2X1 U5714 ( .A(n4140), .B(n4870), .Y(n4887) );
  INVX1 U5715 ( .A(n4887), .Y(n7838) );
  AND2X1 U5716 ( .A(n4164), .B(n4870), .Y(n4899) );
  INVX1 U5717 ( .A(n4899), .Y(n7839) );
  AND2X1 U5718 ( .A(n4188), .B(n4870), .Y(n4911) );
  INVX1 U5719 ( .A(n4911), .Y(n7840) );
  AND2X1 U5720 ( .A(n4134), .B(n4912), .Y(n4926) );
  INVX1 U5721 ( .A(n4926), .Y(n7841) );
  AND2X1 U5722 ( .A(n4158), .B(n4912), .Y(n4938) );
  INVX1 U5723 ( .A(n4938), .Y(n7842) );
  AND2X1 U5724 ( .A(n4182), .B(n4912), .Y(n4950) );
  INVX1 U5725 ( .A(n4950), .Y(n7843) );
  AND2X1 U5726 ( .A(n4136), .B(n4954), .Y(n4969) );
  INVX1 U5727 ( .A(n4969), .Y(n7844) );
  AND2X1 U5728 ( .A(n4160), .B(n4954), .Y(n4981) );
  INVX1 U5729 ( .A(n4981), .Y(n7845) );
  AND2X1 U5730 ( .A(n4184), .B(n4954), .Y(n4993) );
  INVX1 U5731 ( .A(n4993), .Y(n7846) );
  AND2X1 U5732 ( .A(n4130), .B(n4996), .Y(n5008) );
  INVX1 U5733 ( .A(n5008), .Y(n7847) );
  AND2X1 U5734 ( .A(n4154), .B(n4996), .Y(n5020) );
  INVX1 U5735 ( .A(n5020), .Y(n7848) );
  AND2X1 U5736 ( .A(n4178), .B(n4996), .Y(n5032) );
  INVX1 U5737 ( .A(n5032), .Y(n7849) );
  AND2X1 U5738 ( .A(n4132), .B(n5038), .Y(n5051) );
  INVX1 U5739 ( .A(n5051), .Y(n7850) );
  AND2X1 U5740 ( .A(n4156), .B(n5038), .Y(n5063) );
  INVX1 U5741 ( .A(n5063), .Y(n7851) );
  AND2X1 U5742 ( .A(n4180), .B(n5038), .Y(n5075) );
  INVX1 U5743 ( .A(n5075), .Y(n7852) );
  AND2X1 U5744 ( .A(n4150), .B(n5080), .Y(n5102) );
  INVX1 U5745 ( .A(n5102), .Y(n7853) );
  AND2X1 U5746 ( .A(n4174), .B(n5080), .Y(n5114) );
  INVX1 U5747 ( .A(n5114), .Y(n7854) );
  AND2X1 U5748 ( .A(n4128), .B(n5122), .Y(n5133) );
  INVX1 U5749 ( .A(n5133), .Y(n7855) );
  AND2X1 U5750 ( .A(n4152), .B(n5122), .Y(n5145) );
  INVX1 U5751 ( .A(n5145), .Y(n7856) );
  AND2X1 U5752 ( .A(n4176), .B(n5122), .Y(n5157) );
  INVX1 U5753 ( .A(n5157), .Y(n7857) );
  AND2X1 U5754 ( .A(n4138), .B(n5164), .Y(n5180) );
  INVX1 U5755 ( .A(n5180), .Y(n7858) );
  AND2X1 U5756 ( .A(n4162), .B(n5164), .Y(n5192) );
  INVX1 U5757 ( .A(n5192), .Y(n7859) );
  AND2X1 U5758 ( .A(n4186), .B(n5164), .Y(n5204) );
  INVX1 U5759 ( .A(n5204), .Y(n7860) );
  AND2X1 U5760 ( .A(n4140), .B(n5207), .Y(n5224) );
  INVX1 U5761 ( .A(n5224), .Y(n7861) );
  AND2X1 U5762 ( .A(n4164), .B(n5207), .Y(n5236) );
  INVX1 U5763 ( .A(n5236), .Y(n7862) );
  AND2X1 U5764 ( .A(n4188), .B(n5207), .Y(n5248) );
  INVX1 U5765 ( .A(n5248), .Y(n7863) );
  AND2X1 U5766 ( .A(n4134), .B(n5249), .Y(n5263) );
  INVX1 U5767 ( .A(n5263), .Y(n7864) );
  AND2X1 U5768 ( .A(n4158), .B(n5249), .Y(n5275) );
  INVX1 U5769 ( .A(n5275), .Y(n7865) );
  AND2X1 U5770 ( .A(n4182), .B(n5249), .Y(n5287) );
  INVX1 U5771 ( .A(n5287), .Y(n7866) );
  AND2X1 U5772 ( .A(n4136), .B(n5291), .Y(n5306) );
  INVX1 U5773 ( .A(n5306), .Y(n7867) );
  AND2X1 U5774 ( .A(n4160), .B(n5291), .Y(n5318) );
  INVX1 U5775 ( .A(n5318), .Y(n7868) );
  AND2X1 U5776 ( .A(n4184), .B(n5291), .Y(n5330) );
  INVX1 U5777 ( .A(n5330), .Y(n7869) );
  AND2X1 U5778 ( .A(n4130), .B(n5333), .Y(n5345) );
  INVX1 U5779 ( .A(n5345), .Y(n7870) );
  AND2X1 U5780 ( .A(n4154), .B(n5333), .Y(n5357) );
  INVX1 U5781 ( .A(n5357), .Y(n7871) );
  AND2X1 U5782 ( .A(n4178), .B(n5333), .Y(n5369) );
  INVX1 U5783 ( .A(n5369), .Y(n7872) );
  AND2X1 U5784 ( .A(n4132), .B(n5375), .Y(n5388) );
  INVX1 U5785 ( .A(n5388), .Y(n7873) );
  AND2X1 U5786 ( .A(n4156), .B(n5375), .Y(n5400) );
  INVX1 U5787 ( .A(n5400), .Y(n7874) );
  AND2X1 U5788 ( .A(n4180), .B(n5375), .Y(n5412) );
  INVX1 U5789 ( .A(n5412), .Y(n7875) );
  AND2X1 U5790 ( .A(n4150), .B(n5417), .Y(n5439) );
  INVX1 U5791 ( .A(n5439), .Y(n7876) );
  AND2X1 U5792 ( .A(n4174), .B(n5417), .Y(n5451) );
  INVX1 U5793 ( .A(n5451), .Y(n7877) );
  AND2X1 U5794 ( .A(n4128), .B(n5459), .Y(n5470) );
  INVX1 U5795 ( .A(n5470), .Y(n7878) );
  AND2X1 U5796 ( .A(n4152), .B(n5459), .Y(n5482) );
  INVX1 U5797 ( .A(n5482), .Y(n7879) );
  AND2X1 U5798 ( .A(n4176), .B(n5459), .Y(n5494) );
  INVX1 U5799 ( .A(n5494), .Y(n7880) );
  BUFX2 U5800 ( .A(n5503), .Y(n7881) );
  BUFX2 U5801 ( .A(n5506), .Y(n7882) );
  AND2X1 U5802 ( .A(n4112), .B(n4106), .Y(n4111) );
  INVX1 U5803 ( .A(n4111), .Y(n7883) );
  AND2X1 U5804 ( .A(n4122), .B(n4106), .Y(n4121) );
  INVX1 U5805 ( .A(n4121), .Y(n7884) );
  AND2X1 U5806 ( .A(n4110), .B(n4190), .Y(n4192) );
  INVX1 U5807 ( .A(n4192), .Y(n7885) );
  AND2X1 U5808 ( .A(n4120), .B(n4190), .Y(n4197) );
  INVX1 U5809 ( .A(n4197), .Y(n7886) );
  AND2X1 U5810 ( .A(n4116), .B(n4233), .Y(n4238) );
  INVX1 U5811 ( .A(n4238), .Y(n7887) );
  AND2X1 U5812 ( .A(n4126), .B(n4233), .Y(n4243) );
  INVX1 U5813 ( .A(n4243), .Y(n7888) );
  AND2X1 U5814 ( .A(n4114), .B(n4276), .Y(n4280) );
  INVX1 U5815 ( .A(n4280), .Y(n7889) );
  AND2X1 U5816 ( .A(n4124), .B(n4276), .Y(n4285) );
  INVX1 U5817 ( .A(n4285), .Y(n7890) );
  AND2X1 U5818 ( .A(n4136), .B(n4319), .Y(n4334) );
  INVX1 U5819 ( .A(n4334), .Y(n7891) );
  AND2X1 U5820 ( .A(n4160), .B(n4319), .Y(n4346) );
  INVX1 U5821 ( .A(n4346), .Y(n7892) );
  AND2X1 U5822 ( .A(n4184), .B(n4319), .Y(n4358) );
  INVX1 U5823 ( .A(n4358), .Y(n7893) );
  AND2X1 U5824 ( .A(n4134), .B(n4361), .Y(n4375) );
  INVX1 U5825 ( .A(n4375), .Y(n7894) );
  AND2X1 U5826 ( .A(n4158), .B(n4361), .Y(n4387) );
  INVX1 U5827 ( .A(n4387), .Y(n7895) );
  AND2X1 U5828 ( .A(n4182), .B(n4361), .Y(n4399) );
  INVX1 U5829 ( .A(n4399), .Y(n7896) );
  AND2X1 U5830 ( .A(n4140), .B(n4404), .Y(n4421) );
  INVX1 U5831 ( .A(n4421), .Y(n7897) );
  AND2X1 U5832 ( .A(n4164), .B(n4404), .Y(n4433) );
  INVX1 U5833 ( .A(n4433), .Y(n7898) );
  AND2X1 U5834 ( .A(n4188), .B(n4404), .Y(n4445) );
  INVX1 U5835 ( .A(n4445), .Y(n7899) );
  AND2X1 U5836 ( .A(n4138), .B(n4447), .Y(n4463) );
  INVX1 U5837 ( .A(n4463), .Y(n7900) );
  AND2X1 U5838 ( .A(n4162), .B(n4447), .Y(n4475) );
  INVX1 U5839 ( .A(n4475), .Y(n7901) );
  AND2X1 U5840 ( .A(n4186), .B(n4447), .Y(n4487) );
  INVX1 U5841 ( .A(n4487), .Y(n7902) );
  AND2X1 U5842 ( .A(n4128), .B(n4490), .Y(n4501) );
  INVX1 U5843 ( .A(n4501), .Y(n7903) );
  AND2X1 U5844 ( .A(n4152), .B(n4490), .Y(n4513) );
  INVX1 U5845 ( .A(n4513), .Y(n7904) );
  AND2X1 U5846 ( .A(n4176), .B(n4490), .Y(n4525) );
  INVX1 U5847 ( .A(n4525), .Y(n7905) );
  AND2X1 U5848 ( .A(n4150), .B(n4533), .Y(n4555) );
  INVX1 U5849 ( .A(n4555), .Y(n7906) );
  AND2X1 U5850 ( .A(n4174), .B(n4533), .Y(n4567) );
  INVX1 U5851 ( .A(n4567), .Y(n7907) );
  AND2X1 U5852 ( .A(n4132), .B(n4575), .Y(n4588) );
  INVX1 U5853 ( .A(n4588), .Y(n7908) );
  AND2X1 U5854 ( .A(n4156), .B(n4575), .Y(n4600) );
  INVX1 U5855 ( .A(n4600), .Y(n7909) );
  AND2X1 U5856 ( .A(n4180), .B(n4575), .Y(n4612) );
  INVX1 U5857 ( .A(n4612), .Y(n7910) );
  AND2X1 U5858 ( .A(n4130), .B(n4617), .Y(n4629) );
  INVX1 U5859 ( .A(n4629), .Y(n7911) );
  AND2X1 U5860 ( .A(n4154), .B(n4617), .Y(n4641) );
  INVX1 U5861 ( .A(n4641), .Y(n7912) );
  AND2X1 U5862 ( .A(n4178), .B(n4617), .Y(n4653) );
  INVX1 U5863 ( .A(n4653), .Y(n7913) );
  AND2X1 U5864 ( .A(n4112), .B(n4659), .Y(n4662) );
  INVX1 U5865 ( .A(n4662), .Y(n7914) );
  AND2X1 U5866 ( .A(n4122), .B(n4659), .Y(n4667) );
  INVX1 U5867 ( .A(n4667), .Y(n7915) );
  AND2X1 U5868 ( .A(n4110), .B(n4701), .Y(n4703) );
  INVX1 U5869 ( .A(n4703), .Y(n7916) );
  AND2X1 U5870 ( .A(n4120), .B(n4701), .Y(n4708) );
  INVX1 U5871 ( .A(n4708), .Y(n7917) );
  AND2X1 U5872 ( .A(n4116), .B(n4743), .Y(n4748) );
  INVX1 U5873 ( .A(n4748), .Y(n7918) );
  AND2X1 U5874 ( .A(n4126), .B(n4743), .Y(n4753) );
  INVX1 U5875 ( .A(n4753), .Y(n7919) );
  AND2X1 U5876 ( .A(n4114), .B(n4785), .Y(n4789) );
  INVX1 U5877 ( .A(n4789), .Y(n7920) );
  AND2X1 U5878 ( .A(n4124), .B(n4785), .Y(n4794) );
  INVX1 U5879 ( .A(n4794), .Y(n7921) );
  AND2X1 U5880 ( .A(n4136), .B(n4827), .Y(n4842) );
  INVX1 U5881 ( .A(n4842), .Y(n7922) );
  AND2X1 U5882 ( .A(n4160), .B(n4827), .Y(n4854) );
  INVX1 U5883 ( .A(n4854), .Y(n7923) );
  AND2X1 U5884 ( .A(n4184), .B(n4827), .Y(n4866) );
  INVX1 U5885 ( .A(n4866), .Y(n7924) );
  AND2X1 U5886 ( .A(n4134), .B(n4870), .Y(n4884) );
  INVX1 U5887 ( .A(n4884), .Y(n7925) );
  AND2X1 U5888 ( .A(n4158), .B(n4870), .Y(n4896) );
  INVX1 U5889 ( .A(n4896), .Y(n7926) );
  AND2X1 U5890 ( .A(n4182), .B(n4870), .Y(n4908) );
  INVX1 U5891 ( .A(n4908), .Y(n7927) );
  AND2X1 U5892 ( .A(n4140), .B(n4912), .Y(n4929) );
  INVX1 U5893 ( .A(n4929), .Y(n7928) );
  AND2X1 U5894 ( .A(n4164), .B(n4912), .Y(n4941) );
  INVX1 U5895 ( .A(n4941), .Y(n7929) );
  AND2X1 U5896 ( .A(n4188), .B(n4912), .Y(n4953) );
  INVX1 U5897 ( .A(n4953), .Y(n7930) );
  AND2X1 U5898 ( .A(n4138), .B(n4954), .Y(n4970) );
  INVX1 U5899 ( .A(n4970), .Y(n7931) );
  AND2X1 U5900 ( .A(n4162), .B(n4954), .Y(n4982) );
  INVX1 U5901 ( .A(n4982), .Y(n7932) );
  AND2X1 U5902 ( .A(n4186), .B(n4954), .Y(n4994) );
  INVX1 U5903 ( .A(n4994), .Y(n7933) );
  AND2X1 U5904 ( .A(n4128), .B(n4996), .Y(n5007) );
  INVX1 U5905 ( .A(n5007), .Y(n7934) );
  AND2X1 U5906 ( .A(n4152), .B(n4996), .Y(n5019) );
  INVX1 U5907 ( .A(n5019), .Y(n7935) );
  AND2X1 U5908 ( .A(n4176), .B(n4996), .Y(n5031) );
  INVX1 U5909 ( .A(n5031), .Y(n7936) );
  AND2X1 U5910 ( .A(n4150), .B(n5038), .Y(n5060) );
  INVX1 U5911 ( .A(n5060), .Y(n7937) );
  AND2X1 U5912 ( .A(n4174), .B(n5038), .Y(n5072) );
  INVX1 U5913 ( .A(n5072), .Y(n7938) );
  AND2X1 U5914 ( .A(n4132), .B(n5080), .Y(n5093) );
  INVX1 U5915 ( .A(n5093), .Y(n7939) );
  AND2X1 U5916 ( .A(n4156), .B(n5080), .Y(n5105) );
  INVX1 U5917 ( .A(n5105), .Y(n7940) );
  AND2X1 U5918 ( .A(n4180), .B(n5080), .Y(n5117) );
  INVX1 U5919 ( .A(n5117), .Y(n7941) );
  AND2X1 U5920 ( .A(n4130), .B(n5122), .Y(n5134) );
  INVX1 U5921 ( .A(n5134), .Y(n7942) );
  AND2X1 U5922 ( .A(n4154), .B(n5122), .Y(n5146) );
  INVX1 U5923 ( .A(n5146), .Y(n7943) );
  AND2X1 U5924 ( .A(n4178), .B(n5122), .Y(n5158) );
  INVX1 U5925 ( .A(n5158), .Y(n7944) );
  AND2X1 U5926 ( .A(n4136), .B(n5164), .Y(n5179) );
  INVX1 U5927 ( .A(n5179), .Y(n7945) );
  AND2X1 U5928 ( .A(n4160), .B(n5164), .Y(n5191) );
  INVX1 U5929 ( .A(n5191), .Y(n7946) );
  AND2X1 U5930 ( .A(n4184), .B(n5164), .Y(n5203) );
  INVX1 U5931 ( .A(n5203), .Y(n7947) );
  AND2X1 U5932 ( .A(n4134), .B(n5207), .Y(n5221) );
  INVX1 U5933 ( .A(n5221), .Y(n7948) );
  AND2X1 U5934 ( .A(n4158), .B(n5207), .Y(n5233) );
  INVX1 U5935 ( .A(n5233), .Y(n7949) );
  AND2X1 U5936 ( .A(n4182), .B(n5207), .Y(n5245) );
  INVX1 U5937 ( .A(n5245), .Y(n7950) );
  AND2X1 U5938 ( .A(n4140), .B(n5249), .Y(n5266) );
  INVX1 U5939 ( .A(n5266), .Y(n7951) );
  AND2X1 U5940 ( .A(n4164), .B(n5249), .Y(n5278) );
  INVX1 U5941 ( .A(n5278), .Y(n7952) );
  AND2X1 U5942 ( .A(n4188), .B(n5249), .Y(n5290) );
  INVX1 U5943 ( .A(n5290), .Y(n7953) );
  AND2X1 U5944 ( .A(n4138), .B(n5291), .Y(n5307) );
  INVX1 U5945 ( .A(n5307), .Y(n7954) );
  AND2X1 U5946 ( .A(n4162), .B(n5291), .Y(n5319) );
  INVX1 U5947 ( .A(n5319), .Y(n7955) );
  AND2X1 U5948 ( .A(n4186), .B(n5291), .Y(n5331) );
  INVX1 U5949 ( .A(n5331), .Y(n7956) );
  AND2X1 U5950 ( .A(n4128), .B(n5333), .Y(n5344) );
  INVX1 U5951 ( .A(n5344), .Y(n7957) );
  AND2X1 U5952 ( .A(n4152), .B(n5333), .Y(n5356) );
  INVX1 U5953 ( .A(n5356), .Y(n7958) );
  AND2X1 U5954 ( .A(n4176), .B(n5333), .Y(n5368) );
  INVX1 U5955 ( .A(n5368), .Y(n7959) );
  AND2X1 U5956 ( .A(n4150), .B(n5375), .Y(n5397) );
  INVX1 U5957 ( .A(n5397), .Y(n7960) );
  AND2X1 U5958 ( .A(n4174), .B(n5375), .Y(n5409) );
  INVX1 U5959 ( .A(n5409), .Y(n7961) );
  AND2X1 U5960 ( .A(n4132), .B(n5417), .Y(n5430) );
  INVX1 U5961 ( .A(n5430), .Y(n7962) );
  AND2X1 U5962 ( .A(n4156), .B(n5417), .Y(n5442) );
  INVX1 U5963 ( .A(n5442), .Y(n7963) );
  AND2X1 U5964 ( .A(n4180), .B(n5417), .Y(n5454) );
  INVX1 U5965 ( .A(n5454), .Y(n7964) );
  AND2X1 U5966 ( .A(n4130), .B(n5459), .Y(n5471) );
  INVX1 U5967 ( .A(n5471), .Y(n7965) );
  AND2X1 U5968 ( .A(n4154), .B(n5459), .Y(n5483) );
  INVX1 U5969 ( .A(n5483), .Y(n7966) );
  AND2X1 U5970 ( .A(n4178), .B(n5459), .Y(n5495) );
  INVX1 U5971 ( .A(n5495), .Y(n7967) );
  BUFX2 U5972 ( .A(n4104), .Y(n7968) );
  BUFX2 U5973 ( .A(n4275), .Y(n7969) );
  BUFX2 U5974 ( .A(n4403), .Y(n7970) );
  AND2X1 U5975 ( .A(n4062), .B(n8511), .Y(n4083) );
  INVX1 U5976 ( .A(n4083), .Y(n7971) );
  AND2X1 U5977 ( .A(n4110), .B(n4106), .Y(n4109) );
  INVX1 U5978 ( .A(n4109), .Y(n7972) );
  AND2X1 U5979 ( .A(n4120), .B(n4106), .Y(n4119) );
  INVX1 U5980 ( .A(n4119), .Y(n7973) );
  AND2X1 U5981 ( .A(n4112), .B(n4190), .Y(n4193) );
  INVX1 U5982 ( .A(n4193), .Y(n7974) );
  AND2X1 U5983 ( .A(n4122), .B(n4190), .Y(n4198) );
  INVX1 U5984 ( .A(n4198), .Y(n7975) );
  AND2X1 U5985 ( .A(n4114), .B(n4233), .Y(n4237) );
  INVX1 U5986 ( .A(n4237), .Y(n7976) );
  AND2X1 U5987 ( .A(n4124), .B(n4233), .Y(n4242) );
  INVX1 U5988 ( .A(n4242), .Y(n7977) );
  AND2X1 U5989 ( .A(n4116), .B(n4276), .Y(n4281) );
  INVX1 U5990 ( .A(n4281), .Y(n7978) );
  AND2X1 U5991 ( .A(n4126), .B(n4276), .Y(n4286) );
  INVX1 U5992 ( .A(n4286), .Y(n7979) );
  AND2X1 U5993 ( .A(n4134), .B(n4319), .Y(n4333) );
  INVX1 U5994 ( .A(n4333), .Y(n7980) );
  AND2X1 U5995 ( .A(n4158), .B(n4319), .Y(n4345) );
  INVX1 U5996 ( .A(n4345), .Y(n7981) );
  AND2X1 U5997 ( .A(n4182), .B(n4319), .Y(n4357) );
  INVX1 U5998 ( .A(n4357), .Y(n7982) );
  AND2X1 U5999 ( .A(n4136), .B(n4361), .Y(n4376) );
  INVX1 U6000 ( .A(n4376), .Y(n7983) );
  AND2X1 U6001 ( .A(n4160), .B(n4361), .Y(n4388) );
  INVX1 U6002 ( .A(n4388), .Y(n7984) );
  AND2X1 U6003 ( .A(n4184), .B(n4361), .Y(n4400) );
  INVX1 U6004 ( .A(n4400), .Y(n7985) );
  AND2X1 U6005 ( .A(n4138), .B(n4404), .Y(n4420) );
  INVX1 U6006 ( .A(n4420), .Y(n7986) );
  AND2X1 U6007 ( .A(n4162), .B(n4404), .Y(n4432) );
  INVX1 U6008 ( .A(n4432), .Y(n7987) );
  AND2X1 U6009 ( .A(n4186), .B(n4404), .Y(n4444) );
  INVX1 U6010 ( .A(n4444), .Y(n7988) );
  AND2X1 U6011 ( .A(n4140), .B(n4447), .Y(n4464) );
  INVX1 U6012 ( .A(n4464), .Y(n7989) );
  AND2X1 U6013 ( .A(n4164), .B(n4447), .Y(n4476) );
  INVX1 U6014 ( .A(n4476), .Y(n7990) );
  AND2X1 U6015 ( .A(n4188), .B(n4447), .Y(n4488) );
  INVX1 U6016 ( .A(n4488), .Y(n7991) );
  AND2X1 U6017 ( .A(n4150), .B(n4490), .Y(n4512) );
  INVX1 U6018 ( .A(n4512), .Y(n7992) );
  AND2X1 U6019 ( .A(n4174), .B(n4490), .Y(n4524) );
  INVX1 U6020 ( .A(n4524), .Y(n7993) );
  AND2X1 U6021 ( .A(n4128), .B(n4533), .Y(n4544) );
  INVX1 U6022 ( .A(n4544), .Y(n7994) );
  AND2X1 U6023 ( .A(n4152), .B(n4533), .Y(n4556) );
  INVX1 U6024 ( .A(n4556), .Y(n7995) );
  AND2X1 U6025 ( .A(n4176), .B(n4533), .Y(n4568) );
  INVX1 U6026 ( .A(n4568), .Y(n7996) );
  AND2X1 U6027 ( .A(n4130), .B(n4575), .Y(n4587) );
  INVX1 U6028 ( .A(n4587), .Y(n7997) );
  AND2X1 U6029 ( .A(n4154), .B(n4575), .Y(n4599) );
  INVX1 U6030 ( .A(n4599), .Y(n7998) );
  AND2X1 U6031 ( .A(n4178), .B(n4575), .Y(n4611) );
  INVX1 U6032 ( .A(n4611), .Y(n7999) );
  AND2X1 U6033 ( .A(n4132), .B(n4617), .Y(n4630) );
  INVX1 U6034 ( .A(n4630), .Y(n8000) );
  AND2X1 U6035 ( .A(n4156), .B(n4617), .Y(n4642) );
  INVX1 U6036 ( .A(n4642), .Y(n8001) );
  AND2X1 U6037 ( .A(n4180), .B(n4617), .Y(n4654) );
  INVX1 U6038 ( .A(n4654), .Y(n8002) );
  AND2X1 U6039 ( .A(n4110), .B(n4659), .Y(n4661) );
  INVX1 U6040 ( .A(n4661), .Y(n8003) );
  AND2X1 U6041 ( .A(n4120), .B(n4659), .Y(n4666) );
  INVX1 U6042 ( .A(n4666), .Y(n8004) );
  AND2X1 U6043 ( .A(n4112), .B(n4701), .Y(n4704) );
  INVX1 U6044 ( .A(n4704), .Y(n8005) );
  AND2X1 U6045 ( .A(n4122), .B(n4701), .Y(n4709) );
  INVX1 U6046 ( .A(n4709), .Y(n8006) );
  AND2X1 U6047 ( .A(n4114), .B(n4743), .Y(n4747) );
  INVX1 U6048 ( .A(n4747), .Y(n8007) );
  AND2X1 U6049 ( .A(n4124), .B(n4743), .Y(n4752) );
  INVX1 U6050 ( .A(n4752), .Y(n8008) );
  AND2X1 U6051 ( .A(n4116), .B(n4785), .Y(n4790) );
  INVX1 U6052 ( .A(n4790), .Y(n8009) );
  AND2X1 U6053 ( .A(n4126), .B(n4785), .Y(n4795) );
  INVX1 U6054 ( .A(n4795), .Y(n8010) );
  AND2X1 U6055 ( .A(n4134), .B(n4827), .Y(n4841) );
  INVX1 U6056 ( .A(n4841), .Y(n8011) );
  AND2X1 U6057 ( .A(n4158), .B(n4827), .Y(n4853) );
  INVX1 U6058 ( .A(n4853), .Y(n8012) );
  AND2X1 U6059 ( .A(n4182), .B(n4827), .Y(n4865) );
  INVX1 U6060 ( .A(n4865), .Y(n8013) );
  AND2X1 U6061 ( .A(n4136), .B(n4870), .Y(n4885) );
  INVX1 U6062 ( .A(n4885), .Y(n8014) );
  AND2X1 U6063 ( .A(n4160), .B(n4870), .Y(n4897) );
  INVX1 U6064 ( .A(n4897), .Y(n8015) );
  AND2X1 U6065 ( .A(n4184), .B(n4870), .Y(n4909) );
  INVX1 U6066 ( .A(n4909), .Y(n8016) );
  AND2X1 U6067 ( .A(n4138), .B(n4912), .Y(n4928) );
  INVX1 U6068 ( .A(n4928), .Y(n8017) );
  AND2X1 U6069 ( .A(n4162), .B(n4912), .Y(n4940) );
  INVX1 U6070 ( .A(n4940), .Y(n8018) );
  AND2X1 U6071 ( .A(n4186), .B(n4912), .Y(n4952) );
  INVX1 U6072 ( .A(n4952), .Y(n8019) );
  AND2X1 U6073 ( .A(n4140), .B(n4954), .Y(n4971) );
  INVX1 U6074 ( .A(n4971), .Y(n8020) );
  AND2X1 U6075 ( .A(n4164), .B(n4954), .Y(n4983) );
  INVX1 U6076 ( .A(n4983), .Y(n8021) );
  AND2X1 U6077 ( .A(n4188), .B(n4954), .Y(n4995) );
  INVX1 U6078 ( .A(n4995), .Y(n8022) );
  AND2X1 U6079 ( .A(n4150), .B(n4996), .Y(n5018) );
  INVX1 U6080 ( .A(n5018), .Y(n8023) );
  AND2X1 U6081 ( .A(n4174), .B(n4996), .Y(n5030) );
  INVX1 U6082 ( .A(n5030), .Y(n8024) );
  AND2X1 U6083 ( .A(n4128), .B(n5038), .Y(n5049) );
  INVX1 U6084 ( .A(n5049), .Y(n8025) );
  AND2X1 U6085 ( .A(n4152), .B(n5038), .Y(n5061) );
  INVX1 U6086 ( .A(n5061), .Y(n8026) );
  AND2X1 U6087 ( .A(n4176), .B(n5038), .Y(n5073) );
  INVX1 U6088 ( .A(n5073), .Y(n8027) );
  AND2X1 U6089 ( .A(n4130), .B(n5080), .Y(n5092) );
  INVX1 U6090 ( .A(n5092), .Y(n8028) );
  AND2X1 U6091 ( .A(n4154), .B(n5080), .Y(n5104) );
  INVX1 U6092 ( .A(n5104), .Y(n8029) );
  AND2X1 U6093 ( .A(n4178), .B(n5080), .Y(n5116) );
  INVX1 U6094 ( .A(n5116), .Y(n8030) );
  AND2X1 U6095 ( .A(n4132), .B(n5122), .Y(n5135) );
  INVX1 U6096 ( .A(n5135), .Y(n8031) );
  AND2X1 U6097 ( .A(n4156), .B(n5122), .Y(n5147) );
  INVX1 U6098 ( .A(n5147), .Y(n8032) );
  AND2X1 U6099 ( .A(n4180), .B(n5122), .Y(n5159) );
  INVX1 U6100 ( .A(n5159), .Y(n8033) );
  AND2X1 U6101 ( .A(n4134), .B(n5164), .Y(n5178) );
  INVX1 U6102 ( .A(n5178), .Y(n8034) );
  AND2X1 U6103 ( .A(n4158), .B(n5164), .Y(n5190) );
  INVX1 U6104 ( .A(n5190), .Y(n8035) );
  AND2X1 U6105 ( .A(n4182), .B(n5164), .Y(n5202) );
  INVX1 U6106 ( .A(n5202), .Y(n8036) );
  AND2X1 U6107 ( .A(n4136), .B(n5207), .Y(n5222) );
  INVX1 U6108 ( .A(n5222), .Y(n8037) );
  AND2X1 U6109 ( .A(n4160), .B(n5207), .Y(n5234) );
  INVX1 U6110 ( .A(n5234), .Y(n8038) );
  AND2X1 U6111 ( .A(n4184), .B(n5207), .Y(n5246) );
  INVX1 U6112 ( .A(n5246), .Y(n8039) );
  AND2X1 U6113 ( .A(n4138), .B(n5249), .Y(n5265) );
  INVX1 U6114 ( .A(n5265), .Y(n8040) );
  AND2X1 U6115 ( .A(n4162), .B(n5249), .Y(n5277) );
  INVX1 U6116 ( .A(n5277), .Y(n8041) );
  AND2X1 U6117 ( .A(n4186), .B(n5249), .Y(n5289) );
  INVX1 U6118 ( .A(n5289), .Y(n8042) );
  AND2X1 U6119 ( .A(n4140), .B(n5291), .Y(n5308) );
  INVX1 U6120 ( .A(n5308), .Y(n8043) );
  AND2X1 U6121 ( .A(n4164), .B(n5291), .Y(n5320) );
  INVX1 U6122 ( .A(n5320), .Y(n8044) );
  AND2X1 U6123 ( .A(n4188), .B(n5291), .Y(n5332) );
  INVX1 U6124 ( .A(n5332), .Y(n8045) );
  AND2X1 U6125 ( .A(n4150), .B(n5333), .Y(n5355) );
  INVX1 U6126 ( .A(n5355), .Y(n8046) );
  AND2X1 U6127 ( .A(n4174), .B(n5333), .Y(n5367) );
  INVX1 U6128 ( .A(n5367), .Y(n8047) );
  AND2X1 U6129 ( .A(n4128), .B(n5375), .Y(n5386) );
  INVX1 U6130 ( .A(n5386), .Y(n8048) );
  AND2X1 U6131 ( .A(n4152), .B(n5375), .Y(n5398) );
  INVX1 U6132 ( .A(n5398), .Y(n8049) );
  AND2X1 U6133 ( .A(n4176), .B(n5375), .Y(n5410) );
  INVX1 U6134 ( .A(n5410), .Y(n8050) );
  AND2X1 U6135 ( .A(n4130), .B(n5417), .Y(n5429) );
  INVX1 U6136 ( .A(n5429), .Y(n8051) );
  AND2X1 U6137 ( .A(n4154), .B(n5417), .Y(n5441) );
  INVX1 U6138 ( .A(n5441), .Y(n8052) );
  AND2X1 U6139 ( .A(n4178), .B(n5417), .Y(n5453) );
  INVX1 U6140 ( .A(n5453), .Y(n8053) );
  AND2X1 U6141 ( .A(n4132), .B(n5459), .Y(n5472) );
  INVX1 U6142 ( .A(n5472), .Y(n8054) );
  AND2X1 U6143 ( .A(n4156), .B(n5459), .Y(n5484) );
  INVX1 U6144 ( .A(n5484), .Y(n8055) );
  AND2X1 U6145 ( .A(n4180), .B(n5459), .Y(n5496) );
  INVX1 U6146 ( .A(n5496), .Y(n8056) );
  BUFX2 U6147 ( .A(n4096), .Y(n8057) );
  BUFX2 U6148 ( .A(n4095), .Y(n8058) );
  OR2X1 U6149 ( .A(n8518), .B(wr_ptr[4]), .Y(n4097) );
  INVX1 U6150 ( .A(n4097), .Y(n8059) );
  BUFX2 U6151 ( .A(n4232), .Y(n8060) );
  BUFX2 U6152 ( .A(n4446), .Y(n8061) );
  AND2X1 U6153 ( .A(n4148), .B(n4106), .Y(n4147) );
  INVX1 U6154 ( .A(n4147), .Y(n8062) );
  AND2X1 U6155 ( .A(n4172), .B(n4106), .Y(n4171) );
  INVX1 U6156 ( .A(n4171), .Y(n8063) );
  AND2X1 U6157 ( .A(n4108), .B(n4190), .Y(n4191) );
  INVX1 U6158 ( .A(n4191), .Y(n8064) );
  AND2X1 U6159 ( .A(n4146), .B(n4190), .Y(n4210) );
  INVX1 U6160 ( .A(n4210), .Y(n8065) );
  AND2X1 U6161 ( .A(n4170), .B(n4190), .Y(n4222) );
  INVX1 U6162 ( .A(n4222), .Y(n8066) );
  AND2X1 U6163 ( .A(n4144), .B(n4233), .Y(n4252) );
  INVX1 U6164 ( .A(n4252), .Y(n8067) );
  AND2X1 U6165 ( .A(n4168), .B(n4233), .Y(n4264) );
  INVX1 U6166 ( .A(n4264), .Y(n8068) );
  AND2X1 U6167 ( .A(n4142), .B(n4276), .Y(n4294) );
  INVX1 U6168 ( .A(n4294), .Y(n8069) );
  AND2X1 U6169 ( .A(n4166), .B(n4276), .Y(n4306) );
  INVX1 U6170 ( .A(n4306), .Y(n8070) );
  AND2X1 U6171 ( .A(n4132), .B(n4319), .Y(n4332) );
  INVX1 U6172 ( .A(n4332), .Y(n8071) );
  AND2X1 U6173 ( .A(n4156), .B(n4319), .Y(n4344) );
  INVX1 U6174 ( .A(n4344), .Y(n8072) );
  AND2X1 U6175 ( .A(n4180), .B(n4319), .Y(n4356) );
  INVX1 U6176 ( .A(n4356), .Y(n8073) );
  AND2X1 U6177 ( .A(n4130), .B(n4361), .Y(n4373) );
  INVX1 U6178 ( .A(n4373), .Y(n8074) );
  AND2X1 U6179 ( .A(n4154), .B(n4361), .Y(n4385) );
  INVX1 U6180 ( .A(n4385), .Y(n8075) );
  AND2X1 U6181 ( .A(n4178), .B(n4361), .Y(n4397) );
  INVX1 U6182 ( .A(n4397), .Y(n8076) );
  AND2X1 U6183 ( .A(n4128), .B(n4404), .Y(n4415) );
  INVX1 U6184 ( .A(n4415), .Y(n8077) );
  AND2X1 U6185 ( .A(n4152), .B(n4404), .Y(n4427) );
  INVX1 U6186 ( .A(n4427), .Y(n8078) );
  AND2X1 U6187 ( .A(n4176), .B(n4404), .Y(n4439) );
  INVX1 U6188 ( .A(n4439), .Y(n8079) );
  AND2X1 U6189 ( .A(n4150), .B(n4447), .Y(n4469) );
  INVX1 U6190 ( .A(n4469), .Y(n8080) );
  AND2X1 U6191 ( .A(n4174), .B(n4447), .Y(n4481) );
  INVX1 U6192 ( .A(n4481), .Y(n8081) );
  AND2X1 U6193 ( .A(n4140), .B(n4490), .Y(n4507) );
  INVX1 U6194 ( .A(n4507), .Y(n8082) );
  AND2X1 U6195 ( .A(n4164), .B(n4490), .Y(n4519) );
  INVX1 U6196 ( .A(n4519), .Y(n8083) );
  AND2X1 U6197 ( .A(n4188), .B(n4490), .Y(n4531) );
  INVX1 U6198 ( .A(n4531), .Y(n8084) );
  AND2X1 U6199 ( .A(n4138), .B(n4533), .Y(n4549) );
  INVX1 U6200 ( .A(n4549), .Y(n8085) );
  AND2X1 U6201 ( .A(n4162), .B(n4533), .Y(n4561) );
  INVX1 U6202 ( .A(n4561), .Y(n8086) );
  AND2X1 U6203 ( .A(n4186), .B(n4533), .Y(n4573) );
  INVX1 U6204 ( .A(n4573), .Y(n8087) );
  AND2X1 U6205 ( .A(n4136), .B(n4575), .Y(n4590) );
  INVX1 U6206 ( .A(n4590), .Y(n8088) );
  AND2X1 U6207 ( .A(n4160), .B(n4575), .Y(n4602) );
  INVX1 U6208 ( .A(n4602), .Y(n8089) );
  AND2X1 U6209 ( .A(n4184), .B(n4575), .Y(n4614) );
  INVX1 U6210 ( .A(n4614), .Y(n8090) );
  AND2X1 U6211 ( .A(n4134), .B(n4617), .Y(n4631) );
  INVX1 U6212 ( .A(n4631), .Y(n8091) );
  AND2X1 U6213 ( .A(n4158), .B(n4617), .Y(n4643) );
  INVX1 U6214 ( .A(n4643), .Y(n8092) );
  AND2X1 U6215 ( .A(n4182), .B(n4617), .Y(n4655) );
  INVX1 U6216 ( .A(n4655), .Y(n8093) );
  AND2X1 U6217 ( .A(n4148), .B(n4659), .Y(n4680) );
  INVX1 U6218 ( .A(n4680), .Y(n8094) );
  AND2X1 U6219 ( .A(n4172), .B(n4659), .Y(n4692) );
  INVX1 U6220 ( .A(n4692), .Y(n8095) );
  AND2X1 U6221 ( .A(n4108), .B(n4701), .Y(n4702) );
  INVX1 U6222 ( .A(n4702), .Y(n8096) );
  AND2X1 U6223 ( .A(n4146), .B(n4701), .Y(n4721) );
  INVX1 U6224 ( .A(n4721), .Y(n8097) );
  AND2X1 U6225 ( .A(n4170), .B(n4701), .Y(n4733) );
  INVX1 U6226 ( .A(n4733), .Y(n8098) );
  AND2X1 U6227 ( .A(n4144), .B(n4743), .Y(n4762) );
  INVX1 U6228 ( .A(n4762), .Y(n8099) );
  AND2X1 U6229 ( .A(n4168), .B(n4743), .Y(n4774) );
  INVX1 U6230 ( .A(n4774), .Y(n8100) );
  AND2X1 U6231 ( .A(n4142), .B(n4785), .Y(n4803) );
  INVX1 U6232 ( .A(n4803), .Y(n8101) );
  AND2X1 U6233 ( .A(n4166), .B(n4785), .Y(n4815) );
  INVX1 U6234 ( .A(n4815), .Y(n8102) );
  AND2X1 U6235 ( .A(n4132), .B(n4827), .Y(n4840) );
  INVX1 U6236 ( .A(n4840), .Y(n8103) );
  AND2X1 U6237 ( .A(n4156), .B(n4827), .Y(n4852) );
  INVX1 U6238 ( .A(n4852), .Y(n8104) );
  AND2X1 U6239 ( .A(n4180), .B(n4827), .Y(n4864) );
  INVX1 U6240 ( .A(n4864), .Y(n8105) );
  AND2X1 U6241 ( .A(n4130), .B(n4870), .Y(n4882) );
  INVX1 U6242 ( .A(n4882), .Y(n8106) );
  AND2X1 U6243 ( .A(n4154), .B(n4870), .Y(n4894) );
  INVX1 U6244 ( .A(n4894), .Y(n8107) );
  AND2X1 U6245 ( .A(n4178), .B(n4870), .Y(n4906) );
  INVX1 U6246 ( .A(n4906), .Y(n8108) );
  AND2X1 U6247 ( .A(n4128), .B(n4912), .Y(n4923) );
  INVX1 U6248 ( .A(n4923), .Y(n8109) );
  AND2X1 U6249 ( .A(n4152), .B(n4912), .Y(n4935) );
  INVX1 U6250 ( .A(n4935), .Y(n8110) );
  AND2X1 U6251 ( .A(n4176), .B(n4912), .Y(n4947) );
  INVX1 U6252 ( .A(n4947), .Y(n8111) );
  AND2X1 U6253 ( .A(n4150), .B(n4954), .Y(n4976) );
  INVX1 U6254 ( .A(n4976), .Y(n8112) );
  AND2X1 U6255 ( .A(n4174), .B(n4954), .Y(n4988) );
  INVX1 U6256 ( .A(n4988), .Y(n8113) );
  AND2X1 U6257 ( .A(n4140), .B(n4996), .Y(n5013) );
  INVX1 U6258 ( .A(n5013), .Y(n8114) );
  AND2X1 U6259 ( .A(n4164), .B(n4996), .Y(n5025) );
  INVX1 U6260 ( .A(n5025), .Y(n8115) );
  AND2X1 U6261 ( .A(n4188), .B(n4996), .Y(n5037) );
  INVX1 U6262 ( .A(n5037), .Y(n8116) );
  AND2X1 U6263 ( .A(n4138), .B(n5038), .Y(n5054) );
  INVX1 U6264 ( .A(n5054), .Y(n8117) );
  AND2X1 U6265 ( .A(n4162), .B(n5038), .Y(n5066) );
  INVX1 U6266 ( .A(n5066), .Y(n8118) );
  AND2X1 U6267 ( .A(n4186), .B(n5038), .Y(n5078) );
  INVX1 U6268 ( .A(n5078), .Y(n8119) );
  AND2X1 U6269 ( .A(n4136), .B(n5080), .Y(n5095) );
  INVX1 U6270 ( .A(n5095), .Y(n8120) );
  AND2X1 U6271 ( .A(n4160), .B(n5080), .Y(n5107) );
  INVX1 U6272 ( .A(n5107), .Y(n8121) );
  AND2X1 U6273 ( .A(n4184), .B(n5080), .Y(n5119) );
  INVX1 U6274 ( .A(n5119), .Y(n8122) );
  AND2X1 U6275 ( .A(n4134), .B(n5122), .Y(n5136) );
  INVX1 U6276 ( .A(n5136), .Y(n8123) );
  AND2X1 U6277 ( .A(n4158), .B(n5122), .Y(n5148) );
  INVX1 U6278 ( .A(n5148), .Y(n8124) );
  AND2X1 U6279 ( .A(n4182), .B(n5122), .Y(n5160) );
  INVX1 U6280 ( .A(n5160), .Y(n8125) );
  AND2X1 U6281 ( .A(n4132), .B(n5164), .Y(n5177) );
  INVX1 U6282 ( .A(n5177), .Y(n8126) );
  AND2X1 U6283 ( .A(n4156), .B(n5164), .Y(n5189) );
  INVX1 U6284 ( .A(n5189), .Y(n8127) );
  AND2X1 U6285 ( .A(n4180), .B(n5164), .Y(n5201) );
  INVX1 U6286 ( .A(n5201), .Y(n8128) );
  AND2X1 U6287 ( .A(n4130), .B(n5207), .Y(n5219) );
  INVX1 U6288 ( .A(n5219), .Y(n8129) );
  AND2X1 U6289 ( .A(n4154), .B(n5207), .Y(n5231) );
  INVX1 U6290 ( .A(n5231), .Y(n8130) );
  AND2X1 U6291 ( .A(n4178), .B(n5207), .Y(n5243) );
  INVX1 U6292 ( .A(n5243), .Y(n8131) );
  AND2X1 U6293 ( .A(n4128), .B(n5249), .Y(n5260) );
  INVX1 U6294 ( .A(n5260), .Y(n8132) );
  AND2X1 U6295 ( .A(n4152), .B(n5249), .Y(n5272) );
  INVX1 U6296 ( .A(n5272), .Y(n8133) );
  AND2X1 U6297 ( .A(n4176), .B(n5249), .Y(n5284) );
  INVX1 U6298 ( .A(n5284), .Y(n8134) );
  AND2X1 U6299 ( .A(n4150), .B(n5291), .Y(n5313) );
  INVX1 U6300 ( .A(n5313), .Y(n8135) );
  AND2X1 U6301 ( .A(n4174), .B(n5291), .Y(n5325) );
  INVX1 U6302 ( .A(n5325), .Y(n8136) );
  AND2X1 U6303 ( .A(n4140), .B(n5333), .Y(n5350) );
  INVX1 U6304 ( .A(n5350), .Y(n8137) );
  AND2X1 U6305 ( .A(n4164), .B(n5333), .Y(n5362) );
  INVX1 U6306 ( .A(n5362), .Y(n8138) );
  AND2X1 U6307 ( .A(n4188), .B(n5333), .Y(n5374) );
  INVX1 U6308 ( .A(n5374), .Y(n8139) );
  AND2X1 U6309 ( .A(n4138), .B(n5375), .Y(n5391) );
  INVX1 U6310 ( .A(n5391), .Y(n8140) );
  AND2X1 U6311 ( .A(n4162), .B(n5375), .Y(n5403) );
  INVX1 U6312 ( .A(n5403), .Y(n8141) );
  AND2X1 U6313 ( .A(n4186), .B(n5375), .Y(n5415) );
  INVX1 U6314 ( .A(n5415), .Y(n8142) );
  AND2X1 U6315 ( .A(n4136), .B(n5417), .Y(n5432) );
  INVX1 U6316 ( .A(n5432), .Y(n8143) );
  AND2X1 U6317 ( .A(n4160), .B(n5417), .Y(n5444) );
  INVX1 U6318 ( .A(n5444), .Y(n8144) );
  AND2X1 U6319 ( .A(n4184), .B(n5417), .Y(n5456) );
  INVX1 U6320 ( .A(n5456), .Y(n8145) );
  AND2X1 U6321 ( .A(n4134), .B(n5459), .Y(n5473) );
  INVX1 U6322 ( .A(n5473), .Y(n8146) );
  AND2X1 U6323 ( .A(n4158), .B(n5459), .Y(n5485) );
  INVX1 U6324 ( .A(n5485), .Y(n8147) );
  AND2X1 U6325 ( .A(n4182), .B(n5459), .Y(n5497) );
  INVX1 U6326 ( .A(n5497), .Y(n8148) );
  INVX1 U6327 ( .A(n4082), .Y(n8149) );
  INVX1 U6328 ( .A(n4089), .Y(n8150) );
  BUFX2 U6329 ( .A(n5721), .Y(empty_bar) );
  BUFX2 U6330 ( .A(n4489), .Y(n8152) );
  BUFX2 U6331 ( .A(n4105), .Y(n8153) );
  AND2X1 U6332 ( .A(n4108), .B(n4106), .Y(n4107) );
  INVX1 U6333 ( .A(n4107), .Y(n8154) );
  AND2X1 U6334 ( .A(n4146), .B(n4106), .Y(n4145) );
  INVX1 U6335 ( .A(n4145), .Y(n8155) );
  AND2X1 U6336 ( .A(n4170), .B(n4106), .Y(n4169) );
  INVX1 U6337 ( .A(n4169), .Y(n8156) );
  AND2X1 U6338 ( .A(n4148), .B(n4190), .Y(n4211) );
  INVX1 U6339 ( .A(n4211), .Y(n8157) );
  AND2X1 U6340 ( .A(n4172), .B(n4190), .Y(n4223) );
  INVX1 U6341 ( .A(n4223), .Y(n8158) );
  AND2X1 U6342 ( .A(n4142), .B(n4233), .Y(n4251) );
  INVX1 U6343 ( .A(n4251), .Y(n8159) );
  AND2X1 U6344 ( .A(n4166), .B(n4233), .Y(n4263) );
  INVX1 U6345 ( .A(n4263), .Y(n8160) );
  AND2X1 U6346 ( .A(n4144), .B(n4276), .Y(n4295) );
  INVX1 U6347 ( .A(n4295), .Y(n8161) );
  AND2X1 U6348 ( .A(n4168), .B(n4276), .Y(n4307) );
  INVX1 U6349 ( .A(n4307), .Y(n8162) );
  AND2X1 U6350 ( .A(n4130), .B(n4319), .Y(n4331) );
  INVX1 U6351 ( .A(n4331), .Y(n8163) );
  AND2X1 U6352 ( .A(n4154), .B(n4319), .Y(n4343) );
  INVX1 U6353 ( .A(n4343), .Y(n8164) );
  AND2X1 U6354 ( .A(n4178), .B(n4319), .Y(n4355) );
  INVX1 U6355 ( .A(n4355), .Y(n8165) );
  AND2X1 U6356 ( .A(n4132), .B(n4361), .Y(n4374) );
  INVX1 U6357 ( .A(n4374), .Y(n8166) );
  AND2X1 U6358 ( .A(n4156), .B(n4361), .Y(n4386) );
  INVX1 U6359 ( .A(n4386), .Y(n8167) );
  AND2X1 U6360 ( .A(n4180), .B(n4361), .Y(n4398) );
  INVX1 U6361 ( .A(n4398), .Y(n8168) );
  AND2X1 U6362 ( .A(n4150), .B(n4404), .Y(n4426) );
  INVX1 U6363 ( .A(n4426), .Y(n8169) );
  AND2X1 U6364 ( .A(n4174), .B(n4404), .Y(n4438) );
  INVX1 U6365 ( .A(n4438), .Y(n8170) );
  AND2X1 U6366 ( .A(n4128), .B(n4447), .Y(n4458) );
  INVX1 U6367 ( .A(n4458), .Y(n8171) );
  AND2X1 U6368 ( .A(n4152), .B(n4447), .Y(n4470) );
  INVX1 U6369 ( .A(n4470), .Y(n8172) );
  AND2X1 U6370 ( .A(n4176), .B(n4447), .Y(n4482) );
  INVX1 U6371 ( .A(n4482), .Y(n8173) );
  AND2X1 U6372 ( .A(n4138), .B(n4490), .Y(n4506) );
  INVX1 U6373 ( .A(n4506), .Y(n8174) );
  AND2X1 U6374 ( .A(n4162), .B(n4490), .Y(n4518) );
  INVX1 U6375 ( .A(n4518), .Y(n8175) );
  AND2X1 U6376 ( .A(n4186), .B(n4490), .Y(n4530) );
  INVX1 U6377 ( .A(n4530), .Y(n8176) );
  AND2X1 U6378 ( .A(n4140), .B(n4533), .Y(n4550) );
  INVX1 U6379 ( .A(n4550), .Y(n8177) );
  AND2X1 U6380 ( .A(n4164), .B(n4533), .Y(n4562) );
  INVX1 U6381 ( .A(n4562), .Y(n8178) );
  AND2X1 U6382 ( .A(n4188), .B(n4533), .Y(n4574) );
  INVX1 U6383 ( .A(n4574), .Y(n8179) );
  AND2X1 U6384 ( .A(n4134), .B(n4575), .Y(n4589) );
  INVX1 U6385 ( .A(n4589), .Y(n8180) );
  AND2X1 U6386 ( .A(n4158), .B(n4575), .Y(n4601) );
  INVX1 U6387 ( .A(n4601), .Y(n8181) );
  AND2X1 U6388 ( .A(n4182), .B(n4575), .Y(n4613) );
  INVX1 U6389 ( .A(n4613), .Y(n8182) );
  AND2X1 U6390 ( .A(n4136), .B(n4617), .Y(n4632) );
  INVX1 U6391 ( .A(n4632), .Y(n8183) );
  AND2X1 U6392 ( .A(n4160), .B(n4617), .Y(n4644) );
  INVX1 U6393 ( .A(n4644), .Y(n8184) );
  AND2X1 U6394 ( .A(n4184), .B(n4617), .Y(n4656) );
  INVX1 U6395 ( .A(n4656), .Y(n8185) );
  AND2X1 U6396 ( .A(n4108), .B(n4659), .Y(n4660) );
  INVX1 U6397 ( .A(n4660), .Y(n8186) );
  AND2X1 U6398 ( .A(n4146), .B(n4659), .Y(n4679) );
  INVX1 U6399 ( .A(n4679), .Y(n8187) );
  AND2X1 U6400 ( .A(n4170), .B(n4659), .Y(n4691) );
  INVX1 U6401 ( .A(n4691), .Y(n8188) );
  AND2X1 U6402 ( .A(n4148), .B(n4701), .Y(n4722) );
  INVX1 U6403 ( .A(n4722), .Y(n8189) );
  AND2X1 U6404 ( .A(n4172), .B(n4701), .Y(n4734) );
  INVX1 U6405 ( .A(n4734), .Y(n8190) );
  AND2X1 U6406 ( .A(n4142), .B(n4743), .Y(n4761) );
  INVX1 U6407 ( .A(n4761), .Y(n8191) );
  AND2X1 U6408 ( .A(n4166), .B(n4743), .Y(n4773) );
  INVX1 U6409 ( .A(n4773), .Y(n8192) );
  AND2X1 U6410 ( .A(n4144), .B(n4785), .Y(n4804) );
  INVX1 U6411 ( .A(n4804), .Y(n8193) );
  AND2X1 U6412 ( .A(n4168), .B(n4785), .Y(n4816) );
  INVX1 U6413 ( .A(n4816), .Y(n8194) );
  AND2X1 U6414 ( .A(n4130), .B(n4827), .Y(n4839) );
  INVX1 U6415 ( .A(n4839), .Y(n8195) );
  AND2X1 U6416 ( .A(n4154), .B(n4827), .Y(n4851) );
  INVX1 U6417 ( .A(n4851), .Y(n8196) );
  AND2X1 U6418 ( .A(n4178), .B(n4827), .Y(n4863) );
  INVX1 U6419 ( .A(n4863), .Y(n8197) );
  AND2X1 U6420 ( .A(n4132), .B(n4870), .Y(n4883) );
  INVX1 U6421 ( .A(n4883), .Y(n8198) );
  AND2X1 U6422 ( .A(n4156), .B(n4870), .Y(n4895) );
  INVX1 U6423 ( .A(n4895), .Y(n8199) );
  AND2X1 U6424 ( .A(n4180), .B(n4870), .Y(n4907) );
  INVX1 U6425 ( .A(n4907), .Y(n8200) );
  AND2X1 U6426 ( .A(n4150), .B(n4912), .Y(n4934) );
  INVX1 U6427 ( .A(n4934), .Y(n8201) );
  AND2X1 U6428 ( .A(n4174), .B(n4912), .Y(n4946) );
  INVX1 U6429 ( .A(n4946), .Y(n8202) );
  AND2X1 U6430 ( .A(n4128), .B(n4954), .Y(n4965) );
  INVX1 U6431 ( .A(n4965), .Y(n8203) );
  AND2X1 U6432 ( .A(n4152), .B(n4954), .Y(n4977) );
  INVX1 U6433 ( .A(n4977), .Y(n8204) );
  AND2X1 U6434 ( .A(n4176), .B(n4954), .Y(n4989) );
  INVX1 U6435 ( .A(n4989), .Y(n8205) );
  AND2X1 U6436 ( .A(n4138), .B(n4996), .Y(n5012) );
  INVX1 U6437 ( .A(n5012), .Y(n8206) );
  AND2X1 U6438 ( .A(n4162), .B(n4996), .Y(n5024) );
  INVX1 U6439 ( .A(n5024), .Y(n8207) );
  AND2X1 U6440 ( .A(n4186), .B(n4996), .Y(n5036) );
  INVX1 U6441 ( .A(n5036), .Y(n8208) );
  AND2X1 U6442 ( .A(n4140), .B(n5038), .Y(n5055) );
  INVX1 U6443 ( .A(n5055), .Y(n8209) );
  AND2X1 U6444 ( .A(n4164), .B(n5038), .Y(n5067) );
  INVX1 U6445 ( .A(n5067), .Y(n8210) );
  AND2X1 U6446 ( .A(n4188), .B(n5038), .Y(n5079) );
  INVX1 U6447 ( .A(n5079), .Y(n8211) );
  AND2X1 U6448 ( .A(n4134), .B(n5080), .Y(n5094) );
  INVX1 U6449 ( .A(n5094), .Y(n8212) );
  AND2X1 U6450 ( .A(n4158), .B(n5080), .Y(n5106) );
  INVX1 U6451 ( .A(n5106), .Y(n8213) );
  AND2X1 U6452 ( .A(n4182), .B(n5080), .Y(n5118) );
  INVX1 U6453 ( .A(n5118), .Y(n8214) );
  AND2X1 U6454 ( .A(n4136), .B(n5122), .Y(n5137) );
  INVX1 U6455 ( .A(n5137), .Y(n8215) );
  AND2X1 U6456 ( .A(n4160), .B(n5122), .Y(n5149) );
  INVX1 U6457 ( .A(n5149), .Y(n8216) );
  AND2X1 U6458 ( .A(n4184), .B(n5122), .Y(n5161) );
  INVX1 U6459 ( .A(n5161), .Y(n8217) );
  AND2X1 U6460 ( .A(n4130), .B(n5164), .Y(n5176) );
  INVX1 U6461 ( .A(n5176), .Y(n8218) );
  AND2X1 U6462 ( .A(n4154), .B(n5164), .Y(n5188) );
  INVX1 U6463 ( .A(n5188), .Y(n8219) );
  AND2X1 U6464 ( .A(n4178), .B(n5164), .Y(n5200) );
  INVX1 U6465 ( .A(n5200), .Y(n8220) );
  AND2X1 U6466 ( .A(n4132), .B(n5207), .Y(n5220) );
  INVX1 U6467 ( .A(n5220), .Y(n8221) );
  AND2X1 U6468 ( .A(n4156), .B(n5207), .Y(n5232) );
  INVX1 U6469 ( .A(n5232), .Y(n8222) );
  AND2X1 U6470 ( .A(n4180), .B(n5207), .Y(n5244) );
  INVX1 U6471 ( .A(n5244), .Y(n8223) );
  AND2X1 U6472 ( .A(n4150), .B(n5249), .Y(n5271) );
  INVX1 U6473 ( .A(n5271), .Y(n8224) );
  AND2X1 U6474 ( .A(n4174), .B(n5249), .Y(n5283) );
  INVX1 U6475 ( .A(n5283), .Y(n8225) );
  AND2X1 U6476 ( .A(n4128), .B(n5291), .Y(n5302) );
  INVX1 U6477 ( .A(n5302), .Y(n8226) );
  AND2X1 U6478 ( .A(n4152), .B(n5291), .Y(n5314) );
  INVX1 U6479 ( .A(n5314), .Y(n8227) );
  AND2X1 U6480 ( .A(n4176), .B(n5291), .Y(n5326) );
  INVX1 U6481 ( .A(n5326), .Y(n8228) );
  AND2X1 U6482 ( .A(n4138), .B(n5333), .Y(n5349) );
  INVX1 U6483 ( .A(n5349), .Y(n8229) );
  AND2X1 U6484 ( .A(n4162), .B(n5333), .Y(n5361) );
  INVX1 U6485 ( .A(n5361), .Y(n8230) );
  AND2X1 U6486 ( .A(n4186), .B(n5333), .Y(n5373) );
  INVX1 U6487 ( .A(n5373), .Y(n8231) );
  AND2X1 U6488 ( .A(n4140), .B(n5375), .Y(n5392) );
  INVX1 U6489 ( .A(n5392), .Y(n8232) );
  AND2X1 U6490 ( .A(n4164), .B(n5375), .Y(n5404) );
  INVX1 U6491 ( .A(n5404), .Y(n8233) );
  AND2X1 U6492 ( .A(n4188), .B(n5375), .Y(n5416) );
  INVX1 U6493 ( .A(n5416), .Y(n8234) );
  AND2X1 U6494 ( .A(n4134), .B(n5417), .Y(n5431) );
  INVX1 U6495 ( .A(n5431), .Y(n8235) );
  AND2X1 U6496 ( .A(n4158), .B(n5417), .Y(n5443) );
  INVX1 U6497 ( .A(n5443), .Y(n8236) );
  AND2X1 U6498 ( .A(n4182), .B(n5417), .Y(n5455) );
  INVX1 U6499 ( .A(n5455), .Y(n8237) );
  AND2X1 U6500 ( .A(n4136), .B(n5459), .Y(n5474) );
  INVX1 U6501 ( .A(n5474), .Y(n8238) );
  AND2X1 U6502 ( .A(n4160), .B(n5459), .Y(n5486) );
  INVX1 U6503 ( .A(n5486), .Y(n8239) );
  AND2X1 U6504 ( .A(n4184), .B(n5459), .Y(n5498) );
  INVX1 U6505 ( .A(n5498), .Y(n8240) );
  INVX1 U6506 ( .A(n4062), .Y(n8241) );
  BUFX2 U6507 ( .A(n4318), .Y(n8242) );
  BUFX2 U6508 ( .A(n4103), .Y(n8243) );
  AND2X1 U6509 ( .A(n4144), .B(n4106), .Y(n4143) );
  INVX1 U6510 ( .A(n4143), .Y(n8244) );
  AND2X1 U6511 ( .A(n4168), .B(n4106), .Y(n4167) );
  INVX1 U6512 ( .A(n4167), .Y(n8245) );
  AND2X1 U6513 ( .A(n4142), .B(n4190), .Y(n4208) );
  INVX1 U6514 ( .A(n4208), .Y(n8246) );
  AND2X1 U6515 ( .A(n4166), .B(n4190), .Y(n4220) );
  INVX1 U6516 ( .A(n4220), .Y(n8247) );
  AND2X1 U6517 ( .A(n4148), .B(n4233), .Y(n4254) );
  INVX1 U6518 ( .A(n4254), .Y(n8248) );
  AND2X1 U6519 ( .A(n4172), .B(n4233), .Y(n4266) );
  INVX1 U6520 ( .A(n4266), .Y(n8249) );
  AND2X1 U6521 ( .A(n4108), .B(n4276), .Y(n4277) );
  INVX1 U6522 ( .A(n4277), .Y(n8250) );
  AND2X1 U6523 ( .A(n4146), .B(n4276), .Y(n4296) );
  INVX1 U6524 ( .A(n4296), .Y(n8251) );
  AND2X1 U6525 ( .A(n4170), .B(n4276), .Y(n4308) );
  INVX1 U6526 ( .A(n4308), .Y(n8252) );
  AND2X1 U6527 ( .A(n4128), .B(n4319), .Y(n4330) );
  INVX1 U6528 ( .A(n4330), .Y(n8253) );
  AND2X1 U6529 ( .A(n4152), .B(n4319), .Y(n4342) );
  INVX1 U6530 ( .A(n4342), .Y(n8254) );
  AND2X1 U6531 ( .A(n4176), .B(n4319), .Y(n4354) );
  INVX1 U6532 ( .A(n4354), .Y(n8255) );
  AND2X1 U6533 ( .A(n4150), .B(n4361), .Y(n4383) );
  INVX1 U6534 ( .A(n4383), .Y(n8256) );
  AND2X1 U6535 ( .A(n4174), .B(n4361), .Y(n4395) );
  INVX1 U6536 ( .A(n4395), .Y(n8257) );
  AND2X1 U6537 ( .A(n4132), .B(n4404), .Y(n4417) );
  INVX1 U6538 ( .A(n4417), .Y(n8258) );
  AND2X1 U6539 ( .A(n4156), .B(n4404), .Y(n4429) );
  INVX1 U6540 ( .A(n4429), .Y(n8259) );
  AND2X1 U6541 ( .A(n4180), .B(n4404), .Y(n4441) );
  INVX1 U6542 ( .A(n4441), .Y(n8260) );
  AND2X1 U6543 ( .A(n4130), .B(n4447), .Y(n4459) );
  INVX1 U6544 ( .A(n4459), .Y(n8261) );
  AND2X1 U6545 ( .A(n4154), .B(n4447), .Y(n4471) );
  INVX1 U6546 ( .A(n4471), .Y(n8262) );
  AND2X1 U6547 ( .A(n4178), .B(n4447), .Y(n4483) );
  INVX1 U6548 ( .A(n4483), .Y(n8263) );
  AND2X1 U6549 ( .A(n4136), .B(n4490), .Y(n4505) );
  INVX1 U6550 ( .A(n4505), .Y(n8264) );
  AND2X1 U6551 ( .A(n4160), .B(n4490), .Y(n4517) );
  INVX1 U6552 ( .A(n4517), .Y(n8265) );
  AND2X1 U6553 ( .A(n4184), .B(n4490), .Y(n4529) );
  INVX1 U6554 ( .A(n4529), .Y(n8266) );
  AND2X1 U6555 ( .A(n4134), .B(n4533), .Y(n4547) );
  INVX1 U6556 ( .A(n4547), .Y(n8267) );
  AND2X1 U6557 ( .A(n4158), .B(n4533), .Y(n4559) );
  INVX1 U6558 ( .A(n4559), .Y(n8268) );
  AND2X1 U6559 ( .A(n4182), .B(n4533), .Y(n4571) );
  INVX1 U6560 ( .A(n4571), .Y(n8269) );
  AND2X1 U6561 ( .A(n4140), .B(n4575), .Y(n4592) );
  INVX1 U6562 ( .A(n4592), .Y(n8270) );
  AND2X1 U6563 ( .A(n4164), .B(n4575), .Y(n4604) );
  INVX1 U6564 ( .A(n4604), .Y(n8271) );
  AND2X1 U6565 ( .A(n4188), .B(n4575), .Y(n4616) );
  INVX1 U6566 ( .A(n4616), .Y(n8272) );
  AND2X1 U6567 ( .A(n4138), .B(n4617), .Y(n4633) );
  INVX1 U6568 ( .A(n4633), .Y(n8273) );
  AND2X1 U6569 ( .A(n4162), .B(n4617), .Y(n4645) );
  INVX1 U6570 ( .A(n4645), .Y(n8274) );
  AND2X1 U6571 ( .A(n4186), .B(n4617), .Y(n4657) );
  INVX1 U6572 ( .A(n4657), .Y(n8275) );
  AND2X1 U6573 ( .A(n4144), .B(n4659), .Y(n4678) );
  INVX1 U6574 ( .A(n4678), .Y(n8276) );
  AND2X1 U6575 ( .A(n4168), .B(n4659), .Y(n4690) );
  INVX1 U6576 ( .A(n4690), .Y(n8277) );
  AND2X1 U6577 ( .A(n4142), .B(n4701), .Y(n4719) );
  INVX1 U6578 ( .A(n4719), .Y(n8278) );
  AND2X1 U6579 ( .A(n4166), .B(n4701), .Y(n4731) );
  INVX1 U6580 ( .A(n4731), .Y(n8279) );
  AND2X1 U6581 ( .A(n4148), .B(n4743), .Y(n4764) );
  INVX1 U6582 ( .A(n4764), .Y(n8280) );
  AND2X1 U6583 ( .A(n4172), .B(n4743), .Y(n4776) );
  INVX1 U6584 ( .A(n4776), .Y(n8281) );
  AND2X1 U6585 ( .A(n4108), .B(n4785), .Y(n4786) );
  INVX1 U6586 ( .A(n4786), .Y(n8282) );
  AND2X1 U6587 ( .A(n4146), .B(n4785), .Y(n4805) );
  INVX1 U6588 ( .A(n4805), .Y(n8283) );
  AND2X1 U6589 ( .A(n4170), .B(n4785), .Y(n4817) );
  INVX1 U6590 ( .A(n4817), .Y(n8284) );
  AND2X1 U6591 ( .A(n4128), .B(n4827), .Y(n4838) );
  INVX1 U6592 ( .A(n4838), .Y(n8285) );
  AND2X1 U6593 ( .A(n4152), .B(n4827), .Y(n4850) );
  INVX1 U6594 ( .A(n4850), .Y(n8286) );
  AND2X1 U6595 ( .A(n4176), .B(n4827), .Y(n4862) );
  INVX1 U6596 ( .A(n4862), .Y(n8287) );
  AND2X1 U6597 ( .A(n4150), .B(n4870), .Y(n4892) );
  INVX1 U6598 ( .A(n4892), .Y(n8288) );
  AND2X1 U6599 ( .A(n4174), .B(n4870), .Y(n4904) );
  INVX1 U6600 ( .A(n4904), .Y(n8289) );
  AND2X1 U6601 ( .A(n4132), .B(n4912), .Y(n4925) );
  INVX1 U6602 ( .A(n4925), .Y(n8290) );
  AND2X1 U6603 ( .A(n4156), .B(n4912), .Y(n4937) );
  INVX1 U6604 ( .A(n4937), .Y(n8291) );
  AND2X1 U6605 ( .A(n4180), .B(n4912), .Y(n4949) );
  INVX1 U6606 ( .A(n4949), .Y(n8292) );
  AND2X1 U6607 ( .A(n4130), .B(n4954), .Y(n4966) );
  INVX1 U6608 ( .A(n4966), .Y(n8293) );
  AND2X1 U6609 ( .A(n4154), .B(n4954), .Y(n4978) );
  INVX1 U6610 ( .A(n4978), .Y(n8294) );
  AND2X1 U6611 ( .A(n4178), .B(n4954), .Y(n4990) );
  INVX1 U6612 ( .A(n4990), .Y(n8295) );
  AND2X1 U6613 ( .A(n4136), .B(n4996), .Y(n5011) );
  INVX1 U6614 ( .A(n5011), .Y(n8296) );
  AND2X1 U6615 ( .A(n4160), .B(n4996), .Y(n5023) );
  INVX1 U6616 ( .A(n5023), .Y(n8297) );
  AND2X1 U6617 ( .A(n4184), .B(n4996), .Y(n5035) );
  INVX1 U6618 ( .A(n5035), .Y(n8298) );
  AND2X1 U6619 ( .A(n4134), .B(n5038), .Y(n5052) );
  INVX1 U6620 ( .A(n5052), .Y(n8299) );
  AND2X1 U6621 ( .A(n4158), .B(n5038), .Y(n5064) );
  INVX1 U6622 ( .A(n5064), .Y(n8300) );
  AND2X1 U6623 ( .A(n4182), .B(n5038), .Y(n5076) );
  INVX1 U6624 ( .A(n5076), .Y(n8301) );
  AND2X1 U6625 ( .A(n4140), .B(n5080), .Y(n5097) );
  INVX1 U6626 ( .A(n5097), .Y(n8302) );
  AND2X1 U6627 ( .A(n4164), .B(n5080), .Y(n5109) );
  INVX1 U6628 ( .A(n5109), .Y(n8303) );
  AND2X1 U6629 ( .A(n4188), .B(n5080), .Y(n5121) );
  INVX1 U6630 ( .A(n5121), .Y(n8304) );
  AND2X1 U6631 ( .A(n4138), .B(n5122), .Y(n5138) );
  INVX1 U6632 ( .A(n5138), .Y(n8305) );
  AND2X1 U6633 ( .A(n4162), .B(n5122), .Y(n5150) );
  INVX1 U6634 ( .A(n5150), .Y(n8306) );
  AND2X1 U6635 ( .A(n4186), .B(n5122), .Y(n5162) );
  INVX1 U6636 ( .A(n5162), .Y(n8307) );
  AND2X1 U6637 ( .A(n4128), .B(n5164), .Y(n5175) );
  INVX1 U6638 ( .A(n5175), .Y(n8308) );
  AND2X1 U6639 ( .A(n4152), .B(n5164), .Y(n5187) );
  INVX1 U6640 ( .A(n5187), .Y(n8309) );
  AND2X1 U6641 ( .A(n4176), .B(n5164), .Y(n5199) );
  INVX1 U6642 ( .A(n5199), .Y(n8310) );
  AND2X1 U6643 ( .A(n4150), .B(n5207), .Y(n5229) );
  INVX1 U6644 ( .A(n5229), .Y(n8311) );
  AND2X1 U6645 ( .A(n4174), .B(n5207), .Y(n5241) );
  INVX1 U6646 ( .A(n5241), .Y(n8312) );
  AND2X1 U6647 ( .A(n4132), .B(n5249), .Y(n5262) );
  INVX1 U6648 ( .A(n5262), .Y(n8313) );
  AND2X1 U6649 ( .A(n4156), .B(n5249), .Y(n5274) );
  INVX1 U6650 ( .A(n5274), .Y(n8314) );
  AND2X1 U6651 ( .A(n4180), .B(n5249), .Y(n5286) );
  INVX1 U6652 ( .A(n5286), .Y(n8315) );
  AND2X1 U6653 ( .A(n4130), .B(n5291), .Y(n5303) );
  INVX1 U6654 ( .A(n5303), .Y(n8316) );
  AND2X1 U6655 ( .A(n4154), .B(n5291), .Y(n5315) );
  INVX1 U6656 ( .A(n5315), .Y(n8317) );
  AND2X1 U6657 ( .A(n4178), .B(n5291), .Y(n5327) );
  INVX1 U6658 ( .A(n5327), .Y(n8318) );
  AND2X1 U6659 ( .A(n4136), .B(n5333), .Y(n5348) );
  INVX1 U6660 ( .A(n5348), .Y(n8319) );
  AND2X1 U6661 ( .A(n4160), .B(n5333), .Y(n5360) );
  INVX1 U6662 ( .A(n5360), .Y(n8320) );
  AND2X1 U6663 ( .A(n4184), .B(n5333), .Y(n5372) );
  INVX1 U6664 ( .A(n5372), .Y(n8321) );
  AND2X1 U6665 ( .A(n4134), .B(n5375), .Y(n5389) );
  INVX1 U6666 ( .A(n5389), .Y(n8322) );
  AND2X1 U6667 ( .A(n4158), .B(n5375), .Y(n5401) );
  INVX1 U6668 ( .A(n5401), .Y(n8323) );
  AND2X1 U6669 ( .A(n4182), .B(n5375), .Y(n5413) );
  INVX1 U6670 ( .A(n5413), .Y(n8324) );
  AND2X1 U6671 ( .A(n4140), .B(n5417), .Y(n5434) );
  INVX1 U6672 ( .A(n5434), .Y(n8325) );
  AND2X1 U6673 ( .A(n4164), .B(n5417), .Y(n5446) );
  INVX1 U6674 ( .A(n5446), .Y(n8326) );
  AND2X1 U6675 ( .A(n4188), .B(n5417), .Y(n5458) );
  INVX1 U6676 ( .A(n5458), .Y(n8327) );
  AND2X1 U6677 ( .A(n4138), .B(n5459), .Y(n5475) );
  INVX1 U6678 ( .A(n5475), .Y(n8328) );
  AND2X1 U6679 ( .A(n4162), .B(n5459), .Y(n5487) );
  INVX1 U6680 ( .A(n5487), .Y(n8329) );
  AND2X1 U6681 ( .A(n4186), .B(n5459), .Y(n5499) );
  INVX1 U6682 ( .A(n5499), .Y(n8330) );
  BUFX2 U6683 ( .A(n4081), .Y(n8331) );
  AND2X1 U6684 ( .A(n8500), .B(n9831), .Y(n4078) );
  INVX1 U6685 ( .A(n4078), .Y(n8332) );
  BUFX2 U6686 ( .A(n4532), .Y(n8333) );
  BUFX2 U6687 ( .A(n4869), .Y(n8334) );
  AND2X1 U6688 ( .A(n4142), .B(n4106), .Y(n4141) );
  INVX1 U6689 ( .A(n4141), .Y(n8335) );
  AND2X1 U6690 ( .A(n4166), .B(n4106), .Y(n4165) );
  INVX1 U6691 ( .A(n4165), .Y(n8336) );
  AND2X1 U6692 ( .A(n4144), .B(n4190), .Y(n4209) );
  INVX1 U6693 ( .A(n4209), .Y(n8337) );
  AND2X1 U6694 ( .A(n4168), .B(n4190), .Y(n4221) );
  INVX1 U6695 ( .A(n4221), .Y(n8338) );
  AND2X1 U6696 ( .A(n4108), .B(n4233), .Y(n4234) );
  INVX1 U6697 ( .A(n4234), .Y(n8339) );
  AND2X1 U6698 ( .A(n4146), .B(n4233), .Y(n4253) );
  INVX1 U6699 ( .A(n4253), .Y(n8340) );
  AND2X1 U6700 ( .A(n4170), .B(n4233), .Y(n4265) );
  INVX1 U6701 ( .A(n4265), .Y(n8341) );
  AND2X1 U6702 ( .A(n4148), .B(n4276), .Y(n4297) );
  INVX1 U6703 ( .A(n4297), .Y(n8342) );
  AND2X1 U6704 ( .A(n4172), .B(n4276), .Y(n4309) );
  INVX1 U6705 ( .A(n4309), .Y(n8343) );
  AND2X1 U6706 ( .A(n4150), .B(n4319), .Y(n4341) );
  INVX1 U6707 ( .A(n4341), .Y(n8344) );
  AND2X1 U6708 ( .A(n4174), .B(n4319), .Y(n4353) );
  INVX1 U6709 ( .A(n4353), .Y(n8345) );
  AND2X1 U6710 ( .A(n4128), .B(n4361), .Y(n4372) );
  INVX1 U6711 ( .A(n4372), .Y(n8346) );
  AND2X1 U6712 ( .A(n4152), .B(n4361), .Y(n4384) );
  INVX1 U6713 ( .A(n4384), .Y(n8347) );
  AND2X1 U6714 ( .A(n4176), .B(n4361), .Y(n4396) );
  INVX1 U6715 ( .A(n4396), .Y(n8348) );
  AND2X1 U6716 ( .A(n4130), .B(n4404), .Y(n4416) );
  INVX1 U6717 ( .A(n4416), .Y(n8349) );
  AND2X1 U6718 ( .A(n4154), .B(n4404), .Y(n4428) );
  INVX1 U6719 ( .A(n4428), .Y(n8350) );
  AND2X1 U6720 ( .A(n4178), .B(n4404), .Y(n4440) );
  INVX1 U6721 ( .A(n4440), .Y(n8351) );
  AND2X1 U6722 ( .A(n4132), .B(n4447), .Y(n4460) );
  INVX1 U6723 ( .A(n4460), .Y(n8352) );
  AND2X1 U6724 ( .A(n4156), .B(n4447), .Y(n4472) );
  INVX1 U6725 ( .A(n4472), .Y(n8353) );
  AND2X1 U6726 ( .A(n4180), .B(n4447), .Y(n4484) );
  INVX1 U6727 ( .A(n4484), .Y(n8354) );
  AND2X1 U6728 ( .A(n4134), .B(n4490), .Y(n4504) );
  INVX1 U6729 ( .A(n4504), .Y(n8355) );
  AND2X1 U6730 ( .A(n4158), .B(n4490), .Y(n4516) );
  INVX1 U6731 ( .A(n4516), .Y(n8356) );
  AND2X1 U6732 ( .A(n4182), .B(n4490), .Y(n4528) );
  INVX1 U6733 ( .A(n4528), .Y(n8357) );
  AND2X1 U6734 ( .A(n4136), .B(n4533), .Y(n4548) );
  INVX1 U6735 ( .A(n4548), .Y(n8358) );
  AND2X1 U6736 ( .A(n4160), .B(n4533), .Y(n4560) );
  INVX1 U6737 ( .A(n4560), .Y(n8359) );
  AND2X1 U6738 ( .A(n4184), .B(n4533), .Y(n4572) );
  INVX1 U6739 ( .A(n4572), .Y(n8360) );
  AND2X1 U6740 ( .A(n4138), .B(n4575), .Y(n4591) );
  INVX1 U6741 ( .A(n4591), .Y(n8361) );
  AND2X1 U6742 ( .A(n4162), .B(n4575), .Y(n4603) );
  INVX1 U6743 ( .A(n4603), .Y(n8362) );
  AND2X1 U6744 ( .A(n4186), .B(n4575), .Y(n4615) );
  INVX1 U6745 ( .A(n4615), .Y(n8363) );
  AND2X1 U6746 ( .A(n4140), .B(n4617), .Y(n4634) );
  INVX1 U6747 ( .A(n4634), .Y(n8364) );
  AND2X1 U6748 ( .A(n4164), .B(n4617), .Y(n4646) );
  INVX1 U6749 ( .A(n4646), .Y(n8365) );
  AND2X1 U6750 ( .A(n4188), .B(n4617), .Y(n4658) );
  INVX1 U6751 ( .A(n4658), .Y(n8366) );
  AND2X1 U6752 ( .A(n4142), .B(n4659), .Y(n4677) );
  INVX1 U6753 ( .A(n4677), .Y(n8367) );
  AND2X1 U6754 ( .A(n4166), .B(n4659), .Y(n4689) );
  INVX1 U6755 ( .A(n4689), .Y(n8368) );
  AND2X1 U6756 ( .A(n4144), .B(n4701), .Y(n4720) );
  INVX1 U6757 ( .A(n4720), .Y(n8369) );
  AND2X1 U6758 ( .A(n4168), .B(n4701), .Y(n4732) );
  INVX1 U6759 ( .A(n4732), .Y(n8370) );
  AND2X1 U6760 ( .A(n4108), .B(n4743), .Y(n4744) );
  INVX1 U6761 ( .A(n4744), .Y(n8371) );
  AND2X1 U6762 ( .A(n4146), .B(n4743), .Y(n4763) );
  INVX1 U6763 ( .A(n4763), .Y(n8372) );
  AND2X1 U6764 ( .A(n4170), .B(n4743), .Y(n4775) );
  INVX1 U6765 ( .A(n4775), .Y(n8373) );
  AND2X1 U6766 ( .A(n4148), .B(n4785), .Y(n4806) );
  INVX1 U6767 ( .A(n4806), .Y(n8374) );
  AND2X1 U6768 ( .A(n4172), .B(n4785), .Y(n4818) );
  INVX1 U6769 ( .A(n4818), .Y(n8375) );
  AND2X1 U6770 ( .A(n4150), .B(n4827), .Y(n4849) );
  INVX1 U6771 ( .A(n4849), .Y(n8376) );
  AND2X1 U6772 ( .A(n4174), .B(n4827), .Y(n4861) );
  INVX1 U6773 ( .A(n4861), .Y(n8377) );
  AND2X1 U6774 ( .A(n4128), .B(n4870), .Y(n4881) );
  INVX1 U6775 ( .A(n4881), .Y(n8378) );
  AND2X1 U6776 ( .A(n4152), .B(n4870), .Y(n4893) );
  INVX1 U6777 ( .A(n4893), .Y(n8379) );
  AND2X1 U6778 ( .A(n4176), .B(n4870), .Y(n4905) );
  INVX1 U6779 ( .A(n4905), .Y(n8380) );
  AND2X1 U6780 ( .A(n4130), .B(n4912), .Y(n4924) );
  INVX1 U6781 ( .A(n4924), .Y(n8381) );
  AND2X1 U6782 ( .A(n4154), .B(n4912), .Y(n4936) );
  INVX1 U6783 ( .A(n4936), .Y(n8382) );
  AND2X1 U6784 ( .A(n4178), .B(n4912), .Y(n4948) );
  INVX1 U6785 ( .A(n4948), .Y(n8383) );
  AND2X1 U6786 ( .A(n4132), .B(n4954), .Y(n4967) );
  INVX1 U6787 ( .A(n4967), .Y(n8384) );
  AND2X1 U6788 ( .A(n4156), .B(n4954), .Y(n4979) );
  INVX1 U6789 ( .A(n4979), .Y(n8385) );
  AND2X1 U6790 ( .A(n4180), .B(n4954), .Y(n4991) );
  INVX1 U6791 ( .A(n4991), .Y(n8386) );
  AND2X1 U6792 ( .A(n4134), .B(n4996), .Y(n5010) );
  INVX1 U6793 ( .A(n5010), .Y(n8387) );
  AND2X1 U6794 ( .A(n4158), .B(n4996), .Y(n5022) );
  INVX1 U6795 ( .A(n5022), .Y(n8388) );
  AND2X1 U6796 ( .A(n4182), .B(n4996), .Y(n5034) );
  INVX1 U6797 ( .A(n5034), .Y(n8389) );
  AND2X1 U6798 ( .A(n4136), .B(n5038), .Y(n5053) );
  INVX1 U6799 ( .A(n5053), .Y(n8390) );
  AND2X1 U6800 ( .A(n4160), .B(n5038), .Y(n5065) );
  INVX1 U6801 ( .A(n5065), .Y(n8391) );
  AND2X1 U6802 ( .A(n4184), .B(n5038), .Y(n5077) );
  INVX1 U6803 ( .A(n5077), .Y(n8392) );
  AND2X1 U6804 ( .A(n4138), .B(n5080), .Y(n5096) );
  INVX1 U6805 ( .A(n5096), .Y(n8393) );
  AND2X1 U6806 ( .A(n4162), .B(n5080), .Y(n5108) );
  INVX1 U6807 ( .A(n5108), .Y(n8394) );
  AND2X1 U6808 ( .A(n4186), .B(n5080), .Y(n5120) );
  INVX1 U6809 ( .A(n5120), .Y(n8395) );
  AND2X1 U6810 ( .A(n4140), .B(n5122), .Y(n5139) );
  INVX1 U6811 ( .A(n5139), .Y(n8396) );
  AND2X1 U6812 ( .A(n4164), .B(n5122), .Y(n5151) );
  INVX1 U6813 ( .A(n5151), .Y(n8397) );
  AND2X1 U6814 ( .A(n4188), .B(n5122), .Y(n5163) );
  INVX1 U6815 ( .A(n5163), .Y(n8398) );
  AND2X1 U6816 ( .A(n4150), .B(n5164), .Y(n5186) );
  INVX1 U6817 ( .A(n5186), .Y(n8399) );
  AND2X1 U6818 ( .A(n4174), .B(n5164), .Y(n5198) );
  INVX1 U6819 ( .A(n5198), .Y(n8400) );
  AND2X1 U6820 ( .A(n4128), .B(n5207), .Y(n5218) );
  INVX1 U6821 ( .A(n5218), .Y(n8401) );
  AND2X1 U6822 ( .A(n4152), .B(n5207), .Y(n5230) );
  INVX1 U6823 ( .A(n5230), .Y(n8402) );
  AND2X1 U6824 ( .A(n4176), .B(n5207), .Y(n5242) );
  INVX1 U6825 ( .A(n5242), .Y(n8403) );
  AND2X1 U6826 ( .A(n4130), .B(n5249), .Y(n5261) );
  INVX1 U6827 ( .A(n5261), .Y(n8404) );
  AND2X1 U6828 ( .A(n4154), .B(n5249), .Y(n5273) );
  INVX1 U6829 ( .A(n5273), .Y(n8405) );
  AND2X1 U6830 ( .A(n4178), .B(n5249), .Y(n5285) );
  INVX1 U6831 ( .A(n5285), .Y(n8406) );
  AND2X1 U6832 ( .A(n4132), .B(n5291), .Y(n5304) );
  INVX1 U6833 ( .A(n5304), .Y(n8407) );
  AND2X1 U6834 ( .A(n4156), .B(n5291), .Y(n5316) );
  INVX1 U6835 ( .A(n5316), .Y(n8408) );
  AND2X1 U6836 ( .A(n4180), .B(n5291), .Y(n5328) );
  INVX1 U6837 ( .A(n5328), .Y(n8409) );
  AND2X1 U6838 ( .A(n4134), .B(n5333), .Y(n5347) );
  INVX1 U6839 ( .A(n5347), .Y(n8410) );
  AND2X1 U6840 ( .A(n4158), .B(n5333), .Y(n5359) );
  INVX1 U6841 ( .A(n5359), .Y(n8411) );
  AND2X1 U6842 ( .A(n4182), .B(n5333), .Y(n5371) );
  INVX1 U6843 ( .A(n5371), .Y(n8412) );
  AND2X1 U6844 ( .A(n4136), .B(n5375), .Y(n5390) );
  INVX1 U6845 ( .A(n5390), .Y(n8413) );
  AND2X1 U6846 ( .A(n4160), .B(n5375), .Y(n5402) );
  INVX1 U6847 ( .A(n5402), .Y(n8414) );
  AND2X1 U6848 ( .A(n4184), .B(n5375), .Y(n5414) );
  INVX1 U6849 ( .A(n5414), .Y(n8415) );
  AND2X1 U6850 ( .A(n4138), .B(n5417), .Y(n5433) );
  INVX1 U6851 ( .A(n5433), .Y(n8416) );
  AND2X1 U6852 ( .A(n4162), .B(n5417), .Y(n5445) );
  INVX1 U6853 ( .A(n5445), .Y(n8417) );
  AND2X1 U6854 ( .A(n4186), .B(n5417), .Y(n5457) );
  INVX1 U6855 ( .A(n5457), .Y(n8418) );
  AND2X1 U6856 ( .A(n4140), .B(n5459), .Y(n5476) );
  INVX1 U6857 ( .A(n5476), .Y(n8419) );
  AND2X1 U6858 ( .A(n4164), .B(n5459), .Y(n5488) );
  INVX1 U6859 ( .A(n5488), .Y(n8420) );
  AND2X1 U6860 ( .A(n4188), .B(n5459), .Y(n5500) );
  INVX1 U6861 ( .A(n5500), .Y(n8421) );
  AND2X1 U6862 ( .A(n4054), .B(n8514), .Y(n4046) );
  INVX1 U6863 ( .A(n4046), .Y(n8422) );
  AND2X1 U6864 ( .A(n12), .B(n8506), .Y(n5505) );
  INVX1 U6865 ( .A(n5505), .Y(n8423) );
  INVX1 U6866 ( .A(n4076), .Y(n8424) );
  BUFX2 U6867 ( .A(n4189), .Y(n8425) );
  BUFX2 U6868 ( .A(n5206), .Y(n8426) );
  INVX1 U6869 ( .A(n8453), .Y(n8446) );
  INVX1 U6870 ( .A(n8453), .Y(n8445) );
  INVX1 U6871 ( .A(n8453), .Y(n8447) );
  INVX1 U6872 ( .A(n8331), .Y(n8428) );
  INVX1 U6873 ( .A(n8331), .Y(n8427) );
  INVX1 U6874 ( .A(n8453), .Y(n8448) );
  INVX1 U6875 ( .A(n8453), .Y(n8452) );
  INVX1 U6876 ( .A(n8453), .Y(n8451) );
  INVX1 U6877 ( .A(n8453), .Y(n8450) );
  INVX1 U6878 ( .A(n8453), .Y(n8449) );
  INVX1 U6879 ( .A(n8444), .Y(n8438) );
  INVX1 U6880 ( .A(n8444), .Y(n8436) );
  INVX1 U6881 ( .A(n8444), .Y(n8435) );
  INVX1 U6882 ( .A(n8444), .Y(n8437) );
  INVX1 U6883 ( .A(n8444), .Y(n8439) );
  INVX1 U6884 ( .A(n8444), .Y(n8443) );
  INVX1 U6885 ( .A(n8444), .Y(n8442) );
  INVX1 U6886 ( .A(n8444), .Y(n8441) );
  INVX1 U6887 ( .A(n8444), .Y(n8440) );
  INVX1 U6888 ( .A(n8463), .Y(n8457) );
  INVX1 U6889 ( .A(n8463), .Y(n8455) );
  INVX1 U6890 ( .A(n8463), .Y(n8454) );
  INVX1 U6891 ( .A(n8463), .Y(n8456) );
  INVX1 U6892 ( .A(n8463), .Y(n8458) );
  INVX1 U6893 ( .A(n8463), .Y(n8462) );
  INVX1 U6894 ( .A(n8463), .Y(n8461) );
  INVX1 U6895 ( .A(n8463), .Y(n8460) );
  INVX1 U6896 ( .A(n8463), .Y(n8459) );
  INVX1 U6897 ( .A(n8482), .Y(n8489) );
  INVX1 U6898 ( .A(n8482), .Y(n8490) );
  INVX1 U6899 ( .A(n8482), .Y(n8491) );
  INVX1 U6900 ( .A(n8482), .Y(n8488) );
  INVX1 U6901 ( .A(n8499), .Y(n8493) );
  INVX1 U6902 ( .A(n8499), .Y(n8492) );
  INVX1 U6903 ( .A(n8481), .Y(n8475) );
  INVX1 U6904 ( .A(n8481), .Y(n8474) );
  INVX1 U6905 ( .A(n8481), .Y(n8476) );
  INVX1 U6906 ( .A(n8482), .Y(n8485) );
  INVX1 U6907 ( .A(n8482), .Y(n8486) );
  INVX1 U6908 ( .A(n8482), .Y(n8487) );
  INVX1 U6909 ( .A(n8499), .Y(n8497) );
  INVX1 U6910 ( .A(n8499), .Y(n8496) );
  INVX1 U6911 ( .A(n8499), .Y(n8495) );
  INVX1 U6912 ( .A(n8499), .Y(n8494) );
  INVX1 U6913 ( .A(n8481), .Y(n8477) );
  INVX1 U6914 ( .A(n8499), .Y(n8498) );
  INVX1 U6915 ( .A(n8481), .Y(n8480) );
  INVX1 U6916 ( .A(n8481), .Y(n8479) );
  INVX1 U6917 ( .A(n8481), .Y(n8478) );
  INVX1 U6918 ( .A(n8473), .Y(n8467) );
  INVX1 U6919 ( .A(n8473), .Y(n8465) );
  INVX1 U6920 ( .A(n8473), .Y(n8464) );
  INVX1 U6921 ( .A(n8473), .Y(n8466) );
  INVX1 U6922 ( .A(n8482), .Y(n8483) );
  INVX1 U6923 ( .A(n8482), .Y(n8484) );
  INVX1 U6924 ( .A(n8473), .Y(n8468) );
  INVX1 U6925 ( .A(n8473), .Y(n8472) );
  INVX1 U6926 ( .A(n8473), .Y(n8471) );
  INVX1 U6927 ( .A(n8473), .Y(n8470) );
  INVX1 U6928 ( .A(n8473), .Y(n8469) );
  INVX1 U6929 ( .A(n8331), .Y(n8429) );
  INVX1 U6930 ( .A(n8331), .Y(n8430) );
  INVX1 U6931 ( .A(n8502), .Y(n8500) );
  INVX1 U6932 ( .A(n8502), .Y(n8501) );
  INVX1 U6933 ( .A(reset), .Y(n8502) );
  INVX1 U6934 ( .A(n8432), .Y(n8431) );
  INVX1 U6935 ( .A(n1354), .Y(n8499) );
  INVX1 U6936 ( .A(n1359), .Y(n8481) );
  INVX1 U6937 ( .A(n4098), .Y(n8508) );
  INVX1 U6938 ( .A(n8153), .Y(n8509) );
  INVX1 U6939 ( .A(n1362), .Y(n8453) );
  AND2X1 U6940 ( .A(n4074), .B(n8511), .Y(n1362) );
  INVX1 U6941 ( .A(n1363), .Y(n8444) );
  AND2X1 U6942 ( .A(n4075), .B(n8511), .Y(n1363) );
  INVX1 U6943 ( .A(n1361), .Y(n8463) );
  AND2X1 U6944 ( .A(n4073), .B(n8511), .Y(n1361) );
  AND2X1 U6945 ( .A(n8512), .B(n8513), .Y(n4074) );
  INVX1 U6946 ( .A(n8434), .Y(n8433) );
  INVX1 U6947 ( .A(n1374), .Y(n8434) );
  INVX1 U6948 ( .A(n1382), .Y(n8432) );
  INVX1 U6949 ( .A(n7881), .Y(n8505) );
  INVX1 U6950 ( .A(n7115), .Y(n8503) );
  AND2X1 U6951 ( .A(n4054), .B(n15), .Y(n1366) );
  AND2X1 U6952 ( .A(n4062), .B(n16), .Y(n4054) );
  INVX1 U6953 ( .A(put), .Y(n9831) );
  INVX1 U6954 ( .A(wr_ptr[0]), .Y(n8506) );
  INVX1 U6955 ( .A(wr_ptr[3]), .Y(n8518) );
  INVX1 U6956 ( .A(n4100), .Y(n8507) );
  INVX1 U6957 ( .A(wr_ptr[2]), .Y(n8517) );
  INVX1 U6958 ( .A(n1355), .Y(n8482) );
  INVX1 U6959 ( .A(n13), .Y(n8512) );
  INVX1 U6960 ( .A(wr_ptr[4]), .Y(n8515) );
  INVX1 U6961 ( .A(n12), .Y(n8511) );
  INVX1 U6962 ( .A(n15), .Y(n8514) );
  INVX1 U6963 ( .A(n14), .Y(n8513) );
  AND2X1 U6964 ( .A(n4075), .B(n12), .Y(n1354) );
  INVX1 U6965 ( .A(wr_ptr[1]), .Y(n8516) );
  AND2X1 U6966 ( .A(n14), .B(n8512), .Y(n4073) );
  AND2X1 U6967 ( .A(n4074), .B(n12), .Y(n1359) );
  INVX1 U6968 ( .A(n1360), .Y(n8473) );
  AND2X1 U6969 ( .A(n4073), .B(n12), .Y(n1360) );
  AND2X1 U6970 ( .A(n13), .B(n8513), .Y(n4075) );
  INVX1 U6971 ( .A(mem[902]), .Y(n8928) );
  INVX1 U6972 ( .A(mem[738]), .Y(n9092) );
  INVX1 U6973 ( .A(mem[861]), .Y(n8969) );
  INVX1 U6974 ( .A(mem[1230]), .Y(n8600) );
  INVX1 U6975 ( .A(mem[1066]), .Y(n8764) );
  INVX1 U6976 ( .A(mem[1189]), .Y(n8641) );
  INVX1 U6977 ( .A(mem[246]), .Y(n9584) );
  INVX1 U6978 ( .A(mem[82]), .Y(n9748) );
  INVX1 U6979 ( .A(mem[205]), .Y(n9625) );
  INVX1 U6980 ( .A(mem[903]), .Y(n8927) );
  INVX1 U6981 ( .A(mem[739]), .Y(n9091) );
  INVX1 U6982 ( .A(mem[862]), .Y(n8968) );
  INVX1 U6983 ( .A(mem[1231]), .Y(n8599) );
  INVX1 U6984 ( .A(mem[1067]), .Y(n8763) );
  INVX1 U6985 ( .A(mem[1190]), .Y(n8640) );
  INVX1 U6986 ( .A(mem[247]), .Y(n9583) );
  INVX1 U6987 ( .A(mem[83]), .Y(n9747) );
  INVX1 U6988 ( .A(mem[206]), .Y(n9624) );
  INVX1 U6989 ( .A(mem[904]), .Y(n8926) );
  INVX1 U6990 ( .A(mem[740]), .Y(n9090) );
  INVX1 U6991 ( .A(mem[863]), .Y(n8967) );
  INVX1 U6992 ( .A(mem[1232]), .Y(n8598) );
  INVX1 U6993 ( .A(mem[1068]), .Y(n8762) );
  INVX1 U6994 ( .A(mem[1191]), .Y(n8639) );
  INVX1 U6995 ( .A(mem[248]), .Y(n9582) );
  INVX1 U6996 ( .A(mem[84]), .Y(n9746) );
  INVX1 U6997 ( .A(mem[207]), .Y(n9623) );
  INVX1 U6998 ( .A(mem[905]), .Y(n8925) );
  INVX1 U6999 ( .A(mem[741]), .Y(n9089) );
  INVX1 U7000 ( .A(mem[864]), .Y(n8966) );
  INVX1 U7001 ( .A(mem[1233]), .Y(n8597) );
  INVX1 U7002 ( .A(mem[1069]), .Y(n8761) );
  INVX1 U7003 ( .A(mem[1192]), .Y(n8638) );
  INVX1 U7004 ( .A(mem[249]), .Y(n9581) );
  INVX1 U7005 ( .A(mem[85]), .Y(n9745) );
  INVX1 U7006 ( .A(mem[208]), .Y(n9622) );
  INVX1 U7007 ( .A(mem[906]), .Y(n8924) );
  INVX1 U7008 ( .A(mem[742]), .Y(n9088) );
  INVX1 U7009 ( .A(mem[865]), .Y(n8965) );
  INVX1 U7010 ( .A(mem[1234]), .Y(n8596) );
  INVX1 U7011 ( .A(mem[1070]), .Y(n8760) );
  INVX1 U7012 ( .A(mem[1193]), .Y(n8637) );
  INVX1 U7013 ( .A(mem[250]), .Y(n9580) );
  INVX1 U7014 ( .A(mem[86]), .Y(n9744) );
  INVX1 U7015 ( .A(mem[209]), .Y(n9621) );
  INVX1 U7016 ( .A(mem[907]), .Y(n8923) );
  INVX1 U7017 ( .A(mem[743]), .Y(n9087) );
  INVX1 U7018 ( .A(mem[866]), .Y(n8964) );
  INVX1 U7019 ( .A(mem[1235]), .Y(n8595) );
  INVX1 U7020 ( .A(mem[1071]), .Y(n8759) );
  INVX1 U7021 ( .A(mem[1194]), .Y(n8636) );
  INVX1 U7022 ( .A(mem[251]), .Y(n9579) );
  INVX1 U7023 ( .A(mem[87]), .Y(n9743) );
  INVX1 U7024 ( .A(mem[210]), .Y(n9620) );
  INVX1 U7025 ( .A(mem[908]), .Y(n8922) );
  INVX1 U7026 ( .A(mem[744]), .Y(n9086) );
  INVX1 U7027 ( .A(mem[867]), .Y(n8963) );
  INVX1 U7028 ( .A(mem[1236]), .Y(n8594) );
  INVX1 U7029 ( .A(mem[1072]), .Y(n8758) );
  INVX1 U7030 ( .A(mem[1195]), .Y(n8635) );
  INVX1 U7031 ( .A(mem[252]), .Y(n9578) );
  INVX1 U7032 ( .A(mem[88]), .Y(n9742) );
  INVX1 U7033 ( .A(mem[211]), .Y(n9619) );
  INVX1 U7034 ( .A(mem[909]), .Y(n8921) );
  INVX1 U7035 ( .A(mem[745]), .Y(n9085) );
  INVX1 U7036 ( .A(mem[868]), .Y(n8962) );
  INVX1 U7037 ( .A(mem[1237]), .Y(n8593) );
  INVX1 U7038 ( .A(mem[1073]), .Y(n8757) );
  INVX1 U7039 ( .A(mem[1196]), .Y(n8634) );
  INVX1 U7040 ( .A(mem[253]), .Y(n9577) );
  INVX1 U7041 ( .A(mem[89]), .Y(n9741) );
  INVX1 U7042 ( .A(mem[212]), .Y(n9618) );
  INVX1 U7043 ( .A(mem[910]), .Y(n8920) );
  INVX1 U7044 ( .A(mem[746]), .Y(n9084) );
  INVX1 U7045 ( .A(mem[869]), .Y(n8961) );
  INVX1 U7046 ( .A(mem[1238]), .Y(n8592) );
  INVX1 U7047 ( .A(mem[1074]), .Y(n8756) );
  INVX1 U7048 ( .A(mem[1197]), .Y(n8633) );
  INVX1 U7049 ( .A(mem[254]), .Y(n9576) );
  INVX1 U7050 ( .A(mem[90]), .Y(n9740) );
  INVX1 U7051 ( .A(mem[213]), .Y(n9617) );
  INVX1 U7052 ( .A(mem[911]), .Y(n8919) );
  INVX1 U7053 ( .A(mem[747]), .Y(n9083) );
  INVX1 U7054 ( .A(mem[870]), .Y(n8960) );
  INVX1 U7055 ( .A(mem[1239]), .Y(n8591) );
  INVX1 U7056 ( .A(mem[1075]), .Y(n8755) );
  INVX1 U7057 ( .A(mem[1198]), .Y(n8632) );
  INVX1 U7058 ( .A(mem[255]), .Y(n9575) );
  INVX1 U7059 ( .A(mem[91]), .Y(n9739) );
  INVX1 U7060 ( .A(mem[214]), .Y(n9616) );
  INVX1 U7061 ( .A(mem[912]), .Y(n8918) );
  INVX1 U7062 ( .A(mem[748]), .Y(n9082) );
  INVX1 U7063 ( .A(mem[871]), .Y(n8959) );
  INVX1 U7064 ( .A(mem[1240]), .Y(n8590) );
  INVX1 U7065 ( .A(mem[1076]), .Y(n8754) );
  INVX1 U7066 ( .A(mem[1199]), .Y(n8631) );
  INVX1 U7067 ( .A(mem[256]), .Y(n9574) );
  INVX1 U7068 ( .A(mem[92]), .Y(n9738) );
  INVX1 U7069 ( .A(mem[215]), .Y(n9615) );
  INVX1 U7070 ( .A(mem[913]), .Y(n8917) );
  INVX1 U7071 ( .A(mem[749]), .Y(n9081) );
  INVX1 U7072 ( .A(mem[872]), .Y(n8958) );
  INVX1 U7073 ( .A(mem[1241]), .Y(n8589) );
  INVX1 U7074 ( .A(mem[1077]), .Y(n8753) );
  INVX1 U7075 ( .A(mem[1200]), .Y(n8630) );
  INVX1 U7076 ( .A(mem[257]), .Y(n9573) );
  INVX1 U7077 ( .A(mem[93]), .Y(n9737) );
  INVX1 U7078 ( .A(mem[216]), .Y(n9614) );
  INVX1 U7079 ( .A(mem[914]), .Y(n8916) );
  INVX1 U7080 ( .A(mem[750]), .Y(n9080) );
  INVX1 U7081 ( .A(mem[873]), .Y(n8957) );
  INVX1 U7082 ( .A(mem[1242]), .Y(n8588) );
  INVX1 U7083 ( .A(mem[1078]), .Y(n8752) );
  INVX1 U7084 ( .A(mem[1201]), .Y(n8629) );
  INVX1 U7085 ( .A(mem[258]), .Y(n9572) );
  INVX1 U7086 ( .A(mem[94]), .Y(n9736) );
  INVX1 U7087 ( .A(mem[217]), .Y(n9613) );
  INVX1 U7088 ( .A(mem[915]), .Y(n8915) );
  INVX1 U7089 ( .A(mem[751]), .Y(n9079) );
  INVX1 U7090 ( .A(mem[874]), .Y(n8956) );
  INVX1 U7091 ( .A(mem[1243]), .Y(n8587) );
  INVX1 U7092 ( .A(mem[1079]), .Y(n8751) );
  INVX1 U7093 ( .A(mem[1202]), .Y(n8628) );
  INVX1 U7094 ( .A(mem[259]), .Y(n9571) );
  INVX1 U7095 ( .A(mem[95]), .Y(n9735) );
  INVX1 U7096 ( .A(mem[218]), .Y(n9612) );
  INVX1 U7097 ( .A(mem[916]), .Y(n8914) );
  INVX1 U7098 ( .A(mem[752]), .Y(n9078) );
  INVX1 U7099 ( .A(mem[875]), .Y(n8955) );
  INVX1 U7100 ( .A(mem[1244]), .Y(n8586) );
  INVX1 U7101 ( .A(mem[1080]), .Y(n8750) );
  INVX1 U7102 ( .A(mem[1203]), .Y(n8627) );
  INVX1 U7103 ( .A(mem[260]), .Y(n9570) );
  INVX1 U7104 ( .A(mem[96]), .Y(n9734) );
  INVX1 U7105 ( .A(mem[219]), .Y(n9611) );
  INVX1 U7106 ( .A(mem[917]), .Y(n8913) );
  INVX1 U7107 ( .A(mem[753]), .Y(n9077) );
  INVX1 U7108 ( .A(mem[876]), .Y(n8954) );
  INVX1 U7109 ( .A(mem[1245]), .Y(n8585) );
  INVX1 U7110 ( .A(mem[1081]), .Y(n8749) );
  INVX1 U7111 ( .A(mem[1204]), .Y(n8626) );
  INVX1 U7112 ( .A(mem[261]), .Y(n9569) );
  INVX1 U7113 ( .A(mem[97]), .Y(n9733) );
  INVX1 U7114 ( .A(mem[220]), .Y(n9610) );
  INVX1 U7115 ( .A(mem[918]), .Y(n8912) );
  INVX1 U7116 ( .A(mem[754]), .Y(n9076) );
  INVX1 U7117 ( .A(mem[877]), .Y(n8953) );
  INVX1 U7118 ( .A(mem[1246]), .Y(n8584) );
  INVX1 U7119 ( .A(mem[1082]), .Y(n8748) );
  INVX1 U7120 ( .A(mem[1205]), .Y(n8625) );
  INVX1 U7121 ( .A(mem[262]), .Y(n9568) );
  INVX1 U7122 ( .A(mem[98]), .Y(n9732) );
  INVX1 U7123 ( .A(mem[221]), .Y(n9609) );
  INVX1 U7124 ( .A(mem[919]), .Y(n8911) );
  INVX1 U7125 ( .A(mem[755]), .Y(n9075) );
  INVX1 U7126 ( .A(mem[878]), .Y(n8952) );
  INVX1 U7127 ( .A(mem[1247]), .Y(n8583) );
  INVX1 U7128 ( .A(mem[1083]), .Y(n8747) );
  INVX1 U7129 ( .A(mem[1206]), .Y(n8624) );
  INVX1 U7130 ( .A(mem[263]), .Y(n9567) );
  INVX1 U7131 ( .A(mem[99]), .Y(n9731) );
  INVX1 U7132 ( .A(mem[222]), .Y(n9608) );
  INVX1 U7133 ( .A(mem[920]), .Y(n8910) );
  INVX1 U7134 ( .A(mem[756]), .Y(n9074) );
  INVX1 U7135 ( .A(mem[879]), .Y(n8951) );
  INVX1 U7136 ( .A(mem[1248]), .Y(n8582) );
  INVX1 U7137 ( .A(mem[1084]), .Y(n8746) );
  INVX1 U7138 ( .A(mem[1207]), .Y(n8623) );
  INVX1 U7139 ( .A(mem[264]), .Y(n9566) );
  INVX1 U7140 ( .A(mem[100]), .Y(n9730) );
  INVX1 U7141 ( .A(mem[223]), .Y(n9607) );
  INVX1 U7142 ( .A(mem[921]), .Y(n8909) );
  INVX1 U7143 ( .A(mem[757]), .Y(n9073) );
  INVX1 U7144 ( .A(mem[880]), .Y(n8950) );
  INVX1 U7145 ( .A(mem[1249]), .Y(n8581) );
  INVX1 U7146 ( .A(mem[1085]), .Y(n8745) );
  INVX1 U7147 ( .A(mem[1208]), .Y(n8622) );
  INVX1 U7148 ( .A(mem[265]), .Y(n9565) );
  INVX1 U7149 ( .A(mem[101]), .Y(n9729) );
  INVX1 U7150 ( .A(mem[224]), .Y(n9606) );
  INVX1 U7151 ( .A(mem[922]), .Y(n8908) );
  INVX1 U7152 ( .A(mem[758]), .Y(n9072) );
  INVX1 U7153 ( .A(mem[881]), .Y(n8949) );
  INVX1 U7154 ( .A(mem[1250]), .Y(n8580) );
  INVX1 U7155 ( .A(mem[1086]), .Y(n8744) );
  INVX1 U7156 ( .A(mem[1209]), .Y(n8621) );
  INVX1 U7157 ( .A(mem[266]), .Y(n9564) );
  INVX1 U7158 ( .A(mem[102]), .Y(n9728) );
  INVX1 U7159 ( .A(mem[225]), .Y(n9605) );
  INVX1 U7160 ( .A(mem[923]), .Y(n8907) );
  INVX1 U7161 ( .A(mem[759]), .Y(n9071) );
  INVX1 U7162 ( .A(mem[882]), .Y(n8948) );
  INVX1 U7163 ( .A(mem[1251]), .Y(n8579) );
  INVX1 U7164 ( .A(mem[1087]), .Y(n8743) );
  INVX1 U7165 ( .A(mem[1210]), .Y(n8620) );
  INVX1 U7166 ( .A(mem[267]), .Y(n9563) );
  INVX1 U7167 ( .A(mem[103]), .Y(n9727) );
  INVX1 U7168 ( .A(mem[226]), .Y(n9604) );
  INVX1 U7169 ( .A(mem[924]), .Y(n8906) );
  INVX1 U7170 ( .A(mem[760]), .Y(n9070) );
  INVX1 U7171 ( .A(mem[883]), .Y(n8947) );
  INVX1 U7172 ( .A(mem[1252]), .Y(n8578) );
  INVX1 U7173 ( .A(mem[1088]), .Y(n8742) );
  INVX1 U7174 ( .A(mem[1211]), .Y(n8619) );
  INVX1 U7175 ( .A(mem[268]), .Y(n9562) );
  INVX1 U7176 ( .A(mem[104]), .Y(n9726) );
  INVX1 U7177 ( .A(mem[227]), .Y(n9603) );
  INVX1 U7178 ( .A(mem[925]), .Y(n8905) );
  INVX1 U7179 ( .A(mem[761]), .Y(n9069) );
  INVX1 U7180 ( .A(mem[884]), .Y(n8946) );
  INVX1 U7181 ( .A(mem[1253]), .Y(n8577) );
  INVX1 U7182 ( .A(mem[1089]), .Y(n8741) );
  INVX1 U7183 ( .A(mem[1212]), .Y(n8618) );
  INVX1 U7184 ( .A(mem[269]), .Y(n9561) );
  INVX1 U7185 ( .A(mem[105]), .Y(n9725) );
  INVX1 U7186 ( .A(mem[228]), .Y(n9602) );
  INVX1 U7187 ( .A(mem[926]), .Y(n8904) );
  INVX1 U7188 ( .A(mem[762]), .Y(n9068) );
  INVX1 U7189 ( .A(mem[885]), .Y(n8945) );
  INVX1 U7190 ( .A(mem[1254]), .Y(n8576) );
  INVX1 U7191 ( .A(mem[1090]), .Y(n8740) );
  INVX1 U7192 ( .A(mem[1213]), .Y(n8617) );
  INVX1 U7193 ( .A(mem[270]), .Y(n9560) );
  INVX1 U7194 ( .A(mem[106]), .Y(n9724) );
  INVX1 U7195 ( .A(mem[229]), .Y(n9601) );
  INVX1 U7196 ( .A(mem[927]), .Y(n8903) );
  INVX1 U7197 ( .A(mem[763]), .Y(n9067) );
  INVX1 U7198 ( .A(mem[886]), .Y(n8944) );
  INVX1 U7199 ( .A(mem[1255]), .Y(n8575) );
  INVX1 U7200 ( .A(mem[1091]), .Y(n8739) );
  INVX1 U7201 ( .A(mem[1214]), .Y(n8616) );
  INVX1 U7202 ( .A(mem[271]), .Y(n9559) );
  INVX1 U7203 ( .A(mem[107]), .Y(n9723) );
  INVX1 U7204 ( .A(mem[230]), .Y(n9600) );
  INVX1 U7205 ( .A(mem[928]), .Y(n8902) );
  INVX1 U7206 ( .A(mem[764]), .Y(n9066) );
  INVX1 U7207 ( .A(mem[887]), .Y(n8943) );
  INVX1 U7208 ( .A(mem[1256]), .Y(n8574) );
  INVX1 U7209 ( .A(mem[1092]), .Y(n8738) );
  INVX1 U7210 ( .A(mem[1215]), .Y(n8615) );
  INVX1 U7211 ( .A(mem[272]), .Y(n9558) );
  INVX1 U7212 ( .A(mem[108]), .Y(n9722) );
  INVX1 U7213 ( .A(mem[231]), .Y(n9599) );
  INVX1 U7214 ( .A(mem[929]), .Y(n8901) );
  INVX1 U7215 ( .A(mem[765]), .Y(n9065) );
  INVX1 U7216 ( .A(mem[888]), .Y(n8942) );
  INVX1 U7217 ( .A(mem[1257]), .Y(n8573) );
  INVX1 U7218 ( .A(mem[1093]), .Y(n8737) );
  INVX1 U7219 ( .A(mem[1216]), .Y(n8614) );
  INVX1 U7220 ( .A(mem[273]), .Y(n9557) );
  INVX1 U7221 ( .A(mem[109]), .Y(n9721) );
  INVX1 U7222 ( .A(mem[232]), .Y(n9598) );
  INVX1 U7223 ( .A(mem[930]), .Y(n8900) );
  INVX1 U7224 ( .A(mem[766]), .Y(n9064) );
  INVX1 U7225 ( .A(mem[889]), .Y(n8941) );
  INVX1 U7226 ( .A(mem[1258]), .Y(n8572) );
  INVX1 U7227 ( .A(mem[1094]), .Y(n8736) );
  INVX1 U7228 ( .A(mem[1217]), .Y(n8613) );
  INVX1 U7229 ( .A(mem[274]), .Y(n9556) );
  INVX1 U7230 ( .A(mem[110]), .Y(n9720) );
  INVX1 U7231 ( .A(mem[233]), .Y(n9597) );
  INVX1 U7232 ( .A(mem[931]), .Y(n8899) );
  INVX1 U7233 ( .A(mem[767]), .Y(n9063) );
  INVX1 U7234 ( .A(mem[890]), .Y(n8940) );
  INVX1 U7235 ( .A(mem[1259]), .Y(n8571) );
  INVX1 U7236 ( .A(mem[1095]), .Y(n8735) );
  INVX1 U7237 ( .A(mem[1218]), .Y(n8612) );
  INVX1 U7238 ( .A(mem[275]), .Y(n9555) );
  INVX1 U7239 ( .A(mem[111]), .Y(n9719) );
  INVX1 U7240 ( .A(mem[234]), .Y(n9596) );
  INVX1 U7241 ( .A(mem[932]), .Y(n8898) );
  INVX1 U7242 ( .A(mem[768]), .Y(n9062) );
  INVX1 U7243 ( .A(mem[891]), .Y(n8939) );
  INVX1 U7244 ( .A(mem[1260]), .Y(n8570) );
  INVX1 U7245 ( .A(mem[1096]), .Y(n8734) );
  INVX1 U7246 ( .A(mem[1219]), .Y(n8611) );
  INVX1 U7247 ( .A(mem[276]), .Y(n9554) );
  INVX1 U7248 ( .A(mem[112]), .Y(n9718) );
  INVX1 U7249 ( .A(mem[235]), .Y(n9595) );
  INVX1 U7250 ( .A(mem[933]), .Y(n8897) );
  INVX1 U7251 ( .A(mem[769]), .Y(n9061) );
  INVX1 U7252 ( .A(mem[892]), .Y(n8938) );
  INVX1 U7253 ( .A(mem[1261]), .Y(n8569) );
  INVX1 U7254 ( .A(mem[1097]), .Y(n8733) );
  INVX1 U7255 ( .A(mem[1220]), .Y(n8610) );
  INVX1 U7256 ( .A(mem[277]), .Y(n9553) );
  INVX1 U7257 ( .A(mem[113]), .Y(n9717) );
  INVX1 U7258 ( .A(mem[236]), .Y(n9594) );
  INVX1 U7259 ( .A(mem[934]), .Y(n8896) );
  INVX1 U7260 ( .A(mem[770]), .Y(n9060) );
  INVX1 U7261 ( .A(mem[893]), .Y(n8937) );
  INVX1 U7262 ( .A(mem[1262]), .Y(n8568) );
  INVX1 U7263 ( .A(mem[1098]), .Y(n8732) );
  INVX1 U7264 ( .A(mem[1221]), .Y(n8609) );
  INVX1 U7265 ( .A(mem[278]), .Y(n9552) );
  INVX1 U7266 ( .A(mem[114]), .Y(n9716) );
  INVX1 U7267 ( .A(mem[237]), .Y(n9593) );
  INVX1 U7268 ( .A(mem[935]), .Y(n8895) );
  INVX1 U7269 ( .A(mem[771]), .Y(n9059) );
  INVX1 U7270 ( .A(mem[894]), .Y(n8936) );
  INVX1 U7271 ( .A(mem[1263]), .Y(n8567) );
  INVX1 U7272 ( .A(mem[1099]), .Y(n8731) );
  INVX1 U7273 ( .A(mem[1222]), .Y(n8608) );
  INVX1 U7274 ( .A(mem[279]), .Y(n9551) );
  INVX1 U7275 ( .A(mem[115]), .Y(n9715) );
  INVX1 U7276 ( .A(mem[238]), .Y(n9592) );
  INVX1 U7277 ( .A(mem[936]), .Y(n8894) );
  INVX1 U7278 ( .A(mem[772]), .Y(n9058) );
  INVX1 U7279 ( .A(mem[895]), .Y(n8935) );
  INVX1 U7280 ( .A(mem[1264]), .Y(n8566) );
  INVX1 U7281 ( .A(mem[1100]), .Y(n8730) );
  INVX1 U7282 ( .A(mem[1223]), .Y(n8607) );
  INVX1 U7283 ( .A(mem[280]), .Y(n9550) );
  INVX1 U7284 ( .A(mem[116]), .Y(n9714) );
  INVX1 U7285 ( .A(mem[239]), .Y(n9591) );
  INVX1 U7286 ( .A(mem[937]), .Y(n8893) );
  INVX1 U7287 ( .A(mem[773]), .Y(n9057) );
  INVX1 U7288 ( .A(mem[896]), .Y(n8934) );
  INVX1 U7289 ( .A(mem[1265]), .Y(n8565) );
  INVX1 U7290 ( .A(mem[1101]), .Y(n8729) );
  INVX1 U7291 ( .A(mem[1224]), .Y(n8606) );
  INVX1 U7292 ( .A(mem[281]), .Y(n9549) );
  INVX1 U7293 ( .A(mem[117]), .Y(n9713) );
  INVX1 U7294 ( .A(mem[240]), .Y(n9590) );
  INVX1 U7295 ( .A(mem[938]), .Y(n8892) );
  INVX1 U7296 ( .A(mem[774]), .Y(n9056) );
  INVX1 U7297 ( .A(mem[897]), .Y(n8933) );
  INVX1 U7298 ( .A(mem[1266]), .Y(n8564) );
  INVX1 U7299 ( .A(mem[1102]), .Y(n8728) );
  INVX1 U7300 ( .A(mem[1225]), .Y(n8605) );
  INVX1 U7301 ( .A(mem[282]), .Y(n9548) );
  INVX1 U7302 ( .A(mem[118]), .Y(n9712) );
  INVX1 U7303 ( .A(mem[241]), .Y(n9589) );
  INVX1 U7304 ( .A(mem[939]), .Y(n8891) );
  INVX1 U7305 ( .A(mem[775]), .Y(n9055) );
  INVX1 U7306 ( .A(mem[898]), .Y(n8932) );
  INVX1 U7307 ( .A(mem[1267]), .Y(n8563) );
  INVX1 U7308 ( .A(mem[1103]), .Y(n8727) );
  INVX1 U7309 ( .A(mem[1226]), .Y(n8604) );
  INVX1 U7310 ( .A(mem[283]), .Y(n9547) );
  INVX1 U7311 ( .A(mem[119]), .Y(n9711) );
  INVX1 U7312 ( .A(mem[242]), .Y(n9588) );
  INVX1 U7313 ( .A(mem[940]), .Y(n8890) );
  INVX1 U7314 ( .A(mem[776]), .Y(n9054) );
  INVX1 U7315 ( .A(mem[899]), .Y(n8931) );
  INVX1 U7316 ( .A(mem[1268]), .Y(n8562) );
  INVX1 U7317 ( .A(mem[1104]), .Y(n8726) );
  INVX1 U7318 ( .A(mem[1227]), .Y(n8603) );
  INVX1 U7319 ( .A(mem[284]), .Y(n9546) );
  INVX1 U7320 ( .A(mem[120]), .Y(n9710) );
  INVX1 U7321 ( .A(mem[243]), .Y(n9587) );
  INVX1 U7322 ( .A(mem[941]), .Y(n8889) );
  INVX1 U7323 ( .A(mem[777]), .Y(n9053) );
  INVX1 U7324 ( .A(mem[900]), .Y(n8930) );
  INVX1 U7325 ( .A(mem[1269]), .Y(n8561) );
  INVX1 U7326 ( .A(mem[1105]), .Y(n8725) );
  INVX1 U7327 ( .A(mem[1228]), .Y(n8602) );
  INVX1 U7328 ( .A(mem[285]), .Y(n9545) );
  INVX1 U7329 ( .A(mem[121]), .Y(n9709) );
  INVX1 U7330 ( .A(mem[244]), .Y(n9586) );
  INVX1 U7331 ( .A(mem[942]), .Y(n8888) );
  INVX1 U7332 ( .A(mem[778]), .Y(n9052) );
  INVX1 U7333 ( .A(mem[901]), .Y(n8929) );
  INVX1 U7334 ( .A(mem[1270]), .Y(n8560) );
  INVX1 U7335 ( .A(mem[1106]), .Y(n8724) );
  INVX1 U7336 ( .A(mem[1229]), .Y(n8601) );
  INVX1 U7337 ( .A(mem[286]), .Y(n9544) );
  INVX1 U7338 ( .A(mem[122]), .Y(n9708) );
  INVX1 U7339 ( .A(mem[245]), .Y(n9585) );
  INVX1 U7340 ( .A(mem[574]), .Y(n9256) );
  INVX1 U7341 ( .A(mem[410]), .Y(n9420) );
  INVX1 U7342 ( .A(mem[533]), .Y(n9297) );
  INVX1 U7343 ( .A(mem[575]), .Y(n9255) );
  INVX1 U7344 ( .A(mem[411]), .Y(n9419) );
  INVX1 U7345 ( .A(mem[534]), .Y(n9296) );
  INVX1 U7346 ( .A(mem[576]), .Y(n9254) );
  INVX1 U7347 ( .A(mem[412]), .Y(n9418) );
  INVX1 U7348 ( .A(mem[535]), .Y(n9295) );
  INVX1 U7349 ( .A(mem[577]), .Y(n9253) );
  INVX1 U7350 ( .A(mem[413]), .Y(n9417) );
  INVX1 U7351 ( .A(mem[536]), .Y(n9294) );
  INVX1 U7352 ( .A(mem[578]), .Y(n9252) );
  INVX1 U7353 ( .A(mem[414]), .Y(n9416) );
  INVX1 U7354 ( .A(mem[537]), .Y(n9293) );
  INVX1 U7355 ( .A(mem[579]), .Y(n9251) );
  INVX1 U7356 ( .A(mem[415]), .Y(n9415) );
  INVX1 U7357 ( .A(mem[538]), .Y(n9292) );
  INVX1 U7358 ( .A(mem[580]), .Y(n9250) );
  INVX1 U7359 ( .A(mem[416]), .Y(n9414) );
  INVX1 U7360 ( .A(mem[539]), .Y(n9291) );
  INVX1 U7361 ( .A(mem[581]), .Y(n9249) );
  INVX1 U7362 ( .A(mem[417]), .Y(n9413) );
  INVX1 U7363 ( .A(mem[540]), .Y(n9290) );
  INVX1 U7364 ( .A(mem[582]), .Y(n9248) );
  INVX1 U7365 ( .A(mem[418]), .Y(n9412) );
  INVX1 U7366 ( .A(mem[541]), .Y(n9289) );
  INVX1 U7367 ( .A(mem[583]), .Y(n9247) );
  INVX1 U7368 ( .A(mem[419]), .Y(n9411) );
  INVX1 U7369 ( .A(mem[542]), .Y(n9288) );
  INVX1 U7370 ( .A(mem[584]), .Y(n9246) );
  INVX1 U7371 ( .A(mem[420]), .Y(n9410) );
  INVX1 U7372 ( .A(mem[543]), .Y(n9287) );
  INVX1 U7373 ( .A(mem[585]), .Y(n9245) );
  INVX1 U7374 ( .A(mem[421]), .Y(n9409) );
  INVX1 U7375 ( .A(mem[544]), .Y(n9286) );
  INVX1 U7376 ( .A(mem[586]), .Y(n9244) );
  INVX1 U7377 ( .A(mem[422]), .Y(n9408) );
  INVX1 U7378 ( .A(mem[545]), .Y(n9285) );
  INVX1 U7379 ( .A(mem[587]), .Y(n9243) );
  INVX1 U7380 ( .A(mem[423]), .Y(n9407) );
  INVX1 U7381 ( .A(mem[546]), .Y(n9284) );
  INVX1 U7382 ( .A(mem[588]), .Y(n9242) );
  INVX1 U7383 ( .A(mem[424]), .Y(n9406) );
  INVX1 U7384 ( .A(mem[547]), .Y(n9283) );
  INVX1 U7385 ( .A(mem[589]), .Y(n9241) );
  INVX1 U7386 ( .A(mem[425]), .Y(n9405) );
  INVX1 U7387 ( .A(mem[548]), .Y(n9282) );
  INVX1 U7388 ( .A(mem[590]), .Y(n9240) );
  INVX1 U7389 ( .A(mem[426]), .Y(n9404) );
  INVX1 U7390 ( .A(mem[549]), .Y(n9281) );
  INVX1 U7391 ( .A(mem[591]), .Y(n9239) );
  INVX1 U7392 ( .A(mem[427]), .Y(n9403) );
  INVX1 U7393 ( .A(mem[550]), .Y(n9280) );
  INVX1 U7394 ( .A(mem[592]), .Y(n9238) );
  INVX1 U7395 ( .A(mem[428]), .Y(n9402) );
  INVX1 U7396 ( .A(mem[551]), .Y(n9279) );
  INVX1 U7397 ( .A(mem[593]), .Y(n9237) );
  INVX1 U7398 ( .A(mem[429]), .Y(n9401) );
  INVX1 U7399 ( .A(mem[552]), .Y(n9278) );
  INVX1 U7400 ( .A(mem[594]), .Y(n9236) );
  INVX1 U7401 ( .A(mem[430]), .Y(n9400) );
  INVX1 U7402 ( .A(mem[553]), .Y(n9277) );
  INVX1 U7403 ( .A(mem[595]), .Y(n9235) );
  INVX1 U7404 ( .A(mem[431]), .Y(n9399) );
  INVX1 U7405 ( .A(mem[554]), .Y(n9276) );
  INVX1 U7406 ( .A(mem[596]), .Y(n9234) );
  INVX1 U7407 ( .A(mem[432]), .Y(n9398) );
  INVX1 U7408 ( .A(mem[555]), .Y(n9275) );
  INVX1 U7409 ( .A(mem[597]), .Y(n9233) );
  INVX1 U7410 ( .A(mem[433]), .Y(n9397) );
  INVX1 U7411 ( .A(mem[556]), .Y(n9274) );
  INVX1 U7412 ( .A(mem[598]), .Y(n9232) );
  INVX1 U7413 ( .A(mem[434]), .Y(n9396) );
  INVX1 U7414 ( .A(mem[557]), .Y(n9273) );
  INVX1 U7415 ( .A(mem[599]), .Y(n9231) );
  INVX1 U7416 ( .A(mem[435]), .Y(n9395) );
  INVX1 U7417 ( .A(mem[558]), .Y(n9272) );
  INVX1 U7418 ( .A(mem[600]), .Y(n9230) );
  INVX1 U7419 ( .A(mem[436]), .Y(n9394) );
  INVX1 U7420 ( .A(mem[559]), .Y(n9271) );
  INVX1 U7421 ( .A(mem[601]), .Y(n9229) );
  INVX1 U7422 ( .A(mem[437]), .Y(n9393) );
  INVX1 U7423 ( .A(mem[560]), .Y(n9270) );
  INVX1 U7424 ( .A(mem[602]), .Y(n9228) );
  INVX1 U7425 ( .A(mem[438]), .Y(n9392) );
  INVX1 U7426 ( .A(mem[561]), .Y(n9269) );
  INVX1 U7427 ( .A(mem[603]), .Y(n9227) );
  INVX1 U7428 ( .A(mem[439]), .Y(n9391) );
  INVX1 U7429 ( .A(mem[562]), .Y(n9268) );
  INVX1 U7430 ( .A(mem[604]), .Y(n9226) );
  INVX1 U7431 ( .A(mem[440]), .Y(n9390) );
  INVX1 U7432 ( .A(mem[563]), .Y(n9267) );
  INVX1 U7433 ( .A(mem[605]), .Y(n9225) );
  INVX1 U7434 ( .A(mem[441]), .Y(n9389) );
  INVX1 U7435 ( .A(mem[564]), .Y(n9266) );
  INVX1 U7436 ( .A(mem[606]), .Y(n9224) );
  INVX1 U7437 ( .A(mem[442]), .Y(n9388) );
  INVX1 U7438 ( .A(mem[565]), .Y(n9265) );
  INVX1 U7439 ( .A(mem[607]), .Y(n9223) );
  INVX1 U7440 ( .A(mem[443]), .Y(n9387) );
  INVX1 U7441 ( .A(mem[566]), .Y(n9264) );
  INVX1 U7442 ( .A(mem[608]), .Y(n9222) );
  INVX1 U7443 ( .A(mem[444]), .Y(n9386) );
  INVX1 U7444 ( .A(mem[567]), .Y(n9263) );
  INVX1 U7445 ( .A(mem[609]), .Y(n9221) );
  INVX1 U7446 ( .A(mem[445]), .Y(n9385) );
  INVX1 U7447 ( .A(mem[568]), .Y(n9262) );
  INVX1 U7448 ( .A(mem[610]), .Y(n9220) );
  INVX1 U7449 ( .A(mem[446]), .Y(n9384) );
  INVX1 U7450 ( .A(mem[569]), .Y(n9261) );
  INVX1 U7451 ( .A(mem[611]), .Y(n9219) );
  INVX1 U7452 ( .A(mem[447]), .Y(n9383) );
  INVX1 U7453 ( .A(mem[570]), .Y(n9260) );
  INVX1 U7454 ( .A(mem[612]), .Y(n9218) );
  INVX1 U7455 ( .A(mem[448]), .Y(n9382) );
  INVX1 U7456 ( .A(mem[571]), .Y(n9259) );
  INVX1 U7457 ( .A(mem[613]), .Y(n9217) );
  INVX1 U7458 ( .A(mem[449]), .Y(n9381) );
  INVX1 U7459 ( .A(mem[572]), .Y(n9258) );
  INVX1 U7460 ( .A(mem[614]), .Y(n9216) );
  INVX1 U7461 ( .A(mem[450]), .Y(n9380) );
  INVX1 U7462 ( .A(mem[573]), .Y(n9257) );
  INVX1 U7463 ( .A(mem[779]), .Y(n9051) );
  INVX1 U7464 ( .A(mem[656]), .Y(n9174) );
  INVX1 U7465 ( .A(mem[697]), .Y(n9133) );
  INVX1 U7466 ( .A(mem[1107]), .Y(n8723) );
  INVX1 U7467 ( .A(mem[984]), .Y(n8846) );
  INVX1 U7468 ( .A(mem[1025]), .Y(n8805) );
  INVX1 U7469 ( .A(mem[123]), .Y(n9707) );
  INVX1 U7470 ( .A(mem[0]), .Y(n9830) );
  INVX1 U7471 ( .A(mem[41]), .Y(n9789) );
  INVX1 U7472 ( .A(mem[780]), .Y(n9050) );
  INVX1 U7473 ( .A(mem[657]), .Y(n9173) );
  INVX1 U7474 ( .A(mem[698]), .Y(n9132) );
  INVX1 U7475 ( .A(mem[1108]), .Y(n8722) );
  INVX1 U7476 ( .A(mem[985]), .Y(n8845) );
  INVX1 U7477 ( .A(mem[1026]), .Y(n8804) );
  INVX1 U7478 ( .A(mem[124]), .Y(n9706) );
  INVX1 U7479 ( .A(mem[1]), .Y(n9829) );
  INVX1 U7480 ( .A(mem[42]), .Y(n9788) );
  INVX1 U7481 ( .A(mem[781]), .Y(n9049) );
  INVX1 U7482 ( .A(mem[658]), .Y(n9172) );
  INVX1 U7483 ( .A(mem[699]), .Y(n9131) );
  INVX1 U7484 ( .A(mem[1109]), .Y(n8721) );
  INVX1 U7485 ( .A(mem[986]), .Y(n8844) );
  INVX1 U7486 ( .A(mem[1027]), .Y(n8803) );
  INVX1 U7487 ( .A(mem[125]), .Y(n9705) );
  INVX1 U7488 ( .A(mem[2]), .Y(n9828) );
  INVX1 U7489 ( .A(mem[43]), .Y(n9787) );
  INVX1 U7490 ( .A(mem[782]), .Y(n9048) );
  INVX1 U7491 ( .A(mem[659]), .Y(n9171) );
  INVX1 U7492 ( .A(mem[700]), .Y(n9130) );
  INVX1 U7493 ( .A(mem[1110]), .Y(n8720) );
  INVX1 U7494 ( .A(mem[987]), .Y(n8843) );
  INVX1 U7495 ( .A(mem[1028]), .Y(n8802) );
  INVX1 U7496 ( .A(mem[126]), .Y(n9704) );
  INVX1 U7497 ( .A(mem[3]), .Y(n9827) );
  INVX1 U7498 ( .A(mem[44]), .Y(n9786) );
  INVX1 U7499 ( .A(mem[783]), .Y(n9047) );
  INVX1 U7500 ( .A(mem[660]), .Y(n9170) );
  INVX1 U7501 ( .A(mem[701]), .Y(n9129) );
  INVX1 U7502 ( .A(mem[1111]), .Y(n8719) );
  INVX1 U7503 ( .A(mem[988]), .Y(n8842) );
  INVX1 U7504 ( .A(mem[1029]), .Y(n8801) );
  INVX1 U7505 ( .A(mem[127]), .Y(n9703) );
  INVX1 U7506 ( .A(mem[4]), .Y(n9826) );
  INVX1 U7507 ( .A(mem[45]), .Y(n9785) );
  INVX1 U7508 ( .A(mem[784]), .Y(n9046) );
  INVX1 U7509 ( .A(mem[661]), .Y(n9169) );
  INVX1 U7510 ( .A(mem[702]), .Y(n9128) );
  INVX1 U7511 ( .A(mem[1112]), .Y(n8718) );
  INVX1 U7512 ( .A(mem[989]), .Y(n8841) );
  INVX1 U7513 ( .A(mem[1030]), .Y(n8800) );
  INVX1 U7514 ( .A(mem[128]), .Y(n9702) );
  INVX1 U7515 ( .A(mem[5]), .Y(n9825) );
  INVX1 U7516 ( .A(mem[46]), .Y(n9784) );
  INVX1 U7517 ( .A(mem[785]), .Y(n9045) );
  INVX1 U7518 ( .A(mem[662]), .Y(n9168) );
  INVX1 U7519 ( .A(mem[703]), .Y(n9127) );
  INVX1 U7520 ( .A(mem[1113]), .Y(n8717) );
  INVX1 U7521 ( .A(mem[990]), .Y(n8840) );
  INVX1 U7522 ( .A(mem[1031]), .Y(n8799) );
  INVX1 U7523 ( .A(mem[129]), .Y(n9701) );
  INVX1 U7524 ( .A(mem[6]), .Y(n9824) );
  INVX1 U7525 ( .A(mem[47]), .Y(n9783) );
  INVX1 U7526 ( .A(mem[786]), .Y(n9044) );
  INVX1 U7527 ( .A(mem[663]), .Y(n9167) );
  INVX1 U7528 ( .A(mem[704]), .Y(n9126) );
  INVX1 U7529 ( .A(mem[1114]), .Y(n8716) );
  INVX1 U7530 ( .A(mem[991]), .Y(n8839) );
  INVX1 U7531 ( .A(mem[1032]), .Y(n8798) );
  INVX1 U7532 ( .A(mem[130]), .Y(n9700) );
  INVX1 U7533 ( .A(mem[7]), .Y(n9823) );
  INVX1 U7534 ( .A(mem[48]), .Y(n9782) );
  INVX1 U7535 ( .A(mem[787]), .Y(n9043) );
  INVX1 U7536 ( .A(mem[664]), .Y(n9166) );
  INVX1 U7537 ( .A(mem[705]), .Y(n9125) );
  INVX1 U7538 ( .A(mem[1115]), .Y(n8715) );
  INVX1 U7539 ( .A(mem[992]), .Y(n8838) );
  INVX1 U7540 ( .A(mem[1033]), .Y(n8797) );
  INVX1 U7541 ( .A(mem[131]), .Y(n9699) );
  INVX1 U7542 ( .A(mem[8]), .Y(n9822) );
  INVX1 U7543 ( .A(mem[49]), .Y(n9781) );
  INVX1 U7544 ( .A(mem[788]), .Y(n9042) );
  INVX1 U7545 ( .A(mem[665]), .Y(n9165) );
  INVX1 U7546 ( .A(mem[706]), .Y(n9124) );
  INVX1 U7547 ( .A(mem[1116]), .Y(n8714) );
  INVX1 U7548 ( .A(mem[993]), .Y(n8837) );
  INVX1 U7549 ( .A(mem[1034]), .Y(n8796) );
  INVX1 U7550 ( .A(mem[132]), .Y(n9698) );
  INVX1 U7551 ( .A(mem[9]), .Y(n9821) );
  INVX1 U7552 ( .A(mem[50]), .Y(n9780) );
  INVX1 U7553 ( .A(mem[789]), .Y(n9041) );
  INVX1 U7554 ( .A(mem[666]), .Y(n9164) );
  INVX1 U7555 ( .A(mem[707]), .Y(n9123) );
  INVX1 U7556 ( .A(mem[1117]), .Y(n8713) );
  INVX1 U7557 ( .A(mem[994]), .Y(n8836) );
  INVX1 U7558 ( .A(mem[1035]), .Y(n8795) );
  INVX1 U7559 ( .A(mem[133]), .Y(n9697) );
  INVX1 U7560 ( .A(mem[10]), .Y(n9820) );
  INVX1 U7561 ( .A(mem[51]), .Y(n9779) );
  INVX1 U7562 ( .A(mem[790]), .Y(n9040) );
  INVX1 U7563 ( .A(mem[667]), .Y(n9163) );
  INVX1 U7564 ( .A(mem[708]), .Y(n9122) );
  INVX1 U7565 ( .A(mem[1118]), .Y(n8712) );
  INVX1 U7566 ( .A(mem[995]), .Y(n8835) );
  INVX1 U7567 ( .A(mem[1036]), .Y(n8794) );
  INVX1 U7568 ( .A(mem[134]), .Y(n9696) );
  INVX1 U7569 ( .A(mem[11]), .Y(n9819) );
  INVX1 U7570 ( .A(mem[52]), .Y(n9778) );
  INVX1 U7571 ( .A(mem[791]), .Y(n9039) );
  INVX1 U7572 ( .A(mem[668]), .Y(n9162) );
  INVX1 U7573 ( .A(mem[709]), .Y(n9121) );
  INVX1 U7574 ( .A(mem[1119]), .Y(n8711) );
  INVX1 U7575 ( .A(mem[996]), .Y(n8834) );
  INVX1 U7576 ( .A(mem[1037]), .Y(n8793) );
  INVX1 U7577 ( .A(mem[135]), .Y(n9695) );
  INVX1 U7578 ( .A(mem[12]), .Y(n9818) );
  INVX1 U7579 ( .A(mem[53]), .Y(n9777) );
  INVX1 U7580 ( .A(mem[792]), .Y(n9038) );
  INVX1 U7581 ( .A(mem[669]), .Y(n9161) );
  INVX1 U7582 ( .A(mem[710]), .Y(n9120) );
  INVX1 U7583 ( .A(mem[1120]), .Y(n8710) );
  INVX1 U7584 ( .A(mem[997]), .Y(n8833) );
  INVX1 U7585 ( .A(mem[1038]), .Y(n8792) );
  INVX1 U7586 ( .A(mem[136]), .Y(n9694) );
  INVX1 U7587 ( .A(mem[13]), .Y(n9817) );
  INVX1 U7588 ( .A(mem[54]), .Y(n9776) );
  INVX1 U7589 ( .A(mem[793]), .Y(n9037) );
  INVX1 U7590 ( .A(mem[670]), .Y(n9160) );
  INVX1 U7591 ( .A(mem[711]), .Y(n9119) );
  INVX1 U7592 ( .A(mem[1121]), .Y(n8709) );
  INVX1 U7593 ( .A(mem[998]), .Y(n8832) );
  INVX1 U7594 ( .A(mem[1039]), .Y(n8791) );
  INVX1 U7595 ( .A(mem[137]), .Y(n9693) );
  INVX1 U7596 ( .A(mem[14]), .Y(n9816) );
  INVX1 U7597 ( .A(mem[55]), .Y(n9775) );
  INVX1 U7598 ( .A(mem[794]), .Y(n9036) );
  INVX1 U7599 ( .A(mem[671]), .Y(n9159) );
  INVX1 U7600 ( .A(mem[712]), .Y(n9118) );
  INVX1 U7601 ( .A(mem[1122]), .Y(n8708) );
  INVX1 U7602 ( .A(mem[999]), .Y(n8831) );
  INVX1 U7603 ( .A(mem[1040]), .Y(n8790) );
  INVX1 U7604 ( .A(mem[138]), .Y(n9692) );
  INVX1 U7605 ( .A(mem[15]), .Y(n9815) );
  INVX1 U7606 ( .A(mem[56]), .Y(n9774) );
  INVX1 U7607 ( .A(mem[795]), .Y(n9035) );
  INVX1 U7608 ( .A(mem[672]), .Y(n9158) );
  INVX1 U7609 ( .A(mem[713]), .Y(n9117) );
  INVX1 U7610 ( .A(mem[1123]), .Y(n8707) );
  INVX1 U7611 ( .A(mem[1000]), .Y(n8830) );
  INVX1 U7612 ( .A(mem[1041]), .Y(n8789) );
  INVX1 U7613 ( .A(mem[139]), .Y(n9691) );
  INVX1 U7614 ( .A(mem[16]), .Y(n9814) );
  INVX1 U7615 ( .A(mem[57]), .Y(n9773) );
  INVX1 U7616 ( .A(mem[796]), .Y(n9034) );
  INVX1 U7617 ( .A(mem[673]), .Y(n9157) );
  INVX1 U7618 ( .A(mem[714]), .Y(n9116) );
  INVX1 U7619 ( .A(mem[1124]), .Y(n8706) );
  INVX1 U7620 ( .A(mem[1001]), .Y(n8829) );
  INVX1 U7621 ( .A(mem[1042]), .Y(n8788) );
  INVX1 U7622 ( .A(mem[140]), .Y(n9690) );
  INVX1 U7623 ( .A(mem[17]), .Y(n9813) );
  INVX1 U7624 ( .A(mem[58]), .Y(n9772) );
  INVX1 U7625 ( .A(mem[797]), .Y(n9033) );
  INVX1 U7626 ( .A(mem[674]), .Y(n9156) );
  INVX1 U7627 ( .A(mem[715]), .Y(n9115) );
  INVX1 U7628 ( .A(mem[1125]), .Y(n8705) );
  INVX1 U7629 ( .A(mem[1002]), .Y(n8828) );
  INVX1 U7630 ( .A(mem[1043]), .Y(n8787) );
  INVX1 U7631 ( .A(mem[141]), .Y(n9689) );
  INVX1 U7632 ( .A(mem[18]), .Y(n9812) );
  INVX1 U7633 ( .A(mem[59]), .Y(n9771) );
  INVX1 U7634 ( .A(mem[798]), .Y(n9032) );
  INVX1 U7635 ( .A(mem[675]), .Y(n9155) );
  INVX1 U7636 ( .A(mem[716]), .Y(n9114) );
  INVX1 U7637 ( .A(mem[1126]), .Y(n8704) );
  INVX1 U7638 ( .A(mem[1003]), .Y(n8827) );
  INVX1 U7639 ( .A(mem[1044]), .Y(n8786) );
  INVX1 U7640 ( .A(mem[142]), .Y(n9688) );
  INVX1 U7641 ( .A(mem[19]), .Y(n9811) );
  INVX1 U7642 ( .A(mem[60]), .Y(n9770) );
  INVX1 U7643 ( .A(mem[799]), .Y(n9031) );
  INVX1 U7644 ( .A(mem[676]), .Y(n9154) );
  INVX1 U7645 ( .A(mem[717]), .Y(n9113) );
  INVX1 U7646 ( .A(mem[1127]), .Y(n8703) );
  INVX1 U7647 ( .A(mem[1004]), .Y(n8826) );
  INVX1 U7648 ( .A(mem[1045]), .Y(n8785) );
  INVX1 U7649 ( .A(mem[143]), .Y(n9687) );
  INVX1 U7650 ( .A(mem[20]), .Y(n9810) );
  INVX1 U7651 ( .A(mem[61]), .Y(n9769) );
  INVX1 U7652 ( .A(mem[800]), .Y(n9030) );
  INVX1 U7653 ( .A(mem[677]), .Y(n9153) );
  INVX1 U7654 ( .A(mem[718]), .Y(n9112) );
  INVX1 U7655 ( .A(mem[1128]), .Y(n8702) );
  INVX1 U7656 ( .A(mem[1005]), .Y(n8825) );
  INVX1 U7657 ( .A(mem[1046]), .Y(n8784) );
  INVX1 U7658 ( .A(mem[144]), .Y(n9686) );
  INVX1 U7659 ( .A(mem[21]), .Y(n9809) );
  INVX1 U7660 ( .A(mem[62]), .Y(n9768) );
  INVX1 U7661 ( .A(mem[801]), .Y(n9029) );
  INVX1 U7662 ( .A(mem[678]), .Y(n9152) );
  INVX1 U7663 ( .A(mem[719]), .Y(n9111) );
  INVX1 U7664 ( .A(mem[1129]), .Y(n8701) );
  INVX1 U7665 ( .A(mem[1006]), .Y(n8824) );
  INVX1 U7666 ( .A(mem[1047]), .Y(n8783) );
  INVX1 U7667 ( .A(mem[145]), .Y(n9685) );
  INVX1 U7668 ( .A(mem[22]), .Y(n9808) );
  INVX1 U7669 ( .A(mem[63]), .Y(n9767) );
  INVX1 U7670 ( .A(mem[802]), .Y(n9028) );
  INVX1 U7671 ( .A(mem[679]), .Y(n9151) );
  INVX1 U7672 ( .A(mem[720]), .Y(n9110) );
  INVX1 U7673 ( .A(mem[1130]), .Y(n8700) );
  INVX1 U7674 ( .A(mem[1007]), .Y(n8823) );
  INVX1 U7675 ( .A(mem[1048]), .Y(n8782) );
  INVX1 U7676 ( .A(mem[146]), .Y(n9684) );
  INVX1 U7677 ( .A(mem[23]), .Y(n9807) );
  INVX1 U7678 ( .A(mem[64]), .Y(n9766) );
  INVX1 U7679 ( .A(mem[803]), .Y(n9027) );
  INVX1 U7680 ( .A(mem[680]), .Y(n9150) );
  INVX1 U7681 ( .A(mem[721]), .Y(n9109) );
  INVX1 U7682 ( .A(mem[1131]), .Y(n8699) );
  INVX1 U7683 ( .A(mem[1008]), .Y(n8822) );
  INVX1 U7684 ( .A(mem[1049]), .Y(n8781) );
  INVX1 U7685 ( .A(mem[147]), .Y(n9683) );
  INVX1 U7686 ( .A(mem[24]), .Y(n9806) );
  INVX1 U7687 ( .A(mem[65]), .Y(n9765) );
  INVX1 U7688 ( .A(mem[804]), .Y(n9026) );
  INVX1 U7689 ( .A(mem[681]), .Y(n9149) );
  INVX1 U7690 ( .A(mem[722]), .Y(n9108) );
  INVX1 U7691 ( .A(mem[1132]), .Y(n8698) );
  INVX1 U7692 ( .A(mem[1009]), .Y(n8821) );
  INVX1 U7693 ( .A(mem[1050]), .Y(n8780) );
  INVX1 U7694 ( .A(mem[148]), .Y(n9682) );
  INVX1 U7695 ( .A(mem[25]), .Y(n9805) );
  INVX1 U7696 ( .A(mem[66]), .Y(n9764) );
  INVX1 U7697 ( .A(mem[805]), .Y(n9025) );
  INVX1 U7698 ( .A(mem[682]), .Y(n9148) );
  INVX1 U7699 ( .A(mem[723]), .Y(n9107) );
  INVX1 U7700 ( .A(mem[1133]), .Y(n8697) );
  INVX1 U7701 ( .A(mem[1010]), .Y(n8820) );
  INVX1 U7702 ( .A(mem[1051]), .Y(n8779) );
  INVX1 U7703 ( .A(mem[149]), .Y(n9681) );
  INVX1 U7704 ( .A(mem[26]), .Y(n9804) );
  INVX1 U7705 ( .A(mem[67]), .Y(n9763) );
  INVX1 U7706 ( .A(mem[806]), .Y(n9024) );
  INVX1 U7707 ( .A(mem[683]), .Y(n9147) );
  INVX1 U7708 ( .A(mem[724]), .Y(n9106) );
  INVX1 U7709 ( .A(mem[1134]), .Y(n8696) );
  INVX1 U7710 ( .A(mem[1011]), .Y(n8819) );
  INVX1 U7711 ( .A(mem[1052]), .Y(n8778) );
  INVX1 U7712 ( .A(mem[150]), .Y(n9680) );
  INVX1 U7713 ( .A(mem[27]), .Y(n9803) );
  INVX1 U7714 ( .A(mem[68]), .Y(n9762) );
  INVX1 U7715 ( .A(mem[807]), .Y(n9023) );
  INVX1 U7716 ( .A(mem[684]), .Y(n9146) );
  INVX1 U7717 ( .A(mem[725]), .Y(n9105) );
  INVX1 U7718 ( .A(mem[1135]), .Y(n8695) );
  INVX1 U7719 ( .A(mem[1012]), .Y(n8818) );
  INVX1 U7720 ( .A(mem[1053]), .Y(n8777) );
  INVX1 U7721 ( .A(mem[151]), .Y(n9679) );
  INVX1 U7722 ( .A(mem[28]), .Y(n9802) );
  INVX1 U7723 ( .A(mem[69]), .Y(n9761) );
  INVX1 U7724 ( .A(mem[808]), .Y(n9022) );
  INVX1 U7725 ( .A(mem[685]), .Y(n9145) );
  INVX1 U7726 ( .A(mem[726]), .Y(n9104) );
  INVX1 U7727 ( .A(mem[1136]), .Y(n8694) );
  INVX1 U7728 ( .A(mem[1013]), .Y(n8817) );
  INVX1 U7729 ( .A(mem[1054]), .Y(n8776) );
  INVX1 U7730 ( .A(mem[152]), .Y(n9678) );
  INVX1 U7731 ( .A(mem[29]), .Y(n9801) );
  INVX1 U7732 ( .A(mem[70]), .Y(n9760) );
  INVX1 U7733 ( .A(mem[809]), .Y(n9021) );
  INVX1 U7734 ( .A(mem[686]), .Y(n9144) );
  INVX1 U7735 ( .A(mem[727]), .Y(n9103) );
  INVX1 U7736 ( .A(mem[1137]), .Y(n8693) );
  INVX1 U7737 ( .A(mem[1014]), .Y(n8816) );
  INVX1 U7738 ( .A(mem[1055]), .Y(n8775) );
  INVX1 U7739 ( .A(mem[153]), .Y(n9677) );
  INVX1 U7740 ( .A(mem[30]), .Y(n9800) );
  INVX1 U7741 ( .A(mem[71]), .Y(n9759) );
  INVX1 U7742 ( .A(mem[810]), .Y(n9020) );
  INVX1 U7743 ( .A(mem[687]), .Y(n9143) );
  INVX1 U7744 ( .A(mem[728]), .Y(n9102) );
  INVX1 U7745 ( .A(mem[1138]), .Y(n8692) );
  INVX1 U7746 ( .A(mem[1015]), .Y(n8815) );
  INVX1 U7747 ( .A(mem[1056]), .Y(n8774) );
  INVX1 U7748 ( .A(mem[154]), .Y(n9676) );
  INVX1 U7749 ( .A(mem[31]), .Y(n9799) );
  INVX1 U7750 ( .A(mem[72]), .Y(n9758) );
  INVX1 U7751 ( .A(mem[811]), .Y(n9019) );
  INVX1 U7752 ( .A(mem[688]), .Y(n9142) );
  INVX1 U7753 ( .A(mem[729]), .Y(n9101) );
  INVX1 U7754 ( .A(mem[1139]), .Y(n8691) );
  INVX1 U7755 ( .A(mem[1016]), .Y(n8814) );
  INVX1 U7756 ( .A(mem[1057]), .Y(n8773) );
  INVX1 U7757 ( .A(mem[155]), .Y(n9675) );
  INVX1 U7758 ( .A(mem[32]), .Y(n9798) );
  INVX1 U7759 ( .A(mem[73]), .Y(n9757) );
  INVX1 U7760 ( .A(mem[812]), .Y(n9018) );
  INVX1 U7761 ( .A(mem[689]), .Y(n9141) );
  INVX1 U7762 ( .A(mem[730]), .Y(n9100) );
  INVX1 U7763 ( .A(mem[1140]), .Y(n8690) );
  INVX1 U7764 ( .A(mem[1017]), .Y(n8813) );
  INVX1 U7765 ( .A(mem[1058]), .Y(n8772) );
  INVX1 U7766 ( .A(mem[156]), .Y(n9674) );
  INVX1 U7767 ( .A(mem[33]), .Y(n9797) );
  INVX1 U7768 ( .A(mem[74]), .Y(n9756) );
  INVX1 U7769 ( .A(mem[813]), .Y(n9017) );
  INVX1 U7770 ( .A(mem[690]), .Y(n9140) );
  INVX1 U7771 ( .A(mem[731]), .Y(n9099) );
  INVX1 U7772 ( .A(mem[1141]), .Y(n8689) );
  INVX1 U7773 ( .A(mem[1018]), .Y(n8812) );
  INVX1 U7774 ( .A(mem[1059]), .Y(n8771) );
  INVX1 U7775 ( .A(mem[157]), .Y(n9673) );
  INVX1 U7776 ( .A(mem[34]), .Y(n9796) );
  INVX1 U7777 ( .A(mem[75]), .Y(n9755) );
  INVX1 U7778 ( .A(mem[814]), .Y(n9016) );
  INVX1 U7779 ( .A(mem[691]), .Y(n9139) );
  INVX1 U7780 ( .A(mem[732]), .Y(n9098) );
  INVX1 U7781 ( .A(mem[1142]), .Y(n8688) );
  INVX1 U7782 ( .A(mem[1019]), .Y(n8811) );
  INVX1 U7783 ( .A(mem[1060]), .Y(n8770) );
  INVX1 U7784 ( .A(mem[158]), .Y(n9672) );
  INVX1 U7785 ( .A(mem[35]), .Y(n9795) );
  INVX1 U7786 ( .A(mem[76]), .Y(n9754) );
  INVX1 U7787 ( .A(mem[815]), .Y(n9015) );
  INVX1 U7788 ( .A(mem[692]), .Y(n9138) );
  INVX1 U7789 ( .A(mem[733]), .Y(n9097) );
  INVX1 U7790 ( .A(mem[1143]), .Y(n8687) );
  INVX1 U7791 ( .A(mem[1020]), .Y(n8810) );
  INVX1 U7792 ( .A(mem[1061]), .Y(n8769) );
  INVX1 U7793 ( .A(mem[159]), .Y(n9671) );
  INVX1 U7794 ( .A(mem[36]), .Y(n9794) );
  INVX1 U7795 ( .A(mem[77]), .Y(n9753) );
  INVX1 U7796 ( .A(mem[816]), .Y(n9014) );
  INVX1 U7797 ( .A(mem[693]), .Y(n9137) );
  INVX1 U7798 ( .A(mem[734]), .Y(n9096) );
  INVX1 U7799 ( .A(mem[1144]), .Y(n8686) );
  INVX1 U7800 ( .A(mem[1021]), .Y(n8809) );
  INVX1 U7801 ( .A(mem[1062]), .Y(n8768) );
  INVX1 U7802 ( .A(mem[160]), .Y(n9670) );
  INVX1 U7803 ( .A(mem[37]), .Y(n9793) );
  INVX1 U7804 ( .A(mem[78]), .Y(n9752) );
  INVX1 U7805 ( .A(mem[817]), .Y(n9013) );
  INVX1 U7806 ( .A(mem[694]), .Y(n9136) );
  INVX1 U7807 ( .A(mem[735]), .Y(n9095) );
  INVX1 U7808 ( .A(mem[1145]), .Y(n8685) );
  INVX1 U7809 ( .A(mem[1022]), .Y(n8808) );
  INVX1 U7810 ( .A(mem[1063]), .Y(n8767) );
  INVX1 U7811 ( .A(mem[161]), .Y(n9669) );
  INVX1 U7812 ( .A(mem[38]), .Y(n9792) );
  INVX1 U7813 ( .A(mem[79]), .Y(n9751) );
  INVX1 U7814 ( .A(mem[818]), .Y(n9012) );
  INVX1 U7815 ( .A(mem[695]), .Y(n9135) );
  INVX1 U7816 ( .A(mem[736]), .Y(n9094) );
  INVX1 U7817 ( .A(mem[1146]), .Y(n8684) );
  INVX1 U7818 ( .A(mem[1023]), .Y(n8807) );
  INVX1 U7819 ( .A(mem[1064]), .Y(n8766) );
  INVX1 U7820 ( .A(mem[162]), .Y(n9668) );
  INVX1 U7821 ( .A(mem[39]), .Y(n9791) );
  INVX1 U7822 ( .A(mem[80]), .Y(n9750) );
  INVX1 U7823 ( .A(mem[819]), .Y(n9011) );
  INVX1 U7824 ( .A(mem[696]), .Y(n9134) );
  INVX1 U7825 ( .A(mem[737]), .Y(n9093) );
  INVX1 U7826 ( .A(mem[1147]), .Y(n8683) );
  INVX1 U7827 ( .A(mem[1024]), .Y(n8806) );
  INVX1 U7828 ( .A(mem[1065]), .Y(n8765) );
  INVX1 U7829 ( .A(mem[163]), .Y(n9667) );
  INVX1 U7830 ( .A(mem[40]), .Y(n9790) );
  INVX1 U7831 ( .A(mem[81]), .Y(n9749) );
  INVX1 U7832 ( .A(mem[451]), .Y(n9379) );
  INVX1 U7833 ( .A(mem[328]), .Y(n9502) );
  INVX1 U7834 ( .A(mem[369]), .Y(n9461) );
  INVX1 U7835 ( .A(mem[452]), .Y(n9378) );
  INVX1 U7836 ( .A(mem[329]), .Y(n9501) );
  INVX1 U7837 ( .A(mem[370]), .Y(n9460) );
  INVX1 U7838 ( .A(mem[453]), .Y(n9377) );
  INVX1 U7839 ( .A(mem[330]), .Y(n9500) );
  INVX1 U7840 ( .A(mem[371]), .Y(n9459) );
  INVX1 U7841 ( .A(mem[454]), .Y(n9376) );
  INVX1 U7842 ( .A(mem[331]), .Y(n9499) );
  INVX1 U7843 ( .A(mem[372]), .Y(n9458) );
  INVX1 U7844 ( .A(mem[455]), .Y(n9375) );
  INVX1 U7845 ( .A(mem[332]), .Y(n9498) );
  INVX1 U7846 ( .A(mem[373]), .Y(n9457) );
  INVX1 U7847 ( .A(mem[456]), .Y(n9374) );
  INVX1 U7848 ( .A(mem[333]), .Y(n9497) );
  INVX1 U7849 ( .A(mem[374]), .Y(n9456) );
  INVX1 U7850 ( .A(mem[457]), .Y(n9373) );
  INVX1 U7851 ( .A(mem[334]), .Y(n9496) );
  INVX1 U7852 ( .A(mem[375]), .Y(n9455) );
  INVX1 U7853 ( .A(mem[458]), .Y(n9372) );
  INVX1 U7854 ( .A(mem[335]), .Y(n9495) );
  INVX1 U7855 ( .A(mem[376]), .Y(n9454) );
  INVX1 U7856 ( .A(mem[459]), .Y(n9371) );
  INVX1 U7857 ( .A(mem[336]), .Y(n9494) );
  INVX1 U7858 ( .A(mem[377]), .Y(n9453) );
  INVX1 U7859 ( .A(mem[460]), .Y(n9370) );
  INVX1 U7860 ( .A(mem[337]), .Y(n9493) );
  INVX1 U7861 ( .A(mem[378]), .Y(n9452) );
  INVX1 U7862 ( .A(mem[461]), .Y(n9369) );
  INVX1 U7863 ( .A(mem[338]), .Y(n9492) );
  INVX1 U7864 ( .A(mem[379]), .Y(n9451) );
  INVX1 U7865 ( .A(mem[462]), .Y(n9368) );
  INVX1 U7866 ( .A(mem[339]), .Y(n9491) );
  INVX1 U7867 ( .A(mem[380]), .Y(n9450) );
  INVX1 U7868 ( .A(mem[463]), .Y(n9367) );
  INVX1 U7869 ( .A(mem[340]), .Y(n9490) );
  INVX1 U7870 ( .A(mem[381]), .Y(n9449) );
  INVX1 U7871 ( .A(mem[464]), .Y(n9366) );
  INVX1 U7872 ( .A(mem[341]), .Y(n9489) );
  INVX1 U7873 ( .A(mem[382]), .Y(n9448) );
  INVX1 U7874 ( .A(mem[465]), .Y(n9365) );
  INVX1 U7875 ( .A(mem[342]), .Y(n9488) );
  INVX1 U7876 ( .A(mem[383]), .Y(n9447) );
  INVX1 U7877 ( .A(mem[466]), .Y(n9364) );
  INVX1 U7878 ( .A(mem[343]), .Y(n9487) );
  INVX1 U7879 ( .A(mem[384]), .Y(n9446) );
  INVX1 U7880 ( .A(mem[467]), .Y(n9363) );
  INVX1 U7881 ( .A(mem[344]), .Y(n9486) );
  INVX1 U7882 ( .A(mem[385]), .Y(n9445) );
  INVX1 U7883 ( .A(mem[468]), .Y(n9362) );
  INVX1 U7884 ( .A(mem[345]), .Y(n9485) );
  INVX1 U7885 ( .A(mem[386]), .Y(n9444) );
  INVX1 U7886 ( .A(mem[469]), .Y(n9361) );
  INVX1 U7887 ( .A(mem[346]), .Y(n9484) );
  INVX1 U7888 ( .A(mem[387]), .Y(n9443) );
  INVX1 U7889 ( .A(mem[470]), .Y(n9360) );
  INVX1 U7890 ( .A(mem[347]), .Y(n9483) );
  INVX1 U7891 ( .A(mem[388]), .Y(n9442) );
  INVX1 U7892 ( .A(mem[471]), .Y(n9359) );
  INVX1 U7893 ( .A(mem[348]), .Y(n9482) );
  INVX1 U7894 ( .A(mem[389]), .Y(n9441) );
  INVX1 U7895 ( .A(mem[472]), .Y(n9358) );
  INVX1 U7896 ( .A(mem[349]), .Y(n9481) );
  INVX1 U7897 ( .A(mem[390]), .Y(n9440) );
  INVX1 U7898 ( .A(mem[473]), .Y(n9357) );
  INVX1 U7899 ( .A(mem[350]), .Y(n9480) );
  INVX1 U7900 ( .A(mem[391]), .Y(n9439) );
  INVX1 U7901 ( .A(mem[474]), .Y(n9356) );
  INVX1 U7902 ( .A(mem[351]), .Y(n9479) );
  INVX1 U7903 ( .A(mem[392]), .Y(n9438) );
  INVX1 U7904 ( .A(mem[475]), .Y(n9355) );
  INVX1 U7905 ( .A(mem[352]), .Y(n9478) );
  INVX1 U7906 ( .A(mem[393]), .Y(n9437) );
  INVX1 U7907 ( .A(mem[476]), .Y(n9354) );
  INVX1 U7908 ( .A(mem[353]), .Y(n9477) );
  INVX1 U7909 ( .A(mem[394]), .Y(n9436) );
  INVX1 U7910 ( .A(mem[477]), .Y(n9353) );
  INVX1 U7911 ( .A(mem[354]), .Y(n9476) );
  INVX1 U7912 ( .A(mem[395]), .Y(n9435) );
  INVX1 U7913 ( .A(mem[478]), .Y(n9352) );
  INVX1 U7914 ( .A(mem[355]), .Y(n9475) );
  INVX1 U7915 ( .A(mem[396]), .Y(n9434) );
  INVX1 U7916 ( .A(mem[479]), .Y(n9351) );
  INVX1 U7917 ( .A(mem[356]), .Y(n9474) );
  INVX1 U7918 ( .A(mem[397]), .Y(n9433) );
  INVX1 U7919 ( .A(mem[480]), .Y(n9350) );
  INVX1 U7920 ( .A(mem[357]), .Y(n9473) );
  INVX1 U7921 ( .A(mem[398]), .Y(n9432) );
  INVX1 U7922 ( .A(mem[481]), .Y(n9349) );
  INVX1 U7923 ( .A(mem[358]), .Y(n9472) );
  INVX1 U7924 ( .A(mem[399]), .Y(n9431) );
  INVX1 U7925 ( .A(mem[482]), .Y(n9348) );
  INVX1 U7926 ( .A(mem[359]), .Y(n9471) );
  INVX1 U7927 ( .A(mem[400]), .Y(n9430) );
  INVX1 U7928 ( .A(mem[483]), .Y(n9347) );
  INVX1 U7929 ( .A(mem[360]), .Y(n9470) );
  INVX1 U7930 ( .A(mem[401]), .Y(n9429) );
  INVX1 U7931 ( .A(mem[484]), .Y(n9346) );
  INVX1 U7932 ( .A(mem[361]), .Y(n9469) );
  INVX1 U7933 ( .A(mem[402]), .Y(n9428) );
  INVX1 U7934 ( .A(mem[485]), .Y(n9345) );
  INVX1 U7935 ( .A(mem[362]), .Y(n9468) );
  INVX1 U7936 ( .A(mem[403]), .Y(n9427) );
  INVX1 U7937 ( .A(mem[486]), .Y(n9344) );
  INVX1 U7938 ( .A(mem[363]), .Y(n9467) );
  INVX1 U7939 ( .A(mem[404]), .Y(n9426) );
  INVX1 U7940 ( .A(mem[487]), .Y(n9343) );
  INVX1 U7941 ( .A(mem[364]), .Y(n9466) );
  INVX1 U7942 ( .A(mem[405]), .Y(n9425) );
  INVX1 U7943 ( .A(mem[488]), .Y(n9342) );
  INVX1 U7944 ( .A(mem[365]), .Y(n9465) );
  INVX1 U7945 ( .A(mem[406]), .Y(n9424) );
  INVX1 U7946 ( .A(mem[489]), .Y(n9341) );
  INVX1 U7947 ( .A(mem[366]), .Y(n9464) );
  INVX1 U7948 ( .A(mem[407]), .Y(n9423) );
  INVX1 U7949 ( .A(mem[490]), .Y(n9340) );
  INVX1 U7950 ( .A(mem[367]), .Y(n9463) );
  INVX1 U7951 ( .A(mem[408]), .Y(n9422) );
  INVX1 U7952 ( .A(mem[491]), .Y(n9339) );
  INVX1 U7953 ( .A(mem[368]), .Y(n9462) );
  INVX1 U7954 ( .A(mem[409]), .Y(n9421) );
  INVX1 U7955 ( .A(mem[943]), .Y(n8887) );
  INVX1 U7956 ( .A(mem[820]), .Y(n9010) );
  INVX1 U7957 ( .A(mem[1271]), .Y(n8559) );
  INVX1 U7958 ( .A(mem[1148]), .Y(n8682) );
  INVX1 U7959 ( .A(mem[287]), .Y(n9543) );
  INVX1 U7960 ( .A(mem[164]), .Y(n9666) );
  INVX1 U7961 ( .A(mem[944]), .Y(n8886) );
  INVX1 U7962 ( .A(mem[821]), .Y(n9009) );
  INVX1 U7963 ( .A(mem[1272]), .Y(n8558) );
  INVX1 U7964 ( .A(mem[1149]), .Y(n8681) );
  INVX1 U7965 ( .A(mem[288]), .Y(n9542) );
  INVX1 U7966 ( .A(mem[165]), .Y(n9665) );
  INVX1 U7967 ( .A(mem[945]), .Y(n8885) );
  INVX1 U7968 ( .A(mem[822]), .Y(n9008) );
  INVX1 U7969 ( .A(mem[1273]), .Y(n8557) );
  INVX1 U7970 ( .A(mem[1150]), .Y(n8680) );
  INVX1 U7971 ( .A(mem[289]), .Y(n9541) );
  INVX1 U7972 ( .A(mem[166]), .Y(n9664) );
  INVX1 U7973 ( .A(mem[946]), .Y(n8884) );
  INVX1 U7974 ( .A(mem[823]), .Y(n9007) );
  INVX1 U7975 ( .A(mem[1274]), .Y(n8556) );
  INVX1 U7976 ( .A(mem[1151]), .Y(n8679) );
  INVX1 U7977 ( .A(mem[290]), .Y(n9540) );
  INVX1 U7978 ( .A(mem[167]), .Y(n9663) );
  INVX1 U7979 ( .A(mem[947]), .Y(n8883) );
  INVX1 U7980 ( .A(mem[824]), .Y(n9006) );
  INVX1 U7981 ( .A(mem[1275]), .Y(n8555) );
  INVX1 U7982 ( .A(mem[1152]), .Y(n8678) );
  INVX1 U7983 ( .A(mem[291]), .Y(n9539) );
  INVX1 U7984 ( .A(mem[168]), .Y(n9662) );
  INVX1 U7985 ( .A(mem[948]), .Y(n8882) );
  INVX1 U7986 ( .A(mem[825]), .Y(n9005) );
  INVX1 U7987 ( .A(mem[1276]), .Y(n8554) );
  INVX1 U7988 ( .A(mem[1153]), .Y(n8677) );
  INVX1 U7989 ( .A(mem[292]), .Y(n9538) );
  INVX1 U7990 ( .A(mem[169]), .Y(n9661) );
  INVX1 U7991 ( .A(mem[949]), .Y(n8881) );
  INVX1 U7992 ( .A(mem[826]), .Y(n9004) );
  INVX1 U7993 ( .A(mem[1277]), .Y(n8553) );
  INVX1 U7994 ( .A(mem[1154]), .Y(n8676) );
  INVX1 U7995 ( .A(mem[293]), .Y(n9537) );
  INVX1 U7996 ( .A(mem[170]), .Y(n9660) );
  INVX1 U7997 ( .A(mem[950]), .Y(n8880) );
  INVX1 U7998 ( .A(mem[827]), .Y(n9003) );
  INVX1 U7999 ( .A(mem[1278]), .Y(n8552) );
  INVX1 U8000 ( .A(mem[1155]), .Y(n8675) );
  INVX1 U8001 ( .A(mem[294]), .Y(n9536) );
  INVX1 U8002 ( .A(mem[171]), .Y(n9659) );
  INVX1 U8003 ( .A(mem[951]), .Y(n8879) );
  INVX1 U8004 ( .A(mem[828]), .Y(n9002) );
  INVX1 U8005 ( .A(mem[1279]), .Y(n8551) );
  INVX1 U8006 ( .A(mem[1156]), .Y(n8674) );
  INVX1 U8007 ( .A(mem[295]), .Y(n9535) );
  INVX1 U8008 ( .A(mem[172]), .Y(n9658) );
  INVX1 U8009 ( .A(mem[952]), .Y(n8878) );
  INVX1 U8010 ( .A(mem[829]), .Y(n9001) );
  INVX1 U8011 ( .A(mem[1280]), .Y(n8550) );
  INVX1 U8012 ( .A(mem[1157]), .Y(n8673) );
  INVX1 U8013 ( .A(mem[296]), .Y(n9534) );
  INVX1 U8014 ( .A(mem[173]), .Y(n9657) );
  INVX1 U8015 ( .A(mem[953]), .Y(n8877) );
  INVX1 U8016 ( .A(mem[830]), .Y(n9000) );
  INVX1 U8017 ( .A(mem[1281]), .Y(n8549) );
  INVX1 U8018 ( .A(mem[1158]), .Y(n8672) );
  INVX1 U8019 ( .A(mem[297]), .Y(n9533) );
  INVX1 U8020 ( .A(mem[174]), .Y(n9656) );
  INVX1 U8021 ( .A(mem[954]), .Y(n8876) );
  INVX1 U8022 ( .A(mem[831]), .Y(n8999) );
  INVX1 U8023 ( .A(mem[1282]), .Y(n8548) );
  INVX1 U8024 ( .A(mem[1159]), .Y(n8671) );
  INVX1 U8025 ( .A(mem[298]), .Y(n9532) );
  INVX1 U8026 ( .A(mem[175]), .Y(n9655) );
  INVX1 U8027 ( .A(mem[955]), .Y(n8875) );
  INVX1 U8028 ( .A(mem[832]), .Y(n8998) );
  INVX1 U8029 ( .A(mem[1283]), .Y(n8547) );
  INVX1 U8030 ( .A(mem[1160]), .Y(n8670) );
  INVX1 U8031 ( .A(mem[299]), .Y(n9531) );
  INVX1 U8032 ( .A(mem[176]), .Y(n9654) );
  INVX1 U8033 ( .A(mem[956]), .Y(n8874) );
  INVX1 U8034 ( .A(mem[833]), .Y(n8997) );
  INVX1 U8035 ( .A(mem[1284]), .Y(n8546) );
  INVX1 U8036 ( .A(mem[1161]), .Y(n8669) );
  INVX1 U8037 ( .A(mem[300]), .Y(n9530) );
  INVX1 U8038 ( .A(mem[177]), .Y(n9653) );
  INVX1 U8039 ( .A(mem[957]), .Y(n8873) );
  INVX1 U8040 ( .A(mem[834]), .Y(n8996) );
  INVX1 U8041 ( .A(mem[1285]), .Y(n8545) );
  INVX1 U8042 ( .A(mem[1162]), .Y(n8668) );
  INVX1 U8043 ( .A(mem[301]), .Y(n9529) );
  INVX1 U8044 ( .A(mem[178]), .Y(n9652) );
  INVX1 U8045 ( .A(mem[958]), .Y(n8872) );
  INVX1 U8046 ( .A(mem[835]), .Y(n8995) );
  INVX1 U8047 ( .A(mem[1286]), .Y(n8544) );
  INVX1 U8048 ( .A(mem[1163]), .Y(n8667) );
  INVX1 U8049 ( .A(mem[302]), .Y(n9528) );
  INVX1 U8050 ( .A(mem[179]), .Y(n9651) );
  INVX1 U8051 ( .A(mem[959]), .Y(n8871) );
  INVX1 U8052 ( .A(mem[836]), .Y(n8994) );
  INVX1 U8053 ( .A(mem[1287]), .Y(n8543) );
  INVX1 U8054 ( .A(mem[1164]), .Y(n8666) );
  INVX1 U8055 ( .A(mem[303]), .Y(n9527) );
  INVX1 U8056 ( .A(mem[180]), .Y(n9650) );
  INVX1 U8057 ( .A(mem[960]), .Y(n8870) );
  INVX1 U8058 ( .A(mem[837]), .Y(n8993) );
  INVX1 U8059 ( .A(mem[1288]), .Y(n8542) );
  INVX1 U8060 ( .A(mem[1165]), .Y(n8665) );
  INVX1 U8061 ( .A(mem[304]), .Y(n9526) );
  INVX1 U8062 ( .A(mem[181]), .Y(n9649) );
  INVX1 U8063 ( .A(mem[961]), .Y(n8869) );
  INVX1 U8064 ( .A(mem[838]), .Y(n8992) );
  INVX1 U8065 ( .A(mem[1289]), .Y(n8541) );
  INVX1 U8066 ( .A(mem[1166]), .Y(n8664) );
  INVX1 U8067 ( .A(mem[305]), .Y(n9525) );
  INVX1 U8068 ( .A(mem[182]), .Y(n9648) );
  INVX1 U8069 ( .A(mem[962]), .Y(n8868) );
  INVX1 U8070 ( .A(mem[839]), .Y(n8991) );
  INVX1 U8071 ( .A(mem[1290]), .Y(n8540) );
  INVX1 U8072 ( .A(mem[1167]), .Y(n8663) );
  INVX1 U8073 ( .A(mem[306]), .Y(n9524) );
  INVX1 U8074 ( .A(mem[183]), .Y(n9647) );
  INVX1 U8075 ( .A(mem[963]), .Y(n8867) );
  INVX1 U8076 ( .A(mem[840]), .Y(n8990) );
  INVX1 U8077 ( .A(mem[1291]), .Y(n8539) );
  INVX1 U8078 ( .A(mem[1168]), .Y(n8662) );
  INVX1 U8079 ( .A(mem[307]), .Y(n9523) );
  INVX1 U8080 ( .A(mem[184]), .Y(n9646) );
  INVX1 U8081 ( .A(mem[964]), .Y(n8866) );
  INVX1 U8082 ( .A(mem[841]), .Y(n8989) );
  INVX1 U8083 ( .A(mem[1292]), .Y(n8538) );
  INVX1 U8084 ( .A(mem[1169]), .Y(n8661) );
  INVX1 U8085 ( .A(mem[308]), .Y(n9522) );
  INVX1 U8086 ( .A(mem[185]), .Y(n9645) );
  INVX1 U8087 ( .A(mem[965]), .Y(n8865) );
  INVX1 U8088 ( .A(mem[842]), .Y(n8988) );
  INVX1 U8089 ( .A(mem[1293]), .Y(n8537) );
  INVX1 U8090 ( .A(mem[1170]), .Y(n8660) );
  INVX1 U8091 ( .A(mem[309]), .Y(n9521) );
  INVX1 U8092 ( .A(mem[186]), .Y(n9644) );
  INVX1 U8093 ( .A(mem[966]), .Y(n8864) );
  INVX1 U8094 ( .A(mem[843]), .Y(n8987) );
  INVX1 U8095 ( .A(mem[1294]), .Y(n8536) );
  INVX1 U8096 ( .A(mem[1171]), .Y(n8659) );
  INVX1 U8097 ( .A(mem[310]), .Y(n9520) );
  INVX1 U8098 ( .A(mem[187]), .Y(n9643) );
  INVX1 U8099 ( .A(mem[967]), .Y(n8863) );
  INVX1 U8100 ( .A(mem[844]), .Y(n8986) );
  INVX1 U8101 ( .A(mem[1295]), .Y(n8535) );
  INVX1 U8102 ( .A(mem[1172]), .Y(n8658) );
  INVX1 U8103 ( .A(mem[311]), .Y(n9519) );
  INVX1 U8104 ( .A(mem[188]), .Y(n9642) );
  INVX1 U8105 ( .A(mem[968]), .Y(n8862) );
  INVX1 U8106 ( .A(mem[845]), .Y(n8985) );
  INVX1 U8107 ( .A(mem[1296]), .Y(n8534) );
  INVX1 U8108 ( .A(mem[1173]), .Y(n8657) );
  INVX1 U8109 ( .A(mem[312]), .Y(n9518) );
  INVX1 U8110 ( .A(mem[189]), .Y(n9641) );
  INVX1 U8111 ( .A(mem[969]), .Y(n8861) );
  INVX1 U8112 ( .A(mem[846]), .Y(n8984) );
  INVX1 U8113 ( .A(mem[1297]), .Y(n8533) );
  INVX1 U8114 ( .A(mem[1174]), .Y(n8656) );
  INVX1 U8115 ( .A(mem[313]), .Y(n9517) );
  INVX1 U8116 ( .A(mem[190]), .Y(n9640) );
  INVX1 U8117 ( .A(mem[970]), .Y(n8860) );
  INVX1 U8118 ( .A(mem[847]), .Y(n8983) );
  INVX1 U8119 ( .A(mem[1298]), .Y(n8532) );
  INVX1 U8120 ( .A(mem[1175]), .Y(n8655) );
  INVX1 U8121 ( .A(mem[314]), .Y(n9516) );
  INVX1 U8122 ( .A(mem[191]), .Y(n9639) );
  INVX1 U8123 ( .A(mem[971]), .Y(n8859) );
  INVX1 U8124 ( .A(mem[848]), .Y(n8982) );
  INVX1 U8125 ( .A(mem[1299]), .Y(n8531) );
  INVX1 U8126 ( .A(mem[1176]), .Y(n8654) );
  INVX1 U8127 ( .A(mem[315]), .Y(n9515) );
  INVX1 U8128 ( .A(mem[192]), .Y(n9638) );
  INVX1 U8129 ( .A(mem[972]), .Y(n8858) );
  INVX1 U8130 ( .A(mem[849]), .Y(n8981) );
  INVX1 U8131 ( .A(mem[1300]), .Y(n8530) );
  INVX1 U8132 ( .A(mem[1177]), .Y(n8653) );
  INVX1 U8133 ( .A(mem[316]), .Y(n9514) );
  INVX1 U8134 ( .A(mem[193]), .Y(n9637) );
  INVX1 U8135 ( .A(mem[973]), .Y(n8857) );
  INVX1 U8136 ( .A(mem[850]), .Y(n8980) );
  INVX1 U8137 ( .A(mem[1301]), .Y(n8529) );
  INVX1 U8138 ( .A(mem[1178]), .Y(n8652) );
  INVX1 U8139 ( .A(mem[317]), .Y(n9513) );
  INVX1 U8140 ( .A(mem[194]), .Y(n9636) );
  INVX1 U8141 ( .A(mem[974]), .Y(n8856) );
  INVX1 U8142 ( .A(mem[851]), .Y(n8979) );
  INVX1 U8143 ( .A(mem[1302]), .Y(n8528) );
  INVX1 U8144 ( .A(mem[1179]), .Y(n8651) );
  INVX1 U8145 ( .A(mem[318]), .Y(n9512) );
  INVX1 U8146 ( .A(mem[195]), .Y(n9635) );
  INVX1 U8147 ( .A(mem[975]), .Y(n8855) );
  INVX1 U8148 ( .A(mem[852]), .Y(n8978) );
  INVX1 U8149 ( .A(mem[1303]), .Y(n8527) );
  INVX1 U8150 ( .A(mem[1180]), .Y(n8650) );
  INVX1 U8151 ( .A(mem[319]), .Y(n9511) );
  INVX1 U8152 ( .A(mem[196]), .Y(n9634) );
  INVX1 U8153 ( .A(mem[976]), .Y(n8854) );
  INVX1 U8154 ( .A(mem[853]), .Y(n8977) );
  INVX1 U8155 ( .A(mem[1304]), .Y(n8526) );
  INVX1 U8156 ( .A(mem[1181]), .Y(n8649) );
  INVX1 U8157 ( .A(mem[320]), .Y(n9510) );
  INVX1 U8158 ( .A(mem[197]), .Y(n9633) );
  INVX1 U8159 ( .A(mem[977]), .Y(n8853) );
  INVX1 U8160 ( .A(mem[854]), .Y(n8976) );
  INVX1 U8161 ( .A(mem[1305]), .Y(n8525) );
  INVX1 U8162 ( .A(mem[1182]), .Y(n8648) );
  INVX1 U8163 ( .A(mem[321]), .Y(n9509) );
  INVX1 U8164 ( .A(mem[198]), .Y(n9632) );
  INVX1 U8165 ( .A(mem[978]), .Y(n8852) );
  INVX1 U8166 ( .A(mem[855]), .Y(n8975) );
  INVX1 U8167 ( .A(mem[1306]), .Y(n8524) );
  INVX1 U8168 ( .A(mem[1183]), .Y(n8647) );
  INVX1 U8169 ( .A(mem[322]), .Y(n9508) );
  INVX1 U8170 ( .A(mem[199]), .Y(n9631) );
  INVX1 U8171 ( .A(mem[979]), .Y(n8851) );
  INVX1 U8172 ( .A(mem[856]), .Y(n8974) );
  INVX1 U8173 ( .A(mem[1307]), .Y(n8523) );
  INVX1 U8174 ( .A(mem[1184]), .Y(n8646) );
  INVX1 U8175 ( .A(mem[323]), .Y(n9507) );
  INVX1 U8176 ( .A(mem[200]), .Y(n9630) );
  INVX1 U8177 ( .A(mem[980]), .Y(n8850) );
  INVX1 U8178 ( .A(mem[857]), .Y(n8973) );
  INVX1 U8179 ( .A(mem[1308]), .Y(n8522) );
  INVX1 U8180 ( .A(mem[1185]), .Y(n8645) );
  INVX1 U8181 ( .A(mem[324]), .Y(n9506) );
  INVX1 U8182 ( .A(mem[201]), .Y(n9629) );
  INVX1 U8183 ( .A(mem[981]), .Y(n8849) );
  INVX1 U8184 ( .A(mem[858]), .Y(n8972) );
  INVX1 U8185 ( .A(mem[1309]), .Y(n8521) );
  INVX1 U8186 ( .A(mem[1186]), .Y(n8644) );
  INVX1 U8187 ( .A(mem[325]), .Y(n9505) );
  INVX1 U8188 ( .A(mem[202]), .Y(n9628) );
  INVX1 U8189 ( .A(mem[982]), .Y(n8848) );
  INVX1 U8190 ( .A(mem[859]), .Y(n8971) );
  INVX1 U8191 ( .A(mem[1310]), .Y(n8520) );
  INVX1 U8192 ( .A(mem[1187]), .Y(n8643) );
  INVX1 U8193 ( .A(mem[326]), .Y(n9504) );
  INVX1 U8194 ( .A(mem[203]), .Y(n9627) );
  INVX1 U8195 ( .A(mem[983]), .Y(n8847) );
  INVX1 U8196 ( .A(mem[860]), .Y(n8970) );
  INVX1 U8197 ( .A(mem[1311]), .Y(n8519) );
  INVX1 U8198 ( .A(mem[1188]), .Y(n8642) );
  INVX1 U8199 ( .A(mem[327]), .Y(n9503) );
  INVX1 U8200 ( .A(mem[204]), .Y(n9626) );
  INVX1 U8201 ( .A(mem[615]), .Y(n9215) );
  INVX1 U8202 ( .A(mem[492]), .Y(n9338) );
  INVX1 U8203 ( .A(mem[616]), .Y(n9214) );
  INVX1 U8204 ( .A(mem[493]), .Y(n9337) );
  INVX1 U8205 ( .A(mem[617]), .Y(n9213) );
  INVX1 U8206 ( .A(mem[494]), .Y(n9336) );
  INVX1 U8207 ( .A(mem[618]), .Y(n9212) );
  INVX1 U8208 ( .A(mem[495]), .Y(n9335) );
  INVX1 U8209 ( .A(mem[619]), .Y(n9211) );
  INVX1 U8210 ( .A(mem[496]), .Y(n9334) );
  INVX1 U8211 ( .A(mem[620]), .Y(n9210) );
  INVX1 U8212 ( .A(mem[497]), .Y(n9333) );
  INVX1 U8213 ( .A(mem[621]), .Y(n9209) );
  INVX1 U8214 ( .A(mem[498]), .Y(n9332) );
  INVX1 U8215 ( .A(mem[622]), .Y(n9208) );
  INVX1 U8216 ( .A(mem[499]), .Y(n9331) );
  INVX1 U8217 ( .A(mem[623]), .Y(n9207) );
  INVX1 U8218 ( .A(mem[500]), .Y(n9330) );
  INVX1 U8219 ( .A(mem[624]), .Y(n9206) );
  INVX1 U8220 ( .A(mem[501]), .Y(n9329) );
  INVX1 U8221 ( .A(mem[625]), .Y(n9205) );
  INVX1 U8222 ( .A(mem[502]), .Y(n9328) );
  INVX1 U8223 ( .A(mem[626]), .Y(n9204) );
  INVX1 U8224 ( .A(mem[503]), .Y(n9327) );
  INVX1 U8225 ( .A(mem[627]), .Y(n9203) );
  INVX1 U8226 ( .A(mem[504]), .Y(n9326) );
  INVX1 U8227 ( .A(mem[628]), .Y(n9202) );
  INVX1 U8228 ( .A(mem[505]), .Y(n9325) );
  INVX1 U8229 ( .A(mem[629]), .Y(n9201) );
  INVX1 U8230 ( .A(mem[506]), .Y(n9324) );
  INVX1 U8231 ( .A(mem[630]), .Y(n9200) );
  INVX1 U8232 ( .A(mem[507]), .Y(n9323) );
  INVX1 U8233 ( .A(mem[631]), .Y(n9199) );
  INVX1 U8234 ( .A(mem[508]), .Y(n9322) );
  INVX1 U8235 ( .A(mem[632]), .Y(n9198) );
  INVX1 U8236 ( .A(mem[509]), .Y(n9321) );
  INVX1 U8237 ( .A(mem[633]), .Y(n9197) );
  INVX1 U8238 ( .A(mem[510]), .Y(n9320) );
  INVX1 U8239 ( .A(mem[634]), .Y(n9196) );
  INVX1 U8240 ( .A(mem[511]), .Y(n9319) );
  INVX1 U8241 ( .A(mem[635]), .Y(n9195) );
  INVX1 U8242 ( .A(mem[512]), .Y(n9318) );
  INVX1 U8243 ( .A(mem[636]), .Y(n9194) );
  INVX1 U8244 ( .A(mem[513]), .Y(n9317) );
  INVX1 U8245 ( .A(mem[637]), .Y(n9193) );
  INVX1 U8246 ( .A(mem[514]), .Y(n9316) );
  INVX1 U8247 ( .A(mem[638]), .Y(n9192) );
  INVX1 U8248 ( .A(mem[515]), .Y(n9315) );
  INVX1 U8249 ( .A(mem[639]), .Y(n9191) );
  INVX1 U8250 ( .A(mem[516]), .Y(n9314) );
  INVX1 U8251 ( .A(mem[640]), .Y(n9190) );
  INVX1 U8252 ( .A(mem[517]), .Y(n9313) );
  INVX1 U8253 ( .A(mem[641]), .Y(n9189) );
  INVX1 U8254 ( .A(mem[518]), .Y(n9312) );
  INVX1 U8255 ( .A(mem[642]), .Y(n9188) );
  INVX1 U8256 ( .A(mem[519]), .Y(n9311) );
  INVX1 U8257 ( .A(mem[643]), .Y(n9187) );
  INVX1 U8258 ( .A(mem[520]), .Y(n9310) );
  INVX1 U8259 ( .A(mem[644]), .Y(n9186) );
  INVX1 U8260 ( .A(mem[521]), .Y(n9309) );
  INVX1 U8261 ( .A(mem[645]), .Y(n9185) );
  INVX1 U8262 ( .A(mem[522]), .Y(n9308) );
  INVX1 U8263 ( .A(mem[646]), .Y(n9184) );
  INVX1 U8264 ( .A(mem[523]), .Y(n9307) );
  INVX1 U8265 ( .A(mem[647]), .Y(n9183) );
  INVX1 U8266 ( .A(mem[524]), .Y(n9306) );
  INVX1 U8267 ( .A(mem[648]), .Y(n9182) );
  INVX1 U8268 ( .A(mem[525]), .Y(n9305) );
  INVX1 U8269 ( .A(mem[649]), .Y(n9181) );
  INVX1 U8270 ( .A(mem[526]), .Y(n9304) );
  INVX1 U8271 ( .A(mem[650]), .Y(n9180) );
  INVX1 U8272 ( .A(mem[527]), .Y(n9303) );
  INVX1 U8273 ( .A(mem[651]), .Y(n9179) );
  INVX1 U8274 ( .A(mem[528]), .Y(n9302) );
  INVX1 U8275 ( .A(mem[652]), .Y(n9178) );
  INVX1 U8276 ( .A(mem[529]), .Y(n9301) );
  INVX1 U8277 ( .A(mem[653]), .Y(n9177) );
  INVX1 U8278 ( .A(mem[530]), .Y(n9300) );
  INVX1 U8279 ( .A(mem[654]), .Y(n9176) );
  INVX1 U8280 ( .A(mem[531]), .Y(n9299) );
  INVX1 U8281 ( .A(mem[655]), .Y(n9175) );
  INVX1 U8282 ( .A(mem[532]), .Y(n9298) );
  INVX1 U8283 ( .A(n5501), .Y(n8504) );
  INVX1 U8284 ( .A(n16), .Y(n8510) );
  AND2X1 U8285 ( .A(data_in[0]), .B(n8501), .Y(n4188) );
  AND2X1 U8286 ( .A(data_in[3]), .B(n8501), .Y(n4182) );
  AND2X1 U8287 ( .A(data_in[4]), .B(n8501), .Y(n4180) );
  AND2X1 U8288 ( .A(data_in[5]), .B(n8501), .Y(n4178) );
  AND2X1 U8289 ( .A(data_in[6]), .B(n8501), .Y(n4176) );
  AND2X1 U8290 ( .A(data_in[7]), .B(n8501), .Y(n4174) );
  AND2X1 U8291 ( .A(data_in[8]), .B(n8501), .Y(n4172) );
  AND2X1 U8292 ( .A(data_in[9]), .B(n8501), .Y(n4170) );
  AND2X1 U8293 ( .A(data_in[10]), .B(n8501), .Y(n4168) );
  AND2X1 U8294 ( .A(data_in[11]), .B(n8501), .Y(n4166) );
  AND2X1 U8295 ( .A(data_in[12]), .B(n8501), .Y(n4164) );
  AND2X1 U8296 ( .A(data_in[13]), .B(n8501), .Y(n4162) );
  AND2X1 U8297 ( .A(data_in[14]), .B(n8501), .Y(n4160) );
  AND2X1 U8298 ( .A(data_in[15]), .B(n8500), .Y(n4158) );
  AND2X1 U8299 ( .A(data_in[16]), .B(n8501), .Y(n4156) );
  AND2X1 U8300 ( .A(data_in[17]), .B(n8501), .Y(n4154) );
  AND2X1 U8301 ( .A(data_in[18]), .B(n8501), .Y(n4152) );
  AND2X1 U8302 ( .A(data_in[19]), .B(n8501), .Y(n4150) );
  AND2X1 U8303 ( .A(data_in[20]), .B(n8501), .Y(n4148) );
  AND2X1 U8304 ( .A(data_in[21]), .B(n8501), .Y(n4146) );
  AND2X1 U8305 ( .A(data_in[22]), .B(n8501), .Y(n4144) );
  AND2X1 U8306 ( .A(data_in[23]), .B(n8501), .Y(n4142) );
  AND2X1 U8307 ( .A(data_in[24]), .B(n8501), .Y(n4140) );
  AND2X1 U8308 ( .A(data_in[25]), .B(n8501), .Y(n4138) );
  AND2X1 U8309 ( .A(data_in[26]), .B(n8501), .Y(n4136) );
  AND2X1 U8310 ( .A(data_in[27]), .B(n8501), .Y(n4134) );
  AND2X1 U8311 ( .A(data_in[28]), .B(n8501), .Y(n4132) );
  AND2X1 U8312 ( .A(data_in[29]), .B(n8501), .Y(n4130) );
  AND2X1 U8313 ( .A(data_in[1]), .B(n8501), .Y(n4186) );
  AND2X1 U8314 ( .A(data_in[2]), .B(n8501), .Y(n4184) );
  AND2X1 U8315 ( .A(data_in[40]), .B(n8501), .Y(n4108) );
  AND2X1 U8316 ( .A(data_in[30]), .B(n8501), .Y(n4128) );
  AND2X1 U8317 ( .A(data_in[31]), .B(n8501), .Y(n4126) );
  AND2X1 U8318 ( .A(data_in[32]), .B(n8501), .Y(n4124) );
  AND2X1 U8319 ( .A(data_in[33]), .B(n8501), .Y(n4122) );
  AND2X1 U8320 ( .A(data_in[34]), .B(n8501), .Y(n4120) );
  AND2X1 U8321 ( .A(data_in[35]), .B(n8501), .Y(n4118) );
  AND2X1 U8322 ( .A(data_in[36]), .B(n8501), .Y(n4116) );
  AND2X1 U8323 ( .A(data_in[37]), .B(n8501), .Y(n4114) );
  AND2X1 U8324 ( .A(data_in[38]), .B(n8501), .Y(n4112) );
  AND2X1 U8325 ( .A(data_in[39]), .B(n8501), .Y(n4110) );
endmodule


module ddr3_init_engine_DW01_inc_0 ( A, SUM );
  input [18:0] A;
  output [18:0] SUM;

  wire   [18:2] carry;

  HAX1 U1_1_17 ( .A(A[17]), .B(carry[17]), .YC(carry[18]), .YS(SUM[17]) );
  HAX1 U1_1_16 ( .A(A[16]), .B(carry[16]), .YC(carry[17]), .YS(SUM[16]) );
  HAX1 U1_1_15 ( .A(A[15]), .B(carry[15]), .YC(carry[16]), .YS(SUM[15]) );
  HAX1 U1_1_14 ( .A(A[14]), .B(carry[14]), .YC(carry[15]), .YS(SUM[14]) );
  HAX1 U1_1_13 ( .A(A[13]), .B(carry[13]), .YC(carry[14]), .YS(SUM[13]) );
  HAX1 U1_1_12 ( .A(A[12]), .B(carry[12]), .YC(carry[13]), .YS(SUM[12]) );
  HAX1 U1_1_11 ( .A(A[11]), .B(carry[11]), .YC(carry[12]), .YS(SUM[11]) );
  HAX1 U1_1_10 ( .A(A[10]), .B(carry[10]), .YC(carry[11]), .YS(SUM[10]) );
  HAX1 U1_1_9 ( .A(A[9]), .B(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  HAX1 U1_1_8 ( .A(A[8]), .B(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  HAX1 U1_1_7 ( .A(A[7]), .B(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  HAX1 U1_1_6 ( .A(A[6]), .B(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  HAX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry[2]), .YS(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[18]), .B(A[18]), .Y(SUM[18]) );
endmodule


module ddr3_init_engine ( ready, csbar, rasbar, casbar, webar, ba, a, odt, 
        ts_con, cke, clk, resetbar, init, ck, Port15 );
  output [2:0] ba;
  output [13:0] a;
  input clk, resetbar, init, ck;
  output ready, csbar, rasbar, casbar, webar, odt, ts_con, cke;
  inout Port15;
  wire   flag, RESET, INIT, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n216, n55, n56, n57, n58,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n59,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262;
  wire   [18:0] counter;
  assign ba[2] = 1'b0;
  assign a[13] = 1'b0;
  assign a[12] = 1'b0;
  assign a[11] = 1'b0;
  assign a[9] = 1'b0;
  assign a[7] = 1'b0;
  assign a[6] = 1'b0;
  assign a[5] = 1'b0;
  assign a[3] = 1'b0;
  assign a[2] = 1'b0;
  assign a[1] = 1'b0;
  assign a[0] = 1'b0;
  assign odt = 1'b0;
  assign ts_con = 1'b0;

  DFFPOSX1 RESET_reg ( .D(resetbar), .CLK(clk), .Q(RESET) );
  DFFPOSX1 INIT_reg ( .D(init), .CLK(clk), .Q(INIT) );
  DFFPOSX1 flag_reg ( .D(n229), .CLK(clk), .Q(flag) );
  DFFPOSX1 counter_reg_0_ ( .D(n182), .CLK(clk), .Q(counter[0]) );
  DFFPOSX1 counter_reg_1_ ( .D(n181), .CLK(clk), .Q(counter[1]) );
  DFFPOSX1 counter_reg_2_ ( .D(n180), .CLK(clk), .Q(counter[2]) );
  DFFPOSX1 counter_reg_3_ ( .D(n179), .CLK(clk), .Q(counter[3]) );
  DFFPOSX1 counter_reg_4_ ( .D(n178), .CLK(clk), .Q(counter[4]) );
  DFFPOSX1 counter_reg_5_ ( .D(n177), .CLK(clk), .Q(counter[5]) );
  DFFPOSX1 counter_reg_6_ ( .D(n176), .CLK(clk), .Q(counter[6]) );
  DFFPOSX1 counter_reg_7_ ( .D(n175), .CLK(clk), .Q(counter[7]) );
  DFFPOSX1 counter_reg_8_ ( .D(n174), .CLK(clk), .Q(counter[8]) );
  DFFPOSX1 counter_reg_9_ ( .D(n173), .CLK(clk), .Q(counter[9]) );
  DFFPOSX1 counter_reg_10_ ( .D(n172), .CLK(clk), .Q(counter[10]) );
  DFFPOSX1 counter_reg_11_ ( .D(n171), .CLK(clk), .Q(counter[11]) );
  DFFPOSX1 counter_reg_12_ ( .D(n170), .CLK(clk), .Q(counter[12]) );
  DFFPOSX1 counter_reg_13_ ( .D(n169), .CLK(clk), .Q(counter[13]) );
  DFFPOSX1 counter_reg_14_ ( .D(n168), .CLK(clk), .Q(counter[14]) );
  DFFPOSX1 counter_reg_15_ ( .D(n167), .CLK(clk), .Q(counter[15]) );
  DFFPOSX1 counter_reg_16_ ( .D(n166), .CLK(clk), .Q(counter[16]) );
  DFFPOSX1 counter_reg_17_ ( .D(n165), .CLK(clk), .Q(counter[17]) );
  DFFPOSX1 counter_reg_18_ ( .D(n164), .CLK(clk), .Q(counter[18]) );
  DFFPOSX1 ready_reg ( .D(n163), .CLK(clk), .Q(ready) );
  DFFPOSX1 casbar_reg ( .D(n159), .CLK(clk), .Q(casbar) );
  DFFPOSX1 csbar_reg ( .D(n3), .CLK(clk), .Q(csbar) );
  DFFPOSX1 webar_reg ( .D(n161), .CLK(clk), .Q(webar) );
  DFFPOSX1 rasbar_reg ( .D(n4), .CLK(clk), .Q(rasbar) );
  DFFPOSX1 cke_reg ( .D(n158), .CLK(clk), .Q(cke) );
  DFFPOSX1 a_reg_10_ ( .D(n157), .CLK(clk), .Q(a[10]) );
  DFFPOSX1 a_reg_8_ ( .D(n190), .CLK(clk), .Q(a[8]) );
  DFFPOSX1 a_reg_4_ ( .D(n2), .CLK(clk), .Q(a[4]) );
  DFFPOSX1 ba_reg_1_ ( .D(n154), .CLK(clk), .Q(ba[1]) );
  DFFPOSX1 ba_reg_0_ ( .D(n153), .CLK(clk), .Q(ba[0]) );
  OAI21X1 U63 ( .A(n55), .B(n205), .C(n185), .Y(n153) );
  AOI21X1 U66 ( .A(n192), .B(n197), .C(n205), .Y(n60) );
  NAND3X1 U68 ( .A(n63), .B(n64), .C(n42), .Y(n155) );
  OAI21X1 U73 ( .A(n226), .B(n236), .C(n9), .Y(n157) );
  AOI21X1 U75 ( .A(n193), .B(n199), .C(n237), .Y(n71) );
  OAI21X1 U76 ( .A(n211), .B(n193), .C(n220), .Y(n73) );
  OAI21X1 U77 ( .A(n75), .B(n226), .C(n8), .Y(n158) );
  NAND3X1 U79 ( .A(n47), .B(n74), .C(n79), .Y(n77) );
  OAI21X1 U80 ( .A(n240), .B(n48), .C(n7), .Y(n159) );
  OAI21X1 U84 ( .A(n226), .B(n84), .C(n6), .Y(n161) );
  OAI21X1 U86 ( .A(n36), .B(n37), .C(n210), .Y(n84) );
  NAND3X1 U87 ( .A(n198), .B(n45), .C(n204), .Y(n87) );
  NAND3X1 U88 ( .A(n223), .B(n46), .C(n94), .Y(n86) );
  NAND3X1 U91 ( .A(n210), .B(n98), .C(n69), .Y(n82) );
  NAND3X1 U94 ( .A(n240), .B(n199), .C(n100), .Y(n99) );
  NAND3X1 U95 ( .A(n103), .B(n223), .C(n215), .Y(n102) );
  NAND3X1 U96 ( .A(counter[2]), .B(n241), .C(n247), .Y(n96) );
  NAND3X1 U98 ( .A(n112), .B(n217), .C(counter[9]), .Y(n72) );
  NAND3X1 U99 ( .A(n47), .B(counter[1]), .C(n41), .Y(n93) );
  NAND3X1 U102 ( .A(counter[7]), .B(n225), .C(counter[5]), .Y(n107) );
  NAND3X1 U103 ( .A(n252), .B(n253), .C(n250), .Y(n106) );
  NAND3X1 U104 ( .A(n109), .B(n198), .C(n204), .Y(n101) );
  NAND3X1 U105 ( .A(n224), .B(n217), .C(counter[9]), .Y(n89) );
  NAND3X1 U107 ( .A(n225), .B(n246), .C(n40), .Y(n90) );
  OAI21X1 U109 ( .A(n234), .B(n226), .C(n196), .Y(n163) );
  OAI21X1 U111 ( .A(n211), .B(n204), .C(RESET), .Y(n115) );
  NAND3X1 U112 ( .A(n116), .B(n112), .C(counter[12]), .Y(n91) );
  OAI21X1 U113 ( .A(n229), .B(n262), .C(n222), .Y(n164) );
  OAI21X1 U115 ( .A(n230), .B(n261), .C(n213), .Y(n165) );
  OAI21X1 U117 ( .A(n230), .B(n260), .C(n202), .Y(n166) );
  OAI21X1 U119 ( .A(n230), .B(n259), .C(n207), .Y(n167) );
  OAI21X1 U121 ( .A(n229), .B(n258), .C(n195), .Y(n168) );
  OAI21X1 U123 ( .A(n229), .B(n257), .C(n189), .Y(n169) );
  OAI21X1 U125 ( .A(n230), .B(n256), .C(n54), .Y(n170) );
  OAI21X1 U127 ( .A(n229), .B(n255), .C(n184), .Y(n171) );
  OAI21X1 U129 ( .A(n230), .B(n254), .C(n52), .Y(n172) );
  OAI21X1 U131 ( .A(n230), .B(n253), .C(n221), .Y(n173) );
  OAI21X1 U133 ( .A(n229), .B(n252), .C(n201), .Y(n174) );
  OAI21X1 U135 ( .A(n229), .B(n251), .C(n194), .Y(n175) );
  OAI21X1 U137 ( .A(n230), .B(n250), .C(n188), .Y(n176) );
  OAI21X1 U139 ( .A(n229), .B(n249), .C(n59), .Y(n177) );
  OAI21X1 U141 ( .A(n229), .B(n248), .C(n51), .Y(n178) );
  OAI21X1 U143 ( .A(n230), .B(n246), .C(n50), .Y(n179) );
  OAI21X1 U145 ( .A(n230), .B(n243), .C(n49), .Y(n180) );
  OAI21X1 U147 ( .A(n229), .B(n241), .C(n206), .Y(n181) );
  OAI21X1 U149 ( .A(n230), .B(n239), .C(n53), .Y(n182) );
  OAI21X1 U151 ( .A(n233), .B(n214), .C(n226), .Y(n183) );
  AOI21X1 U153 ( .A(n74), .B(n242), .C(n216), .Y(n58) );
  NAND3X1 U154 ( .A(n116), .B(counter[1]), .C(n200), .Y(n68) );
  NOR3X1 U156 ( .A(n246), .B(counter[4]), .C(n209), .Y(n116) );
  NAND3X1 U157 ( .A(counter[9]), .B(counter[6]), .C(n139), .Y(n113) );
  NOR3X1 U158 ( .A(counter[5]), .B(counter[8]), .C(counter[7]), .Y(n139) );
  OAI21X1 U159 ( .A(n100), .B(n211), .C(RESET), .Y(n216) );
  NOR3X1 U161 ( .A(n212), .B(counter[11]), .C(counter[0]), .Y(n141) );
  NAND3X1 U162 ( .A(n260), .B(n261), .C(n257), .Y(n142) );
  NOR3X1 U163 ( .A(n203), .B(n262), .C(n226), .Y(n140) );
  NAND3X1 U165 ( .A(counter[14]), .B(counter[10]), .C(counter[15]), .Y(n143)
         );
  NAND3X1 U167 ( .A(n217), .B(n253), .C(counter[2]), .Y(n144) );
  NAND3X1 U169 ( .A(counter[3]), .B(n225), .C(counter[8]), .Y(n146) );
  NAND3X1 U171 ( .A(n250), .B(n251), .C(n249), .Y(n145) );
  NAND3X1 U173 ( .A(counter[6]), .B(counter[5]), .C(n39), .Y(n147) );
  NAND3X1 U178 ( .A(n249), .B(n250), .C(n38), .Y(n150) );
  NAND3X1 U180 ( .A(counter[7]), .B(counter[8]), .C(n152), .Y(n149) );
  NOR3X1 U181 ( .A(counter[12]), .B(counter[9]), .C(counter[4]), .Y(n152) );
  ddr3_init_engine_DW01_inc_0 add_79 ( .A(counter), .SUM({n28, n27, n26, n25, 
        n24, n23, n22, n21, n20, n19, n18, n17, n16, n15, n14, n13, n12, n11, 
        n10}) );
  OR2X1 U17 ( .A(n31), .B(n34), .Y(n98) );
  AND2X1 U18 ( .A(n55), .B(n197), .Y(n100) );
  AND2X1 U19 ( .A(n192), .B(n43), .Y(n55) );
  AND2X1 U20 ( .A(n45), .B(n208), .Y(n109) );
  AND2X1 U21 ( .A(n46), .B(n193), .Y(n103) );
  OR2X1 U22 ( .A(n218), .B(n219), .Y(n104) );
  OR2X1 U23 ( .A(n32), .B(n33), .Y(n78) );
  AND2X1 U24 ( .A(n183), .B(n214), .Y(n118) );
  AND2X1 U25 ( .A(n208), .B(n215), .Y(n94) );
  AND2X1 U26 ( .A(n74), .B(n5), .Y(n80) );
  AND2X1 U27 ( .A(ba[1]), .B(n220), .Y(n227) );
  OR2X1 U28 ( .A(n43), .B(n205), .Y(n63) );
  AND2X1 U29 ( .A(n64), .B(n191), .Y(n156) );
  AND2X1 U30 ( .A(n1), .B(RESET), .Y(n75) );
  AND2X1 U31 ( .A(n48), .B(RESET), .Y(n88) );
  BUFX2 U32 ( .A(n77), .Y(n1) );
  BUFX2 U33 ( .A(n155), .Y(n2) );
  AND2X1 U34 ( .A(n44), .B(n29), .Y(n162) );
  INVX1 U35 ( .A(n162), .Y(n3) );
  AND2X1 U36 ( .A(n44), .B(n30), .Y(n160) );
  INVX1 U37 ( .A(n160), .Y(n4) );
  BUFX2 U38 ( .A(n99), .Y(n5) );
  AND2X1 U39 ( .A(webar), .B(n88), .Y(n85) );
  INVX1 U40 ( .A(n85), .Y(n6) );
  AND2X1 U41 ( .A(casbar), .B(n48), .Y(n81) );
  INVX1 U42 ( .A(n81), .Y(n7) );
  AND2X1 U43 ( .A(cke), .B(n75), .Y(n76) );
  INVX1 U44 ( .A(n76), .Y(n8) );
  AND2X1 U45 ( .A(a[10]), .B(n237), .Y(n70) );
  INVX1 U46 ( .A(n70), .Y(n9) );
  AND2X1 U47 ( .A(csbar), .B(n88), .Y(n97) );
  INVX1 U48 ( .A(n97), .Y(n29) );
  AND2X1 U49 ( .A(rasbar), .B(n88), .Y(n83) );
  INVX1 U50 ( .A(n83), .Y(n30) );
  BUFX2 U51 ( .A(n101), .Y(n31) );
  BUFX2 U52 ( .A(n106), .Y(n32) );
  BUFX2 U53 ( .A(n107), .Y(n33) );
  BUFX2 U54 ( .A(n102), .Y(n34) );
  BUFX2 U55 ( .A(n60), .Y(n35) );
  BUFX2 U56 ( .A(n86), .Y(n36) );
  BUFX2 U57 ( .A(n87), .Y(n37) );
  OR2X1 U58 ( .A(counter[3]), .B(n187), .Y(n151) );
  INVX1 U59 ( .A(n151), .Y(n38) );
  OR2X1 U60 ( .A(n246), .B(n187), .Y(n148) );
  INVX1 U61 ( .A(n148), .Y(n39) );
  OR2X1 U62 ( .A(n186), .B(n209), .Y(n111) );
  INVX1 U64 ( .A(n111), .Y(n40) );
  OR2X1 U65 ( .A(counter[3]), .B(n243), .Y(n105) );
  INVX1 U67 ( .A(n105), .Y(n41) );
  AND2X1 U69 ( .A(a[4]), .B(n220), .Y(n65) );
  INVX1 U70 ( .A(n65), .Y(n42) );
  AND2X1 U71 ( .A(n112), .B(n245), .Y(n66) );
  INVX1 U72 ( .A(n66), .Y(n43) );
  BUFX2 U74 ( .A(n82), .Y(n44) );
  BUFX2 U78 ( .A(n90), .Y(n45) );
  BUFX2 U81 ( .A(n93), .Y(n46) );
  INVX1 U82 ( .A(n78), .Y(n47) );
  INVX1 U83 ( .A(n80), .Y(n48) );
  AND2X1 U85 ( .A(n12), .B(n231), .Y(n134) );
  INVX1 U89 ( .A(n134), .Y(n49) );
  AND2X1 U90 ( .A(n13), .B(n231), .Y(n133) );
  INVX1 U92 ( .A(n133), .Y(n50) );
  AND2X1 U93 ( .A(n14), .B(n231), .Y(n132) );
  INVX1 U97 ( .A(n132), .Y(n51) );
  AND2X1 U100 ( .A(n20), .B(n232), .Y(n126) );
  INVX1 U101 ( .A(n126), .Y(n52) );
  AND2X1 U106 ( .A(n10), .B(n231), .Y(n136) );
  INVX1 U108 ( .A(n136), .Y(n53) );
  AND2X1 U110 ( .A(n22), .B(n232), .Y(n124) );
  INVX1 U114 ( .A(n124), .Y(n54) );
  AND2X1 U116 ( .A(n15), .B(n231), .Y(n131) );
  INVX1 U118 ( .A(n131), .Y(n59) );
  AND2X1 U120 ( .A(n21), .B(n232), .Y(n125) );
  INVX1 U122 ( .A(n125), .Y(n184) );
  AND2X1 U124 ( .A(ba[0]), .B(n220), .Y(n57) );
  INVX1 U126 ( .A(n57), .Y(n185) );
  AND2X1 U128 ( .A(n243), .B(n241), .Y(n112) );
  INVX1 U130 ( .A(n112), .Y(n186) );
  BUFX2 U132 ( .A(n149), .Y(n187) );
  AND2X1 U134 ( .A(n16), .B(n231), .Y(n130) );
  INVX1 U136 ( .A(n130), .Y(n188) );
  AND2X1 U138 ( .A(n23), .B(n232), .Y(n123) );
  INVX1 U140 ( .A(n123), .Y(n189) );
  INVX1 U142 ( .A(n156), .Y(n190) );
  AND2X1 U144 ( .A(a[8]), .B(n220), .Y(n67) );
  INVX1 U146 ( .A(n67), .Y(n191) );
  OR2X1 U148 ( .A(n205), .B(n199), .Y(n64) );
  AND2X1 U150 ( .A(n247), .B(n224), .Y(n61) );
  INVX1 U152 ( .A(n61), .Y(n192) );
  BUFX2 U155 ( .A(n72), .Y(n193) );
  AND2X1 U160 ( .A(n17), .B(n231), .Y(n129) );
  INVX1 U164 ( .A(n129), .Y(n194) );
  AND2X1 U166 ( .A(n24), .B(n232), .Y(n122) );
  INVX1 U168 ( .A(n122), .Y(n195) );
  AND2X1 U170 ( .A(ready), .B(n234), .Y(n114) );
  INVX1 U172 ( .A(n114), .Y(n196) );
  AND2X1 U174 ( .A(n244), .B(n241), .Y(n62) );
  INVX1 U175 ( .A(n62), .Y(n197) );
  BUFX2 U176 ( .A(n89), .Y(n198) );
  BUFX2 U177 ( .A(n68), .Y(n199) );
  OR2X1 U179 ( .A(counter[12]), .B(n243), .Y(n138) );
  INVX1 U182 ( .A(n138), .Y(n200) );
  AND2X1 U183 ( .A(n18), .B(n231), .Y(n128) );
  INVX1 U184 ( .A(n128), .Y(n201) );
  AND2X1 U185 ( .A(n26), .B(n232), .Y(n120) );
  INVX1 U186 ( .A(n120), .Y(n202) );
  BUFX2 U187 ( .A(n143), .Y(n203) );
  BUFX2 U188 ( .A(n91), .Y(n204) );
  AND2X1 U189 ( .A(n69), .B(n235), .Y(n56) );
  INVX1 U190 ( .A(n56), .Y(n205) );
  AND2X1 U191 ( .A(n11), .B(n231), .Y(n135) );
  INVX1 U192 ( .A(n135), .Y(n206) );
  AND2X1 U193 ( .A(n25), .B(n232), .Y(n121) );
  INVX1 U194 ( .A(n121), .Y(n207) );
  AND2X1 U195 ( .A(n224), .B(n245), .Y(n95) );
  INVX1 U196 ( .A(n95), .Y(n208) );
  BUFX2 U197 ( .A(n113), .Y(n209) );
  INVX1 U198 ( .A(n88), .Y(n210) );
  AND2X1 U199 ( .A(n140), .B(n141), .Y(n74) );
  INVX1 U200 ( .A(n74), .Y(n211) );
  BUFX2 U201 ( .A(n142), .Y(n212) );
  AND2X1 U202 ( .A(n27), .B(n232), .Y(n119) );
  INVX1 U203 ( .A(n119), .Y(n213) );
  AND2X1 U204 ( .A(INIT), .B(n238), .Y(n137) );
  INVX1 U205 ( .A(n137), .Y(n214) );
  BUFX2 U206 ( .A(n96), .Y(n215) );
  INVX1 U207 ( .A(n104), .Y(n217) );
  BUFX2 U208 ( .A(n145), .Y(n218) );
  BUFX2 U209 ( .A(n146), .Y(n219) );
  BUFX2 U210 ( .A(n58), .Y(n220) );
  AND2X1 U211 ( .A(n19), .B(n231), .Y(n127) );
  INVX1 U212 ( .A(n127), .Y(n221) );
  AND2X1 U213 ( .A(n28), .B(n232), .Y(n117) );
  INVX1 U214 ( .A(n117), .Y(n222) );
  AND2X1 U215 ( .A(counter[1]), .B(n244), .Y(n92) );
  INVX1 U216 ( .A(n92), .Y(n223) );
  OR2X1 U217 ( .A(n241), .B(counter[2]), .Y(n110) );
  INVX1 U218 ( .A(n110), .Y(n224) );
  OR2X1 U219 ( .A(n248), .B(counter[12]), .Y(n108) );
  INVX1 U220 ( .A(n108), .Y(n225) );
  AND2X1 U221 ( .A(flag), .B(RESET), .Y(n69) );
  INVX1 U222 ( .A(n69), .Y(n226) );
  BUFX2 U223 ( .A(n118), .Y(n231) );
  BUFX2 U224 ( .A(n118), .Y(n232) );
  INVX1 U225 ( .A(n98), .Y(n240) );
  INVX1 U226 ( .A(n220), .Y(n235) );
  INVX1 U227 ( .A(n73), .Y(n237) );
  INVX1 U228 ( .A(n199), .Y(n242) );
  INVX1 U229 ( .A(RESET), .Y(n233) );
  INVX1 U230 ( .A(flag), .Y(n238) );
  INVX1 U231 ( .A(n115), .Y(n234) );
  INVX1 U232 ( .A(counter[14]), .Y(n258) );
  INVX1 U233 ( .A(counter[15]), .Y(n259) );
  INVX1 U234 ( .A(counter[12]), .Y(n256) );
  INVX1 U235 ( .A(counter[11]), .Y(n255) );
  INVX1 U236 ( .A(counter[10]), .Y(n254) );
  INVX1 U237 ( .A(counter[0]), .Y(n239) );
  INVX1 U238 ( .A(n71), .Y(n236) );
  OR2X1 U239 ( .A(n227), .B(n35), .Y(n154) );
  INVX1 U240 ( .A(counter[1]), .Y(n241) );
  INVX1 U241 ( .A(counter[3]), .Y(n246) );
  INVX1 U242 ( .A(counter[6]), .Y(n250) );
  INVX1 U243 ( .A(counter[9]), .Y(n253) );
  INVX1 U244 ( .A(counter[2]), .Y(n243) );
  INVX1 U245 ( .A(counter[5]), .Y(n249) );
  INVX1 U246 ( .A(counter[8]), .Y(n252) );
  INVX1 U247 ( .A(counter[7]), .Y(n251) );
  INVX1 U248 ( .A(n150), .Y(n247) );
  INVX1 U249 ( .A(counter[4]), .Y(n248) );
  INVX1 U250 ( .A(n144), .Y(n244) );
  INVX1 U251 ( .A(n147), .Y(n245) );
  INVX1 U252 ( .A(counter[18]), .Y(n262) );
  AND2X1 U253 ( .A(n112), .B(counter[3]), .Y(n79) );
  INVX1 U254 ( .A(counter[13]), .Y(n257) );
  INVX1 U255 ( .A(counter[17]), .Y(n261) );
  INVX1 U256 ( .A(counter[16]), .Y(n260) );
  INVX1 U257 ( .A(n183), .Y(n228) );
  INVX1 U258 ( .A(n228), .Y(n229) );
  INVX1 U259 ( .A(n228), .Y(n230) );
endmodule


module SSTL18DDR3DIFF ( PAD, PADN, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD,  PADN;
  wire   n4, n5, n7;

  TBUFX2 b2 ( .A(A), .EN(TS), .Y(PADN) );
  TBUFX2 b1 ( .A(n7), .EN(TS), .Y(PAD) );
  NAND3X1 U4 ( .A(PAD), .B(n5), .C(RI), .Y(n4) );
  INVX1 U1 ( .A(n4), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n7) );
  INVX1 U3 ( .A(PADN), .Y(n5) );
endmodule


module SSTL18DDR3INTERFACE ( ck_pad, ckbar_pad, cke_pad, csbar_pad, rasbar_pad, 
        casbar_pad, webar_pad, ba_pad, a_pad, dm_pad, odt_pad, resetbar_pad, 
        dq_o, dqs_o, dqsbar_o, dq_pad, dqs_pad, dqsbar_pad, ri_i, ts_i, ck_i, 
        cke_i, csbar_i, rasbar_i, casbar_i, webar_i, ba_i, a_i, dq_i, dqs_i, 
        dqsbar_i, dm_i, odt_i, resetbar_i );
  output [2:0] ba_pad;
  output [13:0] a_pad;
  output [1:0] dm_pad;
  output [15:0] dq_o;
  output [1:0] dqs_o;
  output [1:0] dqsbar_o;
  inout [15:0] dq_pad;
  inout [1:0] dqs_pad;
  inout [1:0] dqsbar_pad;
  input [2:0] ba_i;
  input [13:0] a_i;
  input [15:0] dq_i;
  input [1:0] dqs_i;
  input [1:0] dqsbar_i;
  input [1:0] dm_i;
  input ri_i, ts_i, ck_i, cke_i, csbar_i, rasbar_i, casbar_i, webar_i, odt_i,
         resetbar_i;
  output ck_pad, ckbar_pad, cke_pad, csbar_pad, rasbar_pad, casbar_pad,
         webar_pad, odt_pad, resetbar_pad;


  SSTL18DDR3DIFF ck_sstl ( .PAD(ck_pad), .PADN(ckbar_pad), .Z(), .A(ck_i), 
        .RI(1'b0), .TS(1'b1) );
  SSTL18DDR3_45 cke_sstl ( .PAD(cke_pad), .Z(), .A(cke_i), .RI(1'b0), .TS(1'b1) );
  SSTL18DDR3_44 casbar_sstl ( .PAD(casbar_pad), .Z(), .A(casbar_i), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_43 rasbar_sstl ( .PAD(rasbar_pad), .Z(), .A(rasbar_i), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_42 csbar_sstl ( .PAD(csbar_pad), .Z(), .A(csbar_i), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_41 webar_sstl ( .PAD(webar_pad), .Z(), .A(webar_i), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_40 odt_sstl ( .PAD(odt_pad), .Z(), .A(odt_i), .RI(1'b0), .TS(1'b1) );
  SSTL18DDR3_39 resetbar_sstl ( .PAD(resetbar_pad), .Z(), .A(resetbar_i), .RI(
        1'b0), .TS(1'b1) );
  SSTL18DDR3_38 BA_0__sstl_ba ( .PAD(ba_pad[0]), .Z(), .A(ba_i[0]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_37 BA_1__sstl_ba ( .PAD(ba_pad[1]), .Z(), .A(ba_i[1]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_36 BA_2__sstl_ba ( .PAD(ba_pad[2]), .Z(), .A(ba_i[2]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_35 A_0__sstl_a ( .PAD(a_pad[0]), .Z(), .A(a_i[0]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_34 A_1__sstl_a ( .PAD(a_pad[1]), .Z(), .A(a_i[1]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_33 A_2__sstl_a ( .PAD(a_pad[2]), .Z(), .A(a_i[2]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_32 A_3__sstl_a ( .PAD(a_pad[3]), .Z(), .A(a_i[3]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_31 A_4__sstl_a ( .PAD(a_pad[4]), .Z(), .A(a_i[4]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_30 A_5__sstl_a ( .PAD(a_pad[5]), .Z(), .A(a_i[5]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_29 A_6__sstl_a ( .PAD(a_pad[6]), .Z(), .A(a_i[6]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_28 A_7__sstl_a ( .PAD(a_pad[7]), .Z(), .A(a_i[7]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_27 A_8__sstl_a ( .PAD(a_pad[8]), .Z(), .A(a_i[8]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_26 A_9__sstl_a ( .PAD(a_pad[9]), .Z(), .A(a_i[9]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_25 A_10__sstl_a ( .PAD(a_pad[10]), .Z(), .A(a_i[10]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_24 A_11__sstl_a ( .PAD(a_pad[11]), .Z(), .A(a_i[11]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_23 A_12__sstl_a ( .PAD(a_pad[12]), .Z(), .A(a_i[12]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_22 A_13__sstl_a ( .PAD(a_pad[13]), .Z(), .A(a_i[13]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_21 DQ_0__sstl_dq ( .PAD(dq_pad[0]), .Z(dq_o[0]), .A(dq_i[0]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_20 DQ_1__sstl_dq ( .PAD(dq_pad[1]), .Z(dq_o[1]), .A(dq_i[1]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_19 DQ_2__sstl_dq ( .PAD(dq_pad[2]), .Z(dq_o[2]), .A(dq_i[2]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_18 DQ_3__sstl_dq ( .PAD(dq_pad[3]), .Z(dq_o[3]), .A(dq_i[3]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_17 DQ_4__sstl_dq ( .PAD(dq_pad[4]), .Z(dq_o[4]), .A(dq_i[4]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_16 DQ_5__sstl_dq ( .PAD(dq_pad[5]), .Z(dq_o[5]), .A(dq_i[5]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_15 DQ_6__sstl_dq ( .PAD(dq_pad[6]), .Z(dq_o[6]), .A(dq_i[6]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_14 DQ_7__sstl_dq ( .PAD(dq_pad[7]), .Z(dq_o[7]), .A(dq_i[7]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_13 DQ_8__sstl_dq ( .PAD(dq_pad[8]), .Z(dq_o[8]), .A(dq_i[8]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_12 DQ_9__sstl_dq ( .PAD(dq_pad[9]), .Z(dq_o[9]), .A(dq_i[9]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_11 DQ_10__sstl_dq ( .PAD(dq_pad[10]), .Z(dq_o[10]), .A(dq_i[10]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_10 DQ_11__sstl_dq ( .PAD(dq_pad[11]), .Z(dq_o[11]), .A(dq_i[11]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_9 DQ_12__sstl_dq ( .PAD(dq_pad[12]), .Z(dq_o[12]), .A(dq_i[12]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_8 DQ_13__sstl_dq ( .PAD(dq_pad[13]), .Z(dq_o[13]), .A(dq_i[13]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_7 DQ_14__sstl_dq ( .PAD(dq_pad[14]), .Z(dq_o[14]), .A(dq_i[14]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_6 DQ_15__sstl_dq ( .PAD(dq_pad[15]), .Z(dq_o[15]), .A(dq_i[15]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_5 DQS_0__sstl_dqs ( .PAD(dqs_pad[0]), .Z(dqs_o[0]), .A(dqs_i[0]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_4 DQS_1__sstl_dqs ( .PAD(dqs_pad[1]), .Z(dqs_o[1]), .A(dqs_i[1]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_3 DQSBAR_0__sstl_dqsbar ( .PAD(dqsbar_pad[0]), .Z(dqsbar_o[0]), 
        .A(dqsbar_i[0]), .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_2 DQSBAR_1__sstl_dqsbar ( .PAD(dqsbar_pad[1]), .Z(dqsbar_o[1]), 
        .A(dqsbar_i[1]), .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_1 DM_0__sstl_dm ( .PAD(dm_pad[0]), .Z(), .A(dm_i[0]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_0 DM_1__sstl_dm ( .PAD(dm_pad[1]), .Z(), .A(dm_i[1]), .RI(1'b0), 
        .TS(1'b1) );
endmodule


module ddr3_controller ( dout, raddr, fillcount, notfull, ready, ck_pad, 
        ckbar_pad, cke_pad, csbar_pad, rasbar_pad, casbar_pad, webar_pad, 
        ba_pad, a_pad, dm_pad, odt_pad, notempty, resetbar_pad, dq_pad, 
        dqs_pad, dqsbar_pad, clk, resetbar, read, cmd, din, addr, initddr );
  output [15:0] dout;
  output [24:0] raddr;
  output [5:0] fillcount;
  output [2:0] ba_pad;
  output [13:0] a_pad;
  output [1:0] dm_pad;
  inout [15:0] dq_pad;
  inout [1:0] dqs_pad;
  inout [1:0] dqsbar_pad;
  input [2:0] cmd;
  input [15:0] din;
  input [24:0] addr;
  input clk, resetbar, read, initddr;
  output notfull, ready, ck_pad, ckbar_pad, cke_pad, csbar_pad, rasbar_pad,
         casbar_pad, webar_pad, odt_pad, notempty, resetbar_pad;
  wire   ck_i, n6, init_csbar, init_rasbar, init_casbar, init_webar, init_cke,
         csbar_i, rasbar_i, casbar_i, webar_i, n3, n4, n7,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26,
         SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28,
         SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30,
         SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32,
         SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34,
         SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36,
         SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38,
         SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40,
         SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42,
         SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44,
         SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46,
         SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48,
         SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50,
         SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52,
         SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54,
         SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56,
         SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58,
         SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60,
         SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62,
         SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64,
         SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66,
         SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68,
         SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70,
         SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72,
         SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74,
         SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76,
         SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78,
         SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_80,
         SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82,
         SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84,
         SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86,
         SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88,
         SYNOPSYS_UNCONNECTED_89, SYNOPSYS_UNCONNECTED_90,
         SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92,
         SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94,
         SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96,
         SYNOPSYS_UNCONNECTED_97, SYNOPSYS_UNCONNECTED_98,
         SYNOPSYS_UNCONNECTED_99, SYNOPSYS_UNCONNECTED_100,
         SYNOPSYS_UNCONNECTED_101, SYNOPSYS_UNCONNECTED_102,
         SYNOPSYS_UNCONNECTED_103, SYNOPSYS_UNCONNECTED_104,
         SYNOPSYS_UNCONNECTED_105, SYNOPSYS_UNCONNECTED_106,
         SYNOPSYS_UNCONNECTED_107, SYNOPSYS_UNCONNECTED_108,
         SYNOPSYS_UNCONNECTED_109, SYNOPSYS_UNCONNECTED_110,
         SYNOPSYS_UNCONNECTED_111, SYNOPSYS_UNCONNECTED_112,
         SYNOPSYS_UNCONNECTED_113, SYNOPSYS_UNCONNECTED_114,
         SYNOPSYS_UNCONNECTED_115, SYNOPSYS_UNCONNECTED_116,
         SYNOPSYS_UNCONNECTED_117, SYNOPSYS_UNCONNECTED_118;
  wire   [32:0] CMD_data_in;
  wire   [40:0] RETURN_data_in;
  wire   [1:0] init_ba;
  wire   [10:4] init_a;
  wire   [10:4] a_i;
  wire   [1:0] ba_i;
  wire   [15:0] dq_i;
  wire   [1:0] dqs_i;
  wire   [1:0] dqsbar_i;
  wire   [1:0] dm_i;
  assign notfull = 1'b1;

  DFFPOSX1 ck_i_reg ( .D(n3), .CLK(clk), .Q(ck_i) );
  FIFO_DEPTH_P25_WIDTH16 FIFO_IN ( .clk(clk), .reset(resetbar), .data_in(din), 
        .put(1'b0), .get(1'b0), .data_out(dout), .empty_bar(notempty), 
        .full_bar(), .fillcount(fillcount) );
  FIFO_DEPTH_P25_WIDTH33 FIFO_CMD ( .clk(clk), .reset(resetbar), .data_in({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .put(1'b0), 
        .get(1'b0), .data_out({SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, 
        SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, 
        SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, 
        SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10, 
        SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12, 
        SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14, 
        SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16, 
        SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18, 
        SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20, 
        SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22, 
        SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24, 
        SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26, 
        SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28, 
        SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30, 
        SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32, 
        SYNOPSYS_UNCONNECTED_33}), .empty_bar(), .full_bar(), .fillcount({
        SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35, 
        SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37, 
        SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39}) );
  FIFO_DEPTH_P25_WIDTH41 FIFO_RETURN ( .clk(clk), .reset(resetbar), .data_in({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .put(1'b0), .get(1'b0), .data_out({
        SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41, 
        SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_43, 
        SYNOPSYS_UNCONNECTED_44, SYNOPSYS_UNCONNECTED_45, 
        SYNOPSYS_UNCONNECTED_46, SYNOPSYS_UNCONNECTED_47, 
        SYNOPSYS_UNCONNECTED_48, SYNOPSYS_UNCONNECTED_49, 
        SYNOPSYS_UNCONNECTED_50, SYNOPSYS_UNCONNECTED_51, 
        SYNOPSYS_UNCONNECTED_52, SYNOPSYS_UNCONNECTED_53, 
        SYNOPSYS_UNCONNECTED_54, SYNOPSYS_UNCONNECTED_55, 
        SYNOPSYS_UNCONNECTED_56, SYNOPSYS_UNCONNECTED_57, 
        SYNOPSYS_UNCONNECTED_58, SYNOPSYS_UNCONNECTED_59, 
        SYNOPSYS_UNCONNECTED_60, SYNOPSYS_UNCONNECTED_61, 
        SYNOPSYS_UNCONNECTED_62, SYNOPSYS_UNCONNECTED_63, 
        SYNOPSYS_UNCONNECTED_64, SYNOPSYS_UNCONNECTED_65, 
        SYNOPSYS_UNCONNECTED_66, SYNOPSYS_UNCONNECTED_67, 
        SYNOPSYS_UNCONNECTED_68, SYNOPSYS_UNCONNECTED_69, 
        SYNOPSYS_UNCONNECTED_70, SYNOPSYS_UNCONNECTED_71, 
        SYNOPSYS_UNCONNECTED_72, SYNOPSYS_UNCONNECTED_73, 
        SYNOPSYS_UNCONNECTED_74, SYNOPSYS_UNCONNECTED_75, 
        SYNOPSYS_UNCONNECTED_76, SYNOPSYS_UNCONNECTED_77, 
        SYNOPSYS_UNCONNECTED_78, SYNOPSYS_UNCONNECTED_79, 
        SYNOPSYS_UNCONNECTED_80}), .empty_bar(), .full_bar(), .fillcount({
        SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82, 
        SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84, 
        SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86}) );
  ddr3_init_engine XINIT ( .ready(ready), .csbar(init_csbar), .rasbar(
        init_rasbar), .casbar(init_casbar), .webar(init_webar), .ba({
        SYNOPSYS_UNCONNECTED_87, init_ba}), .a({SYNOPSYS_UNCONNECTED_88, 
        SYNOPSYS_UNCONNECTED_89, SYNOPSYS_UNCONNECTED_90, init_a[10], 
        SYNOPSYS_UNCONNECTED_91, init_a[8], SYNOPSYS_UNCONNECTED_92, 
        SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94, init_a[4], 
        SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96, 
        SYNOPSYS_UNCONNECTED_97, SYNOPSYS_UNCONNECTED_98}), .odt(), .ts_con(), 
        .cke(init_cke), .clk(clk), .resetbar(resetbar), .init(initddr), .ck(
        1'b0), .Port15() );
  SSTL18DDR3INTERFACE XSSTL ( .ck_pad(ck_pad), .ckbar_pad(ckbar_pad), 
        .cke_pad(cke_pad), .csbar_pad(csbar_pad), .rasbar_pad(rasbar_pad), 
        .casbar_pad(casbar_pad), .webar_pad(webar_pad), .ba_pad(ba_pad), 
        .a_pad(a_pad), .dm_pad(dm_pad), .odt_pad(odt_pad), .resetbar_pad(
        resetbar_pad), .dq_o({SYNOPSYS_UNCONNECTED_99, 
        SYNOPSYS_UNCONNECTED_100, SYNOPSYS_UNCONNECTED_101, 
        SYNOPSYS_UNCONNECTED_102, SYNOPSYS_UNCONNECTED_103, 
        SYNOPSYS_UNCONNECTED_104, SYNOPSYS_UNCONNECTED_105, 
        SYNOPSYS_UNCONNECTED_106, SYNOPSYS_UNCONNECTED_107, 
        SYNOPSYS_UNCONNECTED_108, SYNOPSYS_UNCONNECTED_109, 
        SYNOPSYS_UNCONNECTED_110, SYNOPSYS_UNCONNECTED_111, 
        SYNOPSYS_UNCONNECTED_112, SYNOPSYS_UNCONNECTED_113, 
        SYNOPSYS_UNCONNECTED_114}), .dqs_o({SYNOPSYS_UNCONNECTED_115, 
        SYNOPSYS_UNCONNECTED_116}), .dqsbar_o({SYNOPSYS_UNCONNECTED_117, 
        SYNOPSYS_UNCONNECTED_118}), .dq_pad(dq_pad), .dqs_pad(dqs_pad), 
        .dqsbar_pad(dqsbar_pad), .ri_i(1'b0), .ts_i(1'b0), .ck_i(ck_i), 
        .cke_i(init_cke), .csbar_i(csbar_i), .rasbar_i(rasbar_i), .casbar_i(
        casbar_i), .webar_i(webar_i), .ba_i({1'b0, ba_i}), .a_i({1'b0, 1'b0, 
        1'b0, a_i[10], 1'b0, a_i[8], 1'b0, 1'b0, 1'b0, a_i[4], 1'b0, 1'b0, 
        1'b0, 1'b0}), .dq_i({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .dqs_i({1'b0, 1'b0}), 
        .dqsbar_i({1'b0, 1'b0}), .dm_i({1'b0, 1'b0}), .odt_i(1'b0), 
        .resetbar_i(1'b0) );
  OR2X1 U27 ( .A(ck_i), .B(n4), .Y(n6) );
  INVX1 U28 ( .A(n6), .Y(n3) );
  INVX1 U29 ( .A(resetbar), .Y(n4) );
  INVX1 U30 ( .A(ready), .Y(n7) );
  AND2X1 U31 ( .A(init_a[10]), .B(n7), .Y(a_i[10]) );
  AND2X1 U32 ( .A(init_a[8]), .B(n7), .Y(a_i[8]) );
  AND2X1 U33 ( .A(init_a[4]), .B(n7), .Y(a_i[4]) );
  AND2X1 U34 ( .A(init_ba[1]), .B(n7), .Y(ba_i[1]) );
  AND2X1 U35 ( .A(init_ba[0]), .B(n7), .Y(ba_i[0]) );
  AND2X1 U36 ( .A(init_webar), .B(n7), .Y(webar_i) );
  AND2X1 U37 ( .A(init_csbar), .B(n7), .Y(csbar_i) );
  AND2X1 U38 ( .A(init_rasbar), .B(n7), .Y(rasbar_i) );
  AND2X1 U39 ( .A(init_casbar), .B(n7), .Y(casbar_i) );
endmodule

