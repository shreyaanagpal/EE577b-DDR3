
module FIFO_2clk_DATA_WIDTH16_FIFO_DEPTH32_PTR_WIDTH6 ( rclk, wclk, reset, we, 
        re, data_in, empty_bar, full_bar, data_out, fillcount );
  input [15:0] data_in;
  output [15:0] data_out;
  output [5:0] fillcount;
  input rclk, wclk, reset, we, re;
  output empty_bar, full_bar;
  wire   n10, n11, n12, n13, n14, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, rd_ptr_bin_5_, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n33, n34, n35, n36, n37, n38, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n88, n89, n90, n91,
         n92, n175, n176, n177, n178, n179, n180, n181, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n1330,
         n1335, n1340, n1345, n1347, n1349, n1351, n1353, n1355, n1357, n1359,
         n1361, n1363, n1365, n1367, n1369, n1371, n1373, n1375, n1377, n1385,
         n1390, n1395, n1400, n1402, n1407, n1415, n1416, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
         n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
         n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
         n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         r301_B_not_0_, r301_B_not_1_, r301_B_not_2_, r301_B_not_3_,
         r301_B_not_4_, r301_B_not_5_, n1, n39, n40, n42, n43, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n87, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n182, n216, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1346, n1368, n1401,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
         n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
         n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
         n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
         n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
         n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
         n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
         n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
         n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
         n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
         n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
         n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
         n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
         n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
         n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
         n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
         n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
         n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
         n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
         n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
         n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
         n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
         n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
         n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
         n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
         n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
         n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
         n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
         n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
         n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
         n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
         n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
         n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
         n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
         n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
         n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
         n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819;
  wire   [5:0] wr_ptr_gray;
  wire   [5:0] wr_ptr_gray_ss;
  wire   [5:0] wr_ptr_gray_s;
  wire   [5:0] rd_ptr_gray;
  wire   [5:0] rd_ptr_gray_ss;
  wire   [5:0] rd_ptr_gray_s;
  wire   [4:0] rd_ptr_bin_ss;
  wire   [5:0] wr_ptr_bin;
  wire   [511:0] fifo;
  wire   [5:2] add_176_carry;
  wire   [5:2] add_158_carry;
  wire   [5:1] r301_carry;

  DFFSR rd_ptr_bin_reg_0_ ( .D(n1418), .CLK(rclk), .R(n5279), .S(1'b1), .Q(n10) );
  DFFSR rd_ptr_bin_reg_5_ ( .D(n1415), .CLK(rclk), .R(n5278), .S(1'b1), .Q(
        rd_ptr_bin_5_) );
  DFFSR rd_ptr_gray_reg_5_ ( .D(n4627), .CLK(rclk), .R(n5278), .S(1'b1), .Q(
        rd_ptr_gray[5]) );
  DFFSR rd_ptr_gray_s_reg_5_ ( .D(n137), .CLK(wclk), .R(n5277), .S(1'b1), .Q(
        rd_ptr_gray_s[5]) );
  DFFSR rd_ptr_gray_ss_reg_5_ ( .D(n134), .CLK(wclk), .R(n5277), .S(1'b1), .Q(
        rd_ptr_gray_ss[5]) );
  DFFSR rd_ptr_gray_reg_4_ ( .D(n15), .CLK(rclk), .R(n5277), .S(1'b1), .Q(
        rd_ptr_gray[4]) );
  DFFSR rd_ptr_gray_s_reg_4_ ( .D(n131), .CLK(wclk), .R(n5277), .S(1'b1), .Q(
        rd_ptr_gray_s[4]) );
  DFFSR rd_ptr_gray_ss_reg_4_ ( .D(n128), .CLK(wclk), .R(n5277), .S(1'b1), .Q(
        rd_ptr_gray_ss[4]) );
  DFFSR wr_ptr_bin_reg_5_ ( .D(n1407), .CLK(wclk), .R(n5280), .S(1'b1), .Q(
        wr_ptr_bin[5]) );
  DFFSR wr_ptr_gray_reg_5_ ( .D(n4630), .CLK(wclk), .R(n5280), .S(1'b1), .Q(
        wr_ptr_gray[5]) );
  DFFSR wr_ptr_gray_s_reg_5_ ( .D(n125), .CLK(rclk), .R(n5280), .S(1'b1), .Q(
        wr_ptr_gray_s[5]) );
  DFFSR wr_ptr_gray_ss_reg_5_ ( .D(n122), .CLK(rclk), .R(n5280), .S(1'b1), .Q(
        wr_ptr_gray_ss[5]) );
  DFFSR wr_ptr_bin_reg_1_ ( .D(n1400), .CLK(wclk), .R(n5281), .S(1'b1), .Q(
        wr_ptr_bin[1]) );
  DFFSR wr_ptr_gray_reg_0_ ( .D(n24), .CLK(wclk), .R(n5281), .S(1'b1), .Q(
        wr_ptr_gray[0]) );
  DFFSR wr_ptr_gray_s_reg_0_ ( .D(n119), .CLK(rclk), .R(n5281), .S(1'b1), .Q(
        wr_ptr_gray_s[0]) );
  DFFSR wr_ptr_gray_ss_reg_0_ ( .D(n116), .CLK(rclk), .R(n5281), .S(1'b1), .Q(
        wr_ptr_gray_ss[0]) );
  DFFSR wr_ptr_bin_reg_2_ ( .D(n1395), .CLK(wclk), .R(n5281), .S(1'b1), .Q(
        wr_ptr_bin[2]) );
  DFFSR wr_ptr_gray_reg_1_ ( .D(n861), .CLK(wclk), .R(n5281), .S(1'b1), .Q(
        wr_ptr_gray[1]) );
  DFFSR wr_ptr_gray_s_reg_1_ ( .D(n113), .CLK(rclk), .R(n5281), .S(1'b1), .Q(
        wr_ptr_gray_s[1]) );
  DFFSR wr_ptr_gray_ss_reg_1_ ( .D(n110), .CLK(rclk), .R(n5281), .S(1'b1), .Q(
        wr_ptr_gray_ss[1]) );
  DFFSR wr_ptr_bin_reg_3_ ( .D(n1390), .CLK(wclk), .R(n5281), .S(1'b1), .Q(
        wr_ptr_bin[3]) );
  DFFSR wr_ptr_gray_reg_2_ ( .D(n22), .CLK(wclk), .R(n5281), .S(1'b1), .Q(
        wr_ptr_gray[2]) );
  DFFSR wr_ptr_gray_s_reg_2_ ( .D(n107), .CLK(rclk), .R(n5281), .S(1'b1), .Q(
        wr_ptr_gray_s[2]) );
  DFFSR wr_ptr_gray_ss_reg_2_ ( .D(n104), .CLK(rclk), .R(n5280), .S(1'b1), .Q(
        wr_ptr_gray_ss[2]) );
  DFFSR wr_ptr_bin_reg_4_ ( .D(n1385), .CLK(wclk), .R(n5280), .S(1'b1), .Q(
        wr_ptr_bin[4]) );
  DFFSR wr_ptr_gray_reg_3_ ( .D(n21), .CLK(wclk), .R(n5279), .S(1'b1), .Q(
        wr_ptr_gray[3]) );
  DFFSR wr_ptr_gray_s_reg_3_ ( .D(n101), .CLK(rclk), .R(n5279), .S(1'b1), .Q(
        wr_ptr_gray_s[3]) );
  DFFSR wr_ptr_gray_ss_reg_3_ ( .D(n98), .CLK(rclk), .R(n5279), .S(1'b1), .Q(
        wr_ptr_gray_ss[3]) );
  DFFSR wr_ptr_gray_reg_4_ ( .D(n20), .CLK(wclk), .R(n5279), .S(1'b1), .Q(
        wr_ptr_gray[4]) );
  DFFSR wr_ptr_gray_s_reg_4_ ( .D(n95), .CLK(rclk), .R(n5279), .S(1'b1), .Q(
        wr_ptr_gray_s[4]) );
  DFFSR wr_ptr_gray_ss_reg_4_ ( .D(n87), .CLK(rclk), .R(n5279), .S(1'b1), .Q(
        wr_ptr_gray_ss[4]) );
  DFFSR data_out_reg_0_ ( .D(n1377), .CLK(rclk), .R(n5277), .S(1'b1), .Q(n5837) );
  DFFSR data_out_reg_1_ ( .D(n1375), .CLK(rclk), .R(n5277), .S(1'b1), .Q(n5836) );
  DFFSR data_out_reg_2_ ( .D(n1373), .CLK(rclk), .R(n5277), .S(1'b1), .Q(n5835) );
  DFFSR data_out_reg_3_ ( .D(n1371), .CLK(rclk), .R(n5277), .S(1'b1), .Q(n5834) );
  DFFSR data_out_reg_5_ ( .D(n1367), .CLK(rclk), .R(n5276), .S(1'b1), .Q(n5832) );
  DFFSR data_out_reg_6_ ( .D(n1365), .CLK(rclk), .R(n5276), .S(1'b1), .Q(n5831) );
  DFFSR data_out_reg_7_ ( .D(n1363), .CLK(rclk), .R(n5276), .S(1'b1), .Q(n5830) );
  DFFSR data_out_reg_8_ ( .D(n1361), .CLK(rclk), .R(n5276), .S(1'b1), .Q(n5829) );
  DFFSR data_out_reg_9_ ( .D(n1359), .CLK(rclk), .R(n5276), .S(1'b1), .Q(n5828) );
  DFFSR data_out_reg_10_ ( .D(n1357), .CLK(rclk), .R(n5276), .S(1'b1), .Q(
        n5827) );
  DFFSR data_out_reg_11_ ( .D(n1355), .CLK(rclk), .R(n5276), .S(1'b1), .Q(
        n5826) );
  DFFSR data_out_reg_12_ ( .D(n1353), .CLK(rclk), .R(n5276), .S(1'b1), .Q(
        n5825) );
  DFFSR data_out_reg_13_ ( .D(n1351), .CLK(rclk), .R(n5276), .S(1'b1), .Q(
        n5824) );
  DFFSR data_out_reg_14_ ( .D(n1349), .CLK(rclk), .R(n5276), .S(1'b1), .Q(
        n5823) );
  DFFSR rd_ptr_bin_reg_1_ ( .D(n1345), .CLK(rclk), .R(n5279), .S(1'b1), .Q(n11) );
  DFFSR rd_ptr_gray_reg_0_ ( .D(n19), .CLK(rclk), .R(n5279), .S(1'b1), .Q(
        rd_ptr_gray[0]) );
  DFFSR rd_ptr_gray_s_reg_0_ ( .D(n68), .CLK(wclk), .R(n5279), .S(1'b1), .Q(
        rd_ptr_gray_s[0]) );
  DFFSR rd_ptr_gray_ss_reg_0_ ( .D(n65), .CLK(wclk), .R(n5278), .S(1'b1), .Q(
        rd_ptr_gray_ss[0]) );
  DFFSR rd_ptr_bin_reg_2_ ( .D(n1340), .CLK(rclk), .R(n5278), .S(1'b1), .Q(n12) );
  DFFSR rd_ptr_gray_reg_1_ ( .D(n18), .CLK(rclk), .R(n5278), .S(1'b1), .Q(
        rd_ptr_gray[1]) );
  DFFSR rd_ptr_gray_s_reg_1_ ( .D(n62), .CLK(wclk), .R(n5278), .S(1'b1), .Q(
        rd_ptr_gray_s[1]) );
  DFFSR rd_ptr_gray_ss_reg_1_ ( .D(n59), .CLK(wclk), .R(n5278), .S(1'b1), .Q(
        rd_ptr_gray_ss[1]) );
  DFFSR rd_ptr_bin_reg_3_ ( .D(n1335), .CLK(rclk), .R(n5278), .S(1'b1), .Q(n13) );
  DFFSR rd_ptr_gray_reg_2_ ( .D(n17), .CLK(rclk), .R(n5278), .S(1'b1), .Q(
        rd_ptr_gray[2]) );
  DFFSR rd_ptr_gray_s_reg_2_ ( .D(n56), .CLK(wclk), .R(n5278), .S(1'b1), .Q(
        rd_ptr_gray_s[2]) );
  DFFSR rd_ptr_gray_ss_reg_2_ ( .D(n53), .CLK(wclk), .R(n5278), .S(1'b1), .Q(
        rd_ptr_gray_ss[2]) );
  DFFSR rd_ptr_bin_reg_4_ ( .D(n1330), .CLK(rclk), .R(n5278), .S(1'b1), .Q(n14) );
  DFFSR rd_ptr_gray_reg_3_ ( .D(n16), .CLK(rclk), .R(n5277), .S(1'b1), .Q(
        rd_ptr_gray[3]) );
  DFFSR rd_ptr_gray_s_reg_3_ ( .D(n50), .CLK(wclk), .R(n5277), .S(1'b1), .Q(
        rd_ptr_gray_s[3]) );
  DFFSR rd_ptr_gray_ss_reg_3_ ( .D(n47), .CLK(wclk), .R(n5277), .S(1'b1), .Q(
        rd_ptr_gray_ss[3]) );
  XOR2X1 U7 ( .A(rd_ptr_bin_ss[4]), .B(n3051), .Y(rd_ptr_bin_ss[3]) );
  XOR2X1 U8 ( .A(n4601), .B(n39), .Y(rd_ptr_bin_ss[4]) );
  OAI21X1 U9 ( .A(n175), .B(n176), .C(n3033), .Y(n1330) );
  INVX1 U11 ( .A(n4652), .Y(n176) );
  OAI21X1 U12 ( .A(n175), .B(n178), .C(n3030), .Y(n1335) );
  INVX1 U14 ( .A(n4751), .Y(n178) );
  OAI21X1 U15 ( .A(n175), .B(n180), .C(n3027), .Y(n1340) );
  OAI21X1 U17 ( .A(n175), .B(n5293), .C(n3024), .Y(n1345) );
  INVX1 U19 ( .A(n847), .Y(n1347) );
  INVX1 U21 ( .A(n186), .Y(n1349) );
  AOI22X1 U22 ( .A(data_out[14]), .B(n4649), .C(n72), .D(n175), .Y(n186) );
  INVX1 U23 ( .A(n834), .Y(n1351) );
  INVX1 U25 ( .A(n188), .Y(n1353) );
  AOI22X1 U26 ( .A(data_out[12]), .B(n4649), .C(n74), .D(n175), .Y(n188) );
  INVX1 U27 ( .A(n189), .Y(n1355) );
  AOI22X1 U28 ( .A(data_out[11]), .B(n4649), .C(n75), .D(n175), .Y(n189) );
  INVX1 U29 ( .A(n821), .Y(n1357) );
  INVX1 U31 ( .A(n191), .Y(n1359) );
  AOI22X1 U32 ( .A(data_out[9]), .B(n4649), .C(n77), .D(n175), .Y(n191) );
  INVX1 U33 ( .A(n192), .Y(n1361) );
  AOI22X1 U34 ( .A(data_out[8]), .B(n4649), .C(n78), .D(n175), .Y(n192) );
  INVX1 U35 ( .A(n171), .Y(n1363) );
  INVX1 U37 ( .A(n194), .Y(n1365) );
  AOI22X1 U38 ( .A(data_out[6]), .B(n4649), .C(n80), .D(n175), .Y(n194) );
  INVX1 U39 ( .A(n195), .Y(n1367) );
  AOI22X1 U40 ( .A(data_out[5]), .B(n4649), .C(n81), .D(n175), .Y(n195) );
  INVX1 U41 ( .A(n158), .Y(n1369) );
  INVX1 U43 ( .A(n197), .Y(n1371) );
  AOI22X1 U44 ( .A(data_out[3]), .B(n4649), .C(n83), .D(n175), .Y(n197) );
  INVX1 U45 ( .A(n198), .Y(n1373) );
  AOI22X1 U46 ( .A(data_out[2]), .B(n4649), .C(n84), .D(n175), .Y(n198) );
  INVX1 U47 ( .A(n145), .Y(n1375) );
  INVX1 U49 ( .A(n200), .Y(n1377) );
  AOI22X1 U50 ( .A(data_out[0]), .B(n4649), .C(n86), .D(n175), .Y(n200) );
  OAI21X1 U51 ( .A(n201), .B(n202), .C(n3022), .Y(n1385) );
  OAI21X1 U53 ( .A(n201), .B(n204), .C(n3020), .Y(n1390) );
  OAI21X1 U55 ( .A(n201), .B(n206), .C(n3017), .Y(n1395) );
  OAI21X1 U57 ( .A(n201), .B(n208), .C(n3014), .Y(n1400) );
  OAI21X1 U59 ( .A(n201), .B(n210), .C(n3011), .Y(n1402) );
  OAI21X1 U61 ( .A(n201), .B(n212), .C(n3008), .Y(n1407) );
  INVX1 U63 ( .A(n4630), .Y(n212) );
  OAI21X1 U64 ( .A(n175), .B(n214), .C(n3005), .Y(n1415) );
  INVX1 U66 ( .A(reset), .Y(n1416) );
  OAI21X1 U67 ( .A(n175), .B(n5314), .C(n3002), .Y(n1418) );
  INVX1 U69 ( .A(n4649), .Y(n175) );
  OAI21X1 U71 ( .A(n4655), .B(n219), .C(n2999), .Y(n1419) );
  OAI21X1 U73 ( .A(n4655), .B(n221), .C(n2996), .Y(n1420) );
  OAI21X1 U75 ( .A(n4655), .B(n223), .C(n2993), .Y(n1421) );
  OAI21X1 U77 ( .A(n4655), .B(n225), .C(n2990), .Y(n1422) );
  OAI21X1 U79 ( .A(n4655), .B(n227), .C(n2987), .Y(n1423) );
  OAI21X1 U81 ( .A(n4655), .B(n229), .C(n2984), .Y(n1424) );
  OAI21X1 U83 ( .A(n4655), .B(n231), .C(n2981), .Y(n1425) );
  OAI21X1 U85 ( .A(n4655), .B(n233), .C(n2978), .Y(n1426) );
  OAI21X1 U87 ( .A(n4655), .B(n235), .C(n2975), .Y(n1427) );
  OAI21X1 U89 ( .A(n4655), .B(n237), .C(n2972), .Y(n1428) );
  OAI21X1 U91 ( .A(n4655), .B(n239), .C(n2969), .Y(n1429) );
  OAI21X1 U93 ( .A(n4655), .B(n241), .C(n2966), .Y(n1430) );
  OAI21X1 U95 ( .A(n4655), .B(n243), .C(n2963), .Y(n1431) );
  OAI21X1 U97 ( .A(n4655), .B(n245), .C(n2960), .Y(n1432) );
  OAI21X1 U99 ( .A(n4655), .B(n247), .C(n2957), .Y(n1433) );
  OAI21X1 U101 ( .A(n4655), .B(n249), .C(n2954), .Y(n1434) );
  OAI21X1 U104 ( .A(n219), .B(n4748), .C(n2951), .Y(n1435) );
  OAI21X1 U106 ( .A(n221), .B(n4748), .C(n2948), .Y(n1436) );
  OAI21X1 U108 ( .A(n223), .B(n4748), .C(n2945), .Y(n1437) );
  OAI21X1 U110 ( .A(n225), .B(n4748), .C(n2942), .Y(n1438) );
  OAI21X1 U112 ( .A(n227), .B(n4748), .C(n2939), .Y(n1439) );
  OAI21X1 U114 ( .A(n229), .B(n4748), .C(n2936), .Y(n1440) );
  OAI21X1 U116 ( .A(n231), .B(n4748), .C(n2933), .Y(n1441) );
  OAI21X1 U118 ( .A(n233), .B(n4748), .C(n2930), .Y(n1442) );
  OAI21X1 U120 ( .A(n235), .B(n4748), .C(n2927), .Y(n1443) );
  OAI21X1 U122 ( .A(n237), .B(n4748), .C(n2924), .Y(n1444) );
  OAI21X1 U124 ( .A(n239), .B(n4748), .C(n2921), .Y(n1445) );
  OAI21X1 U126 ( .A(n241), .B(n4748), .C(n2918), .Y(n1446) );
  OAI21X1 U128 ( .A(n243), .B(n4748), .C(n2915), .Y(n1447) );
  OAI21X1 U130 ( .A(n245), .B(n4748), .C(n2912), .Y(n1448) );
  OAI21X1 U132 ( .A(n247), .B(n4748), .C(n2909), .Y(n1449) );
  OAI21X1 U134 ( .A(n249), .B(n4748), .C(n2906), .Y(n1450) );
  OAI21X1 U137 ( .A(n219), .B(n4745), .C(n2903), .Y(n1451) );
  OAI21X1 U139 ( .A(n221), .B(n4745), .C(n2900), .Y(n1452) );
  OAI21X1 U141 ( .A(n223), .B(n4745), .C(n2897), .Y(n1453) );
  OAI21X1 U143 ( .A(n225), .B(n4745), .C(n2894), .Y(n1454) );
  OAI21X1 U145 ( .A(n227), .B(n4745), .C(n2891), .Y(n1455) );
  OAI21X1 U147 ( .A(n229), .B(n4745), .C(n2888), .Y(n1456) );
  OAI21X1 U149 ( .A(n231), .B(n4745), .C(n2885), .Y(n1457) );
  OAI21X1 U151 ( .A(n233), .B(n4745), .C(n2882), .Y(n1458) );
  OAI21X1 U153 ( .A(n235), .B(n4745), .C(n2879), .Y(n1459) );
  OAI21X1 U155 ( .A(n237), .B(n4745), .C(n2876), .Y(n1460) );
  OAI21X1 U157 ( .A(n239), .B(n4745), .C(n2873), .Y(n1461) );
  OAI21X1 U159 ( .A(n241), .B(n4745), .C(n2870), .Y(n1462) );
  OAI21X1 U161 ( .A(n243), .B(n4745), .C(n2867), .Y(n1463) );
  OAI21X1 U163 ( .A(n245), .B(n4745), .C(n2864), .Y(n1464) );
  OAI21X1 U165 ( .A(n247), .B(n4745), .C(n2861), .Y(n1465) );
  OAI21X1 U167 ( .A(n249), .B(n4745), .C(n2858), .Y(n1466) );
  OAI21X1 U170 ( .A(n219), .B(n4742), .C(n2855), .Y(n1467) );
  OAI21X1 U172 ( .A(n221), .B(n4742), .C(n2852), .Y(n1468) );
  OAI21X1 U174 ( .A(n223), .B(n4742), .C(n2849), .Y(n1469) );
  OAI21X1 U176 ( .A(n225), .B(n4742), .C(n2846), .Y(n1470) );
  OAI21X1 U178 ( .A(n227), .B(n4742), .C(n2843), .Y(n1471) );
  OAI21X1 U180 ( .A(n229), .B(n4742), .C(n2840), .Y(n1472) );
  OAI21X1 U182 ( .A(n231), .B(n4742), .C(n2837), .Y(n1473) );
  OAI21X1 U184 ( .A(n233), .B(n4742), .C(n2834), .Y(n1474) );
  OAI21X1 U186 ( .A(n235), .B(n4742), .C(n2831), .Y(n1475) );
  OAI21X1 U188 ( .A(n237), .B(n4742), .C(n2828), .Y(n1476) );
  OAI21X1 U190 ( .A(n239), .B(n4742), .C(n2825), .Y(n1477) );
  OAI21X1 U192 ( .A(n241), .B(n4742), .C(n2822), .Y(n1478) );
  OAI21X1 U194 ( .A(n243), .B(n4742), .C(n2819), .Y(n1479) );
  OAI21X1 U196 ( .A(n245), .B(n4742), .C(n2816), .Y(n1480) );
  OAI21X1 U198 ( .A(n247), .B(n4742), .C(n2813), .Y(n1481) );
  OAI21X1 U200 ( .A(n249), .B(n4742), .C(n2810), .Y(n1482) );
  OAI21X1 U203 ( .A(n219), .B(n4739), .C(n2807), .Y(n1483) );
  OAI21X1 U205 ( .A(n221), .B(n4739), .C(n2804), .Y(n1484) );
  OAI21X1 U207 ( .A(n223), .B(n4739), .C(n2801), .Y(n1485) );
  OAI21X1 U209 ( .A(n225), .B(n4739), .C(n2798), .Y(n1486) );
  OAI21X1 U211 ( .A(n227), .B(n4739), .C(n2795), .Y(n1487) );
  OAI21X1 U213 ( .A(n229), .B(n4739), .C(n2792), .Y(n1488) );
  OAI21X1 U215 ( .A(n231), .B(n4739), .C(n2789), .Y(n1489) );
  OAI21X1 U217 ( .A(n233), .B(n4739), .C(n2786), .Y(n1490) );
  OAI21X1 U219 ( .A(n235), .B(n4739), .C(n2783), .Y(n1491) );
  OAI21X1 U221 ( .A(n237), .B(n4739), .C(n2780), .Y(n1492) );
  OAI21X1 U223 ( .A(n239), .B(n4739), .C(n2777), .Y(n1493) );
  OAI21X1 U225 ( .A(n241), .B(n4739), .C(n2774), .Y(n1494) );
  OAI21X1 U227 ( .A(n243), .B(n4739), .C(n2771), .Y(n1495) );
  OAI21X1 U229 ( .A(n245), .B(n4739), .C(n2768), .Y(n1496) );
  OAI21X1 U231 ( .A(n247), .B(n4739), .C(n2765), .Y(n1497) );
  OAI21X1 U233 ( .A(n249), .B(n4739), .C(n2762), .Y(n1498) );
  OAI21X1 U236 ( .A(n219), .B(n4736), .C(n2759), .Y(n1499) );
  OAI21X1 U238 ( .A(n221), .B(n4736), .C(n2756), .Y(n1500) );
  OAI21X1 U240 ( .A(n223), .B(n4736), .C(n2753), .Y(n1501) );
  OAI21X1 U242 ( .A(n225), .B(n4736), .C(n2750), .Y(n1502) );
  OAI21X1 U244 ( .A(n227), .B(n4736), .C(n2747), .Y(n1503) );
  OAI21X1 U246 ( .A(n229), .B(n4736), .C(n2744), .Y(n1504) );
  OAI21X1 U248 ( .A(n231), .B(n4736), .C(n2741), .Y(n1505) );
  OAI21X1 U250 ( .A(n233), .B(n4736), .C(n2738), .Y(n1506) );
  OAI21X1 U252 ( .A(n235), .B(n4736), .C(n2735), .Y(n1507) );
  OAI21X1 U254 ( .A(n237), .B(n4736), .C(n2732), .Y(n1508) );
  OAI21X1 U256 ( .A(n239), .B(n4736), .C(n2729), .Y(n1509) );
  OAI21X1 U258 ( .A(n241), .B(n4736), .C(n2726), .Y(n1510) );
  OAI21X1 U260 ( .A(n243), .B(n4736), .C(n2723), .Y(n1511) );
  OAI21X1 U262 ( .A(n245), .B(n4736), .C(n2720), .Y(n1512) );
  OAI21X1 U264 ( .A(n247), .B(n4736), .C(n2717), .Y(n1513) );
  OAI21X1 U266 ( .A(n249), .B(n4736), .C(n2714), .Y(n1514) );
  OAI21X1 U269 ( .A(n219), .B(n4733), .C(n2711), .Y(n1515) );
  OAI21X1 U271 ( .A(n221), .B(n4733), .C(n2708), .Y(n1516) );
  OAI21X1 U273 ( .A(n223), .B(n4733), .C(n2705), .Y(n1517) );
  OAI21X1 U275 ( .A(n225), .B(n4733), .C(n2702), .Y(n1518) );
  OAI21X1 U277 ( .A(n227), .B(n4733), .C(n2699), .Y(n1519) );
  OAI21X1 U279 ( .A(n229), .B(n4733), .C(n2696), .Y(n1520) );
  OAI21X1 U281 ( .A(n231), .B(n4733), .C(n2693), .Y(n1521) );
  OAI21X1 U283 ( .A(n233), .B(n4733), .C(n2690), .Y(n1522) );
  OAI21X1 U285 ( .A(n235), .B(n4733), .C(n2687), .Y(n1523) );
  OAI21X1 U287 ( .A(n237), .B(n4733), .C(n2684), .Y(n1524) );
  OAI21X1 U289 ( .A(n239), .B(n4733), .C(n2681), .Y(n1525) );
  OAI21X1 U291 ( .A(n241), .B(n4733), .C(n2678), .Y(n1526) );
  OAI21X1 U293 ( .A(n243), .B(n4733), .C(n2675), .Y(n1527) );
  OAI21X1 U295 ( .A(n245), .B(n4733), .C(n2672), .Y(n1528) );
  OAI21X1 U297 ( .A(n247), .B(n4733), .C(n2669), .Y(n1529) );
  OAI21X1 U299 ( .A(n249), .B(n4733), .C(n2666), .Y(n1530) );
  OAI21X1 U302 ( .A(n219), .B(n4730), .C(n2663), .Y(n1531) );
  OAI21X1 U304 ( .A(n221), .B(n4730), .C(n2660), .Y(n1532) );
  OAI21X1 U306 ( .A(n223), .B(n4730), .C(n2657), .Y(n1533) );
  OAI21X1 U308 ( .A(n225), .B(n4730), .C(n2654), .Y(n1534) );
  OAI21X1 U310 ( .A(n227), .B(n4730), .C(n2651), .Y(n1535) );
  OAI21X1 U312 ( .A(n229), .B(n4730), .C(n2648), .Y(n1536) );
  OAI21X1 U314 ( .A(n231), .B(n4730), .C(n2645), .Y(n1537) );
  OAI21X1 U316 ( .A(n233), .B(n4730), .C(n2642), .Y(n1538) );
  OAI21X1 U318 ( .A(n235), .B(n4730), .C(n2639), .Y(n1539) );
  OAI21X1 U320 ( .A(n237), .B(n4730), .C(n2636), .Y(n1540) );
  OAI21X1 U322 ( .A(n239), .B(n4730), .C(n2633), .Y(n1541) );
  OAI21X1 U324 ( .A(n241), .B(n4730), .C(n2630), .Y(n1542) );
  OAI21X1 U326 ( .A(n243), .B(n4730), .C(n2627), .Y(n1543) );
  OAI21X1 U328 ( .A(n245), .B(n4730), .C(n2624), .Y(n1544) );
  OAI21X1 U330 ( .A(n247), .B(n4730), .C(n2621), .Y(n1545) );
  OAI21X1 U332 ( .A(n249), .B(n4730), .C(n2618), .Y(n1546) );
  INVX1 U335 ( .A(n379), .Y(n252) );
  NAND3X1 U336 ( .A(n204), .B(n202), .C(n201), .Y(n379) );
  OAI21X1 U337 ( .A(n219), .B(n4727), .C(n2615), .Y(n1547) );
  OAI21X1 U339 ( .A(n221), .B(n4727), .C(n2612), .Y(n1548) );
  OAI21X1 U341 ( .A(n223), .B(n4727), .C(n2609), .Y(n1549) );
  OAI21X1 U343 ( .A(n225), .B(n4727), .C(n2606), .Y(n1550) );
  OAI21X1 U345 ( .A(n227), .B(n4727), .C(n2603), .Y(n1551) );
  OAI21X1 U347 ( .A(n229), .B(n4727), .C(n2600), .Y(n1552) );
  OAI21X1 U349 ( .A(n231), .B(n4727), .C(n2597), .Y(n1553) );
  OAI21X1 U351 ( .A(n233), .B(n4727), .C(n2594), .Y(n1554) );
  OAI21X1 U353 ( .A(n235), .B(n4727), .C(n2591), .Y(n1555) );
  OAI21X1 U355 ( .A(n237), .B(n4727), .C(n2588), .Y(n1556) );
  OAI21X1 U357 ( .A(n239), .B(n4727), .C(n2585), .Y(n1557) );
  OAI21X1 U359 ( .A(n241), .B(n4727), .C(n2582), .Y(n1558) );
  OAI21X1 U361 ( .A(n243), .B(n4727), .C(n2579), .Y(n1559) );
  OAI21X1 U363 ( .A(n245), .B(n4727), .C(n2576), .Y(n1560) );
  OAI21X1 U365 ( .A(n247), .B(n4727), .C(n2573), .Y(n1561) );
  OAI21X1 U367 ( .A(n249), .B(n4727), .C(n2570), .Y(n1562) );
  OAI21X1 U370 ( .A(n219), .B(n4724), .C(n2567), .Y(n1563) );
  OAI21X1 U372 ( .A(n221), .B(n4724), .C(n2564), .Y(n1564) );
  OAI21X1 U374 ( .A(n223), .B(n4724), .C(n2561), .Y(n1565) );
  OAI21X1 U376 ( .A(n225), .B(n4724), .C(n2558), .Y(n1566) );
  OAI21X1 U378 ( .A(n227), .B(n4724), .C(n2555), .Y(n1567) );
  OAI21X1 U380 ( .A(n229), .B(n4724), .C(n2552), .Y(n1568) );
  OAI21X1 U382 ( .A(n231), .B(n4724), .C(n2549), .Y(n1569) );
  OAI21X1 U384 ( .A(n233), .B(n4724), .C(n2546), .Y(n1570) );
  OAI21X1 U386 ( .A(n235), .B(n4724), .C(n2543), .Y(n1571) );
  OAI21X1 U388 ( .A(n237), .B(n4724), .C(n2540), .Y(n1572) );
  OAI21X1 U390 ( .A(n239), .B(n4724), .C(n2537), .Y(n1573) );
  OAI21X1 U392 ( .A(n241), .B(n4724), .C(n2534), .Y(n1574) );
  OAI21X1 U394 ( .A(n243), .B(n4724), .C(n2531), .Y(n1575) );
  OAI21X1 U396 ( .A(n245), .B(n4724), .C(n2528), .Y(n1576) );
  OAI21X1 U398 ( .A(n247), .B(n4724), .C(n2525), .Y(n1577) );
  OAI21X1 U400 ( .A(n249), .B(n4724), .C(n2522), .Y(n1578) );
  OAI21X1 U403 ( .A(n219), .B(n4721), .C(n2519), .Y(n1579) );
  OAI21X1 U405 ( .A(n221), .B(n4721), .C(n2516), .Y(n1580) );
  OAI21X1 U407 ( .A(n223), .B(n4721), .C(n2513), .Y(n1581) );
  OAI21X1 U409 ( .A(n225), .B(n4721), .C(n2510), .Y(n1582) );
  OAI21X1 U411 ( .A(n227), .B(n4721), .C(n2507), .Y(n1583) );
  OAI21X1 U413 ( .A(n229), .B(n4721), .C(n2504), .Y(n1584) );
  OAI21X1 U415 ( .A(n231), .B(n4721), .C(n2501), .Y(n1585) );
  OAI21X1 U417 ( .A(n233), .B(n4721), .C(n2498), .Y(n1586) );
  OAI21X1 U419 ( .A(n235), .B(n4721), .C(n2495), .Y(n1587) );
  OAI21X1 U421 ( .A(n237), .B(n4721), .C(n2492), .Y(n1588) );
  OAI21X1 U423 ( .A(n239), .B(n4721), .C(n2489), .Y(n1589) );
  OAI21X1 U425 ( .A(n241), .B(n4721), .C(n2486), .Y(n1590) );
  OAI21X1 U427 ( .A(n243), .B(n4721), .C(n2483), .Y(n1591) );
  OAI21X1 U429 ( .A(n245), .B(n4721), .C(n2480), .Y(n1592) );
  OAI21X1 U431 ( .A(n247), .B(n4721), .C(n2477), .Y(n1593) );
  OAI21X1 U433 ( .A(n249), .B(n4721), .C(n2474), .Y(n1594) );
  OAI21X1 U436 ( .A(n219), .B(n4718), .C(n2471), .Y(n1595) );
  OAI21X1 U438 ( .A(n221), .B(n4718), .C(n2468), .Y(n1596) );
  OAI21X1 U440 ( .A(n223), .B(n4718), .C(n2465), .Y(n1597) );
  OAI21X1 U442 ( .A(n225), .B(n4718), .C(n2462), .Y(n1598) );
  OAI21X1 U444 ( .A(n227), .B(n4718), .C(n2459), .Y(n1599) );
  OAI21X1 U446 ( .A(n229), .B(n4718), .C(n2456), .Y(n1600) );
  OAI21X1 U448 ( .A(n231), .B(n4718), .C(n2453), .Y(n1601) );
  OAI21X1 U450 ( .A(n233), .B(n4718), .C(n2450), .Y(n1602) );
  OAI21X1 U452 ( .A(n235), .B(n4718), .C(n2447), .Y(n1603) );
  OAI21X1 U454 ( .A(n237), .B(n4718), .C(n2444), .Y(n1604) );
  OAI21X1 U456 ( .A(n239), .B(n4718), .C(n2441), .Y(n1605) );
  OAI21X1 U458 ( .A(n241), .B(n4718), .C(n2438), .Y(n1606) );
  OAI21X1 U460 ( .A(n243), .B(n4718), .C(n2435), .Y(n1607) );
  OAI21X1 U462 ( .A(n245), .B(n4718), .C(n2432), .Y(n1608) );
  OAI21X1 U464 ( .A(n247), .B(n4718), .C(n2429), .Y(n1609) );
  OAI21X1 U466 ( .A(n249), .B(n4718), .C(n2426), .Y(n1610) );
  OAI21X1 U469 ( .A(n219), .B(n4715), .C(n2423), .Y(n1611) );
  OAI21X1 U471 ( .A(n221), .B(n4715), .C(n2420), .Y(n1612) );
  OAI21X1 U473 ( .A(n223), .B(n4715), .C(n2417), .Y(n1613) );
  OAI21X1 U475 ( .A(n225), .B(n4715), .C(n2414), .Y(n1614) );
  OAI21X1 U477 ( .A(n227), .B(n4715), .C(n2411), .Y(n1615) );
  OAI21X1 U479 ( .A(n229), .B(n4715), .C(n2408), .Y(n1616) );
  OAI21X1 U481 ( .A(n231), .B(n4715), .C(n2405), .Y(n1617) );
  OAI21X1 U483 ( .A(n233), .B(n4715), .C(n2402), .Y(n1618) );
  OAI21X1 U485 ( .A(n235), .B(n4715), .C(n2399), .Y(n1619) );
  OAI21X1 U487 ( .A(n237), .B(n4715), .C(n2396), .Y(n1620) );
  OAI21X1 U489 ( .A(n239), .B(n4715), .C(n2393), .Y(n1621) );
  OAI21X1 U491 ( .A(n241), .B(n4715), .C(n2390), .Y(n1622) );
  OAI21X1 U493 ( .A(n243), .B(n4715), .C(n2387), .Y(n1623) );
  OAI21X1 U495 ( .A(n245), .B(n4715), .C(n2384), .Y(n1624) );
  OAI21X1 U497 ( .A(n247), .B(n4715), .C(n2381), .Y(n1625) );
  OAI21X1 U499 ( .A(n249), .B(n4715), .C(n2378), .Y(n1626) );
  OAI21X1 U502 ( .A(n219), .B(n4712), .C(n2375), .Y(n1627) );
  OAI21X1 U504 ( .A(n221), .B(n4712), .C(n2372), .Y(n1628) );
  OAI21X1 U506 ( .A(n223), .B(n4712), .C(n2369), .Y(n1629) );
  OAI21X1 U508 ( .A(n225), .B(n4712), .C(n2366), .Y(n1630) );
  OAI21X1 U510 ( .A(n227), .B(n4712), .C(n2363), .Y(n1631) );
  OAI21X1 U512 ( .A(n229), .B(n4712), .C(n2360), .Y(n1632) );
  OAI21X1 U514 ( .A(n231), .B(n4712), .C(n2357), .Y(n1633) );
  OAI21X1 U516 ( .A(n233), .B(n4712), .C(n2354), .Y(n1634) );
  OAI21X1 U518 ( .A(n235), .B(n4712), .C(n2351), .Y(n1635) );
  OAI21X1 U520 ( .A(n237), .B(n4712), .C(n2348), .Y(n1636) );
  OAI21X1 U522 ( .A(n239), .B(n4712), .C(n2345), .Y(n1637) );
  OAI21X1 U524 ( .A(n241), .B(n4712), .C(n2342), .Y(n1638) );
  OAI21X1 U526 ( .A(n243), .B(n4712), .C(n2339), .Y(n1639) );
  OAI21X1 U528 ( .A(n245), .B(n4712), .C(n2336), .Y(n1640) );
  OAI21X1 U530 ( .A(n247), .B(n4712), .C(n2333), .Y(n1641) );
  OAI21X1 U532 ( .A(n249), .B(n4712), .C(n2330), .Y(n1642) );
  OAI21X1 U535 ( .A(n219), .B(n4709), .C(n2327), .Y(n1643) );
  OAI21X1 U537 ( .A(n221), .B(n4709), .C(n2324), .Y(n1644) );
  OAI21X1 U539 ( .A(n223), .B(n4709), .C(n2321), .Y(n1645) );
  OAI21X1 U541 ( .A(n225), .B(n4709), .C(n2318), .Y(n1646) );
  OAI21X1 U543 ( .A(n227), .B(n4709), .C(n2315), .Y(n1647) );
  OAI21X1 U545 ( .A(n229), .B(n4709), .C(n2312), .Y(n1648) );
  OAI21X1 U547 ( .A(n231), .B(n4709), .C(n2309), .Y(n1649) );
  OAI21X1 U549 ( .A(n233), .B(n4709), .C(n2306), .Y(n1650) );
  OAI21X1 U551 ( .A(n235), .B(n4709), .C(n2303), .Y(n1651) );
  OAI21X1 U553 ( .A(n237), .B(n4709), .C(n2300), .Y(n1652) );
  OAI21X1 U555 ( .A(n239), .B(n4709), .C(n2297), .Y(n1653) );
  OAI21X1 U557 ( .A(n241), .B(n4709), .C(n2294), .Y(n1654) );
  OAI21X1 U559 ( .A(n243), .B(n4709), .C(n2291), .Y(n1655) );
  OAI21X1 U561 ( .A(n245), .B(n4709), .C(n2288), .Y(n1656) );
  OAI21X1 U563 ( .A(n247), .B(n4709), .C(n2285), .Y(n1657) );
  OAI21X1 U565 ( .A(n249), .B(n4709), .C(n2282), .Y(n1658) );
  OAI21X1 U568 ( .A(n219), .B(n4706), .C(n2279), .Y(n1659) );
  OAI21X1 U570 ( .A(n221), .B(n4706), .C(n2276), .Y(n1660) );
  OAI21X1 U572 ( .A(n223), .B(n4706), .C(n2273), .Y(n1661) );
  OAI21X1 U574 ( .A(n225), .B(n4706), .C(n2270), .Y(n1662) );
  OAI21X1 U576 ( .A(n227), .B(n4706), .C(n2267), .Y(n1663) );
  OAI21X1 U578 ( .A(n229), .B(n4706), .C(n2264), .Y(n1664) );
  OAI21X1 U580 ( .A(n231), .B(n4706), .C(n2261), .Y(n1665) );
  OAI21X1 U582 ( .A(n233), .B(n4706), .C(n2258), .Y(n1666) );
  OAI21X1 U584 ( .A(n235), .B(n4706), .C(n2255), .Y(n1667) );
  OAI21X1 U586 ( .A(n237), .B(n4706), .C(n2252), .Y(n1668) );
  OAI21X1 U588 ( .A(n239), .B(n4706), .C(n2249), .Y(n1669) );
  OAI21X1 U590 ( .A(n241), .B(n4706), .C(n2246), .Y(n1670) );
  OAI21X1 U592 ( .A(n243), .B(n4706), .C(n2243), .Y(n1671) );
  OAI21X1 U594 ( .A(n245), .B(n4706), .C(n2240), .Y(n1672) );
  OAI21X1 U596 ( .A(n247), .B(n4706), .C(n2237), .Y(n1673) );
  OAI21X1 U598 ( .A(n249), .B(n4706), .C(n2234), .Y(n1674) );
  INVX1 U601 ( .A(n517), .Y(n397) );
  NAND3X1 U602 ( .A(n201), .B(n202), .C(n4642), .Y(n517) );
  INVX1 U603 ( .A(n4639), .Y(n202) );
  OAI21X1 U604 ( .A(n219), .B(n4703), .C(n2231), .Y(n1675) );
  OAI21X1 U606 ( .A(n221), .B(n4703), .C(n2228), .Y(n1676) );
  OAI21X1 U608 ( .A(n223), .B(n4703), .C(n2225), .Y(n1677) );
  OAI21X1 U610 ( .A(n225), .B(n4703), .C(n2222), .Y(n1678) );
  OAI21X1 U612 ( .A(n227), .B(n4703), .C(n2219), .Y(n1679) );
  OAI21X1 U614 ( .A(n229), .B(n4703), .C(n2216), .Y(n1680) );
  OAI21X1 U616 ( .A(n231), .B(n4703), .C(n2213), .Y(n1681) );
  OAI21X1 U618 ( .A(n233), .B(n4703), .C(n2210), .Y(n1682) );
  OAI21X1 U620 ( .A(n235), .B(n4703), .C(n2207), .Y(n1683) );
  OAI21X1 U622 ( .A(n237), .B(n4703), .C(n2204), .Y(n1684) );
  OAI21X1 U624 ( .A(n239), .B(n4703), .C(n2201), .Y(n1685) );
  OAI21X1 U626 ( .A(n241), .B(n4703), .C(n2198), .Y(n1686) );
  OAI21X1 U628 ( .A(n243), .B(n4703), .C(n2195), .Y(n1687) );
  OAI21X1 U630 ( .A(n245), .B(n4703), .C(n2192), .Y(n1688) );
  OAI21X1 U632 ( .A(n247), .B(n4703), .C(n2189), .Y(n1689) );
  OAI21X1 U634 ( .A(n249), .B(n4703), .C(n2186), .Y(n1690) );
  OAI21X1 U637 ( .A(n219), .B(n4700), .C(n2183), .Y(n1691) );
  OAI21X1 U639 ( .A(n221), .B(n4700), .C(n2180), .Y(n1692) );
  OAI21X1 U641 ( .A(n223), .B(n4700), .C(n2177), .Y(n1693) );
  OAI21X1 U643 ( .A(n225), .B(n4700), .C(n2174), .Y(n1694) );
  OAI21X1 U645 ( .A(n227), .B(n4700), .C(n2171), .Y(n1695) );
  OAI21X1 U647 ( .A(n229), .B(n4700), .C(n2168), .Y(n1696) );
  OAI21X1 U649 ( .A(n231), .B(n4700), .C(n2165), .Y(n1697) );
  OAI21X1 U651 ( .A(n233), .B(n4700), .C(n2162), .Y(n1698) );
  OAI21X1 U653 ( .A(n235), .B(n4700), .C(n2159), .Y(n1699) );
  OAI21X1 U655 ( .A(n237), .B(n4700), .C(n2156), .Y(n1700) );
  OAI21X1 U657 ( .A(n239), .B(n4700), .C(n2153), .Y(n1701) );
  OAI21X1 U659 ( .A(n241), .B(n4700), .C(n2150), .Y(n1702) );
  OAI21X1 U661 ( .A(n243), .B(n4700), .C(n2147), .Y(n1703) );
  OAI21X1 U663 ( .A(n245), .B(n4700), .C(n2144), .Y(n1704) );
  OAI21X1 U665 ( .A(n247), .B(n4700), .C(n2141), .Y(n1705) );
  OAI21X1 U667 ( .A(n249), .B(n4700), .C(n2138), .Y(n1706) );
  OAI21X1 U670 ( .A(n219), .B(n4697), .C(n2135), .Y(n1707) );
  OAI21X1 U672 ( .A(n221), .B(n4697), .C(n2132), .Y(n1708) );
  OAI21X1 U674 ( .A(n223), .B(n4697), .C(n2129), .Y(n1709) );
  OAI21X1 U676 ( .A(n225), .B(n4697), .C(n2126), .Y(n1710) );
  OAI21X1 U678 ( .A(n227), .B(n4697), .C(n2123), .Y(n1711) );
  OAI21X1 U680 ( .A(n229), .B(n4697), .C(n2120), .Y(n1712) );
  OAI21X1 U682 ( .A(n231), .B(n4697), .C(n2117), .Y(n1713) );
  OAI21X1 U684 ( .A(n233), .B(n4697), .C(n2114), .Y(n1714) );
  OAI21X1 U686 ( .A(n235), .B(n4697), .C(n2111), .Y(n1715) );
  OAI21X1 U688 ( .A(n237), .B(n4697), .C(n2108), .Y(n1716) );
  OAI21X1 U690 ( .A(n239), .B(n4697), .C(n2105), .Y(n1717) );
  OAI21X1 U692 ( .A(n241), .B(n4697), .C(n2102), .Y(n1718) );
  OAI21X1 U694 ( .A(n243), .B(n4697), .C(n2099), .Y(n1719) );
  OAI21X1 U696 ( .A(n245), .B(n4697), .C(n2096), .Y(n1720) );
  OAI21X1 U698 ( .A(n247), .B(n4697), .C(n2093), .Y(n1721) );
  OAI21X1 U700 ( .A(n249), .B(n4697), .C(n2090), .Y(n1722) );
  OAI21X1 U703 ( .A(n219), .B(n4694), .C(n2087), .Y(n1723) );
  OAI21X1 U705 ( .A(n221), .B(n4694), .C(n2084), .Y(n1724) );
  OAI21X1 U707 ( .A(n223), .B(n4694), .C(n2081), .Y(n1725) );
  OAI21X1 U709 ( .A(n225), .B(n4694), .C(n2078), .Y(n1726) );
  OAI21X1 U711 ( .A(n227), .B(n4694), .C(n2075), .Y(n1727) );
  OAI21X1 U713 ( .A(n229), .B(n4694), .C(n2072), .Y(n1728) );
  OAI21X1 U715 ( .A(n231), .B(n4694), .C(n2069), .Y(n1729) );
  OAI21X1 U717 ( .A(n233), .B(n4694), .C(n2066), .Y(n1730) );
  OAI21X1 U719 ( .A(n235), .B(n4694), .C(n2063), .Y(n1731) );
  OAI21X1 U721 ( .A(n237), .B(n4694), .C(n2060), .Y(n1732) );
  OAI21X1 U723 ( .A(n239), .B(n4694), .C(n2057), .Y(n1733) );
  OAI21X1 U725 ( .A(n241), .B(n4694), .C(n2054), .Y(n1734) );
  OAI21X1 U727 ( .A(n243), .B(n4694), .C(n2051), .Y(n1735) );
  OAI21X1 U729 ( .A(n245), .B(n4694), .C(n2048), .Y(n1736) );
  OAI21X1 U731 ( .A(n247), .B(n4694), .C(n2045), .Y(n1737) );
  OAI21X1 U733 ( .A(n249), .B(n4694), .C(n2042), .Y(n1738) );
  OAI21X1 U736 ( .A(n219), .B(n4691), .C(n2039), .Y(n1739) );
  OAI21X1 U738 ( .A(n221), .B(n4691), .C(n2036), .Y(n1740) );
  OAI21X1 U740 ( .A(n223), .B(n4691), .C(n2033), .Y(n1741) );
  OAI21X1 U742 ( .A(n225), .B(n4691), .C(n2030), .Y(n1742) );
  OAI21X1 U744 ( .A(n227), .B(n4691), .C(n2027), .Y(n1743) );
  OAI21X1 U746 ( .A(n229), .B(n4691), .C(n2024), .Y(n1744) );
  OAI21X1 U748 ( .A(n231), .B(n4691), .C(n2021), .Y(n1745) );
  OAI21X1 U750 ( .A(n233), .B(n4691), .C(n2018), .Y(n1746) );
  OAI21X1 U752 ( .A(n235), .B(n4691), .C(n2015), .Y(n1747) );
  OAI21X1 U754 ( .A(n237), .B(n4691), .C(n2012), .Y(n1748) );
  OAI21X1 U756 ( .A(n239), .B(n4691), .C(n2009), .Y(n1749) );
  OAI21X1 U758 ( .A(n241), .B(n4691), .C(n2006), .Y(n1750) );
  OAI21X1 U760 ( .A(n243), .B(n4691), .C(n2003), .Y(n1751) );
  OAI21X1 U762 ( .A(n245), .B(n4691), .C(n2000), .Y(n1752) );
  OAI21X1 U764 ( .A(n247), .B(n4691), .C(n1997), .Y(n1753) );
  OAI21X1 U766 ( .A(n249), .B(n4691), .C(n1994), .Y(n1754) );
  OAI21X1 U769 ( .A(n219), .B(n4688), .C(n1991), .Y(n1755) );
  OAI21X1 U771 ( .A(n221), .B(n4688), .C(n1988), .Y(n1756) );
  OAI21X1 U773 ( .A(n223), .B(n4688), .C(n1985), .Y(n1757) );
  OAI21X1 U775 ( .A(n225), .B(n4688), .C(n1982), .Y(n1758) );
  OAI21X1 U777 ( .A(n227), .B(n4688), .C(n1979), .Y(n1759) );
  OAI21X1 U779 ( .A(n229), .B(n4688), .C(n1976), .Y(n1760) );
  OAI21X1 U781 ( .A(n231), .B(n4688), .C(n1973), .Y(n1761) );
  OAI21X1 U783 ( .A(n233), .B(n4688), .C(n1970), .Y(n1762) );
  OAI21X1 U785 ( .A(n235), .B(n4688), .C(n1967), .Y(n1763) );
  OAI21X1 U787 ( .A(n237), .B(n4688), .C(n1964), .Y(n1764) );
  OAI21X1 U789 ( .A(n239), .B(n4688), .C(n1961), .Y(n1765) );
  OAI21X1 U791 ( .A(n241), .B(n4688), .C(n1958), .Y(n1766) );
  OAI21X1 U793 ( .A(n243), .B(n4688), .C(n1955), .Y(n1767) );
  OAI21X1 U795 ( .A(n245), .B(n4688), .C(n1952), .Y(n1768) );
  OAI21X1 U797 ( .A(n247), .B(n4688), .C(n1949), .Y(n1769) );
  OAI21X1 U799 ( .A(n249), .B(n4688), .C(n1946), .Y(n1770) );
  OAI21X1 U802 ( .A(n219), .B(n4685), .C(n1943), .Y(n1771) );
  OAI21X1 U804 ( .A(n221), .B(n4685), .C(n1940), .Y(n1772) );
  OAI21X1 U806 ( .A(n223), .B(n4685), .C(n1937), .Y(n1773) );
  OAI21X1 U808 ( .A(n225), .B(n4685), .C(n1934), .Y(n1774) );
  OAI21X1 U810 ( .A(n227), .B(n4685), .C(n1931), .Y(n1775) );
  OAI21X1 U812 ( .A(n229), .B(n4685), .C(n1346), .Y(n1776) );
  OAI21X1 U814 ( .A(n231), .B(n4685), .C(n1323), .Y(n1777) );
  OAI21X1 U816 ( .A(n233), .B(n4685), .C(n1320), .Y(n1778) );
  OAI21X1 U818 ( .A(n235), .B(n4685), .C(n1317), .Y(n1779) );
  OAI21X1 U820 ( .A(n237), .B(n4685), .C(n1314), .Y(n1780) );
  OAI21X1 U822 ( .A(n239), .B(n4685), .C(n1311), .Y(n1781) );
  OAI21X1 U824 ( .A(n241), .B(n4685), .C(n1308), .Y(n1782) );
  OAI21X1 U826 ( .A(n243), .B(n4685), .C(n1305), .Y(n1783) );
  OAI21X1 U828 ( .A(n245), .B(n4685), .C(n1302), .Y(n1784) );
  OAI21X1 U830 ( .A(n247), .B(n4685), .C(n1299), .Y(n1785) );
  OAI21X1 U832 ( .A(n249), .B(n4685), .C(n1296), .Y(n1786) );
  OAI21X1 U835 ( .A(n219), .B(n4682), .C(n1293), .Y(n1787) );
  OAI21X1 U837 ( .A(n221), .B(n4682), .C(n1290), .Y(n1788) );
  OAI21X1 U839 ( .A(n223), .B(n4682), .C(n1287), .Y(n1789) );
  OAI21X1 U841 ( .A(n225), .B(n4682), .C(n1284), .Y(n1790) );
  OAI21X1 U843 ( .A(n227), .B(n4682), .C(n1281), .Y(n1791) );
  OAI21X1 U845 ( .A(n229), .B(n4682), .C(n1278), .Y(n1792) );
  OAI21X1 U847 ( .A(n231), .B(n4682), .C(n1275), .Y(n1793) );
  OAI21X1 U849 ( .A(n233), .B(n4682), .C(n1272), .Y(n1794) );
  OAI21X1 U851 ( .A(n235), .B(n4682), .C(n1269), .Y(n1795) );
  OAI21X1 U853 ( .A(n237), .B(n4682), .C(n1266), .Y(n1796) );
  OAI21X1 U855 ( .A(n239), .B(n4682), .C(n1263), .Y(n1797) );
  OAI21X1 U857 ( .A(n241), .B(n4682), .C(n1260), .Y(n1798) );
  OAI21X1 U859 ( .A(n243), .B(n4682), .C(n1257), .Y(n1799) );
  OAI21X1 U861 ( .A(n245), .B(n4682), .C(n1254), .Y(n1800) );
  OAI21X1 U863 ( .A(n247), .B(n4682), .C(n1251), .Y(n1801) );
  OAI21X1 U865 ( .A(n249), .B(n4682), .C(n1248), .Y(n1802) );
  INVX1 U868 ( .A(n655), .Y(n535) );
  NAND3X1 U869 ( .A(n201), .B(n204), .C(n4639), .Y(n655) );
  INVX1 U870 ( .A(n4642), .Y(n204) );
  OAI21X1 U871 ( .A(n219), .B(n4679), .C(n1245), .Y(n1803) );
  OAI21X1 U873 ( .A(n221), .B(n4679), .C(n1242), .Y(n1804) );
  OAI21X1 U875 ( .A(n223), .B(n4679), .C(n1239), .Y(n1805) );
  OAI21X1 U877 ( .A(n225), .B(n4679), .C(n1236), .Y(n1806) );
  OAI21X1 U879 ( .A(n227), .B(n4679), .C(n1233), .Y(n1807) );
  OAI21X1 U881 ( .A(n229), .B(n4679), .C(n1230), .Y(n1808) );
  OAI21X1 U883 ( .A(n231), .B(n4679), .C(n1227), .Y(n1809) );
  OAI21X1 U885 ( .A(n233), .B(n4679), .C(n1224), .Y(n1810) );
  OAI21X1 U887 ( .A(n235), .B(n4679), .C(n1221), .Y(n1811) );
  OAI21X1 U889 ( .A(n237), .B(n4679), .C(n1218), .Y(n1812) );
  OAI21X1 U891 ( .A(n239), .B(n4679), .C(n1215), .Y(n1813) );
  OAI21X1 U893 ( .A(n241), .B(n4679), .C(n1212), .Y(n1814) );
  OAI21X1 U895 ( .A(n243), .B(n4679), .C(n1209), .Y(n1815) );
  OAI21X1 U897 ( .A(n245), .B(n4679), .C(n1206), .Y(n1816) );
  OAI21X1 U899 ( .A(n247), .B(n4679), .C(n1203), .Y(n1817) );
  OAI21X1 U901 ( .A(n249), .B(n4679), .C(n1200), .Y(n1818) );
  NOR3X1 U904 ( .A(n4633), .B(n4636), .C(n4645), .Y(n251) );
  OAI21X1 U905 ( .A(n219), .B(n4676), .C(n1197), .Y(n1819) );
  OAI21X1 U907 ( .A(n221), .B(n4676), .C(n1194), .Y(n1820) );
  OAI21X1 U909 ( .A(n223), .B(n4676), .C(n1191), .Y(n1821) );
  OAI21X1 U911 ( .A(n225), .B(n4676), .C(n1188), .Y(n1822) );
  OAI21X1 U913 ( .A(n227), .B(n4676), .C(n1185), .Y(n1823) );
  OAI21X1 U915 ( .A(n229), .B(n4676), .C(n1182), .Y(n1824) );
  OAI21X1 U917 ( .A(n231), .B(n4676), .C(n1179), .Y(n1825) );
  OAI21X1 U919 ( .A(n233), .B(n4676), .C(n1176), .Y(n1826) );
  OAI21X1 U921 ( .A(n235), .B(n4676), .C(n1173), .Y(n1827) );
  OAI21X1 U923 ( .A(n237), .B(n4676), .C(n1170), .Y(n1828) );
  OAI21X1 U925 ( .A(n239), .B(n4676), .C(n1167), .Y(n1829) );
  OAI21X1 U927 ( .A(n241), .B(n4676), .C(n1164), .Y(n1830) );
  OAI21X1 U929 ( .A(n243), .B(n4676), .C(n1161), .Y(n1831) );
  OAI21X1 U931 ( .A(n245), .B(n4676), .C(n1158), .Y(n1832) );
  OAI21X1 U933 ( .A(n247), .B(n4676), .C(n1155), .Y(n1833) );
  OAI21X1 U935 ( .A(n249), .B(n4676), .C(n1152), .Y(n1834) );
  NOR3X1 U938 ( .A(n4633), .B(n4636), .C(n210), .Y(n270) );
  OAI21X1 U939 ( .A(n219), .B(n4673), .C(n1149), .Y(n1835) );
  OAI21X1 U941 ( .A(n221), .B(n4673), .C(n1146), .Y(n1836) );
  OAI21X1 U943 ( .A(n223), .B(n4673), .C(n1143), .Y(n1837) );
  OAI21X1 U945 ( .A(n225), .B(n4673), .C(n1140), .Y(n1838) );
  OAI21X1 U947 ( .A(n227), .B(n4673), .C(n1137), .Y(n1839) );
  OAI21X1 U949 ( .A(n229), .B(n4673), .C(n1134), .Y(n1840) );
  OAI21X1 U951 ( .A(n231), .B(n4673), .C(n1131), .Y(n1841) );
  OAI21X1 U953 ( .A(n233), .B(n4673), .C(n1128), .Y(n1842) );
  OAI21X1 U955 ( .A(n235), .B(n4673), .C(n1125), .Y(n1843) );
  OAI21X1 U957 ( .A(n237), .B(n4673), .C(n1122), .Y(n1844) );
  OAI21X1 U959 ( .A(n239), .B(n4673), .C(n1119), .Y(n1845) );
  OAI21X1 U961 ( .A(n241), .B(n4673), .C(n1116), .Y(n1846) );
  OAI21X1 U963 ( .A(n243), .B(n4673), .C(n1113), .Y(n1847) );
  OAI21X1 U965 ( .A(n245), .B(n4673), .C(n1110), .Y(n1848) );
  OAI21X1 U967 ( .A(n247), .B(n4673), .C(n1107), .Y(n1849) );
  OAI21X1 U969 ( .A(n249), .B(n4673), .C(n1104), .Y(n1850) );
  OAI21X1 U973 ( .A(n219), .B(n4670), .C(n1101), .Y(n1851) );
  OAI21X1 U975 ( .A(n221), .B(n4670), .C(n1098), .Y(n1852) );
  OAI21X1 U977 ( .A(n223), .B(n4670), .C(n1095), .Y(n1853) );
  OAI21X1 U979 ( .A(n225), .B(n4670), .C(n1092), .Y(n1854) );
  OAI21X1 U981 ( .A(n227), .B(n4670), .C(n1089), .Y(n1855) );
  OAI21X1 U983 ( .A(n229), .B(n4670), .C(n1086), .Y(n1856) );
  OAI21X1 U985 ( .A(n231), .B(n4670), .C(n1083), .Y(n1857) );
  OAI21X1 U987 ( .A(n233), .B(n4670), .C(n1080), .Y(n1858) );
  OAI21X1 U989 ( .A(n235), .B(n4670), .C(n1077), .Y(n1859) );
  OAI21X1 U991 ( .A(n237), .B(n4670), .C(n1074), .Y(n1860) );
  OAI21X1 U993 ( .A(n239), .B(n4670), .C(n1071), .Y(n1861) );
  OAI21X1 U995 ( .A(n241), .B(n4670), .C(n1068), .Y(n1862) );
  OAI21X1 U997 ( .A(n243), .B(n4670), .C(n1065), .Y(n1863) );
  OAI21X1 U999 ( .A(n245), .B(n4670), .C(n1062), .Y(n1864) );
  OAI21X1 U1001 ( .A(n247), .B(n4670), .C(n1059), .Y(n1865) );
  OAI21X1 U1003 ( .A(n249), .B(n4670), .C(n1056), .Y(n1866) );
  OAI21X1 U1007 ( .A(n219), .B(n4667), .C(n1053), .Y(n1867) );
  OAI21X1 U1009 ( .A(n221), .B(n4667), .C(n1050), .Y(n1868) );
  OAI21X1 U1011 ( .A(n223), .B(n4667), .C(n1047), .Y(n1869) );
  OAI21X1 U1013 ( .A(n225), .B(n4667), .C(n1044), .Y(n1870) );
  OAI21X1 U1015 ( .A(n227), .B(n4667), .C(n1041), .Y(n1871) );
  OAI21X1 U1017 ( .A(n229), .B(n4667), .C(n1038), .Y(n1872) );
  OAI21X1 U1019 ( .A(n231), .B(n4667), .C(n1035), .Y(n1873) );
  OAI21X1 U1021 ( .A(n233), .B(n4667), .C(n1032), .Y(n1874) );
  OAI21X1 U1023 ( .A(n235), .B(n4667), .C(n1029), .Y(n1875) );
  OAI21X1 U1025 ( .A(n237), .B(n4667), .C(n1026), .Y(n1876) );
  OAI21X1 U1027 ( .A(n239), .B(n4667), .C(n1023), .Y(n1877) );
  OAI21X1 U1029 ( .A(n241), .B(n4667), .C(n1020), .Y(n1878) );
  OAI21X1 U1031 ( .A(n243), .B(n4667), .C(n1017), .Y(n1879) );
  OAI21X1 U1033 ( .A(n245), .B(n4667), .C(n1014), .Y(n1880) );
  OAI21X1 U1035 ( .A(n247), .B(n4667), .C(n1011), .Y(n1881) );
  OAI21X1 U1037 ( .A(n249), .B(n4667), .C(n1008), .Y(n1882) );
  OAI21X1 U1041 ( .A(n219), .B(n4664), .C(n1005), .Y(n1883) );
  OAI21X1 U1043 ( .A(n221), .B(n4664), .C(n1002), .Y(n1884) );
  OAI21X1 U1045 ( .A(n223), .B(n4664), .C(n999), .Y(n1885) );
  OAI21X1 U1047 ( .A(n225), .B(n4664), .C(n996), .Y(n1886) );
  OAI21X1 U1049 ( .A(n227), .B(n4664), .C(n993), .Y(n1887) );
  OAI21X1 U1051 ( .A(n229), .B(n4664), .C(n990), .Y(n1888) );
  OAI21X1 U1053 ( .A(n231), .B(n4664), .C(n987), .Y(n1889) );
  OAI21X1 U1055 ( .A(n233), .B(n4664), .C(n984), .Y(n1890) );
  OAI21X1 U1057 ( .A(n235), .B(n4664), .C(n981), .Y(n1891) );
  OAI21X1 U1059 ( .A(n237), .B(n4664), .C(n978), .Y(n1892) );
  OAI21X1 U1061 ( .A(n239), .B(n4664), .C(n975), .Y(n1893) );
  OAI21X1 U1063 ( .A(n241), .B(n4664), .C(n972), .Y(n1894) );
  OAI21X1 U1065 ( .A(n243), .B(n4664), .C(n969), .Y(n1895) );
  OAI21X1 U1067 ( .A(n245), .B(n4664), .C(n966), .Y(n1896) );
  OAI21X1 U1069 ( .A(n247), .B(n4664), .C(n963), .Y(n1897) );
  OAI21X1 U1071 ( .A(n249), .B(n4664), .C(n960), .Y(n1898) );
  OAI21X1 U1075 ( .A(n219), .B(n4661), .C(n957), .Y(n1899) );
  OAI21X1 U1077 ( .A(n221), .B(n4661), .C(n954), .Y(n1900) );
  OAI21X1 U1079 ( .A(n223), .B(n4661), .C(n951), .Y(n1901) );
  OAI21X1 U1081 ( .A(n225), .B(n4661), .C(n948), .Y(n1902) );
  OAI21X1 U1083 ( .A(n227), .B(n4661), .C(n945), .Y(n1903) );
  OAI21X1 U1085 ( .A(n229), .B(n4661), .C(n942), .Y(n1904) );
  OAI21X1 U1087 ( .A(n231), .B(n4661), .C(n939), .Y(n1905) );
  OAI21X1 U1089 ( .A(n233), .B(n4661), .C(n936), .Y(n1906) );
  OAI21X1 U1091 ( .A(n235), .B(n4661), .C(n933), .Y(n1907) );
  OAI21X1 U1093 ( .A(n237), .B(n4661), .C(n930), .Y(n1908) );
  OAI21X1 U1095 ( .A(n239), .B(n4661), .C(n927), .Y(n1909) );
  OAI21X1 U1097 ( .A(n241), .B(n4661), .C(n924), .Y(n1910) );
  OAI21X1 U1099 ( .A(n243), .B(n4661), .C(n921), .Y(n1911) );
  OAI21X1 U1101 ( .A(n245), .B(n4661), .C(n918), .Y(n1912) );
  OAI21X1 U1103 ( .A(n247), .B(n4661), .C(n915), .Y(n1913) );
  OAI21X1 U1105 ( .A(n249), .B(n4661), .C(n912), .Y(n1914) );
  NOR3X1 U1108 ( .A(n206), .B(n4646), .C(n208), .Y(n360) );
  OAI21X1 U1109 ( .A(n219), .B(n4658), .C(n909), .Y(n1915) );
  INVX1 U1111 ( .A(data_in[15]), .Y(n219) );
  OAI21X1 U1112 ( .A(n221), .B(n4658), .C(n906), .Y(n1916) );
  INVX1 U1114 ( .A(data_in[14]), .Y(n221) );
  OAI21X1 U1115 ( .A(n223), .B(n4658), .C(n903), .Y(n1917) );
  INVX1 U1117 ( .A(data_in[13]), .Y(n223) );
  OAI21X1 U1118 ( .A(n225), .B(n4658), .C(n900), .Y(n1918) );
  INVX1 U1120 ( .A(data_in[12]), .Y(n225) );
  OAI21X1 U1121 ( .A(n227), .B(n4658), .C(n897), .Y(n1919) );
  INVX1 U1123 ( .A(data_in[11]), .Y(n227) );
  OAI21X1 U1124 ( .A(n229), .B(n4658), .C(n894), .Y(n1920) );
  INVX1 U1126 ( .A(data_in[10]), .Y(n229) );
  OAI21X1 U1127 ( .A(n231), .B(n4658), .C(n891), .Y(n1921) );
  INVX1 U1129 ( .A(data_in[9]), .Y(n231) );
  OAI21X1 U1130 ( .A(n233), .B(n4658), .C(n888), .Y(n1922) );
  INVX1 U1132 ( .A(data_in[8]), .Y(n233) );
  OAI21X1 U1133 ( .A(n235), .B(n4658), .C(n885), .Y(n1923) );
  INVX1 U1135 ( .A(data_in[7]), .Y(n235) );
  OAI21X1 U1136 ( .A(n237), .B(n4658), .C(n882), .Y(n1924) );
  INVX1 U1138 ( .A(data_in[6]), .Y(n237) );
  OAI21X1 U1139 ( .A(n239), .B(n4658), .C(n879), .Y(n1925) );
  INVX1 U1141 ( .A(data_in[5]), .Y(n239) );
  OAI21X1 U1142 ( .A(n241), .B(n4658), .C(n876), .Y(n1926) );
  INVX1 U1144 ( .A(data_in[4]), .Y(n241) );
  OAI21X1 U1145 ( .A(n243), .B(n4658), .C(n873), .Y(n1927) );
  INVX1 U1147 ( .A(data_in[3]), .Y(n243) );
  OAI21X1 U1148 ( .A(n245), .B(n4658), .C(n870), .Y(n1928) );
  INVX1 U1150 ( .A(data_in[2]), .Y(n245) );
  OAI21X1 U1151 ( .A(n247), .B(n4658), .C(n867), .Y(n1929) );
  INVX1 U1153 ( .A(data_in[1]), .Y(n247) );
  OAI21X1 U1154 ( .A(n249), .B(n4658), .C(n864), .Y(n1930) );
  NOR3X1 U1157 ( .A(n208), .B(n206), .C(n210), .Y(n378) );
  INVX1 U1158 ( .A(n4645), .Y(n210) );
  INVX1 U1159 ( .A(n795), .Y(n673) );
  NAND3X1 U1160 ( .A(n4639), .B(n201), .C(n4642), .Y(n795) );
  INVX1 U1162 ( .A(data_in[0]), .Y(n249) );
  XOR2X1 U1163 ( .A(n4633), .B(n4645), .Y(n24) );
  INVX1 U1166 ( .A(n4636), .Y(n206) );
  INVX1 U1168 ( .A(n4633), .Y(n208) );
  XOR2X1 U1169 ( .A(n4642), .B(n4636), .Y(n22) );
  XOR2X1 U1170 ( .A(n4639), .B(n4642), .Y(n21) );
  XOR2X1 U1171 ( .A(n4630), .B(n4639), .Y(n20) );
  XOR2X1 U1172 ( .A(n5285), .B(n5298), .Y(n19) );
  XOR2X1 U1173 ( .A(n5275), .B(n5285), .Y(n18) );
  XOR2X1 U1174 ( .A(n4751), .B(n5275), .Y(n17) );
  XOR2X1 U1175 ( .A(n4652), .B(n4751), .Y(n16) );
  XOR2X1 U1176 ( .A(n4627), .B(n4652), .Y(n15) );
  NAND3X1 U1177 ( .A(n3036), .B(fillcount[5]), .C(n797), .Y(n5821) );
  NOR3X1 U1178 ( .A(fillcount[2]), .B(fillcount[4]), .C(fillcount[3]), .Y(n797) );
  NAND3X1 U1180 ( .A(n140), .B(n799), .C(n3042), .Y(n5820) );
  XOR2X1 U1182 ( .A(n4652), .B(n803), .Y(n802) );
  XOR2X1 U1183 ( .A(n4751), .B(n804), .Y(n801) );
  XOR2X1 U1184 ( .A(n214), .B(n4609), .Y(n799) );
  INVX1 U1185 ( .A(n4627), .Y(n214) );
  AOI22X1 U1186 ( .A(n805), .B(n143), .C(n807), .D(n3039), .Y(n798) );
  NAND3X1 U1187 ( .A(n809), .B(n180), .C(n810), .Y(n808) );
  XOR2X1 U1188 ( .A(n5319), .B(n811), .Y(n810) );
  INVX1 U1190 ( .A(n5275), .Y(n180) );
  XOR2X1 U1191 ( .A(n4624), .B(n5295), .Y(n809) );
  NAND3X1 U1193 ( .A(n812), .B(n813), .C(n5275), .Y(n806) );
  XOR2X1 U1194 ( .A(n4624), .B(n5285), .Y(n813) );
  XOR2X1 U1195 ( .A(n5298), .B(n811), .Y(n812) );
  XOR2X1 U1196 ( .A(n4624), .B(n3060), .Y(n811) );
  INVX1 U1197 ( .A(n807), .Y(n805) );
  XNOR2X1 U1198 ( .A(n804), .B(n3048), .Y(n807) );
  XOR2X1 U1199 ( .A(n803), .B(n3057), .Y(n804) );
  XOR2X1 U1200 ( .A(n4609), .B(n3054), .Y(n803) );
  HAX1 add_176_U1_1_1 ( .A(n5285), .B(n5313), .YC(add_176_carry[2]), .YS(n88)
         );
  HAX1 add_176_U1_1_2 ( .A(n5275), .B(add_176_carry[2]), .YC(add_176_carry[3]), 
        .YS(n89) );
  HAX1 add_176_U1_1_3 ( .A(n4751), .B(add_176_carry[3]), .YC(add_176_carry[4]), 
        .YS(n90) );
  HAX1 add_176_U1_1_4 ( .A(n4652), .B(add_176_carry[4]), .YC(add_176_carry[5]), 
        .YS(n91) );
  HAX1 add_158_U1_1_1 ( .A(n4633), .B(n4646), .YC(add_158_carry[2]), .YS(n34)
         );
  HAX1 add_158_U1_1_2 ( .A(n4636), .B(add_158_carry[2]), .YC(add_158_carry[3]), 
        .YS(n35) );
  HAX1 add_158_U1_1_3 ( .A(n4642), .B(add_158_carry[3]), .YC(add_158_carry[4]), 
        .YS(n36) );
  HAX1 add_158_U1_1_4 ( .A(n4639), .B(add_158_carry[4]), .YC(add_158_carry[5]), 
        .YS(n37) );
  FAX1 r301_U2_1 ( .A(n4633), .B(r301_B_not_1_), .C(r301_carry[1]), .YC(
        r301_carry[2]), .YS(fillcount[1]) );
  FAX1 r301_U2_2 ( .A(n4636), .B(r301_B_not_2_), .C(r301_carry[2]), .YC(
        r301_carry[3]), .YS(fillcount[2]) );
  FAX1 r301_U2_3 ( .A(n4642), .B(r301_B_not_3_), .C(r301_carry[3]), .YC(
        r301_carry[4]), .YS(fillcount[3]) );
  FAX1 r301_U2_4 ( .A(n4639), .B(r301_B_not_4_), .C(r301_carry[4]), .YC(
        r301_carry[5]), .YS(fillcount[4]) );
  FAX1 r301_U2_5 ( .A(n4630), .B(r301_B_not_5_), .C(r301_carry[5]), .YC(), 
        .YS(fillcount[5]) );
  DFFSR fifo_reg_0__15_ ( .D(n1419), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[511]) );
  DFFSR fifo_reg_0__14_ ( .D(n1420), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[510]) );
  DFFSR fifo_reg_0__13_ ( .D(n1421), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[509]) );
  DFFSR fifo_reg_0__12_ ( .D(n1422), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[508]) );
  DFFSR fifo_reg_0__11_ ( .D(n1423), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[507]) );
  DFFSR fifo_reg_0__10_ ( .D(n1424), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[506]) );
  DFFSR fifo_reg_0__9_ ( .D(n1425), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[505]) );
  DFFSR fifo_reg_0__8_ ( .D(n1426), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[504]) );
  DFFSR fifo_reg_0__7_ ( .D(n1427), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[503]) );
  DFFSR fifo_reg_0__6_ ( .D(n1428), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[502]) );
  DFFSR fifo_reg_0__5_ ( .D(n1429), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[501]) );
  DFFSR fifo_reg_0__4_ ( .D(n1430), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[500]) );
  DFFSR fifo_reg_0__3_ ( .D(n1431), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[499]) );
  DFFSR fifo_reg_0__2_ ( .D(n1432), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[498]) );
  DFFSR fifo_reg_0__1_ ( .D(n1433), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[497]) );
  DFFSR fifo_reg_0__0_ ( .D(n1434), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[496]) );
  DFFSR fifo_reg_7__15_ ( .D(n1531), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[399]) );
  DFFSR fifo_reg_7__14_ ( .D(n1532), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[398]) );
  DFFSR fifo_reg_7__13_ ( .D(n1533), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[397]) );
  DFFSR fifo_reg_7__12_ ( .D(n1534), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[396]) );
  DFFSR fifo_reg_7__11_ ( .D(n1535), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[395]) );
  DFFSR fifo_reg_7__10_ ( .D(n1536), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[394]) );
  DFFSR fifo_reg_7__9_ ( .D(n1537), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[393]) );
  DFFSR fifo_reg_7__8_ ( .D(n1538), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[392]) );
  DFFSR fifo_reg_7__7_ ( .D(n1539), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[391]) );
  DFFSR fifo_reg_7__6_ ( .D(n1540), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[390]) );
  DFFSR fifo_reg_7__5_ ( .D(n1541), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[389]) );
  DFFSR fifo_reg_7__4_ ( .D(n1542), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[388]) );
  DFFSR fifo_reg_7__3_ ( .D(n1543), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[387]) );
  DFFSR fifo_reg_7__2_ ( .D(n1544), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[386]) );
  DFFSR fifo_reg_7__1_ ( .D(n1545), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[385]) );
  DFFSR fifo_reg_7__0_ ( .D(n1546), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[384]) );
  DFFSR fifo_reg_6__15_ ( .D(n1515), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[415]) );
  DFFSR fifo_reg_6__14_ ( .D(n1516), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[414]) );
  DFFSR fifo_reg_6__13_ ( .D(n1517), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[413]) );
  DFFSR fifo_reg_6__12_ ( .D(n1518), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[412]) );
  DFFSR fifo_reg_6__11_ ( .D(n1519), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[411]) );
  DFFSR fifo_reg_6__10_ ( .D(n1520), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[410]) );
  DFFSR fifo_reg_6__9_ ( .D(n1521), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[409]) );
  DFFSR fifo_reg_6__8_ ( .D(n1522), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[408]) );
  DFFSR fifo_reg_6__7_ ( .D(n1523), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[407]) );
  DFFSR fifo_reg_6__6_ ( .D(n1524), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[406]) );
  DFFSR fifo_reg_6__5_ ( .D(n1525), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[405]) );
  DFFSR fifo_reg_6__4_ ( .D(n1526), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[404]) );
  DFFSR fifo_reg_6__3_ ( .D(n1527), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[403]) );
  DFFSR fifo_reg_6__2_ ( .D(n1528), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[402]) );
  DFFSR fifo_reg_6__1_ ( .D(n1529), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[401]) );
  DFFSR fifo_reg_6__0_ ( .D(n1530), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[400]) );
  DFFSR fifo_reg_5__15_ ( .D(n1499), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[431]) );
  DFFSR fifo_reg_5__14_ ( .D(n1500), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[430]) );
  DFFSR fifo_reg_5__13_ ( .D(n1501), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[429]) );
  DFFSR fifo_reg_5__12_ ( .D(n1502), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[428]) );
  DFFSR fifo_reg_5__11_ ( .D(n1503), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[427]) );
  DFFSR fifo_reg_5__10_ ( .D(n1504), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[426]) );
  DFFSR fifo_reg_5__9_ ( .D(n1505), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[425]) );
  DFFSR fifo_reg_5__8_ ( .D(n1506), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[424]) );
  DFFSR fifo_reg_5__7_ ( .D(n1507), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[423]) );
  DFFSR fifo_reg_5__6_ ( .D(n1508), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[422]) );
  DFFSR fifo_reg_5__5_ ( .D(n1509), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[421]) );
  DFFSR fifo_reg_5__4_ ( .D(n1510), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[420]) );
  DFFSR fifo_reg_5__3_ ( .D(n1511), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[419]) );
  DFFSR fifo_reg_5__2_ ( .D(n1512), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[418]) );
  DFFSR fifo_reg_5__1_ ( .D(n1513), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[417]) );
  DFFSR fifo_reg_5__0_ ( .D(n1514), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[416]) );
  DFFSR fifo_reg_4__15_ ( .D(n1483), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[447]) );
  DFFSR fifo_reg_4__14_ ( .D(n1484), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[446]) );
  DFFSR fifo_reg_4__13_ ( .D(n1485), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[445]) );
  DFFSR fifo_reg_4__12_ ( .D(n1486), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[444]) );
  DFFSR fifo_reg_4__11_ ( .D(n1487), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[443]) );
  DFFSR fifo_reg_4__10_ ( .D(n1488), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[442]) );
  DFFSR fifo_reg_4__9_ ( .D(n1489), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[441]) );
  DFFSR fifo_reg_4__8_ ( .D(n1490), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[440]) );
  DFFSR fifo_reg_4__7_ ( .D(n1491), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[439]) );
  DFFSR fifo_reg_4__6_ ( .D(n1492), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[438]) );
  DFFSR fifo_reg_4__5_ ( .D(n1493), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[437]) );
  DFFSR fifo_reg_4__4_ ( .D(n1494), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[436]) );
  DFFSR fifo_reg_4__3_ ( .D(n1495), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[435]) );
  DFFSR fifo_reg_4__2_ ( .D(n1496), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[434]) );
  DFFSR fifo_reg_4__1_ ( .D(n1497), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[433]) );
  DFFSR fifo_reg_4__0_ ( .D(n1498), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[432]) );
  DFFSR fifo_reg_3__15_ ( .D(n1467), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[463]) );
  DFFSR fifo_reg_3__14_ ( .D(n1468), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[462]) );
  DFFSR fifo_reg_3__13_ ( .D(n1469), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[461]) );
  DFFSR fifo_reg_3__12_ ( .D(n1470), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[460]) );
  DFFSR fifo_reg_3__11_ ( .D(n1471), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[459]) );
  DFFSR fifo_reg_3__10_ ( .D(n1472), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[458]) );
  DFFSR fifo_reg_3__9_ ( .D(n1473), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[457]) );
  DFFSR fifo_reg_3__8_ ( .D(n1474), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[456]) );
  DFFSR fifo_reg_3__7_ ( .D(n1475), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[455]) );
  DFFSR fifo_reg_3__6_ ( .D(n1476), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[454]) );
  DFFSR fifo_reg_3__5_ ( .D(n1477), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[453]) );
  DFFSR fifo_reg_3__4_ ( .D(n1478), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[452]) );
  DFFSR fifo_reg_3__3_ ( .D(n1479), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[451]) );
  DFFSR fifo_reg_3__2_ ( .D(n1480), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[450]) );
  DFFSR fifo_reg_3__1_ ( .D(n1481), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[449]) );
  DFFSR fifo_reg_3__0_ ( .D(n1482), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[448]) );
  DFFSR fifo_reg_2__15_ ( .D(n1451), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[479]) );
  DFFSR fifo_reg_2__14_ ( .D(n1452), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[478]) );
  DFFSR fifo_reg_2__13_ ( .D(n1453), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[477]) );
  DFFSR fifo_reg_2__12_ ( .D(n1454), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[476]) );
  DFFSR fifo_reg_2__11_ ( .D(n1455), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[475]) );
  DFFSR fifo_reg_2__10_ ( .D(n1456), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[474]) );
  DFFSR fifo_reg_2__9_ ( .D(n1457), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[473]) );
  DFFSR fifo_reg_2__8_ ( .D(n1458), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[472]) );
  DFFSR fifo_reg_2__7_ ( .D(n1459), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[471]) );
  DFFSR fifo_reg_2__6_ ( .D(n1460), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[470]) );
  DFFSR fifo_reg_2__5_ ( .D(n1461), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[469]) );
  DFFSR fifo_reg_2__4_ ( .D(n1462), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[468]) );
  DFFSR fifo_reg_2__3_ ( .D(n1463), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[467]) );
  DFFSR fifo_reg_2__2_ ( .D(n1464), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[466]) );
  DFFSR fifo_reg_2__1_ ( .D(n1465), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[465]) );
  DFFSR fifo_reg_2__0_ ( .D(n1466), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[464]) );
  DFFSR fifo_reg_1__15_ ( .D(n1435), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[495]) );
  DFFSR fifo_reg_1__14_ ( .D(n1436), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[494]) );
  DFFSR fifo_reg_1__13_ ( .D(n1437), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[493]) );
  DFFSR fifo_reg_1__12_ ( .D(n1438), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[492]) );
  DFFSR fifo_reg_1__11_ ( .D(n1439), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[491]) );
  DFFSR fifo_reg_1__10_ ( .D(n1440), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[490]) );
  DFFSR fifo_reg_1__9_ ( .D(n1441), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[489]) );
  DFFSR fifo_reg_1__8_ ( .D(n1442), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[488]) );
  DFFSR fifo_reg_1__7_ ( .D(n1443), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[487]) );
  DFFSR fifo_reg_1__6_ ( .D(n1444), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[486]) );
  DFFSR fifo_reg_1__5_ ( .D(n1445), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[485]) );
  DFFSR fifo_reg_1__4_ ( .D(n1446), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[484]) );
  DFFSR fifo_reg_1__3_ ( .D(n1447), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[483]) );
  DFFSR fifo_reg_1__2_ ( .D(n1448), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[482]) );
  DFFSR fifo_reg_1__1_ ( .D(n1449), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[481]) );
  DFFSR fifo_reg_1__0_ ( .D(n1450), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[480]) );
  DFFSR fifo_reg_25__15_ ( .D(n1819), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[111]) );
  DFFSR fifo_reg_25__14_ ( .D(n1820), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[110]) );
  DFFSR fifo_reg_25__13_ ( .D(n1821), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[109]) );
  DFFSR fifo_reg_25__12_ ( .D(n1822), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[108]) );
  DFFSR fifo_reg_25__11_ ( .D(n1823), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[107]) );
  DFFSR fifo_reg_25__10_ ( .D(n1824), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[106]) );
  DFFSR fifo_reg_25__9_ ( .D(n1825), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[105]) );
  DFFSR fifo_reg_25__8_ ( .D(n1826), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[104]) );
  DFFSR fifo_reg_25__7_ ( .D(n1827), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[103]) );
  DFFSR fifo_reg_25__6_ ( .D(n1828), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[102]) );
  DFFSR fifo_reg_25__5_ ( .D(n1829), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[101]) );
  DFFSR fifo_reg_25__4_ ( .D(n1830), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[100]) );
  DFFSR fifo_reg_25__3_ ( .D(n1831), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[99]) );
  DFFSR fifo_reg_25__2_ ( .D(n1832), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[98]) );
  DFFSR fifo_reg_25__1_ ( .D(n1833), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[97]) );
  DFFSR fifo_reg_25__0_ ( .D(n1834), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[96]) );
  DFFSR fifo_reg_24__15_ ( .D(n1803), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[127]) );
  DFFSR fifo_reg_24__14_ ( .D(n1804), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[126]) );
  DFFSR fifo_reg_24__13_ ( .D(n1805), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[125]) );
  DFFSR fifo_reg_24__12_ ( .D(n1806), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[124]) );
  DFFSR fifo_reg_24__11_ ( .D(n1807), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[123]) );
  DFFSR fifo_reg_24__10_ ( .D(n1808), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[122]) );
  DFFSR fifo_reg_24__9_ ( .D(n1809), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[121]) );
  DFFSR fifo_reg_24__8_ ( .D(n1810), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[120]) );
  DFFSR fifo_reg_24__7_ ( .D(n1811), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[119]) );
  DFFSR fifo_reg_24__6_ ( .D(n1812), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[118]) );
  DFFSR fifo_reg_24__5_ ( .D(n1813), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[117]) );
  DFFSR fifo_reg_24__4_ ( .D(n1814), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[116]) );
  DFFSR fifo_reg_24__3_ ( .D(n1815), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[115]) );
  DFFSR fifo_reg_24__2_ ( .D(n1816), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[114]) );
  DFFSR fifo_reg_24__1_ ( .D(n1817), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[113]) );
  DFFSR fifo_reg_24__0_ ( .D(n1818), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[112]) );
  DFFSR fifo_reg_31__15_ ( .D(n1915), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[15]) );
  DFFSR fifo_reg_31__14_ ( .D(n1916), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[14]) );
  DFFSR fifo_reg_31__13_ ( .D(n1917), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[13]) );
  DFFSR fifo_reg_31__12_ ( .D(n1918), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[12]) );
  DFFSR fifo_reg_31__11_ ( .D(n1919), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[11]) );
  DFFSR fifo_reg_31__10_ ( .D(n1920), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[10]) );
  DFFSR fifo_reg_31__9_ ( .D(n1921), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[9]) );
  DFFSR fifo_reg_31__8_ ( .D(n1922), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[8]) );
  DFFSR fifo_reg_31__7_ ( .D(n1923), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[7]) );
  DFFSR fifo_reg_31__6_ ( .D(n1924), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[6]) );
  DFFSR fifo_reg_31__5_ ( .D(n1925), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[5]) );
  DFFSR fifo_reg_31__4_ ( .D(n1926), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[4]) );
  DFFSR fifo_reg_31__3_ ( .D(n1927), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[3]) );
  DFFSR fifo_reg_31__2_ ( .D(n1928), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[2]) );
  DFFSR fifo_reg_31__1_ ( .D(n1929), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[1]) );
  DFFSR fifo_reg_31__0_ ( .D(n1930), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[0]) );
  DFFSR fifo_reg_30__15_ ( .D(n1899), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[31]) );
  DFFSR fifo_reg_30__14_ ( .D(n1900), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[30]) );
  DFFSR fifo_reg_30__13_ ( .D(n1901), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[29]) );
  DFFSR fifo_reg_30__12_ ( .D(n1902), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[28]) );
  DFFSR fifo_reg_30__11_ ( .D(n1903), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[27]) );
  DFFSR fifo_reg_30__10_ ( .D(n1904), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[26]) );
  DFFSR fifo_reg_30__9_ ( .D(n1905), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[25]) );
  DFFSR fifo_reg_30__8_ ( .D(n1906), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[24]) );
  DFFSR fifo_reg_30__7_ ( .D(n1907), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[23]) );
  DFFSR fifo_reg_30__6_ ( .D(n1908), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[22]) );
  DFFSR fifo_reg_30__5_ ( .D(n1909), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[21]) );
  DFFSR fifo_reg_30__4_ ( .D(n1910), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[20]) );
  DFFSR fifo_reg_30__3_ ( .D(n1911), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[19]) );
  DFFSR fifo_reg_30__2_ ( .D(n1912), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[18]) );
  DFFSR fifo_reg_30__1_ ( .D(n1913), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[17]) );
  DFFSR fifo_reg_30__0_ ( .D(n1914), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[16]) );
  DFFSR fifo_reg_28__15_ ( .D(n1867), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[63]) );
  DFFSR fifo_reg_28__14_ ( .D(n1868), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[62]) );
  DFFSR fifo_reg_28__13_ ( .D(n1869), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[61]) );
  DFFSR fifo_reg_28__12_ ( .D(n1870), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[60]) );
  DFFSR fifo_reg_28__11_ ( .D(n1871), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[59]) );
  DFFSR fifo_reg_28__10_ ( .D(n1872), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[58]) );
  DFFSR fifo_reg_28__9_ ( .D(n1873), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[57]) );
  DFFSR fifo_reg_28__8_ ( .D(n1874), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[56]) );
  DFFSR fifo_reg_28__7_ ( .D(n1875), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[55]) );
  DFFSR fifo_reg_28__6_ ( .D(n1876), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[54]) );
  DFFSR fifo_reg_28__5_ ( .D(n1877), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[53]) );
  DFFSR fifo_reg_28__4_ ( .D(n1878), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[52]) );
  DFFSR fifo_reg_28__3_ ( .D(n1879), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[51]) );
  DFFSR fifo_reg_28__2_ ( .D(n1880), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[50]) );
  DFFSR fifo_reg_28__1_ ( .D(n1881), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[49]) );
  DFFSR fifo_reg_28__0_ ( .D(n1882), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[48]) );
  DFFSR fifo_reg_26__15_ ( .D(n1835), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[95]) );
  DFFSR fifo_reg_26__14_ ( .D(n1836), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[94]) );
  DFFSR fifo_reg_26__13_ ( .D(n1837), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[93]) );
  DFFSR fifo_reg_26__12_ ( .D(n1838), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[92]) );
  DFFSR fifo_reg_26__11_ ( .D(n1839), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[91]) );
  DFFSR fifo_reg_26__10_ ( .D(n1840), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[90]) );
  DFFSR fifo_reg_26__9_ ( .D(n1841), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[89]) );
  DFFSR fifo_reg_26__8_ ( .D(n1842), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[88]) );
  DFFSR fifo_reg_26__7_ ( .D(n1843), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[87]) );
  DFFSR fifo_reg_26__6_ ( .D(n1844), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[86]) );
  DFFSR fifo_reg_26__5_ ( .D(n1845), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[85]) );
  DFFSR fifo_reg_26__4_ ( .D(n1846), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[84]) );
  DFFSR fifo_reg_26__3_ ( .D(n1847), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[83]) );
  DFFSR fifo_reg_26__2_ ( .D(n1848), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[82]) );
  DFFSR fifo_reg_26__1_ ( .D(n1849), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[81]) );
  DFFSR fifo_reg_26__0_ ( .D(n1850), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[80]) );
  DFFSR fifo_reg_29__15_ ( .D(n1883), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[47]) );
  DFFSR fifo_reg_29__14_ ( .D(n1884), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[46]) );
  DFFSR fifo_reg_29__13_ ( .D(n1885), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[45]) );
  DFFSR fifo_reg_29__12_ ( .D(n1886), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[44]) );
  DFFSR fifo_reg_29__11_ ( .D(n1887), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[43]) );
  DFFSR fifo_reg_29__10_ ( .D(n1888), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[42]) );
  DFFSR fifo_reg_29__9_ ( .D(n1889), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[41]) );
  DFFSR fifo_reg_29__8_ ( .D(n1890), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[40]) );
  DFFSR fifo_reg_29__7_ ( .D(n1891), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[39]) );
  DFFSR fifo_reg_29__6_ ( .D(n1892), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[38]) );
  DFFSR fifo_reg_29__5_ ( .D(n1893), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[37]) );
  DFFSR fifo_reg_29__4_ ( .D(n1894), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[36]) );
  DFFSR fifo_reg_29__3_ ( .D(n1895), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[35]) );
  DFFSR fifo_reg_29__2_ ( .D(n1896), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[34]) );
  DFFSR fifo_reg_29__1_ ( .D(n1897), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[33]) );
  DFFSR fifo_reg_29__0_ ( .D(n1898), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[32]) );
  DFFSR fifo_reg_27__15_ ( .D(n1851), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[79]) );
  DFFSR fifo_reg_27__14_ ( .D(n1852), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[78]) );
  DFFSR fifo_reg_27__13_ ( .D(n1853), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[77]) );
  DFFSR fifo_reg_27__12_ ( .D(n1854), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[76]) );
  DFFSR fifo_reg_27__11_ ( .D(n1855), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[75]) );
  DFFSR fifo_reg_27__10_ ( .D(n1856), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[74]) );
  DFFSR fifo_reg_27__9_ ( .D(n1857), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[73]) );
  DFFSR fifo_reg_27__8_ ( .D(n1858), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[72]) );
  DFFSR fifo_reg_27__7_ ( .D(n1859), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[71]) );
  DFFSR fifo_reg_27__6_ ( .D(n1860), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[70]) );
  DFFSR fifo_reg_27__5_ ( .D(n1861), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[69]) );
  DFFSR fifo_reg_27__4_ ( .D(n1862), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[68]) );
  DFFSR fifo_reg_27__3_ ( .D(n1863), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[67]) );
  DFFSR fifo_reg_27__2_ ( .D(n1864), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[66]) );
  DFFSR fifo_reg_27__1_ ( .D(n1865), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[65]) );
  DFFSR fifo_reg_27__0_ ( .D(n1866), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[64]) );
  DFFSR fifo_reg_9__15_ ( .D(n1563), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[367]) );
  DFFSR fifo_reg_9__14_ ( .D(n1564), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[366]) );
  DFFSR fifo_reg_9__13_ ( .D(n1565), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[365]) );
  DFFSR fifo_reg_9__12_ ( .D(n1566), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[364]) );
  DFFSR fifo_reg_9__11_ ( .D(n1567), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[363]) );
  DFFSR fifo_reg_9__10_ ( .D(n1568), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[362]) );
  DFFSR fifo_reg_9__9_ ( .D(n1569), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[361]) );
  DFFSR fifo_reg_9__8_ ( .D(n1570), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[360]) );
  DFFSR fifo_reg_9__7_ ( .D(n1571), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[359]) );
  DFFSR fifo_reg_9__6_ ( .D(n1572), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[358]) );
  DFFSR fifo_reg_9__5_ ( .D(n1573), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[357]) );
  DFFSR fifo_reg_9__4_ ( .D(n1574), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[356]) );
  DFFSR fifo_reg_9__3_ ( .D(n1575), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[355]) );
  DFFSR fifo_reg_9__2_ ( .D(n1576), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[354]) );
  DFFSR fifo_reg_9__1_ ( .D(n1577), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[353]) );
  DFFSR fifo_reg_9__0_ ( .D(n1578), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[352]) );
  DFFSR fifo_reg_8__15_ ( .D(n1547), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[383]) );
  DFFSR fifo_reg_8__14_ ( .D(n1548), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[382]) );
  DFFSR fifo_reg_8__13_ ( .D(n1549), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[381]) );
  DFFSR fifo_reg_8__12_ ( .D(n1550), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[380]) );
  DFFSR fifo_reg_8__11_ ( .D(n1551), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[379]) );
  DFFSR fifo_reg_8__10_ ( .D(n1552), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[378]) );
  DFFSR fifo_reg_8__9_ ( .D(n1553), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[377]) );
  DFFSR fifo_reg_8__8_ ( .D(n1554), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[376]) );
  DFFSR fifo_reg_8__7_ ( .D(n1555), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[375]) );
  DFFSR fifo_reg_8__6_ ( .D(n1556), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[374]) );
  DFFSR fifo_reg_8__5_ ( .D(n1557), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[373]) );
  DFFSR fifo_reg_8__4_ ( .D(n1558), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[372]) );
  DFFSR fifo_reg_8__3_ ( .D(n1559), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[371]) );
  DFFSR fifo_reg_8__2_ ( .D(n1560), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[370]) );
  DFFSR fifo_reg_8__1_ ( .D(n1561), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[369]) );
  DFFSR fifo_reg_8__0_ ( .D(n1562), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[368]) );
  DFFSR fifo_reg_17__15_ ( .D(n1691), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[239]) );
  DFFSR fifo_reg_17__14_ ( .D(n1692), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[238]) );
  DFFSR fifo_reg_17__13_ ( .D(n1693), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[237]) );
  DFFSR fifo_reg_17__12_ ( .D(n1694), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[236]) );
  DFFSR fifo_reg_17__11_ ( .D(n1695), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[235]) );
  DFFSR fifo_reg_17__10_ ( .D(n1696), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[234]) );
  DFFSR fifo_reg_17__9_ ( .D(n1697), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[233]) );
  DFFSR fifo_reg_17__8_ ( .D(n1698), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[232]) );
  DFFSR fifo_reg_17__7_ ( .D(n1699), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[231]) );
  DFFSR fifo_reg_17__6_ ( .D(n1700), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[230]) );
  DFFSR fifo_reg_17__5_ ( .D(n1701), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[229]) );
  DFFSR fifo_reg_17__4_ ( .D(n1702), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[228]) );
  DFFSR fifo_reg_17__3_ ( .D(n1703), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[227]) );
  DFFSR fifo_reg_17__2_ ( .D(n1704), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[226]) );
  DFFSR fifo_reg_17__1_ ( .D(n1705), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[225]) );
  DFFSR fifo_reg_17__0_ ( .D(n1706), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[224]) );
  DFFSR fifo_reg_16__15_ ( .D(n1675), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[255]) );
  DFFSR fifo_reg_16__14_ ( .D(n1676), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[254]) );
  DFFSR fifo_reg_16__13_ ( .D(n1677), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[253]) );
  DFFSR fifo_reg_16__12_ ( .D(n1678), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[252]) );
  DFFSR fifo_reg_16__11_ ( .D(n1679), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[251]) );
  DFFSR fifo_reg_16__10_ ( .D(n1680), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[250]) );
  DFFSR fifo_reg_16__9_ ( .D(n1681), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[249]) );
  DFFSR fifo_reg_16__8_ ( .D(n1682), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[248]) );
  DFFSR fifo_reg_16__7_ ( .D(n1683), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[247]) );
  DFFSR fifo_reg_16__6_ ( .D(n1684), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[246]) );
  DFFSR fifo_reg_16__5_ ( .D(n1685), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[245]) );
  DFFSR fifo_reg_16__4_ ( .D(n1686), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[244]) );
  DFFSR fifo_reg_16__3_ ( .D(n1687), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[243]) );
  DFFSR fifo_reg_16__2_ ( .D(n1688), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[242]) );
  DFFSR fifo_reg_16__1_ ( .D(n1689), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[241]) );
  DFFSR fifo_reg_16__0_ ( .D(n1690), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[240]) );
  DFFSR fifo_reg_15__15_ ( .D(n1659), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[271]) );
  DFFSR fifo_reg_15__14_ ( .D(n1660), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[270]) );
  DFFSR fifo_reg_15__13_ ( .D(n1661), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[269]) );
  DFFSR fifo_reg_15__12_ ( .D(n1662), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[268]) );
  DFFSR fifo_reg_15__11_ ( .D(n1663), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[267]) );
  DFFSR fifo_reg_15__10_ ( .D(n1664), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[266]) );
  DFFSR fifo_reg_15__9_ ( .D(n1665), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[265]) );
  DFFSR fifo_reg_15__8_ ( .D(n1666), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[264]) );
  DFFSR fifo_reg_15__7_ ( .D(n1667), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[263]) );
  DFFSR fifo_reg_15__6_ ( .D(n1668), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[262]) );
  DFFSR fifo_reg_15__5_ ( .D(n1669), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[261]) );
  DFFSR fifo_reg_15__4_ ( .D(n1670), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[260]) );
  DFFSR fifo_reg_15__3_ ( .D(n1671), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[259]) );
  DFFSR fifo_reg_15__2_ ( .D(n1672), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[258]) );
  DFFSR fifo_reg_15__1_ ( .D(n1673), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[257]) );
  DFFSR fifo_reg_15__0_ ( .D(n1674), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[256]) );
  DFFSR fifo_reg_14__15_ ( .D(n1643), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[287]) );
  DFFSR fifo_reg_14__14_ ( .D(n1644), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[286]) );
  DFFSR fifo_reg_14__13_ ( .D(n1645), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[285]) );
  DFFSR fifo_reg_14__12_ ( .D(n1646), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[284]) );
  DFFSR fifo_reg_14__11_ ( .D(n1647), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[283]) );
  DFFSR fifo_reg_14__10_ ( .D(n1648), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[282]) );
  DFFSR fifo_reg_14__9_ ( .D(n1649), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[281]) );
  DFFSR fifo_reg_14__8_ ( .D(n1650), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[280]) );
  DFFSR fifo_reg_14__7_ ( .D(n1651), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[279]) );
  DFFSR fifo_reg_14__6_ ( .D(n1652), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[278]) );
  DFFSR fifo_reg_14__5_ ( .D(n1653), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[277]) );
  DFFSR fifo_reg_14__4_ ( .D(n1654), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[276]) );
  DFFSR fifo_reg_14__3_ ( .D(n1655), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[275]) );
  DFFSR fifo_reg_14__2_ ( .D(n1656), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[274]) );
  DFFSR fifo_reg_14__1_ ( .D(n1657), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[273]) );
  DFFSR fifo_reg_14__0_ ( .D(n1658), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[272]) );
  DFFSR fifo_reg_23__15_ ( .D(n1787), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[143]) );
  DFFSR fifo_reg_23__14_ ( .D(n1788), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[142]) );
  DFFSR fifo_reg_23__13_ ( .D(n1789), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[141]) );
  DFFSR fifo_reg_23__12_ ( .D(n1790), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[140]) );
  DFFSR fifo_reg_23__11_ ( .D(n1791), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[139]) );
  DFFSR fifo_reg_23__10_ ( .D(n1792), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[138]) );
  DFFSR fifo_reg_23__9_ ( .D(n1793), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[137]) );
  DFFSR fifo_reg_23__8_ ( .D(n1794), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[136]) );
  DFFSR fifo_reg_23__7_ ( .D(n1795), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[135]) );
  DFFSR fifo_reg_23__6_ ( .D(n1796), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[134]) );
  DFFSR fifo_reg_23__5_ ( .D(n1797), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[133]) );
  DFFSR fifo_reg_23__4_ ( .D(n1798), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[132]) );
  DFFSR fifo_reg_23__3_ ( .D(n1799), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[131]) );
  DFFSR fifo_reg_23__2_ ( .D(n1800), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[130]) );
  DFFSR fifo_reg_23__1_ ( .D(n1801), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[129]) );
  DFFSR fifo_reg_23__0_ ( .D(n1802), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[128]) );
  DFFSR fifo_reg_22__15_ ( .D(n1771), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[159]) );
  DFFSR fifo_reg_22__14_ ( .D(n1772), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[158]) );
  DFFSR fifo_reg_22__13_ ( .D(n1773), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[157]) );
  DFFSR fifo_reg_22__12_ ( .D(n1774), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[156]) );
  DFFSR fifo_reg_22__11_ ( .D(n1775), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[155]) );
  DFFSR fifo_reg_22__10_ ( .D(n1776), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[154]) );
  DFFSR fifo_reg_22__9_ ( .D(n1777), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[153]) );
  DFFSR fifo_reg_22__8_ ( .D(n1778), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[152]) );
  DFFSR fifo_reg_22__7_ ( .D(n1779), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[151]) );
  DFFSR fifo_reg_22__6_ ( .D(n1780), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[150]) );
  DFFSR fifo_reg_22__5_ ( .D(n1781), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[149]) );
  DFFSR fifo_reg_22__4_ ( .D(n1782), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[148]) );
  DFFSR fifo_reg_22__3_ ( .D(n1783), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[147]) );
  DFFSR fifo_reg_22__2_ ( .D(n1784), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[146]) );
  DFFSR fifo_reg_22__1_ ( .D(n1785), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[145]) );
  DFFSR fifo_reg_22__0_ ( .D(n1786), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[144]) );
  DFFSR fifo_reg_12__15_ ( .D(n1611), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[319]) );
  DFFSR fifo_reg_12__14_ ( .D(n1612), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[318]) );
  DFFSR fifo_reg_12__13_ ( .D(n1613), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[317]) );
  DFFSR fifo_reg_12__12_ ( .D(n1614), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[316]) );
  DFFSR fifo_reg_12__11_ ( .D(n1615), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[315]) );
  DFFSR fifo_reg_12__10_ ( .D(n1616), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[314]) );
  DFFSR fifo_reg_12__9_ ( .D(n1617), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[313]) );
  DFFSR fifo_reg_12__8_ ( .D(n1618), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[312]) );
  DFFSR fifo_reg_12__7_ ( .D(n1619), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[311]) );
  DFFSR fifo_reg_12__6_ ( .D(n1620), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[310]) );
  DFFSR fifo_reg_12__5_ ( .D(n1621), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[309]) );
  DFFSR fifo_reg_12__4_ ( .D(n1622), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[308]) );
  DFFSR fifo_reg_12__3_ ( .D(n1623), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[307]) );
  DFFSR fifo_reg_12__2_ ( .D(n1624), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[306]) );
  DFFSR fifo_reg_12__1_ ( .D(n1625), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[305]) );
  DFFSR fifo_reg_12__0_ ( .D(n1626), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[304]) );
  DFFSR fifo_reg_10__15_ ( .D(n1579), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[351]) );
  DFFSR fifo_reg_10__14_ ( .D(n1580), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[350]) );
  DFFSR fifo_reg_10__13_ ( .D(n1581), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[349]) );
  DFFSR fifo_reg_10__12_ ( .D(n1582), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[348]) );
  DFFSR fifo_reg_10__11_ ( .D(n1583), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[347]) );
  DFFSR fifo_reg_10__10_ ( .D(n1584), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[346]) );
  DFFSR fifo_reg_10__9_ ( .D(n1585), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[345]) );
  DFFSR fifo_reg_10__8_ ( .D(n1586), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[344]) );
  DFFSR fifo_reg_10__7_ ( .D(n1587), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[343]) );
  DFFSR fifo_reg_10__6_ ( .D(n1588), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[342]) );
  DFFSR fifo_reg_10__5_ ( .D(n1589), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[341]) );
  DFFSR fifo_reg_10__4_ ( .D(n1590), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[340]) );
  DFFSR fifo_reg_10__3_ ( .D(n1591), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[339]) );
  DFFSR fifo_reg_10__2_ ( .D(n1592), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[338]) );
  DFFSR fifo_reg_10__1_ ( .D(n1593), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[337]) );
  DFFSR fifo_reg_10__0_ ( .D(n1594), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[336]) );
  DFFSR fifo_reg_20__15_ ( .D(n1739), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[191]) );
  DFFSR fifo_reg_20__14_ ( .D(n1740), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[190]) );
  DFFSR fifo_reg_20__13_ ( .D(n1741), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[189]) );
  DFFSR fifo_reg_20__12_ ( .D(n1742), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[188]) );
  DFFSR fifo_reg_20__11_ ( .D(n1743), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[187]) );
  DFFSR fifo_reg_20__10_ ( .D(n1744), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[186]) );
  DFFSR fifo_reg_20__9_ ( .D(n1745), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[185]) );
  DFFSR fifo_reg_20__8_ ( .D(n1746), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[184]) );
  DFFSR fifo_reg_20__7_ ( .D(n1747), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[183]) );
  DFFSR fifo_reg_20__6_ ( .D(n1748), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[182]) );
  DFFSR fifo_reg_20__5_ ( .D(n1749), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[181]) );
  DFFSR fifo_reg_20__4_ ( .D(n1750), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[180]) );
  DFFSR fifo_reg_20__3_ ( .D(n1751), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[179]) );
  DFFSR fifo_reg_20__2_ ( .D(n1752), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[178]) );
  DFFSR fifo_reg_20__1_ ( .D(n1753), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[177]) );
  DFFSR fifo_reg_20__0_ ( .D(n1754), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[176]) );
  DFFSR fifo_reg_18__15_ ( .D(n1707), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[223]) );
  DFFSR fifo_reg_18__14_ ( .D(n1708), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[222]) );
  DFFSR fifo_reg_18__13_ ( .D(n1709), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[221]) );
  DFFSR fifo_reg_18__12_ ( .D(n1710), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[220]) );
  DFFSR fifo_reg_18__11_ ( .D(n1711), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[219]) );
  DFFSR fifo_reg_18__10_ ( .D(n1712), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[218]) );
  DFFSR fifo_reg_18__9_ ( .D(n1713), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[217]) );
  DFFSR fifo_reg_18__8_ ( .D(n1714), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[216]) );
  DFFSR fifo_reg_18__7_ ( .D(n1715), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[215]) );
  DFFSR fifo_reg_18__6_ ( .D(n1716), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[214]) );
  DFFSR fifo_reg_18__5_ ( .D(n1717), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[213]) );
  DFFSR fifo_reg_18__4_ ( .D(n1718), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[212]) );
  DFFSR fifo_reg_18__3_ ( .D(n1719), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[211]) );
  DFFSR fifo_reg_18__2_ ( .D(n1720), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[210]) );
  DFFSR fifo_reg_18__1_ ( .D(n1721), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[209]) );
  DFFSR fifo_reg_18__0_ ( .D(n1722), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[208]) );
  DFFSR fifo_reg_13__15_ ( .D(n1627), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[303]) );
  DFFSR fifo_reg_13__14_ ( .D(n1628), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[302]) );
  DFFSR fifo_reg_13__13_ ( .D(n1629), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[301]) );
  DFFSR fifo_reg_13__12_ ( .D(n1630), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[300]) );
  DFFSR fifo_reg_13__11_ ( .D(n1631), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[299]) );
  DFFSR fifo_reg_13__10_ ( .D(n1632), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[298]) );
  DFFSR fifo_reg_13__9_ ( .D(n1633), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[297]) );
  DFFSR fifo_reg_13__8_ ( .D(n1634), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[296]) );
  DFFSR fifo_reg_13__7_ ( .D(n1635), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[295]) );
  DFFSR fifo_reg_13__6_ ( .D(n1636), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[294]) );
  DFFSR fifo_reg_13__5_ ( .D(n1637), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[293]) );
  DFFSR fifo_reg_13__4_ ( .D(n1638), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[292]) );
  DFFSR fifo_reg_13__3_ ( .D(n1639), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[291]) );
  DFFSR fifo_reg_13__2_ ( .D(n1640), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[290]) );
  DFFSR fifo_reg_13__1_ ( .D(n1641), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[289]) );
  DFFSR fifo_reg_13__0_ ( .D(n1642), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[288]) );
  DFFSR fifo_reg_11__15_ ( .D(n1595), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[335]) );
  DFFSR fifo_reg_11__14_ ( .D(n1596), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[334]) );
  DFFSR fifo_reg_11__13_ ( .D(n1597), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[333]) );
  DFFSR fifo_reg_11__12_ ( .D(n1598), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[332]) );
  DFFSR fifo_reg_11__11_ ( .D(n1599), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[331]) );
  DFFSR fifo_reg_11__10_ ( .D(n1600), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[330]) );
  DFFSR fifo_reg_11__9_ ( .D(n1601), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[329]) );
  DFFSR fifo_reg_11__8_ ( .D(n1602), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[328]) );
  DFFSR fifo_reg_11__7_ ( .D(n1603), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[327]) );
  DFFSR fifo_reg_11__6_ ( .D(n1604), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[326]) );
  DFFSR fifo_reg_11__5_ ( .D(n1605), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[325]) );
  DFFSR fifo_reg_11__4_ ( .D(n1606), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[324]) );
  DFFSR fifo_reg_11__3_ ( .D(n1607), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[323]) );
  DFFSR fifo_reg_11__2_ ( .D(n1608), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[322]) );
  DFFSR fifo_reg_11__1_ ( .D(n1609), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[321]) );
  DFFSR fifo_reg_11__0_ ( .D(n1610), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[320]) );
  DFFSR fifo_reg_21__15_ ( .D(n1755), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[175]) );
  DFFSR fifo_reg_21__14_ ( .D(n1756), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[174]) );
  DFFSR fifo_reg_21__13_ ( .D(n1757), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[173]) );
  DFFSR fifo_reg_21__12_ ( .D(n1758), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[172]) );
  DFFSR fifo_reg_21__11_ ( .D(n1759), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[171]) );
  DFFSR fifo_reg_21__10_ ( .D(n1760), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[170]) );
  DFFSR fifo_reg_21__9_ ( .D(n1761), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[169]) );
  DFFSR fifo_reg_21__8_ ( .D(n1762), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[168]) );
  DFFSR fifo_reg_21__7_ ( .D(n1763), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[167]) );
  DFFSR fifo_reg_21__6_ ( .D(n1764), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[166]) );
  DFFSR fifo_reg_21__5_ ( .D(n1765), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[165]) );
  DFFSR fifo_reg_21__4_ ( .D(n1766), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[164]) );
  DFFSR fifo_reg_21__3_ ( .D(n1767), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[163]) );
  DFFSR fifo_reg_21__2_ ( .D(n1768), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[162]) );
  DFFSR fifo_reg_21__1_ ( .D(n1769), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[161]) );
  DFFSR fifo_reg_21__0_ ( .D(n1770), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[160]) );
  DFFSR fifo_reg_19__15_ ( .D(n1723), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[207]) );
  DFFSR fifo_reg_19__14_ ( .D(n1724), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[206]) );
  DFFSR fifo_reg_19__13_ ( .D(n1725), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[205]) );
  DFFSR fifo_reg_19__12_ ( .D(n1726), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[204]) );
  DFFSR fifo_reg_19__11_ ( .D(n1727), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[203]) );
  DFFSR fifo_reg_19__10_ ( .D(n1728), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[202]) );
  DFFSR fifo_reg_19__9_ ( .D(n1729), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[201]) );
  DFFSR fifo_reg_19__8_ ( .D(n1730), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[200]) );
  DFFSR fifo_reg_19__7_ ( .D(n1731), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[199]) );
  DFFSR fifo_reg_19__6_ ( .D(n1732), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[198]) );
  DFFSR fifo_reg_19__5_ ( .D(n1733), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[197]) );
  DFFSR fifo_reg_19__4_ ( .D(n1734), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[196]) );
  DFFSR fifo_reg_19__3_ ( .D(n1735), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[195]) );
  DFFSR fifo_reg_19__2_ ( .D(n1736), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[194]) );
  DFFSR fifo_reg_19__1_ ( .D(n1737), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        fifo[193]) );
  DFFSR fifo_reg_19__0_ ( .D(n1738), .CLK(wclk), .R(n4754), .S(1'b1), .Q(
        fifo[192]) );
  DFFSR wr_ptr_bin_reg_0_ ( .D(n1402), .CLK(wclk), .R(n4755), .S(1'b1), .Q(
        wr_ptr_bin[0]) );
  DFFSR data_out_reg_15_ ( .D(n1347), .CLK(rclk), .R(n4754), .S(1'b1), .Q(
        n5822) );
  DFFSR data_out_reg_4_ ( .D(n1369), .CLK(rclk), .R(n4755), .S(1'b1), .Q(n5833) );
  OR2X1 U3 ( .A(n4645), .B(r301_B_not_0_), .Y(n5819) );
  INVX1 U4 ( .A(n5819), .Y(n1) );
  BUFX2 U5 ( .A(n5833), .Y(data_out[4]) );
  BUFX2 U6 ( .A(n5822), .Y(data_out[15]) );
  BUFX2 U10 ( .A(n5824), .Y(data_out[13]) );
  BUFX2 U13 ( .A(n5827), .Y(data_out[10]) );
  BUFX2 U16 ( .A(n5830), .Y(data_out[7]) );
  BUFX2 U18 ( .A(n5836), .Y(data_out[1]) );
  BUFX2 U20 ( .A(n5823), .Y(data_out[14]) );
  BUFX2 U24 ( .A(n5825), .Y(data_out[12]) );
  BUFX2 U30 ( .A(n5826), .Y(data_out[11]) );
  BUFX2 U36 ( .A(n5828), .Y(data_out[9]) );
  BUFX2 U42 ( .A(n5829), .Y(data_out[8]) );
  BUFX2 U48 ( .A(n5831), .Y(data_out[6]) );
  BUFX2 U52 ( .A(n5832), .Y(data_out[5]) );
  BUFX2 U54 ( .A(n5834), .Y(data_out[3]) );
  BUFX2 U56 ( .A(n5835), .Y(data_out[2]) );
  BUFX2 U58 ( .A(n5837), .Y(data_out[0]) );
  BUFX2 U60 ( .A(rd_ptr_gray_ss[4]), .Y(n39) );
  INVX1 U62 ( .A(n42), .Y(n40) );
  INVX1 U65 ( .A(n40), .Y(empty_bar) );
  BUFX2 U68 ( .A(n5820), .Y(n42) );
  INVX1 U70 ( .A(n45), .Y(n43) );
  INVX1 U72 ( .A(n43), .Y(full_bar) );
  BUFX2 U74 ( .A(n5821), .Y(n45) );
  INVX1 U76 ( .A(n48), .Y(n46) );
  INVX1 U78 ( .A(n46), .Y(n47) );
  BUFX2 U80 ( .A(rd_ptr_gray_s[3]), .Y(n48) );
  INVX1 U82 ( .A(n51), .Y(n49) );
  INVX1 U84 ( .A(n49), .Y(n50) );
  BUFX2 U86 ( .A(rd_ptr_gray[3]), .Y(n51) );
  INVX1 U88 ( .A(n54), .Y(n52) );
  INVX1 U90 ( .A(n52), .Y(n53) );
  BUFX2 U92 ( .A(rd_ptr_gray_s[2]), .Y(n54) );
  INVX1 U94 ( .A(n57), .Y(n55) );
  INVX1 U96 ( .A(n55), .Y(n56) );
  BUFX2 U98 ( .A(rd_ptr_gray[2]), .Y(n57) );
  INVX1 U100 ( .A(n60), .Y(n58) );
  INVX1 U102 ( .A(n58), .Y(n59) );
  BUFX2 U103 ( .A(rd_ptr_gray_s[1]), .Y(n60) );
  INVX1 U105 ( .A(n63), .Y(n61) );
  INVX1 U107 ( .A(n61), .Y(n62) );
  BUFX2 U109 ( .A(rd_ptr_gray[1]), .Y(n63) );
  INVX1 U111 ( .A(n66), .Y(n64) );
  INVX1 U113 ( .A(n64), .Y(n65) );
  BUFX2 U115 ( .A(rd_ptr_gray_s[0]), .Y(n66) );
  INVX1 U117 ( .A(n69), .Y(n67) );
  INVX1 U119 ( .A(n67), .Y(n68) );
  BUFX2 U121 ( .A(rd_ptr_gray[0]), .Y(n69) );
  INVX1 U123 ( .A(n93), .Y(n70) );
  INVX1 U125 ( .A(n70), .Y(n87) );
  BUFX2 U127 ( .A(wr_ptr_gray_s[4]), .Y(n93) );
  INVX1 U129 ( .A(n96), .Y(n94) );
  INVX1 U131 ( .A(n94), .Y(n95) );
  BUFX2 U133 ( .A(wr_ptr_gray[4]), .Y(n96) );
  INVX1 U135 ( .A(n99), .Y(n97) );
  INVX1 U136 ( .A(n97), .Y(n98) );
  BUFX2 U138 ( .A(wr_ptr_gray_s[3]), .Y(n99) );
  INVX1 U140 ( .A(n102), .Y(n100) );
  INVX1 U142 ( .A(n100), .Y(n101) );
  BUFX2 U144 ( .A(wr_ptr_gray[3]), .Y(n102) );
  INVX1 U146 ( .A(n105), .Y(n103) );
  INVX1 U148 ( .A(n103), .Y(n104) );
  BUFX2 U150 ( .A(wr_ptr_gray_s[2]), .Y(n105) );
  INVX1 U152 ( .A(n108), .Y(n106) );
  INVX1 U154 ( .A(n106), .Y(n107) );
  BUFX2 U156 ( .A(wr_ptr_gray[2]), .Y(n108) );
  INVX1 U158 ( .A(n111), .Y(n109) );
  INVX1 U160 ( .A(n109), .Y(n110) );
  BUFX2 U162 ( .A(wr_ptr_gray_s[1]), .Y(n111) );
  INVX1 U164 ( .A(n114), .Y(n112) );
  INVX1 U166 ( .A(n112), .Y(n113) );
  BUFX2 U168 ( .A(wr_ptr_gray[1]), .Y(n114) );
  INVX1 U169 ( .A(n117), .Y(n115) );
  INVX1 U171 ( .A(n115), .Y(n116) );
  BUFX2 U173 ( .A(wr_ptr_gray_s[0]), .Y(n117) );
  INVX1 U175 ( .A(n120), .Y(n118) );
  INVX1 U177 ( .A(n118), .Y(n119) );
  BUFX2 U179 ( .A(wr_ptr_gray[0]), .Y(n120) );
  INVX1 U181 ( .A(n123), .Y(n121) );
  INVX1 U183 ( .A(n121), .Y(n122) );
  BUFX2 U185 ( .A(wr_ptr_gray_s[5]), .Y(n123) );
  INVX1 U187 ( .A(n126), .Y(n124) );
  INVX1 U189 ( .A(n124), .Y(n125) );
  BUFX2 U191 ( .A(wr_ptr_gray[5]), .Y(n126) );
  INVX1 U193 ( .A(n129), .Y(n127) );
  INVX1 U195 ( .A(n127), .Y(n128) );
  BUFX2 U197 ( .A(rd_ptr_gray_s[4]), .Y(n129) );
  INVX1 U199 ( .A(n132), .Y(n130) );
  INVX1 U201 ( .A(n130), .Y(n131) );
  BUFX2 U202 ( .A(rd_ptr_gray[4]), .Y(n132) );
  INVX1 U204 ( .A(n135), .Y(n133) );
  INVX1 U206 ( .A(n133), .Y(n134) );
  BUFX2 U208 ( .A(rd_ptr_gray_s[5]), .Y(n135) );
  INVX1 U210 ( .A(n138), .Y(n136) );
  INVX1 U212 ( .A(n136), .Y(n137) );
  BUFX2 U214 ( .A(rd_ptr_gray[5]), .Y(n138) );
  INVX1 U216 ( .A(n141), .Y(n139) );
  INVX1 U218 ( .A(n139), .Y(n140) );
  BUFX2 U220 ( .A(n798), .Y(n141) );
  INVX1 U222 ( .A(n144), .Y(n142) );
  INVX1 U224 ( .A(n142), .Y(n143) );
  BUFX2 U226 ( .A(n806), .Y(n144) );
  OR2X1 U228 ( .A(n147), .B(n150), .Y(n199) );
  INVX1 U230 ( .A(n199), .Y(n145) );
  INVX1 U232 ( .A(n148), .Y(n146) );
  INVX1 U234 ( .A(n146), .Y(n147) );
  OR2X1 U235 ( .A(n154), .B(n155), .Y(n152) );
  INVX1 U237 ( .A(n152), .Y(n148) );
  INVX1 U239 ( .A(n151), .Y(n149) );
  INVX1 U241 ( .A(n149), .Y(n150) );
  OR2X1 U243 ( .A(n156), .B(n157), .Y(n153) );
  INVX1 U245 ( .A(n153), .Y(n151) );
  INVX1 U247 ( .A(n4649), .Y(n154) );
  INVX1 U249 ( .A(data_out[1]), .Y(n155) );
  INVX1 U251 ( .A(n175), .Y(n156) );
  INVX1 U253 ( .A(n85), .Y(n157) );
  INVX1 U255 ( .A(n5804), .Y(n85) );
  OR2X1 U257 ( .A(n160), .B(n163), .Y(n196) );
  INVX1 U259 ( .A(n196), .Y(n158) );
  INVX1 U261 ( .A(n161), .Y(n159) );
  INVX1 U263 ( .A(n159), .Y(n160) );
  OR2X1 U265 ( .A(n167), .B(n168), .Y(n165) );
  INVX1 U267 ( .A(n165), .Y(n161) );
  INVX1 U268 ( .A(n164), .Y(n162) );
  INVX1 U270 ( .A(n162), .Y(n163) );
  OR2X1 U272 ( .A(n169), .B(n170), .Y(n166) );
  INVX1 U274 ( .A(n166), .Y(n164) );
  INVX1 U276 ( .A(n4649), .Y(n167) );
  INVX1 U278 ( .A(data_out[4]), .Y(n168) );
  INVX1 U280 ( .A(n175), .Y(n169) );
  INVX1 U282 ( .A(n82), .Y(n170) );
  INVX1 U284 ( .A(n5807), .Y(n82) );
  OR2X1 U286 ( .A(n173), .B(n216), .Y(n193) );
  INVX1 U288 ( .A(n193), .Y(n171) );
  INVX1 U290 ( .A(n174), .Y(n172) );
  INVX1 U292 ( .A(n172), .Y(n173) );
  OR2X1 U294 ( .A(n817), .B(n818), .Y(n815) );
  INVX1 U296 ( .A(n815), .Y(n174) );
  INVX1 U298 ( .A(n814), .Y(n182) );
  INVX1 U300 ( .A(n182), .Y(n216) );
  OR2X1 U301 ( .A(n819), .B(n820), .Y(n816) );
  INVX1 U303 ( .A(n816), .Y(n814) );
  INVX1 U305 ( .A(n4649), .Y(n817) );
  INVX1 U307 ( .A(data_out[7]), .Y(n818) );
  INVX1 U309 ( .A(n175), .Y(n819) );
  INVX1 U311 ( .A(n79), .Y(n820) );
  INVX1 U313 ( .A(n5810), .Y(n79) );
  OR2X1 U315 ( .A(n823), .B(n826), .Y(n190) );
  INVX1 U317 ( .A(n190), .Y(n821) );
  INVX1 U319 ( .A(n824), .Y(n822) );
  INVX1 U321 ( .A(n822), .Y(n823) );
  OR2X1 U323 ( .A(n830), .B(n831), .Y(n828) );
  INVX1 U325 ( .A(n828), .Y(n824) );
  INVX1 U327 ( .A(n827), .Y(n825) );
  INVX1 U329 ( .A(n825), .Y(n826) );
  OR2X1 U331 ( .A(n832), .B(n833), .Y(n829) );
  INVX1 U333 ( .A(n829), .Y(n827) );
  INVX1 U334 ( .A(n4649), .Y(n830) );
  INVX1 U338 ( .A(data_out[10]), .Y(n831) );
  INVX1 U340 ( .A(n175), .Y(n832) );
  INVX1 U342 ( .A(n76), .Y(n833) );
  INVX1 U344 ( .A(n5813), .Y(n76) );
  OR2X1 U346 ( .A(n836), .B(n839), .Y(n187) );
  INVX1 U348 ( .A(n187), .Y(n834) );
  INVX1 U350 ( .A(n837), .Y(n835) );
  INVX1 U352 ( .A(n835), .Y(n836) );
  OR2X1 U354 ( .A(n843), .B(n844), .Y(n841) );
  INVX1 U356 ( .A(n841), .Y(n837) );
  INVX1 U358 ( .A(n840), .Y(n838) );
  INVX1 U360 ( .A(n838), .Y(n839) );
  OR2X1 U362 ( .A(n845), .B(n846), .Y(n842) );
  INVX1 U364 ( .A(n842), .Y(n840) );
  INVX1 U366 ( .A(n4649), .Y(n843) );
  INVX1 U368 ( .A(data_out[13]), .Y(n844) );
  INVX1 U369 ( .A(n175), .Y(n845) );
  INVX1 U371 ( .A(n73), .Y(n846) );
  INVX1 U373 ( .A(n5816), .Y(n73) );
  OR2X1 U375 ( .A(n849), .B(n852), .Y(n184) );
  INVX1 U377 ( .A(n184), .Y(n847) );
  INVX1 U379 ( .A(n850), .Y(n848) );
  INVX1 U381 ( .A(n848), .Y(n849) );
  OR2X1 U383 ( .A(n856), .B(n857), .Y(n854) );
  INVX1 U385 ( .A(n854), .Y(n850) );
  INVX1 U387 ( .A(n853), .Y(n851) );
  INVX1 U389 ( .A(n851), .Y(n852) );
  OR2X1 U391 ( .A(n858), .B(n859), .Y(n855) );
  INVX1 U393 ( .A(n855), .Y(n853) );
  INVX1 U395 ( .A(n4649), .Y(n856) );
  INVX1 U397 ( .A(data_out[15]), .Y(n857) );
  INVX1 U399 ( .A(n175), .Y(n858) );
  INVX1 U401 ( .A(n71), .Y(n859) );
  INVX1 U402 ( .A(n5818), .Y(n71) );
  AND2X1 U404 ( .A(n673), .B(n4621), .Y(n691) );
  AND2X1 U406 ( .A(n673), .B(n4618), .Y(n709) );
  AND2X1 U408 ( .A(n673), .B(n4615), .Y(n726) );
  AND2X1 U410 ( .A(n673), .B(n4612), .Y(n744) );
  AND2X1 U412 ( .A(n673), .B(n360), .Y(n761) );
  AND2X1 U414 ( .A(n673), .B(n251), .Y(n656) );
  AND2X1 U416 ( .A(n673), .B(n270), .Y(n674) );
  AND2X1 U418 ( .A(n535), .B(n251), .Y(n518) );
  AND2X1 U420 ( .A(n535), .B(n270), .Y(n536) );
  AND2X1 U422 ( .A(n535), .B(n4621), .Y(n553) );
  AND2X1 U424 ( .A(n535), .B(n4618), .Y(n570) );
  AND2X1 U426 ( .A(n535), .B(n4615), .Y(n587) );
  AND2X1 U428 ( .A(n535), .B(n4612), .Y(n604) );
  AND2X1 U430 ( .A(n535), .B(n360), .Y(n621) );
  AND2X1 U432 ( .A(n397), .B(n251), .Y(n380) );
  AND2X1 U434 ( .A(n397), .B(n270), .Y(n398) );
  AND2X1 U435 ( .A(n397), .B(n4621), .Y(n415) );
  AND2X1 U437 ( .A(n397), .B(n4618), .Y(n432) );
  AND2X1 U439 ( .A(n397), .B(n4615), .Y(n449) );
  AND2X1 U441 ( .A(n397), .B(n4612), .Y(n466) );
  AND2X1 U443 ( .A(n397), .B(n360), .Y(n483) );
  AND2X1 U445 ( .A(n270), .B(n252), .Y(n253) );
  AND2X1 U447 ( .A(n4621), .B(n252), .Y(n271) );
  AND2X1 U449 ( .A(n4618), .B(n252), .Y(n289) );
  AND2X1 U451 ( .A(n4615), .B(n252), .Y(n307) );
  AND2X1 U453 ( .A(n4612), .B(n252), .Y(n325) );
  AND2X1 U455 ( .A(n360), .B(n252), .Y(n343) );
  INVX1 U457 ( .A(n862), .Y(n860) );
  INVX1 U459 ( .A(n860), .Y(n861) );
  AND2X1 U461 ( .A(n4606), .B(n4603), .Y(n23) );
  INVX1 U463 ( .A(n23), .Y(n862) );
  INVX1 U465 ( .A(n865), .Y(n863) );
  INVX1 U467 ( .A(n863), .Y(n864) );
  AND2X1 U468 ( .A(n4311), .B(n4658), .Y(n794) );
  INVX1 U470 ( .A(n794), .Y(n865) );
  INVX1 U472 ( .A(n868), .Y(n866) );
  INVX1 U474 ( .A(n866), .Y(n867) );
  AND2X1 U476 ( .A(n4314), .B(n4658), .Y(n793) );
  INVX1 U478 ( .A(n793), .Y(n868) );
  INVX1 U480 ( .A(n871), .Y(n869) );
  INVX1 U482 ( .A(n869), .Y(n870) );
  AND2X1 U484 ( .A(n4317), .B(n4658), .Y(n792) );
  INVX1 U486 ( .A(n792), .Y(n871) );
  INVX1 U488 ( .A(n874), .Y(n872) );
  INVX1 U490 ( .A(n872), .Y(n873) );
  AND2X1 U492 ( .A(n4320), .B(n4658), .Y(n791) );
  INVX1 U494 ( .A(n791), .Y(n874) );
  INVX1 U496 ( .A(n877), .Y(n875) );
  INVX1 U498 ( .A(n875), .Y(n876) );
  AND2X1 U500 ( .A(n4323), .B(n4658), .Y(n790) );
  INVX1 U501 ( .A(n790), .Y(n877) );
  INVX1 U503 ( .A(n880), .Y(n878) );
  INVX1 U505 ( .A(n878), .Y(n879) );
  AND2X1 U507 ( .A(n4326), .B(n4658), .Y(n789) );
  INVX1 U509 ( .A(n789), .Y(n880) );
  INVX1 U511 ( .A(n883), .Y(n881) );
  INVX1 U513 ( .A(n881), .Y(n882) );
  AND2X1 U515 ( .A(n4329), .B(n4658), .Y(n788) );
  INVX1 U517 ( .A(n788), .Y(n883) );
  INVX1 U519 ( .A(n886), .Y(n884) );
  INVX1 U521 ( .A(n884), .Y(n885) );
  AND2X1 U523 ( .A(n4332), .B(n4658), .Y(n787) );
  INVX1 U525 ( .A(n787), .Y(n886) );
  INVX1 U527 ( .A(n889), .Y(n887) );
  INVX1 U529 ( .A(n887), .Y(n888) );
  AND2X1 U531 ( .A(n4335), .B(n4658), .Y(n786) );
  INVX1 U533 ( .A(n786), .Y(n889) );
  INVX1 U534 ( .A(n892), .Y(n890) );
  INVX1 U536 ( .A(n890), .Y(n891) );
  AND2X1 U538 ( .A(n4338), .B(n4658), .Y(n785) );
  INVX1 U540 ( .A(n785), .Y(n892) );
  INVX1 U542 ( .A(n895), .Y(n893) );
  INVX1 U544 ( .A(n893), .Y(n894) );
  AND2X1 U546 ( .A(n4341), .B(n4658), .Y(n784) );
  INVX1 U548 ( .A(n784), .Y(n895) );
  INVX1 U550 ( .A(n898), .Y(n896) );
  INVX1 U552 ( .A(n896), .Y(n897) );
  AND2X1 U554 ( .A(n4344), .B(n4658), .Y(n783) );
  INVX1 U556 ( .A(n783), .Y(n898) );
  INVX1 U558 ( .A(n901), .Y(n899) );
  INVX1 U560 ( .A(n899), .Y(n900) );
  AND2X1 U562 ( .A(n4347), .B(n4658), .Y(n782) );
  INVX1 U564 ( .A(n782), .Y(n901) );
  INVX1 U566 ( .A(n904), .Y(n902) );
  INVX1 U567 ( .A(n902), .Y(n903) );
  AND2X1 U569 ( .A(n4350), .B(n4658), .Y(n781) );
  INVX1 U571 ( .A(n781), .Y(n904) );
  INVX1 U573 ( .A(n907), .Y(n905) );
  INVX1 U575 ( .A(n905), .Y(n906) );
  AND2X1 U577 ( .A(n4353), .B(n4658), .Y(n780) );
  INVX1 U579 ( .A(n780), .Y(n907) );
  INVX1 U581 ( .A(n910), .Y(n908) );
  INVX1 U583 ( .A(n908), .Y(n909) );
  AND2X1 U585 ( .A(n4356), .B(n4658), .Y(n779) );
  INVX1 U587 ( .A(n779), .Y(n910) );
  INVX1 U589 ( .A(n913), .Y(n911) );
  INVX1 U591 ( .A(n911), .Y(n912) );
  AND2X1 U593 ( .A(n3543), .B(n4661), .Y(n777) );
  INVX1 U595 ( .A(n777), .Y(n913) );
  INVX1 U597 ( .A(n916), .Y(n914) );
  INVX1 U599 ( .A(n914), .Y(n915) );
  AND2X1 U600 ( .A(n3546), .B(n4661), .Y(n776) );
  INVX1 U605 ( .A(n776), .Y(n916) );
  INVX1 U607 ( .A(n919), .Y(n917) );
  INVX1 U609 ( .A(n917), .Y(n918) );
  AND2X1 U611 ( .A(n3549), .B(n4661), .Y(n775) );
  INVX1 U613 ( .A(n775), .Y(n919) );
  INVX1 U615 ( .A(n922), .Y(n920) );
  INVX1 U617 ( .A(n920), .Y(n921) );
  AND2X1 U619 ( .A(n3552), .B(n4661), .Y(n774) );
  INVX1 U621 ( .A(n774), .Y(n922) );
  INVX1 U623 ( .A(n925), .Y(n923) );
  INVX1 U625 ( .A(n923), .Y(n924) );
  AND2X1 U627 ( .A(n3555), .B(n4661), .Y(n773) );
  INVX1 U629 ( .A(n773), .Y(n925) );
  INVX1 U631 ( .A(n928), .Y(n926) );
  INVX1 U633 ( .A(n926), .Y(n927) );
  AND2X1 U635 ( .A(n3558), .B(n4661), .Y(n772) );
  INVX1 U636 ( .A(n772), .Y(n928) );
  INVX1 U638 ( .A(n931), .Y(n929) );
  INVX1 U640 ( .A(n929), .Y(n930) );
  AND2X1 U642 ( .A(n3561), .B(n4661), .Y(n771) );
  INVX1 U644 ( .A(n771), .Y(n931) );
  INVX1 U646 ( .A(n934), .Y(n932) );
  INVX1 U648 ( .A(n932), .Y(n933) );
  AND2X1 U650 ( .A(n3564), .B(n4661), .Y(n770) );
  INVX1 U652 ( .A(n770), .Y(n934) );
  INVX1 U654 ( .A(n937), .Y(n935) );
  INVX1 U656 ( .A(n935), .Y(n936) );
  AND2X1 U658 ( .A(n3567), .B(n4661), .Y(n769) );
  INVX1 U660 ( .A(n769), .Y(n937) );
  INVX1 U662 ( .A(n940), .Y(n938) );
  INVX1 U664 ( .A(n938), .Y(n939) );
  AND2X1 U666 ( .A(n3570), .B(n4661), .Y(n768) );
  INVX1 U668 ( .A(n768), .Y(n940) );
  INVX1 U669 ( .A(n943), .Y(n941) );
  INVX1 U671 ( .A(n941), .Y(n942) );
  AND2X1 U673 ( .A(n3573), .B(n4661), .Y(n767) );
  INVX1 U675 ( .A(n767), .Y(n943) );
  INVX1 U677 ( .A(n946), .Y(n944) );
  INVX1 U679 ( .A(n944), .Y(n945) );
  AND2X1 U681 ( .A(n3576), .B(n4661), .Y(n766) );
  INVX1 U683 ( .A(n766), .Y(n946) );
  INVX1 U685 ( .A(n949), .Y(n947) );
  INVX1 U687 ( .A(n947), .Y(n948) );
  AND2X1 U689 ( .A(n3579), .B(n4661), .Y(n765) );
  INVX1 U691 ( .A(n765), .Y(n949) );
  INVX1 U693 ( .A(n952), .Y(n950) );
  INVX1 U695 ( .A(n950), .Y(n951) );
  AND2X1 U697 ( .A(n3582), .B(n4661), .Y(n764) );
  INVX1 U699 ( .A(n764), .Y(n952) );
  INVX1 U701 ( .A(n955), .Y(n953) );
  INVX1 U702 ( .A(n953), .Y(n954) );
  AND2X1 U704 ( .A(n3585), .B(n4661), .Y(n763) );
  INVX1 U706 ( .A(n763), .Y(n955) );
  INVX1 U708 ( .A(n958), .Y(n956) );
  INVX1 U710 ( .A(n956), .Y(n957) );
  AND2X1 U712 ( .A(n3588), .B(n4661), .Y(n762) );
  INVX1 U714 ( .A(n762), .Y(n958) );
  INVX1 U716 ( .A(n961), .Y(n959) );
  INVX1 U718 ( .A(n959), .Y(n960) );
  AND2X1 U720 ( .A(n4263), .B(n4664), .Y(n760) );
  INVX1 U722 ( .A(n760), .Y(n961) );
  INVX1 U724 ( .A(n964), .Y(n962) );
  INVX1 U726 ( .A(n962), .Y(n963) );
  AND2X1 U728 ( .A(n4266), .B(n4664), .Y(n759) );
  INVX1 U730 ( .A(n759), .Y(n964) );
  INVX1 U732 ( .A(n967), .Y(n965) );
  INVX1 U734 ( .A(n965), .Y(n966) );
  AND2X1 U735 ( .A(n4269), .B(n4664), .Y(n758) );
  INVX1 U737 ( .A(n758), .Y(n967) );
  INVX1 U739 ( .A(n970), .Y(n968) );
  INVX1 U741 ( .A(n968), .Y(n969) );
  AND2X1 U743 ( .A(n4272), .B(n4664), .Y(n757) );
  INVX1 U745 ( .A(n757), .Y(n970) );
  INVX1 U747 ( .A(n973), .Y(n971) );
  INVX1 U749 ( .A(n971), .Y(n972) );
  AND2X1 U751 ( .A(n4275), .B(n4664), .Y(n756) );
  INVX1 U753 ( .A(n756), .Y(n973) );
  INVX1 U755 ( .A(n976), .Y(n974) );
  INVX1 U757 ( .A(n974), .Y(n975) );
  AND2X1 U759 ( .A(n4278), .B(n4664), .Y(n755) );
  INVX1 U761 ( .A(n755), .Y(n976) );
  INVX1 U763 ( .A(n979), .Y(n977) );
  INVX1 U765 ( .A(n977), .Y(n978) );
  AND2X1 U767 ( .A(n4281), .B(n4664), .Y(n754) );
  INVX1 U768 ( .A(n754), .Y(n979) );
  INVX1 U770 ( .A(n982), .Y(n980) );
  INVX1 U772 ( .A(n980), .Y(n981) );
  AND2X1 U774 ( .A(n4284), .B(n4664), .Y(n753) );
  INVX1 U776 ( .A(n753), .Y(n982) );
  INVX1 U778 ( .A(n985), .Y(n983) );
  INVX1 U780 ( .A(n983), .Y(n984) );
  AND2X1 U782 ( .A(n4287), .B(n4664), .Y(n752) );
  INVX1 U784 ( .A(n752), .Y(n985) );
  INVX1 U786 ( .A(n988), .Y(n986) );
  INVX1 U788 ( .A(n986), .Y(n987) );
  AND2X1 U790 ( .A(n4290), .B(n4664), .Y(n751) );
  INVX1 U792 ( .A(n751), .Y(n988) );
  INVX1 U794 ( .A(n991), .Y(n989) );
  INVX1 U796 ( .A(n989), .Y(n990) );
  AND2X1 U798 ( .A(n4293), .B(n4664), .Y(n750) );
  INVX1 U800 ( .A(n750), .Y(n991) );
  INVX1 U801 ( .A(n994), .Y(n992) );
  INVX1 U803 ( .A(n992), .Y(n993) );
  AND2X1 U805 ( .A(n4296), .B(n4664), .Y(n749) );
  INVX1 U807 ( .A(n749), .Y(n994) );
  INVX1 U809 ( .A(n997), .Y(n995) );
  INVX1 U811 ( .A(n995), .Y(n996) );
  AND2X1 U813 ( .A(n4299), .B(n4664), .Y(n748) );
  INVX1 U815 ( .A(n748), .Y(n997) );
  INVX1 U817 ( .A(n1000), .Y(n998) );
  INVX1 U819 ( .A(n998), .Y(n999) );
  AND2X1 U821 ( .A(n4302), .B(n4664), .Y(n747) );
  INVX1 U823 ( .A(n747), .Y(n1000) );
  INVX1 U825 ( .A(n1003), .Y(n1001) );
  INVX1 U827 ( .A(n1001), .Y(n1002) );
  AND2X1 U829 ( .A(n4305), .B(n4664), .Y(n746) );
  INVX1 U831 ( .A(n746), .Y(n1003) );
  INVX1 U833 ( .A(n1006), .Y(n1004) );
  INVX1 U834 ( .A(n1004), .Y(n1005) );
  AND2X1 U836 ( .A(n4308), .B(n4664), .Y(n745) );
  INVX1 U838 ( .A(n745), .Y(n1006) );
  INVX1 U840 ( .A(n1009), .Y(n1007) );
  INVX1 U842 ( .A(n1007), .Y(n1008) );
  AND2X1 U844 ( .A(n3495), .B(n4667), .Y(n742) );
  INVX1 U846 ( .A(n742), .Y(n1009) );
  INVX1 U848 ( .A(n1012), .Y(n1010) );
  INVX1 U850 ( .A(n1010), .Y(n1011) );
  AND2X1 U852 ( .A(n3498), .B(n4667), .Y(n741) );
  INVX1 U854 ( .A(n741), .Y(n1012) );
  INVX1 U856 ( .A(n1015), .Y(n1013) );
  INVX1 U858 ( .A(n1013), .Y(n1014) );
  AND2X1 U860 ( .A(n3501), .B(n4667), .Y(n740) );
  INVX1 U862 ( .A(n740), .Y(n1015) );
  INVX1 U864 ( .A(n1018), .Y(n1016) );
  INVX1 U866 ( .A(n1016), .Y(n1017) );
  AND2X1 U867 ( .A(n3504), .B(n4667), .Y(n739) );
  INVX1 U872 ( .A(n739), .Y(n1018) );
  INVX1 U874 ( .A(n1021), .Y(n1019) );
  INVX1 U876 ( .A(n1019), .Y(n1020) );
  AND2X1 U878 ( .A(n3507), .B(n4667), .Y(n738) );
  INVX1 U880 ( .A(n738), .Y(n1021) );
  INVX1 U882 ( .A(n1024), .Y(n1022) );
  INVX1 U884 ( .A(n1022), .Y(n1023) );
  AND2X1 U886 ( .A(n3510), .B(n4667), .Y(n737) );
  INVX1 U888 ( .A(n737), .Y(n1024) );
  INVX1 U890 ( .A(n1027), .Y(n1025) );
  INVX1 U892 ( .A(n1025), .Y(n1026) );
  AND2X1 U894 ( .A(n3513), .B(n4667), .Y(n736) );
  INVX1 U896 ( .A(n736), .Y(n1027) );
  INVX1 U898 ( .A(n1030), .Y(n1028) );
  INVX1 U900 ( .A(n1028), .Y(n1029) );
  AND2X1 U902 ( .A(n3516), .B(n4667), .Y(n735) );
  INVX1 U903 ( .A(n735), .Y(n1030) );
  INVX1 U906 ( .A(n1033), .Y(n1031) );
  INVX1 U908 ( .A(n1031), .Y(n1032) );
  AND2X1 U910 ( .A(n3519), .B(n4667), .Y(n734) );
  INVX1 U912 ( .A(n734), .Y(n1033) );
  INVX1 U914 ( .A(n1036), .Y(n1034) );
  INVX1 U916 ( .A(n1034), .Y(n1035) );
  AND2X1 U918 ( .A(n3522), .B(n4667), .Y(n733) );
  INVX1 U920 ( .A(n733), .Y(n1036) );
  INVX1 U922 ( .A(n1039), .Y(n1037) );
  INVX1 U924 ( .A(n1037), .Y(n1038) );
  AND2X1 U926 ( .A(n3525), .B(n4667), .Y(n732) );
  INVX1 U928 ( .A(n732), .Y(n1039) );
  INVX1 U930 ( .A(n1042), .Y(n1040) );
  INVX1 U932 ( .A(n1040), .Y(n1041) );
  AND2X1 U934 ( .A(n3528), .B(n4667), .Y(n731) );
  INVX1 U936 ( .A(n731), .Y(n1042) );
  INVX1 U937 ( .A(n1045), .Y(n1043) );
  INVX1 U940 ( .A(n1043), .Y(n1044) );
  AND2X1 U942 ( .A(n3531), .B(n4667), .Y(n730) );
  INVX1 U944 ( .A(n730), .Y(n1045) );
  INVX1 U946 ( .A(n1048), .Y(n1046) );
  INVX1 U948 ( .A(n1046), .Y(n1047) );
  AND2X1 U950 ( .A(n3534), .B(n4667), .Y(n729) );
  INVX1 U952 ( .A(n729), .Y(n1048) );
  INVX1 U954 ( .A(n1051), .Y(n1049) );
  INVX1 U956 ( .A(n1049), .Y(n1050) );
  AND2X1 U958 ( .A(n3537), .B(n4667), .Y(n728) );
  INVX1 U960 ( .A(n728), .Y(n1051) );
  INVX1 U962 ( .A(n1054), .Y(n1052) );
  INVX1 U964 ( .A(n1052), .Y(n1053) );
  AND2X1 U966 ( .A(n3540), .B(n4667), .Y(n727) );
  INVX1 U968 ( .A(n727), .Y(n1054) );
  INVX1 U970 ( .A(n1057), .Y(n1055) );
  INVX1 U971 ( .A(n1055), .Y(n1056) );
  AND2X1 U972 ( .A(n4215), .B(n4670), .Y(n725) );
  INVX1 U974 ( .A(n725), .Y(n1057) );
  INVX1 U976 ( .A(n1060), .Y(n1058) );
  INVX1 U978 ( .A(n1058), .Y(n1059) );
  AND2X1 U980 ( .A(n4218), .B(n4670), .Y(n724) );
  INVX1 U982 ( .A(n724), .Y(n1060) );
  INVX1 U984 ( .A(n1063), .Y(n1061) );
  INVX1 U986 ( .A(n1061), .Y(n1062) );
  AND2X1 U988 ( .A(n4221), .B(n4670), .Y(n723) );
  INVX1 U990 ( .A(n723), .Y(n1063) );
  INVX1 U992 ( .A(n1066), .Y(n1064) );
  INVX1 U994 ( .A(n1064), .Y(n1065) );
  AND2X1 U996 ( .A(n4224), .B(n4670), .Y(n722) );
  INVX1 U998 ( .A(n722), .Y(n1066) );
  INVX1 U1000 ( .A(n1069), .Y(n1067) );
  INVX1 U1002 ( .A(n1067), .Y(n1068) );
  AND2X1 U1004 ( .A(n4227), .B(n4670), .Y(n721) );
  INVX1 U1005 ( .A(n721), .Y(n1069) );
  INVX1 U1006 ( .A(n1072), .Y(n1070) );
  INVX1 U1008 ( .A(n1070), .Y(n1071) );
  AND2X1 U1010 ( .A(n4230), .B(n4670), .Y(n720) );
  INVX1 U1012 ( .A(n720), .Y(n1072) );
  INVX1 U1014 ( .A(n1075), .Y(n1073) );
  INVX1 U1016 ( .A(n1073), .Y(n1074) );
  AND2X1 U1018 ( .A(n4233), .B(n4670), .Y(n719) );
  INVX1 U1020 ( .A(n719), .Y(n1075) );
  INVX1 U1022 ( .A(n1078), .Y(n1076) );
  INVX1 U1024 ( .A(n1076), .Y(n1077) );
  AND2X1 U1026 ( .A(n4236), .B(n4670), .Y(n718) );
  INVX1 U1028 ( .A(n718), .Y(n1078) );
  INVX1 U1030 ( .A(n1081), .Y(n1079) );
  INVX1 U1032 ( .A(n1079), .Y(n1080) );
  AND2X1 U1034 ( .A(n4239), .B(n4670), .Y(n717) );
  INVX1 U1036 ( .A(n717), .Y(n1081) );
  INVX1 U1038 ( .A(n1084), .Y(n1082) );
  INVX1 U1039 ( .A(n1082), .Y(n1083) );
  AND2X1 U1040 ( .A(n4242), .B(n4670), .Y(n716) );
  INVX1 U1042 ( .A(n716), .Y(n1084) );
  INVX1 U1044 ( .A(n1087), .Y(n1085) );
  INVX1 U1046 ( .A(n1085), .Y(n1086) );
  AND2X1 U1048 ( .A(n4245), .B(n4670), .Y(n715) );
  INVX1 U1050 ( .A(n715), .Y(n1087) );
  INVX1 U1052 ( .A(n1090), .Y(n1088) );
  INVX1 U1054 ( .A(n1088), .Y(n1089) );
  AND2X1 U1056 ( .A(n4248), .B(n4670), .Y(n714) );
  INVX1 U1058 ( .A(n714), .Y(n1090) );
  INVX1 U1060 ( .A(n1093), .Y(n1091) );
  INVX1 U1062 ( .A(n1091), .Y(n1092) );
  AND2X1 U1064 ( .A(n4251), .B(n4670), .Y(n713) );
  INVX1 U1066 ( .A(n713), .Y(n1093) );
  INVX1 U1068 ( .A(n1096), .Y(n1094) );
  INVX1 U1070 ( .A(n1094), .Y(n1095) );
  AND2X1 U1072 ( .A(n4254), .B(n4670), .Y(n712) );
  INVX1 U1073 ( .A(n712), .Y(n1096) );
  INVX1 U1074 ( .A(n1099), .Y(n1097) );
  INVX1 U1076 ( .A(n1097), .Y(n1098) );
  AND2X1 U1078 ( .A(n4257), .B(n4670), .Y(n711) );
  INVX1 U1080 ( .A(n711), .Y(n1099) );
  INVX1 U1082 ( .A(n1102), .Y(n1100) );
  INVX1 U1084 ( .A(n1100), .Y(n1101) );
  AND2X1 U1086 ( .A(n4260), .B(n4670), .Y(n710) );
  INVX1 U1088 ( .A(n710), .Y(n1102) );
  INVX1 U1090 ( .A(n1105), .Y(n1103) );
  INVX1 U1092 ( .A(n1103), .Y(n1104) );
  AND2X1 U1094 ( .A(n3447), .B(n4673), .Y(n707) );
  INVX1 U1096 ( .A(n707), .Y(n1105) );
  INVX1 U1098 ( .A(n1108), .Y(n1106) );
  INVX1 U1100 ( .A(n1106), .Y(n1107) );
  AND2X1 U1102 ( .A(n3450), .B(n4673), .Y(n706) );
  INVX1 U1104 ( .A(n706), .Y(n1108) );
  INVX1 U1106 ( .A(n1111), .Y(n1109) );
  INVX1 U1107 ( .A(n1109), .Y(n1110) );
  AND2X1 U1110 ( .A(n3453), .B(n4673), .Y(n705) );
  INVX1 U1113 ( .A(n705), .Y(n1111) );
  INVX1 U1116 ( .A(n1114), .Y(n1112) );
  INVX1 U1119 ( .A(n1112), .Y(n1113) );
  AND2X1 U1122 ( .A(n3456), .B(n4673), .Y(n704) );
  INVX1 U1125 ( .A(n704), .Y(n1114) );
  INVX1 U1128 ( .A(n1117), .Y(n1115) );
  INVX1 U1131 ( .A(n1115), .Y(n1116) );
  AND2X1 U1134 ( .A(n3459), .B(n4673), .Y(n703) );
  INVX1 U1137 ( .A(n703), .Y(n1117) );
  INVX1 U1140 ( .A(n1120), .Y(n1118) );
  INVX1 U1143 ( .A(n1118), .Y(n1119) );
  AND2X1 U1146 ( .A(n3462), .B(n4673), .Y(n702) );
  INVX1 U1149 ( .A(n702), .Y(n1120) );
  INVX1 U1152 ( .A(n1123), .Y(n1121) );
  INVX1 U1155 ( .A(n1121), .Y(n1122) );
  AND2X1 U1156 ( .A(n3465), .B(n4673), .Y(n701) );
  INVX1 U1161 ( .A(n701), .Y(n1123) );
  INVX1 U1164 ( .A(n1126), .Y(n1124) );
  INVX1 U1165 ( .A(n1124), .Y(n1125) );
  AND2X1 U1167 ( .A(n3468), .B(n4673), .Y(n700) );
  INVX1 U1179 ( .A(n700), .Y(n1126) );
  INVX1 U1181 ( .A(n1129), .Y(n1127) );
  INVX1 U1189 ( .A(n1127), .Y(n1128) );
  AND2X1 U1192 ( .A(n3471), .B(n4673), .Y(n699) );
  INVX1 U1201 ( .A(n699), .Y(n1129) );
  INVX1 U1202 ( .A(n1132), .Y(n1130) );
  INVX1 U1203 ( .A(n1130), .Y(n1131) );
  AND2X1 U1204 ( .A(n3474), .B(n4673), .Y(n698) );
  INVX1 U1205 ( .A(n698), .Y(n1132) );
  INVX1 U1206 ( .A(n1135), .Y(n1133) );
  INVX1 U1207 ( .A(n1133), .Y(n1134) );
  AND2X1 U1208 ( .A(n3477), .B(n4673), .Y(n697) );
  INVX1 U1209 ( .A(n697), .Y(n1135) );
  INVX1 U1210 ( .A(n1138), .Y(n1136) );
  INVX1 U1211 ( .A(n1136), .Y(n1137) );
  AND2X1 U1212 ( .A(n3480), .B(n4673), .Y(n696) );
  INVX1 U1213 ( .A(n696), .Y(n1138) );
  INVX1 U1214 ( .A(n1141), .Y(n1139) );
  INVX1 U1215 ( .A(n1139), .Y(n1140) );
  AND2X1 U1216 ( .A(n3483), .B(n4673), .Y(n695) );
  INVX1 U1217 ( .A(n695), .Y(n1141) );
  INVX1 U1218 ( .A(n1144), .Y(n1142) );
  INVX1 U1219 ( .A(n1142), .Y(n1143) );
  AND2X1 U1220 ( .A(n3486), .B(n4673), .Y(n694) );
  INVX1 U1221 ( .A(n694), .Y(n1144) );
  INVX1 U1222 ( .A(n1147), .Y(n1145) );
  INVX1 U1223 ( .A(n1145), .Y(n1146) );
  AND2X1 U1224 ( .A(n3489), .B(n4673), .Y(n693) );
  INVX1 U1225 ( .A(n693), .Y(n1147) );
  INVX1 U1226 ( .A(n1150), .Y(n1148) );
  INVX1 U1227 ( .A(n1148), .Y(n1149) );
  AND2X1 U1228 ( .A(n3492), .B(n4673), .Y(n692) );
  INVX1 U1229 ( .A(n692), .Y(n1150) );
  INVX1 U1230 ( .A(n1153), .Y(n1151) );
  INVX1 U1231 ( .A(n1151), .Y(n1152) );
  AND2X1 U1232 ( .A(n4359), .B(n4676), .Y(n690) );
  INVX1 U1233 ( .A(n690), .Y(n1153) );
  INVX1 U1234 ( .A(n1156), .Y(n1154) );
  INVX1 U1235 ( .A(n1154), .Y(n1155) );
  AND2X1 U1236 ( .A(n4362), .B(n4676), .Y(n689) );
  INVX1 U1237 ( .A(n689), .Y(n1156) );
  INVX1 U1238 ( .A(n1159), .Y(n1157) );
  INVX1 U1239 ( .A(n1157), .Y(n1158) );
  AND2X1 U1240 ( .A(n4365), .B(n4676), .Y(n688) );
  INVX1 U1241 ( .A(n688), .Y(n1159) );
  INVX1 U1242 ( .A(n1162), .Y(n1160) );
  INVX1 U1243 ( .A(n1160), .Y(n1161) );
  AND2X1 U1244 ( .A(n4368), .B(n4676), .Y(n687) );
  INVX1 U1245 ( .A(n687), .Y(n1162) );
  INVX1 U1246 ( .A(n1165), .Y(n1163) );
  INVX1 U1247 ( .A(n1163), .Y(n1164) );
  AND2X1 U1248 ( .A(n4371), .B(n4676), .Y(n686) );
  INVX1 U1249 ( .A(n686), .Y(n1165) );
  INVX1 U1250 ( .A(n1168), .Y(n1166) );
  INVX1 U1251 ( .A(n1166), .Y(n1167) );
  AND2X1 U1252 ( .A(n4374), .B(n4676), .Y(n685) );
  INVX1 U1253 ( .A(n685), .Y(n1168) );
  INVX1 U1254 ( .A(n1171), .Y(n1169) );
  INVX1 U1255 ( .A(n1169), .Y(n1170) );
  AND2X1 U1256 ( .A(n4377), .B(n4676), .Y(n684) );
  INVX1 U1257 ( .A(n684), .Y(n1171) );
  INVX1 U1258 ( .A(n1174), .Y(n1172) );
  INVX1 U1259 ( .A(n1172), .Y(n1173) );
  AND2X1 U1260 ( .A(n4380), .B(n4676), .Y(n683) );
  INVX1 U1261 ( .A(n683), .Y(n1174) );
  INVX1 U1262 ( .A(n1177), .Y(n1175) );
  INVX1 U1263 ( .A(n1175), .Y(n1176) );
  AND2X1 U1264 ( .A(n4383), .B(n4676), .Y(n682) );
  INVX1 U1265 ( .A(n682), .Y(n1177) );
  INVX1 U1266 ( .A(n1180), .Y(n1178) );
  INVX1 U1267 ( .A(n1178), .Y(n1179) );
  AND2X1 U1268 ( .A(n4386), .B(n4676), .Y(n681) );
  INVX1 U1269 ( .A(n681), .Y(n1180) );
  INVX1 U1270 ( .A(n1183), .Y(n1181) );
  INVX1 U1271 ( .A(n1181), .Y(n1182) );
  AND2X1 U1272 ( .A(n4389), .B(n4676), .Y(n680) );
  INVX1 U1273 ( .A(n680), .Y(n1183) );
  INVX1 U1274 ( .A(n1186), .Y(n1184) );
  INVX1 U1275 ( .A(n1184), .Y(n1185) );
  AND2X1 U1276 ( .A(n4392), .B(n4676), .Y(n679) );
  INVX1 U1277 ( .A(n679), .Y(n1186) );
  INVX1 U1278 ( .A(n1189), .Y(n1187) );
  INVX1 U1279 ( .A(n1187), .Y(n1188) );
  AND2X1 U1280 ( .A(n4395), .B(n4676), .Y(n678) );
  INVX1 U1281 ( .A(n678), .Y(n1189) );
  INVX1 U1282 ( .A(n1192), .Y(n1190) );
  INVX1 U1283 ( .A(n1190), .Y(n1191) );
  AND2X1 U1284 ( .A(n4398), .B(n4676), .Y(n677) );
  INVX1 U1285 ( .A(n677), .Y(n1192) );
  INVX1 U1286 ( .A(n1195), .Y(n1193) );
  INVX1 U1287 ( .A(n1193), .Y(n1194) );
  AND2X1 U1288 ( .A(n4401), .B(n4676), .Y(n676) );
  INVX1 U1289 ( .A(n676), .Y(n1195) );
  INVX1 U1290 ( .A(n1198), .Y(n1196) );
  INVX1 U1291 ( .A(n1196), .Y(n1197) );
  AND2X1 U1292 ( .A(n4404), .B(n4676), .Y(n675) );
  INVX1 U1293 ( .A(n675), .Y(n1198) );
  INVX1 U1294 ( .A(n1201), .Y(n1199) );
  INVX1 U1295 ( .A(n1199), .Y(n1200) );
  AND2X1 U1296 ( .A(n3591), .B(n4679), .Y(n672) );
  INVX1 U1297 ( .A(n672), .Y(n1201) );
  INVX1 U1298 ( .A(n1204), .Y(n1202) );
  INVX1 U1299 ( .A(n1202), .Y(n1203) );
  AND2X1 U1300 ( .A(n3594), .B(n4679), .Y(n671) );
  INVX1 U1301 ( .A(n671), .Y(n1204) );
  INVX1 U1302 ( .A(n1207), .Y(n1205) );
  INVX1 U1303 ( .A(n1205), .Y(n1206) );
  AND2X1 U1304 ( .A(n3597), .B(n4679), .Y(n670) );
  INVX1 U1305 ( .A(n670), .Y(n1207) );
  INVX1 U1306 ( .A(n1210), .Y(n1208) );
  INVX1 U1307 ( .A(n1208), .Y(n1209) );
  AND2X1 U1308 ( .A(n3600), .B(n4679), .Y(n669) );
  INVX1 U1309 ( .A(n669), .Y(n1210) );
  INVX1 U1310 ( .A(n1213), .Y(n1211) );
  INVX1 U1311 ( .A(n1211), .Y(n1212) );
  AND2X1 U1312 ( .A(n3603), .B(n4679), .Y(n668) );
  INVX1 U1313 ( .A(n668), .Y(n1213) );
  INVX1 U1314 ( .A(n1216), .Y(n1214) );
  INVX1 U1315 ( .A(n1214), .Y(n1215) );
  AND2X1 U1316 ( .A(n3606), .B(n4679), .Y(n667) );
  INVX1 U1317 ( .A(n667), .Y(n1216) );
  INVX1 U1318 ( .A(n1219), .Y(n1217) );
  INVX1 U1319 ( .A(n1217), .Y(n1218) );
  AND2X1 U1320 ( .A(n3609), .B(n4679), .Y(n666) );
  INVX1 U1321 ( .A(n666), .Y(n1219) );
  INVX1 U1322 ( .A(n1222), .Y(n1220) );
  INVX1 U1323 ( .A(n1220), .Y(n1221) );
  AND2X1 U1324 ( .A(n3612), .B(n4679), .Y(n665) );
  INVX1 U1325 ( .A(n665), .Y(n1222) );
  INVX1 U1326 ( .A(n1225), .Y(n1223) );
  INVX1 U1327 ( .A(n1223), .Y(n1224) );
  AND2X1 U1328 ( .A(n3615), .B(n4679), .Y(n664) );
  INVX1 U1329 ( .A(n664), .Y(n1225) );
  INVX1 U1330 ( .A(n1228), .Y(n1226) );
  INVX1 U1331 ( .A(n1226), .Y(n1227) );
  AND2X1 U1332 ( .A(n3618), .B(n4679), .Y(n663) );
  INVX1 U1333 ( .A(n663), .Y(n1228) );
  INVX1 U1334 ( .A(n1231), .Y(n1229) );
  INVX1 U1335 ( .A(n1229), .Y(n1230) );
  AND2X1 U1336 ( .A(n3621), .B(n4679), .Y(n662) );
  INVX1 U1337 ( .A(n662), .Y(n1231) );
  INVX1 U1338 ( .A(n1234), .Y(n1232) );
  INVX1 U1339 ( .A(n1232), .Y(n1233) );
  AND2X1 U1340 ( .A(n3624), .B(n4679), .Y(n661) );
  INVX1 U1341 ( .A(n661), .Y(n1234) );
  INVX1 U1342 ( .A(n1237), .Y(n1235) );
  INVX1 U1343 ( .A(n1235), .Y(n1236) );
  AND2X1 U1344 ( .A(n3627), .B(n4679), .Y(n660) );
  INVX1 U1345 ( .A(n660), .Y(n1237) );
  INVX1 U1346 ( .A(n1240), .Y(n1238) );
  INVX1 U1347 ( .A(n1238), .Y(n1239) );
  AND2X1 U1348 ( .A(n3630), .B(n4679), .Y(n659) );
  INVX1 U1349 ( .A(n659), .Y(n1240) );
  INVX1 U1350 ( .A(n1243), .Y(n1241) );
  INVX1 U1351 ( .A(n1241), .Y(n1242) );
  AND2X1 U1352 ( .A(n3633), .B(n4679), .Y(n658) );
  INVX1 U1353 ( .A(n658), .Y(n1243) );
  INVX1 U1354 ( .A(n1246), .Y(n1244) );
  INVX1 U1355 ( .A(n1244), .Y(n1245) );
  AND2X1 U1356 ( .A(n3636), .B(n4679), .Y(n657) );
  INVX1 U1357 ( .A(n657), .Y(n1246) );
  INVX1 U1358 ( .A(n1249), .Y(n1247) );
  INVX1 U1359 ( .A(n1247), .Y(n1248) );
  AND2X1 U1360 ( .A(n4023), .B(n4682), .Y(n654) );
  INVX1 U1361 ( .A(n654), .Y(n1249) );
  INVX1 U1362 ( .A(n1252), .Y(n1250) );
  INVX1 U1363 ( .A(n1250), .Y(n1251) );
  AND2X1 U1364 ( .A(n4026), .B(n4682), .Y(n653) );
  INVX1 U1365 ( .A(n653), .Y(n1252) );
  INVX1 U1366 ( .A(n1255), .Y(n1253) );
  INVX1 U1367 ( .A(n1253), .Y(n1254) );
  AND2X1 U1368 ( .A(n4029), .B(n4682), .Y(n652) );
  INVX1 U1369 ( .A(n652), .Y(n1255) );
  INVX1 U1370 ( .A(n1258), .Y(n1256) );
  INVX1 U1371 ( .A(n1256), .Y(n1257) );
  AND2X1 U1372 ( .A(n4032), .B(n4682), .Y(n651) );
  INVX1 U1373 ( .A(n651), .Y(n1258) );
  INVX1 U1374 ( .A(n1261), .Y(n1259) );
  INVX1 U1375 ( .A(n1259), .Y(n1260) );
  AND2X1 U1376 ( .A(n4035), .B(n4682), .Y(n650) );
  INVX1 U1377 ( .A(n650), .Y(n1261) );
  INVX1 U1378 ( .A(n1264), .Y(n1262) );
  INVX1 U1379 ( .A(n1262), .Y(n1263) );
  AND2X1 U1380 ( .A(n4038), .B(n4682), .Y(n649) );
  INVX1 U1381 ( .A(n649), .Y(n1264) );
  INVX1 U1382 ( .A(n1267), .Y(n1265) );
  INVX1 U1383 ( .A(n1265), .Y(n1266) );
  AND2X1 U1384 ( .A(n4041), .B(n4682), .Y(n648) );
  INVX1 U1385 ( .A(n648), .Y(n1267) );
  INVX1 U1386 ( .A(n1270), .Y(n1268) );
  INVX1 U1387 ( .A(n1268), .Y(n1269) );
  AND2X1 U1388 ( .A(n4044), .B(n4682), .Y(n647) );
  INVX1 U1389 ( .A(n647), .Y(n1270) );
  INVX1 U1390 ( .A(n1273), .Y(n1271) );
  INVX1 U1391 ( .A(n1271), .Y(n1272) );
  AND2X1 U1392 ( .A(n4047), .B(n4682), .Y(n646) );
  INVX1 U1393 ( .A(n646), .Y(n1273) );
  INVX1 U1394 ( .A(n1276), .Y(n1274) );
  INVX1 U1395 ( .A(n1274), .Y(n1275) );
  AND2X1 U1396 ( .A(n4050), .B(n4682), .Y(n645) );
  INVX1 U1397 ( .A(n645), .Y(n1276) );
  INVX1 U1398 ( .A(n1279), .Y(n1277) );
  INVX1 U1399 ( .A(n1277), .Y(n1278) );
  AND2X1 U1400 ( .A(n4053), .B(n4682), .Y(n644) );
  INVX1 U1401 ( .A(n644), .Y(n1279) );
  INVX1 U1402 ( .A(n1282), .Y(n1280) );
  INVX1 U1403 ( .A(n1280), .Y(n1281) );
  AND2X1 U1404 ( .A(n4056), .B(n4682), .Y(n643) );
  INVX1 U1405 ( .A(n643), .Y(n1282) );
  INVX1 U1406 ( .A(n1285), .Y(n1283) );
  INVX1 U1407 ( .A(n1283), .Y(n1284) );
  AND2X1 U1408 ( .A(n4059), .B(n4682), .Y(n642) );
  INVX1 U1409 ( .A(n642), .Y(n1285) );
  INVX1 U1410 ( .A(n1288), .Y(n1286) );
  INVX1 U1411 ( .A(n1286), .Y(n1287) );
  AND2X1 U1412 ( .A(n4062), .B(n4682), .Y(n641) );
  INVX1 U1413 ( .A(n641), .Y(n1288) );
  INVX1 U1414 ( .A(n1291), .Y(n1289) );
  INVX1 U1415 ( .A(n1289), .Y(n1290) );
  AND2X1 U1416 ( .A(n4065), .B(n4682), .Y(n640) );
  INVX1 U1417 ( .A(n640), .Y(n1291) );
  INVX1 U1418 ( .A(n1294), .Y(n1292) );
  INVX1 U1419 ( .A(n1292), .Y(n1293) );
  AND2X1 U1420 ( .A(n4068), .B(n4682), .Y(n639) );
  INVX1 U1421 ( .A(n639), .Y(n1294) );
  INVX1 U1422 ( .A(n1297), .Y(n1295) );
  INVX1 U1423 ( .A(n1295), .Y(n1296) );
  AND2X1 U1424 ( .A(n3255), .B(n4685), .Y(n637) );
  INVX1 U1425 ( .A(n637), .Y(n1297) );
  INVX1 U1426 ( .A(n1300), .Y(n1298) );
  INVX1 U1427 ( .A(n1298), .Y(n1299) );
  AND2X1 U1428 ( .A(n3258), .B(n4685), .Y(n636) );
  INVX1 U1429 ( .A(n636), .Y(n1300) );
  INVX1 U1430 ( .A(n1303), .Y(n1301) );
  INVX1 U1431 ( .A(n1301), .Y(n1302) );
  AND2X1 U1432 ( .A(n3261), .B(n4685), .Y(n635) );
  INVX1 U1433 ( .A(n635), .Y(n1303) );
  INVX1 U1434 ( .A(n1306), .Y(n1304) );
  INVX1 U1435 ( .A(n1304), .Y(n1305) );
  AND2X1 U1436 ( .A(n3264), .B(n4685), .Y(n634) );
  INVX1 U1437 ( .A(n634), .Y(n1306) );
  INVX1 U1438 ( .A(n1309), .Y(n1307) );
  INVX1 U1439 ( .A(n1307), .Y(n1308) );
  AND2X1 U1440 ( .A(n3267), .B(n4685), .Y(n633) );
  INVX1 U1441 ( .A(n633), .Y(n1309) );
  INVX1 U1442 ( .A(n1312), .Y(n1310) );
  INVX1 U1443 ( .A(n1310), .Y(n1311) );
  AND2X1 U1444 ( .A(n3270), .B(n4685), .Y(n632) );
  INVX1 U1445 ( .A(n632), .Y(n1312) );
  INVX1 U1446 ( .A(n1315), .Y(n1313) );
  INVX1 U1447 ( .A(n1313), .Y(n1314) );
  AND2X1 U1448 ( .A(n3273), .B(n4685), .Y(n631) );
  INVX1 U1449 ( .A(n631), .Y(n1315) );
  INVX1 U1450 ( .A(n1318), .Y(n1316) );
  INVX1 U1451 ( .A(n1316), .Y(n1317) );
  AND2X1 U1452 ( .A(n3276), .B(n4685), .Y(n630) );
  INVX1 U1453 ( .A(n630), .Y(n1318) );
  INVX1 U1454 ( .A(n1321), .Y(n1319) );
  INVX1 U1455 ( .A(n1319), .Y(n1320) );
  AND2X1 U1456 ( .A(n3279), .B(n4685), .Y(n629) );
  INVX1 U1457 ( .A(n629), .Y(n1321) );
  INVX1 U1458 ( .A(n1324), .Y(n1322) );
  INVX1 U1459 ( .A(n1322), .Y(n1323) );
  AND2X1 U1460 ( .A(n3282), .B(n4685), .Y(n628) );
  INVX1 U1461 ( .A(n628), .Y(n1324) );
  INVX1 U1462 ( .A(n1368), .Y(n1325) );
  INVX1 U1463 ( .A(n1325), .Y(n1346) );
  AND2X1 U1464 ( .A(n3285), .B(n4685), .Y(n627) );
  INVX1 U1465 ( .A(n627), .Y(n1368) );
  INVX1 U1466 ( .A(n1932), .Y(n1401) );
  INVX1 U1467 ( .A(n1401), .Y(n1931) );
  AND2X1 U1468 ( .A(n3288), .B(n4685), .Y(n626) );
  INVX1 U1469 ( .A(n626), .Y(n1932) );
  INVX1 U1470 ( .A(n1935), .Y(n1933) );
  INVX1 U1471 ( .A(n1933), .Y(n1934) );
  AND2X1 U1472 ( .A(n3291), .B(n4685), .Y(n625) );
  INVX1 U1473 ( .A(n625), .Y(n1935) );
  INVX1 U1474 ( .A(n1938), .Y(n1936) );
  INVX1 U1475 ( .A(n1936), .Y(n1937) );
  AND2X1 U1476 ( .A(n3294), .B(n4685), .Y(n624) );
  INVX1 U1477 ( .A(n624), .Y(n1938) );
  INVX1 U1478 ( .A(n1941), .Y(n1939) );
  INVX1 U1479 ( .A(n1939), .Y(n1940) );
  AND2X1 U1480 ( .A(n3297), .B(n4685), .Y(n623) );
  INVX1 U1481 ( .A(n623), .Y(n1941) );
  INVX1 U1482 ( .A(n1944), .Y(n1942) );
  INVX1 U1483 ( .A(n1942), .Y(n1943) );
  AND2X1 U1484 ( .A(n3300), .B(n4685), .Y(n622) );
  INVX1 U1485 ( .A(n622), .Y(n1944) );
  INVX1 U1486 ( .A(n1947), .Y(n1945) );
  INVX1 U1487 ( .A(n1945), .Y(n1946) );
  AND2X1 U1488 ( .A(n3879), .B(n4688), .Y(n620) );
  INVX1 U1489 ( .A(n620), .Y(n1947) );
  INVX1 U1490 ( .A(n1950), .Y(n1948) );
  INVX1 U1491 ( .A(n1948), .Y(n1949) );
  AND2X1 U1492 ( .A(n3882), .B(n4688), .Y(n619) );
  INVX1 U1493 ( .A(n619), .Y(n1950) );
  INVX1 U1494 ( .A(n1953), .Y(n1951) );
  INVX1 U1495 ( .A(n1951), .Y(n1952) );
  AND2X1 U1496 ( .A(n3885), .B(n4688), .Y(n618) );
  INVX1 U1497 ( .A(n618), .Y(n1953) );
  INVX1 U1498 ( .A(n1956), .Y(n1954) );
  INVX1 U1499 ( .A(n1954), .Y(n1955) );
  AND2X1 U1500 ( .A(n3888), .B(n4688), .Y(n617) );
  INVX1 U1501 ( .A(n617), .Y(n1956) );
  INVX1 U1502 ( .A(n1959), .Y(n1957) );
  INVX1 U1503 ( .A(n1957), .Y(n1958) );
  AND2X1 U1504 ( .A(n3891), .B(n4688), .Y(n616) );
  INVX1 U1505 ( .A(n616), .Y(n1959) );
  INVX1 U1506 ( .A(n1962), .Y(n1960) );
  INVX1 U1507 ( .A(n1960), .Y(n1961) );
  AND2X1 U1508 ( .A(n3894), .B(n4688), .Y(n615) );
  INVX1 U1509 ( .A(n615), .Y(n1962) );
  INVX1 U1510 ( .A(n1965), .Y(n1963) );
  INVX1 U1511 ( .A(n1963), .Y(n1964) );
  AND2X1 U1512 ( .A(n3897), .B(n4688), .Y(n614) );
  INVX1 U1513 ( .A(n614), .Y(n1965) );
  INVX1 U1514 ( .A(n1968), .Y(n1966) );
  INVX1 U1515 ( .A(n1966), .Y(n1967) );
  AND2X1 U1516 ( .A(n3900), .B(n4688), .Y(n613) );
  INVX1 U1517 ( .A(n613), .Y(n1968) );
  INVX1 U1518 ( .A(n1971), .Y(n1969) );
  INVX1 U1519 ( .A(n1969), .Y(n1970) );
  AND2X1 U1520 ( .A(n3903), .B(n4688), .Y(n612) );
  INVX1 U1521 ( .A(n612), .Y(n1971) );
  INVX1 U1522 ( .A(n1974), .Y(n1972) );
  INVX1 U1523 ( .A(n1972), .Y(n1973) );
  AND2X1 U1524 ( .A(n3906), .B(n4688), .Y(n611) );
  INVX1 U1525 ( .A(n611), .Y(n1974) );
  INVX1 U1526 ( .A(n1977), .Y(n1975) );
  INVX1 U1527 ( .A(n1975), .Y(n1976) );
  AND2X1 U1528 ( .A(n3909), .B(n4688), .Y(n610) );
  INVX1 U1529 ( .A(n610), .Y(n1977) );
  INVX1 U1530 ( .A(n1980), .Y(n1978) );
  INVX1 U1531 ( .A(n1978), .Y(n1979) );
  AND2X1 U1532 ( .A(n3912), .B(n4688), .Y(n609) );
  INVX1 U1533 ( .A(n609), .Y(n1980) );
  INVX1 U1534 ( .A(n1983), .Y(n1981) );
  INVX1 U1535 ( .A(n1981), .Y(n1982) );
  AND2X1 U1536 ( .A(n3915), .B(n4688), .Y(n608) );
  INVX1 U1537 ( .A(n608), .Y(n1983) );
  INVX1 U1538 ( .A(n1986), .Y(n1984) );
  INVX1 U1539 ( .A(n1984), .Y(n1985) );
  AND2X1 U1540 ( .A(n3918), .B(n4688), .Y(n607) );
  INVX1 U1541 ( .A(n607), .Y(n1986) );
  INVX1 U1542 ( .A(n1989), .Y(n1987) );
  INVX1 U1543 ( .A(n1987), .Y(n1988) );
  AND2X1 U1544 ( .A(n3921), .B(n4688), .Y(n606) );
  INVX1 U1545 ( .A(n606), .Y(n1989) );
  INVX1 U1546 ( .A(n1992), .Y(n1990) );
  INVX1 U1547 ( .A(n1990), .Y(n1991) );
  AND2X1 U1548 ( .A(n3924), .B(n4688), .Y(n605) );
  INVX1 U1549 ( .A(n605), .Y(n1992) );
  INVX1 U1550 ( .A(n1995), .Y(n1993) );
  INVX1 U1551 ( .A(n1993), .Y(n1994) );
  AND2X1 U1552 ( .A(n3111), .B(n4691), .Y(n603) );
  INVX1 U1553 ( .A(n603), .Y(n1995) );
  INVX1 U1554 ( .A(n1998), .Y(n1996) );
  INVX1 U1555 ( .A(n1996), .Y(n1997) );
  AND2X1 U1556 ( .A(n3114), .B(n4691), .Y(n602) );
  INVX1 U1557 ( .A(n602), .Y(n1998) );
  INVX1 U1558 ( .A(n2001), .Y(n1999) );
  INVX1 U1559 ( .A(n1999), .Y(n2000) );
  AND2X1 U1560 ( .A(n3117), .B(n4691), .Y(n601) );
  INVX1 U1561 ( .A(n601), .Y(n2001) );
  INVX1 U1562 ( .A(n2004), .Y(n2002) );
  INVX1 U1563 ( .A(n2002), .Y(n2003) );
  AND2X1 U1564 ( .A(n3120), .B(n4691), .Y(n600) );
  INVX1 U1565 ( .A(n600), .Y(n2004) );
  INVX1 U1566 ( .A(n2007), .Y(n2005) );
  INVX1 U1567 ( .A(n2005), .Y(n2006) );
  AND2X1 U1568 ( .A(n3123), .B(n4691), .Y(n599) );
  INVX1 U1569 ( .A(n599), .Y(n2007) );
  INVX1 U1570 ( .A(n2010), .Y(n2008) );
  INVX1 U1571 ( .A(n2008), .Y(n2009) );
  AND2X1 U1572 ( .A(n3126), .B(n4691), .Y(n598) );
  INVX1 U1573 ( .A(n598), .Y(n2010) );
  INVX1 U1574 ( .A(n2013), .Y(n2011) );
  INVX1 U1575 ( .A(n2011), .Y(n2012) );
  AND2X1 U1576 ( .A(n3129), .B(n4691), .Y(n597) );
  INVX1 U1577 ( .A(n597), .Y(n2013) );
  INVX1 U1578 ( .A(n2016), .Y(n2014) );
  INVX1 U1579 ( .A(n2014), .Y(n2015) );
  AND2X1 U1580 ( .A(n3132), .B(n4691), .Y(n596) );
  INVX1 U1581 ( .A(n596), .Y(n2016) );
  INVX1 U1582 ( .A(n2019), .Y(n2017) );
  INVX1 U1583 ( .A(n2017), .Y(n2018) );
  AND2X1 U1584 ( .A(n3135), .B(n4691), .Y(n595) );
  INVX1 U1585 ( .A(n595), .Y(n2019) );
  INVX1 U1586 ( .A(n2022), .Y(n2020) );
  INVX1 U1587 ( .A(n2020), .Y(n2021) );
  AND2X1 U1588 ( .A(n3138), .B(n4691), .Y(n594) );
  INVX1 U1589 ( .A(n594), .Y(n2022) );
  INVX1 U1590 ( .A(n2025), .Y(n2023) );
  INVX1 U1591 ( .A(n2023), .Y(n2024) );
  AND2X1 U1592 ( .A(n3141), .B(n4691), .Y(n593) );
  INVX1 U1593 ( .A(n593), .Y(n2025) );
  INVX1 U1594 ( .A(n2028), .Y(n2026) );
  INVX1 U1595 ( .A(n2026), .Y(n2027) );
  AND2X1 U1596 ( .A(n3144), .B(n4691), .Y(n592) );
  INVX1 U1597 ( .A(n592), .Y(n2028) );
  INVX1 U1598 ( .A(n2031), .Y(n2029) );
  INVX1 U1599 ( .A(n2029), .Y(n2030) );
  AND2X1 U1600 ( .A(n3147), .B(n4691), .Y(n591) );
  INVX1 U1601 ( .A(n591), .Y(n2031) );
  INVX1 U1602 ( .A(n2034), .Y(n2032) );
  INVX1 U1603 ( .A(n2032), .Y(n2033) );
  AND2X1 U1604 ( .A(n3150), .B(n4691), .Y(n590) );
  INVX1 U1605 ( .A(n590), .Y(n2034) );
  INVX1 U1606 ( .A(n2037), .Y(n2035) );
  INVX1 U1607 ( .A(n2035), .Y(n2036) );
  AND2X1 U1608 ( .A(n3153), .B(n4691), .Y(n589) );
  INVX1 U1609 ( .A(n589), .Y(n2037) );
  INVX1 U1610 ( .A(n2040), .Y(n2038) );
  INVX1 U1611 ( .A(n2038), .Y(n2039) );
  AND2X1 U1612 ( .A(n3156), .B(n4691), .Y(n588) );
  INVX1 U1613 ( .A(n588), .Y(n2040) );
  INVX1 U1614 ( .A(n2043), .Y(n2041) );
  INVX1 U1615 ( .A(n2041), .Y(n2042) );
  AND2X1 U1616 ( .A(n3831), .B(n4694), .Y(n586) );
  INVX1 U1617 ( .A(n586), .Y(n2043) );
  INVX1 U1618 ( .A(n2046), .Y(n2044) );
  INVX1 U1619 ( .A(n2044), .Y(n2045) );
  AND2X1 U1620 ( .A(n3834), .B(n4694), .Y(n585) );
  INVX1 U1621 ( .A(n585), .Y(n2046) );
  INVX1 U1622 ( .A(n2049), .Y(n2047) );
  INVX1 U1623 ( .A(n2047), .Y(n2048) );
  AND2X1 U1624 ( .A(n3837), .B(n4694), .Y(n584) );
  INVX1 U1625 ( .A(n584), .Y(n2049) );
  INVX1 U1626 ( .A(n2052), .Y(n2050) );
  INVX1 U1627 ( .A(n2050), .Y(n2051) );
  AND2X1 U1628 ( .A(n3840), .B(n4694), .Y(n583) );
  INVX1 U1629 ( .A(n583), .Y(n2052) );
  INVX1 U1630 ( .A(n2055), .Y(n2053) );
  INVX1 U1631 ( .A(n2053), .Y(n2054) );
  AND2X1 U1632 ( .A(n3843), .B(n4694), .Y(n582) );
  INVX1 U1633 ( .A(n582), .Y(n2055) );
  INVX1 U1634 ( .A(n2058), .Y(n2056) );
  INVX1 U1635 ( .A(n2056), .Y(n2057) );
  AND2X1 U1636 ( .A(n3846), .B(n4694), .Y(n581) );
  INVX1 U1637 ( .A(n581), .Y(n2058) );
  INVX1 U1638 ( .A(n2061), .Y(n2059) );
  INVX1 U1639 ( .A(n2059), .Y(n2060) );
  AND2X1 U1640 ( .A(n3849), .B(n4694), .Y(n580) );
  INVX1 U1641 ( .A(n580), .Y(n2061) );
  INVX1 U1642 ( .A(n2064), .Y(n2062) );
  INVX1 U1643 ( .A(n2062), .Y(n2063) );
  AND2X1 U1644 ( .A(n3852), .B(n4694), .Y(n579) );
  INVX1 U1645 ( .A(n579), .Y(n2064) );
  INVX1 U1646 ( .A(n2067), .Y(n2065) );
  INVX1 U1647 ( .A(n2065), .Y(n2066) );
  AND2X1 U1648 ( .A(n3855), .B(n4694), .Y(n578) );
  INVX1 U1649 ( .A(n578), .Y(n2067) );
  INVX1 U1650 ( .A(n2070), .Y(n2068) );
  INVX1 U1651 ( .A(n2068), .Y(n2069) );
  AND2X1 U1652 ( .A(n3858), .B(n4694), .Y(n577) );
  INVX1 U1653 ( .A(n577), .Y(n2070) );
  INVX1 U1654 ( .A(n2073), .Y(n2071) );
  INVX1 U1655 ( .A(n2071), .Y(n2072) );
  AND2X1 U1656 ( .A(n3861), .B(n4694), .Y(n576) );
  INVX1 U1657 ( .A(n576), .Y(n2073) );
  INVX1 U1658 ( .A(n2076), .Y(n2074) );
  INVX1 U1659 ( .A(n2074), .Y(n2075) );
  AND2X1 U1660 ( .A(n3864), .B(n4694), .Y(n575) );
  INVX1 U1661 ( .A(n575), .Y(n2076) );
  INVX1 U1662 ( .A(n2079), .Y(n2077) );
  INVX1 U1663 ( .A(n2077), .Y(n2078) );
  AND2X1 U1664 ( .A(n3867), .B(n4694), .Y(n574) );
  INVX1 U1665 ( .A(n574), .Y(n2079) );
  INVX1 U1666 ( .A(n2082), .Y(n2080) );
  INVX1 U1667 ( .A(n2080), .Y(n2081) );
  AND2X1 U1668 ( .A(n3870), .B(n4694), .Y(n573) );
  INVX1 U1669 ( .A(n573), .Y(n2082) );
  INVX1 U1670 ( .A(n2085), .Y(n2083) );
  INVX1 U1671 ( .A(n2083), .Y(n2084) );
  AND2X1 U1672 ( .A(n3873), .B(n4694), .Y(n572) );
  INVX1 U1673 ( .A(n572), .Y(n2085) );
  INVX1 U1674 ( .A(n2088), .Y(n2086) );
  INVX1 U1675 ( .A(n2086), .Y(n2087) );
  AND2X1 U1676 ( .A(n3876), .B(n4694), .Y(n571) );
  INVX1 U1677 ( .A(n571), .Y(n2088) );
  INVX1 U1678 ( .A(n2091), .Y(n2089) );
  INVX1 U1679 ( .A(n2089), .Y(n2090) );
  AND2X1 U1680 ( .A(n3063), .B(n4697), .Y(n569) );
  INVX1 U1681 ( .A(n569), .Y(n2091) );
  INVX1 U1682 ( .A(n2094), .Y(n2092) );
  INVX1 U1683 ( .A(n2092), .Y(n2093) );
  AND2X1 U1684 ( .A(n3066), .B(n4697), .Y(n568) );
  INVX1 U1685 ( .A(n568), .Y(n2094) );
  INVX1 U1686 ( .A(n2097), .Y(n2095) );
  INVX1 U1687 ( .A(n2095), .Y(n2096) );
  AND2X1 U1688 ( .A(n3069), .B(n4697), .Y(n567) );
  INVX1 U1689 ( .A(n567), .Y(n2097) );
  INVX1 U1690 ( .A(n2100), .Y(n2098) );
  INVX1 U1691 ( .A(n2098), .Y(n2099) );
  AND2X1 U1692 ( .A(n3072), .B(n4697), .Y(n566) );
  INVX1 U1693 ( .A(n566), .Y(n2100) );
  INVX1 U1694 ( .A(n2103), .Y(n2101) );
  INVX1 U1695 ( .A(n2101), .Y(n2102) );
  AND2X1 U1696 ( .A(n3075), .B(n4697), .Y(n565) );
  INVX1 U1697 ( .A(n565), .Y(n2103) );
  INVX1 U1698 ( .A(n2106), .Y(n2104) );
  INVX1 U1699 ( .A(n2104), .Y(n2105) );
  AND2X1 U1700 ( .A(n3078), .B(n4697), .Y(n564) );
  INVX1 U1701 ( .A(n564), .Y(n2106) );
  INVX1 U1702 ( .A(n2109), .Y(n2107) );
  INVX1 U1703 ( .A(n2107), .Y(n2108) );
  AND2X1 U1704 ( .A(n3081), .B(n4697), .Y(n563) );
  INVX1 U1705 ( .A(n563), .Y(n2109) );
  INVX1 U1706 ( .A(n2112), .Y(n2110) );
  INVX1 U1707 ( .A(n2110), .Y(n2111) );
  AND2X1 U1708 ( .A(n3084), .B(n4697), .Y(n562) );
  INVX1 U1709 ( .A(n562), .Y(n2112) );
  INVX1 U1710 ( .A(n2115), .Y(n2113) );
  INVX1 U1711 ( .A(n2113), .Y(n2114) );
  AND2X1 U1712 ( .A(n3087), .B(n4697), .Y(n561) );
  INVX1 U1729 ( .A(n561), .Y(n2115) );
  INVX1 U1740 ( .A(n2118), .Y(n2116) );
  INVX1 U1764 ( .A(n2116), .Y(n2117) );
  AND2X1 U1777 ( .A(n3090), .B(n4697), .Y(n560) );
  INVX1 U1778 ( .A(n560), .Y(n2118) );
  INVX1 U1779 ( .A(n2121), .Y(n2119) );
  INVX1 U1780 ( .A(n2119), .Y(n2120) );
  AND2X1 U1781 ( .A(n3093), .B(n4697), .Y(n559) );
  INVX1 U1782 ( .A(n559), .Y(n2121) );
  INVX1 U1783 ( .A(n2124), .Y(n2122) );
  INVX1 U1784 ( .A(n2122), .Y(n2123) );
  AND2X1 U1785 ( .A(n3096), .B(n4697), .Y(n558) );
  INVX1 U1786 ( .A(n558), .Y(n2124) );
  INVX1 U1787 ( .A(n2127), .Y(n2125) );
  INVX1 U1788 ( .A(n2125), .Y(n2126) );
  AND2X1 U1789 ( .A(n3099), .B(n4697), .Y(n557) );
  INVX1 U1790 ( .A(n557), .Y(n2127) );
  INVX1 U1791 ( .A(n2130), .Y(n2128) );
  INVX1 U1792 ( .A(n2128), .Y(n2129) );
  AND2X1 U1793 ( .A(n3102), .B(n4697), .Y(n556) );
  INVX1 U1794 ( .A(n556), .Y(n2130) );
  INVX1 U1795 ( .A(n2133), .Y(n2131) );
  INVX1 U1796 ( .A(n2131), .Y(n2132) );
  AND2X1 U1797 ( .A(n3105), .B(n4697), .Y(n555) );
  INVX1 U1798 ( .A(n555), .Y(n2133) );
  INVX1 U1799 ( .A(n2136), .Y(n2134) );
  INVX1 U1800 ( .A(n2134), .Y(n2135) );
  AND2X1 U1801 ( .A(n3108), .B(n4697), .Y(n554) );
  INVX1 U1802 ( .A(n554), .Y(n2136) );
  INVX1 U1803 ( .A(n2139), .Y(n2137) );
  INVX1 U1804 ( .A(n2137), .Y(n2138) );
  AND2X1 U1805 ( .A(n4119), .B(n4700), .Y(n552) );
  INVX1 U1806 ( .A(n552), .Y(n2139) );
  INVX1 U1807 ( .A(n2142), .Y(n2140) );
  INVX1 U1808 ( .A(n2140), .Y(n2141) );
  AND2X1 U1809 ( .A(n4122), .B(n4700), .Y(n551) );
  INVX1 U1810 ( .A(n551), .Y(n2142) );
  INVX1 U1811 ( .A(n2145), .Y(n2143) );
  INVX1 U1812 ( .A(n2143), .Y(n2144) );
  AND2X1 U1813 ( .A(n4125), .B(n4700), .Y(n550) );
  INVX1 U1814 ( .A(n550), .Y(n2145) );
  INVX1 U1815 ( .A(n2148), .Y(n2146) );
  INVX1 U1816 ( .A(n2146), .Y(n2147) );
  AND2X1 U1817 ( .A(n4128), .B(n4700), .Y(n549) );
  INVX1 U1818 ( .A(n549), .Y(n2148) );
  INVX1 U1819 ( .A(n2151), .Y(n2149) );
  INVX1 U1820 ( .A(n2149), .Y(n2150) );
  AND2X1 U1821 ( .A(n4131), .B(n4700), .Y(n548) );
  INVX1 U1822 ( .A(n548), .Y(n2151) );
  INVX1 U1823 ( .A(n2154), .Y(n2152) );
  INVX1 U1824 ( .A(n2152), .Y(n2153) );
  AND2X1 U1825 ( .A(n4134), .B(n4700), .Y(n547) );
  INVX1 U1826 ( .A(n547), .Y(n2154) );
  INVX1 U1827 ( .A(n2157), .Y(n2155) );
  INVX1 U1828 ( .A(n2155), .Y(n2156) );
  AND2X1 U1829 ( .A(n4137), .B(n4700), .Y(n546) );
  INVX1 U1830 ( .A(n546), .Y(n2157) );
  INVX1 U1831 ( .A(n2160), .Y(n2158) );
  INVX1 U1832 ( .A(n2158), .Y(n2159) );
  AND2X1 U1833 ( .A(n4140), .B(n4700), .Y(n545) );
  INVX1 U1834 ( .A(n545), .Y(n2160) );
  INVX1 U1835 ( .A(n2163), .Y(n2161) );
  INVX1 U1836 ( .A(n2161), .Y(n2162) );
  AND2X1 U1837 ( .A(n4143), .B(n4700), .Y(n544) );
  INVX1 U1838 ( .A(n544), .Y(n2163) );
  INVX1 U1839 ( .A(n2166), .Y(n2164) );
  INVX1 U1840 ( .A(n2164), .Y(n2165) );
  AND2X1 U1841 ( .A(n4146), .B(n4700), .Y(n543) );
  INVX1 U1842 ( .A(n543), .Y(n2166) );
  INVX1 U1843 ( .A(n2169), .Y(n2167) );
  INVX1 U1844 ( .A(n2167), .Y(n2168) );
  AND2X1 U1845 ( .A(n4149), .B(n4700), .Y(n542) );
  INVX1 U1846 ( .A(n542), .Y(n2169) );
  INVX1 U1847 ( .A(n2172), .Y(n2170) );
  INVX1 U1848 ( .A(n2170), .Y(n2171) );
  AND2X1 U1849 ( .A(n4152), .B(n4700), .Y(n541) );
  INVX1 U1850 ( .A(n541), .Y(n2172) );
  INVX1 U1851 ( .A(n2175), .Y(n2173) );
  INVX1 U1852 ( .A(n2173), .Y(n2174) );
  AND2X1 U1853 ( .A(n4155), .B(n4700), .Y(n540) );
  INVX1 U1854 ( .A(n540), .Y(n2175) );
  INVX1 U1855 ( .A(n2178), .Y(n2176) );
  INVX1 U1856 ( .A(n2176), .Y(n2177) );
  AND2X1 U1857 ( .A(n4158), .B(n4700), .Y(n539) );
  INVX1 U1858 ( .A(n539), .Y(n2178) );
  INVX1 U1859 ( .A(n2181), .Y(n2179) );
  INVX1 U1860 ( .A(n2179), .Y(n2180) );
  AND2X1 U1861 ( .A(n4161), .B(n4700), .Y(n538) );
  INVX1 U1862 ( .A(n538), .Y(n2181) );
  INVX1 U1863 ( .A(n2184), .Y(n2182) );
  INVX1 U1864 ( .A(n2182), .Y(n2183) );
  AND2X1 U1865 ( .A(n4164), .B(n4700), .Y(n537) );
  INVX1 U1866 ( .A(n537), .Y(n2184) );
  INVX1 U1867 ( .A(n2187), .Y(n2185) );
  INVX1 U1868 ( .A(n2185), .Y(n2186) );
  AND2X1 U1869 ( .A(n3351), .B(n4703), .Y(n534) );
  INVX1 U1870 ( .A(n534), .Y(n2187) );
  INVX1 U1871 ( .A(n2190), .Y(n2188) );
  INVX1 U1872 ( .A(n2188), .Y(n2189) );
  AND2X1 U1873 ( .A(n3354), .B(n4703), .Y(n533) );
  INVX1 U1874 ( .A(n533), .Y(n2190) );
  INVX1 U1875 ( .A(n2193), .Y(n2191) );
  INVX1 U1876 ( .A(n2191), .Y(n2192) );
  AND2X1 U1877 ( .A(n3357), .B(n4703), .Y(n532) );
  INVX1 U1878 ( .A(n532), .Y(n2193) );
  INVX1 U1879 ( .A(n2196), .Y(n2194) );
  INVX1 U1880 ( .A(n2194), .Y(n2195) );
  AND2X1 U1881 ( .A(n3360), .B(n4703), .Y(n531) );
  INVX1 U1882 ( .A(n531), .Y(n2196) );
  INVX1 U1883 ( .A(n2199), .Y(n2197) );
  INVX1 U1884 ( .A(n2197), .Y(n2198) );
  AND2X1 U1885 ( .A(n3363), .B(n4703), .Y(n530) );
  INVX1 U1886 ( .A(n530), .Y(n2199) );
  INVX1 U1887 ( .A(n2202), .Y(n2200) );
  INVX1 U1888 ( .A(n2200), .Y(n2201) );
  AND2X1 U1889 ( .A(n3366), .B(n4703), .Y(n529) );
  INVX1 U1890 ( .A(n529), .Y(n2202) );
  INVX1 U1891 ( .A(n2205), .Y(n2203) );
  INVX1 U1892 ( .A(n2203), .Y(n2204) );
  AND2X1 U1893 ( .A(n3369), .B(n4703), .Y(n528) );
  INVX1 U1894 ( .A(n528), .Y(n2205) );
  INVX1 U1895 ( .A(n2208), .Y(n2206) );
  INVX1 U1896 ( .A(n2206), .Y(n2207) );
  AND2X1 U1897 ( .A(n3372), .B(n4703), .Y(n527) );
  INVX1 U1898 ( .A(n527), .Y(n2208) );
  INVX1 U1899 ( .A(n2211), .Y(n2209) );
  INVX1 U1900 ( .A(n2209), .Y(n2210) );
  AND2X1 U1901 ( .A(n3375), .B(n4703), .Y(n526) );
  INVX1 U1902 ( .A(n526), .Y(n2211) );
  INVX1 U1903 ( .A(n2214), .Y(n2212) );
  INVX1 U1904 ( .A(n2212), .Y(n2213) );
  AND2X1 U1905 ( .A(n3378), .B(n4703), .Y(n525) );
  INVX1 U1906 ( .A(n525), .Y(n2214) );
  INVX1 U1907 ( .A(n2217), .Y(n2215) );
  INVX1 U1908 ( .A(n2215), .Y(n2216) );
  AND2X1 U1909 ( .A(n3381), .B(n4703), .Y(n524) );
  INVX1 U1910 ( .A(n524), .Y(n2217) );
  INVX1 U1911 ( .A(n2220), .Y(n2218) );
  INVX1 U1912 ( .A(n2218), .Y(n2219) );
  AND2X1 U1913 ( .A(n3384), .B(n4703), .Y(n523) );
  INVX1 U1914 ( .A(n523), .Y(n2220) );
  INVX1 U1915 ( .A(n2223), .Y(n2221) );
  INVX1 U1916 ( .A(n2221), .Y(n2222) );
  AND2X1 U1917 ( .A(n3387), .B(n4703), .Y(n522) );
  INVX1 U1918 ( .A(n522), .Y(n2223) );
  INVX1 U1919 ( .A(n2226), .Y(n2224) );
  INVX1 U1920 ( .A(n2224), .Y(n2225) );
  AND2X1 U1921 ( .A(n3390), .B(n4703), .Y(n521) );
  INVX1 U1922 ( .A(n521), .Y(n2226) );
  INVX1 U1923 ( .A(n2229), .Y(n2227) );
  INVX1 U1924 ( .A(n2227), .Y(n2228) );
  AND2X1 U1925 ( .A(n3393), .B(n4703), .Y(n520) );
  INVX1 U1926 ( .A(n520), .Y(n2229) );
  INVX1 U1927 ( .A(n2232), .Y(n2230) );
  INVX1 U1928 ( .A(n2230), .Y(n2231) );
  AND2X1 U1929 ( .A(n3396), .B(n4703), .Y(n519) );
  INVX1 U1930 ( .A(n519), .Y(n2232) );
  INVX1 U1931 ( .A(n2235), .Y(n2233) );
  INVX1 U1932 ( .A(n2233), .Y(n2234) );
  AND2X1 U1933 ( .A(n4071), .B(n4706), .Y(n516) );
  INVX1 U1934 ( .A(n516), .Y(n2235) );
  INVX1 U1935 ( .A(n2238), .Y(n2236) );
  INVX1 U1936 ( .A(n2236), .Y(n2237) );
  AND2X1 U1937 ( .A(n4074), .B(n4706), .Y(n515) );
  INVX1 U1938 ( .A(n515), .Y(n2238) );
  INVX1 U1939 ( .A(n2241), .Y(n2239) );
  INVX1 U1940 ( .A(n2239), .Y(n2240) );
  AND2X1 U1941 ( .A(n4077), .B(n4706), .Y(n514) );
  INVX1 U1942 ( .A(n514), .Y(n2241) );
  INVX1 U1943 ( .A(n2244), .Y(n2242) );
  INVX1 U1944 ( .A(n2242), .Y(n2243) );
  AND2X1 U1945 ( .A(n4080), .B(n4706), .Y(n513) );
  INVX1 U1946 ( .A(n513), .Y(n2244) );
  INVX1 U1947 ( .A(n2247), .Y(n2245) );
  INVX1 U1948 ( .A(n2245), .Y(n2246) );
  AND2X1 U1949 ( .A(n4083), .B(n4706), .Y(n512) );
  INVX1 U1950 ( .A(n512), .Y(n2247) );
  INVX1 U1951 ( .A(n2250), .Y(n2248) );
  INVX1 U1952 ( .A(n2248), .Y(n2249) );
  AND2X1 U1953 ( .A(n4086), .B(n4706), .Y(n511) );
  INVX1 U1954 ( .A(n511), .Y(n2250) );
  INVX1 U1955 ( .A(n2253), .Y(n2251) );
  INVX1 U1956 ( .A(n2251), .Y(n2252) );
  AND2X1 U1957 ( .A(n4089), .B(n4706), .Y(n510) );
  INVX1 U1958 ( .A(n510), .Y(n2253) );
  INVX1 U1959 ( .A(n2256), .Y(n2254) );
  INVX1 U1960 ( .A(n2254), .Y(n2255) );
  AND2X1 U1961 ( .A(n4092), .B(n4706), .Y(n509) );
  INVX1 U1962 ( .A(n509), .Y(n2256) );
  INVX1 U1963 ( .A(n2259), .Y(n2257) );
  INVX1 U1964 ( .A(n2257), .Y(n2258) );
  AND2X1 U1965 ( .A(n4095), .B(n4706), .Y(n508) );
  INVX1 U1966 ( .A(n508), .Y(n2259) );
  INVX1 U1967 ( .A(n2262), .Y(n2260) );
  INVX1 U1968 ( .A(n2260), .Y(n2261) );
  AND2X1 U1969 ( .A(n4098), .B(n4706), .Y(n507) );
  INVX1 U1970 ( .A(n507), .Y(n2262) );
  INVX1 U1971 ( .A(n2265), .Y(n2263) );
  INVX1 U1972 ( .A(n2263), .Y(n2264) );
  AND2X1 U1973 ( .A(n4101), .B(n4706), .Y(n506) );
  INVX1 U1974 ( .A(n506), .Y(n2265) );
  INVX1 U1975 ( .A(n2268), .Y(n2266) );
  INVX1 U1976 ( .A(n2266), .Y(n2267) );
  AND2X1 U1977 ( .A(n4104), .B(n4706), .Y(n505) );
  INVX1 U1978 ( .A(n505), .Y(n2268) );
  INVX1 U1979 ( .A(n2271), .Y(n2269) );
  INVX1 U1980 ( .A(n2269), .Y(n2270) );
  AND2X1 U1981 ( .A(n4107), .B(n4706), .Y(n504) );
  INVX1 U1982 ( .A(n504), .Y(n2271) );
  INVX1 U1983 ( .A(n2274), .Y(n2272) );
  INVX1 U1984 ( .A(n2272), .Y(n2273) );
  AND2X1 U1985 ( .A(n4110), .B(n4706), .Y(n503) );
  INVX1 U1986 ( .A(n503), .Y(n2274) );
  INVX1 U1987 ( .A(n2277), .Y(n2275) );
  INVX1 U1988 ( .A(n2275), .Y(n2276) );
  AND2X1 U1989 ( .A(n4113), .B(n4706), .Y(n502) );
  INVX1 U1990 ( .A(n502), .Y(n2277) );
  INVX1 U1991 ( .A(n2280), .Y(n2278) );
  INVX1 U1992 ( .A(n2278), .Y(n2279) );
  AND2X1 U1993 ( .A(n4116), .B(n4706), .Y(n501) );
  INVX1 U1994 ( .A(n501), .Y(n2280) );
  INVX1 U1995 ( .A(n2283), .Y(n2281) );
  INVX1 U1996 ( .A(n2281), .Y(n2282) );
  AND2X1 U1997 ( .A(n3303), .B(n4709), .Y(n499) );
  INVX1 U1998 ( .A(n499), .Y(n2283) );
  INVX1 U1999 ( .A(n2286), .Y(n2284) );
  INVX1 U2000 ( .A(n2284), .Y(n2285) );
  AND2X1 U2001 ( .A(n3306), .B(n4709), .Y(n498) );
  INVX1 U2002 ( .A(n498), .Y(n2286) );
  INVX1 U2003 ( .A(n2289), .Y(n2287) );
  INVX1 U2004 ( .A(n2287), .Y(n2288) );
  AND2X1 U2005 ( .A(n3309), .B(n4709), .Y(n497) );
  INVX1 U2006 ( .A(n497), .Y(n2289) );
  INVX1 U2007 ( .A(n2292), .Y(n2290) );
  INVX1 U2008 ( .A(n2290), .Y(n2291) );
  AND2X1 U2009 ( .A(n3312), .B(n4709), .Y(n496) );
  INVX1 U2010 ( .A(n496), .Y(n2292) );
  INVX1 U2011 ( .A(n2295), .Y(n2293) );
  INVX1 U2012 ( .A(n2293), .Y(n2294) );
  AND2X1 U2013 ( .A(n3315), .B(n4709), .Y(n495) );
  INVX1 U2014 ( .A(n495), .Y(n2295) );
  INVX1 U2015 ( .A(n2298), .Y(n2296) );
  INVX1 U2016 ( .A(n2296), .Y(n2297) );
  AND2X1 U2017 ( .A(n3318), .B(n4709), .Y(n494) );
  INVX1 U2018 ( .A(n494), .Y(n2298) );
  INVX1 U2019 ( .A(n2301), .Y(n2299) );
  INVX1 U2020 ( .A(n2299), .Y(n2300) );
  AND2X1 U2021 ( .A(n3321), .B(n4709), .Y(n493) );
  INVX1 U2022 ( .A(n493), .Y(n2301) );
  INVX1 U2023 ( .A(n2304), .Y(n2302) );
  INVX1 U2024 ( .A(n2302), .Y(n2303) );
  AND2X1 U2025 ( .A(n3324), .B(n4709), .Y(n492) );
  INVX1 U2026 ( .A(n492), .Y(n2304) );
  INVX1 U2027 ( .A(n2307), .Y(n2305) );
  INVX1 U2028 ( .A(n2305), .Y(n2306) );
  AND2X1 U2029 ( .A(n3327), .B(n4709), .Y(n491) );
  INVX1 U2030 ( .A(n491), .Y(n2307) );
  INVX1 U2031 ( .A(n2310), .Y(n2308) );
  INVX1 U2032 ( .A(n2308), .Y(n2309) );
  AND2X1 U2033 ( .A(n3330), .B(n4709), .Y(n490) );
  INVX1 U2034 ( .A(n490), .Y(n2310) );
  INVX1 U2035 ( .A(n2313), .Y(n2311) );
  INVX1 U2036 ( .A(n2311), .Y(n2312) );
  AND2X1 U2037 ( .A(n3333), .B(n4709), .Y(n489) );
  INVX1 U2038 ( .A(n489), .Y(n2313) );
  INVX1 U2039 ( .A(n2316), .Y(n2314) );
  INVX1 U2040 ( .A(n2314), .Y(n2315) );
  AND2X1 U2041 ( .A(n3336), .B(n4709), .Y(n488) );
  INVX1 U2042 ( .A(n488), .Y(n2316) );
  INVX1 U2043 ( .A(n2319), .Y(n2317) );
  INVX1 U2044 ( .A(n2317), .Y(n2318) );
  AND2X1 U2045 ( .A(n3339), .B(n4709), .Y(n487) );
  INVX1 U2046 ( .A(n487), .Y(n2319) );
  INVX1 U2047 ( .A(n2322), .Y(n2320) );
  INVX1 U2048 ( .A(n2320), .Y(n2321) );
  AND2X1 U2049 ( .A(n3342), .B(n4709), .Y(n486) );
  INVX1 U2050 ( .A(n486), .Y(n2322) );
  INVX1 U2051 ( .A(n2325), .Y(n2323) );
  INVX1 U2052 ( .A(n2323), .Y(n2324) );
  AND2X1 U2053 ( .A(n3345), .B(n4709), .Y(n485) );
  INVX1 U2054 ( .A(n485), .Y(n2325) );
  INVX1 U2055 ( .A(n2328), .Y(n2326) );
  INVX1 U2056 ( .A(n2326), .Y(n2327) );
  AND2X1 U2057 ( .A(n3348), .B(n4709), .Y(n484) );
  INVX1 U2058 ( .A(n484), .Y(n2328) );
  INVX1 U2059 ( .A(n2331), .Y(n2329) );
  INVX1 U2060 ( .A(n2329), .Y(n2330) );
  AND2X1 U2061 ( .A(n3975), .B(n4712), .Y(n482) );
  INVX1 U2062 ( .A(n482), .Y(n2331) );
  INVX1 U2063 ( .A(n2334), .Y(n2332) );
  INVX1 U2064 ( .A(n2332), .Y(n2333) );
  AND2X1 U2065 ( .A(n3978), .B(n4712), .Y(n481) );
  INVX1 U2066 ( .A(n481), .Y(n2334) );
  INVX1 U2067 ( .A(n2337), .Y(n2335) );
  INVX1 U2068 ( .A(n2335), .Y(n2336) );
  AND2X1 U2069 ( .A(n3981), .B(n4712), .Y(n480) );
  INVX1 U2070 ( .A(n480), .Y(n2337) );
  INVX1 U2071 ( .A(n2340), .Y(n2338) );
  INVX1 U2072 ( .A(n2338), .Y(n2339) );
  AND2X1 U2073 ( .A(n3984), .B(n4712), .Y(n479) );
  INVX1 U2074 ( .A(n479), .Y(n2340) );
  INVX1 U2075 ( .A(n2343), .Y(n2341) );
  INVX1 U2076 ( .A(n2341), .Y(n2342) );
  AND2X1 U2077 ( .A(n3987), .B(n4712), .Y(n478) );
  INVX1 U2078 ( .A(n478), .Y(n2343) );
  INVX1 U2079 ( .A(n2346), .Y(n2344) );
  INVX1 U2080 ( .A(n2344), .Y(n2345) );
  AND2X1 U2081 ( .A(n3990), .B(n4712), .Y(n477) );
  INVX1 U2082 ( .A(n477), .Y(n2346) );
  INVX1 U2083 ( .A(n2349), .Y(n2347) );
  INVX1 U2084 ( .A(n2347), .Y(n2348) );
  AND2X1 U2085 ( .A(n3993), .B(n4712), .Y(n476) );
  INVX1 U2086 ( .A(n476), .Y(n2349) );
  INVX1 U2087 ( .A(n2352), .Y(n2350) );
  INVX1 U2088 ( .A(n2350), .Y(n2351) );
  AND2X1 U2089 ( .A(n3996), .B(n4712), .Y(n475) );
  INVX1 U2090 ( .A(n475), .Y(n2352) );
  INVX1 U2091 ( .A(n2355), .Y(n2353) );
  INVX1 U2092 ( .A(n2353), .Y(n2354) );
  AND2X1 U2093 ( .A(n3999), .B(n4712), .Y(n474) );
  INVX1 U2094 ( .A(n474), .Y(n2355) );
  INVX1 U2095 ( .A(n2358), .Y(n2356) );
  INVX1 U2096 ( .A(n2356), .Y(n2357) );
  AND2X1 U2097 ( .A(n4002), .B(n4712), .Y(n473) );
  INVX1 U2098 ( .A(n473), .Y(n2358) );
  INVX1 U2099 ( .A(n2361), .Y(n2359) );
  INVX1 U2100 ( .A(n2359), .Y(n2360) );
  AND2X1 U2101 ( .A(n4005), .B(n4712), .Y(n472) );
  INVX1 U2102 ( .A(n472), .Y(n2361) );
  INVX1 U2103 ( .A(n2364), .Y(n2362) );
  INVX1 U2104 ( .A(n2362), .Y(n2363) );
  AND2X1 U2105 ( .A(n4008), .B(n4712), .Y(n471) );
  INVX1 U2106 ( .A(n471), .Y(n2364) );
  INVX1 U2107 ( .A(n2367), .Y(n2365) );
  INVX1 U2108 ( .A(n2365), .Y(n2366) );
  AND2X1 U2109 ( .A(n4011), .B(n4712), .Y(n470) );
  INVX1 U2110 ( .A(n470), .Y(n2367) );
  INVX1 U2111 ( .A(n2370), .Y(n2368) );
  INVX1 U2112 ( .A(n2368), .Y(n2369) );
  AND2X1 U2113 ( .A(n4014), .B(n4712), .Y(n469) );
  INVX1 U2114 ( .A(n469), .Y(n2370) );
  INVX1 U2115 ( .A(n2373), .Y(n2371) );
  INVX1 U2116 ( .A(n2371), .Y(n2372) );
  AND2X1 U2117 ( .A(n4017), .B(n4712), .Y(n468) );
  INVX1 U2118 ( .A(n468), .Y(n2373) );
  INVX1 U2119 ( .A(n2376), .Y(n2374) );
  INVX1 U2120 ( .A(n2374), .Y(n2375) );
  AND2X1 U2121 ( .A(n4020), .B(n4712), .Y(n467) );
  INVX1 U2122 ( .A(n467), .Y(n2376) );
  INVX1 U2123 ( .A(n2379), .Y(n2377) );
  INVX1 U2124 ( .A(n2377), .Y(n2378) );
  AND2X1 U2125 ( .A(n3207), .B(n4715), .Y(n465) );
  INVX1 U2126 ( .A(n465), .Y(n2379) );
  INVX1 U2127 ( .A(n2382), .Y(n2380) );
  INVX1 U2128 ( .A(n2380), .Y(n2381) );
  AND2X1 U2129 ( .A(n3210), .B(n4715), .Y(n464) );
  INVX1 U2130 ( .A(n464), .Y(n2382) );
  INVX1 U2131 ( .A(n2385), .Y(n2383) );
  INVX1 U2132 ( .A(n2383), .Y(n2384) );
  AND2X1 U2133 ( .A(n3213), .B(n4715), .Y(n463) );
  INVX1 U2134 ( .A(n463), .Y(n2385) );
  INVX1 U2135 ( .A(n2388), .Y(n2386) );
  INVX1 U2136 ( .A(n2386), .Y(n2387) );
  AND2X1 U2137 ( .A(n3216), .B(n4715), .Y(n462) );
  INVX1 U2138 ( .A(n462), .Y(n2388) );
  INVX1 U2139 ( .A(n2391), .Y(n2389) );
  INVX1 U2140 ( .A(n2389), .Y(n2390) );
  AND2X1 U2141 ( .A(n3219), .B(n4715), .Y(n461) );
  INVX1 U2142 ( .A(n461), .Y(n2391) );
  INVX1 U2143 ( .A(n2394), .Y(n2392) );
  INVX1 U2144 ( .A(n2392), .Y(n2393) );
  AND2X1 U2145 ( .A(n3222), .B(n4715), .Y(n460) );
  INVX1 U2146 ( .A(n460), .Y(n2394) );
  INVX1 U2147 ( .A(n2397), .Y(n2395) );
  INVX1 U2148 ( .A(n2395), .Y(n2396) );
  AND2X1 U2149 ( .A(n3225), .B(n4715), .Y(n459) );
  INVX1 U2150 ( .A(n459), .Y(n2397) );
  INVX1 U2151 ( .A(n2400), .Y(n2398) );
  INVX1 U2152 ( .A(n2398), .Y(n2399) );
  AND2X1 U2153 ( .A(n3228), .B(n4715), .Y(n458) );
  INVX1 U2154 ( .A(n458), .Y(n2400) );
  INVX1 U2155 ( .A(n2403), .Y(n2401) );
  INVX1 U2156 ( .A(n2401), .Y(n2402) );
  AND2X1 U2157 ( .A(n3231), .B(n4715), .Y(n457) );
  INVX1 U2158 ( .A(n457), .Y(n2403) );
  INVX1 U2159 ( .A(n2406), .Y(n2404) );
  INVX1 U2160 ( .A(n2404), .Y(n2405) );
  AND2X1 U2161 ( .A(n3234), .B(n4715), .Y(n456) );
  INVX1 U2162 ( .A(n456), .Y(n2406) );
  INVX1 U2163 ( .A(n2409), .Y(n2407) );
  INVX1 U2164 ( .A(n2407), .Y(n2408) );
  AND2X1 U2165 ( .A(n3237), .B(n4715), .Y(n455) );
  INVX1 U2166 ( .A(n455), .Y(n2409) );
  INVX1 U2167 ( .A(n2412), .Y(n2410) );
  INVX1 U2168 ( .A(n2410), .Y(n2411) );
  AND2X1 U2169 ( .A(n3240), .B(n4715), .Y(n454) );
  INVX1 U2170 ( .A(n454), .Y(n2412) );
  INVX1 U2171 ( .A(n2415), .Y(n2413) );
  INVX1 U2172 ( .A(n2413), .Y(n2414) );
  AND2X1 U2173 ( .A(n3243), .B(n4715), .Y(n453) );
  INVX1 U2174 ( .A(n453), .Y(n2415) );
  INVX1 U2175 ( .A(n2418), .Y(n2416) );
  INVX1 U2176 ( .A(n2416), .Y(n2417) );
  AND2X1 U2177 ( .A(n3246), .B(n4715), .Y(n452) );
  INVX1 U2178 ( .A(n452), .Y(n2418) );
  INVX1 U2179 ( .A(n2421), .Y(n2419) );
  INVX1 U2180 ( .A(n2419), .Y(n2420) );
  AND2X1 U2181 ( .A(n3249), .B(n4715), .Y(n451) );
  INVX1 U2182 ( .A(n451), .Y(n2421) );
  INVX1 U2183 ( .A(n2424), .Y(n2422) );
  INVX1 U2184 ( .A(n2422), .Y(n2423) );
  AND2X1 U2185 ( .A(n3252), .B(n4715), .Y(n450) );
  INVX1 U2186 ( .A(n450), .Y(n2424) );
  INVX1 U2187 ( .A(n2427), .Y(n2425) );
  INVX1 U2188 ( .A(n2425), .Y(n2426) );
  AND2X1 U2189 ( .A(n3927), .B(n4718), .Y(n448) );
  INVX1 U2190 ( .A(n448), .Y(n2427) );
  INVX1 U2191 ( .A(n2430), .Y(n2428) );
  INVX1 U2192 ( .A(n2428), .Y(n2429) );
  AND2X1 U2193 ( .A(n3930), .B(n4718), .Y(n447) );
  INVX1 U2194 ( .A(n447), .Y(n2430) );
  INVX1 U2195 ( .A(n2433), .Y(n2431) );
  INVX1 U2196 ( .A(n2431), .Y(n2432) );
  AND2X1 U2197 ( .A(n3933), .B(n4718), .Y(n446) );
  INVX1 U2198 ( .A(n446), .Y(n2433) );
  INVX1 U2199 ( .A(n2436), .Y(n2434) );
  INVX1 U2200 ( .A(n2434), .Y(n2435) );
  AND2X1 U2201 ( .A(n3936), .B(n4718), .Y(n445) );
  INVX1 U2202 ( .A(n445), .Y(n2436) );
  INVX1 U2203 ( .A(n2439), .Y(n2437) );
  INVX1 U2204 ( .A(n2437), .Y(n2438) );
  AND2X1 U2205 ( .A(n3939), .B(n4718), .Y(n444) );
  INVX1 U2206 ( .A(n444), .Y(n2439) );
  INVX1 U2207 ( .A(n2442), .Y(n2440) );
  INVX1 U2208 ( .A(n2440), .Y(n2441) );
  AND2X1 U2209 ( .A(n3942), .B(n4718), .Y(n443) );
  INVX1 U2210 ( .A(n443), .Y(n2442) );
  INVX1 U2211 ( .A(n2445), .Y(n2443) );
  INVX1 U2212 ( .A(n2443), .Y(n2444) );
  AND2X1 U2213 ( .A(n3945), .B(n4718), .Y(n442) );
  INVX1 U2214 ( .A(n442), .Y(n2445) );
  INVX1 U2215 ( .A(n2448), .Y(n2446) );
  INVX1 U2216 ( .A(n2446), .Y(n2447) );
  AND2X1 U2217 ( .A(n3948), .B(n4718), .Y(n441) );
  INVX1 U2218 ( .A(n441), .Y(n2448) );
  INVX1 U2219 ( .A(n2451), .Y(n2449) );
  INVX1 U2220 ( .A(n2449), .Y(n2450) );
  AND2X1 U2221 ( .A(n3951), .B(n4718), .Y(n440) );
  INVX1 U2222 ( .A(n440), .Y(n2451) );
  INVX1 U2223 ( .A(n2454), .Y(n2452) );
  INVX1 U2224 ( .A(n2452), .Y(n2453) );
  AND2X1 U2225 ( .A(n3954), .B(n4718), .Y(n439) );
  INVX1 U2226 ( .A(n439), .Y(n2454) );
  INVX1 U2227 ( .A(n2457), .Y(n2455) );
  INVX1 U2228 ( .A(n2455), .Y(n2456) );
  AND2X1 U2229 ( .A(n3957), .B(n4718), .Y(n438) );
  INVX1 U2230 ( .A(n438), .Y(n2457) );
  INVX1 U2231 ( .A(n2460), .Y(n2458) );
  INVX1 U2232 ( .A(n2458), .Y(n2459) );
  AND2X1 U2233 ( .A(n3960), .B(n4718), .Y(n437) );
  INVX1 U2234 ( .A(n437), .Y(n2460) );
  INVX1 U2235 ( .A(n2463), .Y(n2461) );
  INVX1 U2236 ( .A(n2461), .Y(n2462) );
  AND2X1 U2237 ( .A(n3963), .B(n4718), .Y(n436) );
  INVX1 U2238 ( .A(n436), .Y(n2463) );
  INVX1 U2239 ( .A(n2466), .Y(n2464) );
  INVX1 U2240 ( .A(n2464), .Y(n2465) );
  AND2X1 U2241 ( .A(n3966), .B(n4718), .Y(n435) );
  INVX1 U2242 ( .A(n435), .Y(n2466) );
  INVX1 U2243 ( .A(n2469), .Y(n2467) );
  INVX1 U2244 ( .A(n2467), .Y(n2468) );
  AND2X1 U2245 ( .A(n3969), .B(n4718), .Y(n434) );
  INVX1 U2246 ( .A(n434), .Y(n2469) );
  INVX1 U2247 ( .A(n2472), .Y(n2470) );
  INVX1 U2248 ( .A(n2470), .Y(n2471) );
  AND2X1 U2249 ( .A(n3972), .B(n4718), .Y(n433) );
  INVX1 U2250 ( .A(n433), .Y(n2472) );
  INVX1 U2251 ( .A(n2475), .Y(n2473) );
  INVX1 U2252 ( .A(n2473), .Y(n2474) );
  AND2X1 U2253 ( .A(n3159), .B(n4721), .Y(n431) );
  INVX1 U2254 ( .A(n431), .Y(n2475) );
  INVX1 U2255 ( .A(n2478), .Y(n2476) );
  INVX1 U2256 ( .A(n2476), .Y(n2477) );
  AND2X1 U2257 ( .A(n3162), .B(n4721), .Y(n430) );
  INVX1 U2258 ( .A(n430), .Y(n2478) );
  INVX1 U2259 ( .A(n2481), .Y(n2479) );
  INVX1 U2260 ( .A(n2479), .Y(n2480) );
  AND2X1 U2261 ( .A(n3165), .B(n4721), .Y(n429) );
  INVX1 U2262 ( .A(n429), .Y(n2481) );
  INVX1 U2263 ( .A(n2484), .Y(n2482) );
  INVX1 U2264 ( .A(n2482), .Y(n2483) );
  AND2X1 U2265 ( .A(n3168), .B(n4721), .Y(n428) );
  INVX1 U2266 ( .A(n428), .Y(n2484) );
  INVX1 U2267 ( .A(n2487), .Y(n2485) );
  INVX1 U2268 ( .A(n2485), .Y(n2486) );
  AND2X1 U2269 ( .A(n3171), .B(n4721), .Y(n427) );
  INVX1 U2270 ( .A(n427), .Y(n2487) );
  INVX1 U2271 ( .A(n2490), .Y(n2488) );
  INVX1 U2272 ( .A(n2488), .Y(n2489) );
  AND2X1 U2273 ( .A(n3174), .B(n4721), .Y(n426) );
  INVX1 U2274 ( .A(n426), .Y(n2490) );
  INVX1 U2275 ( .A(n2493), .Y(n2491) );
  INVX1 U2276 ( .A(n2491), .Y(n2492) );
  AND2X1 U2277 ( .A(n3177), .B(n4721), .Y(n425) );
  INVX1 U2278 ( .A(n425), .Y(n2493) );
  INVX1 U2279 ( .A(n2496), .Y(n2494) );
  INVX1 U2280 ( .A(n2494), .Y(n2495) );
  AND2X1 U2281 ( .A(n3180), .B(n4721), .Y(n424) );
  INVX1 U2282 ( .A(n424), .Y(n2496) );
  INVX1 U2283 ( .A(n2499), .Y(n2497) );
  INVX1 U2284 ( .A(n2497), .Y(n2498) );
  AND2X1 U2285 ( .A(n3183), .B(n4721), .Y(n423) );
  INVX1 U2286 ( .A(n423), .Y(n2499) );
  INVX1 U2287 ( .A(n2502), .Y(n2500) );
  INVX1 U2288 ( .A(n2500), .Y(n2501) );
  AND2X1 U2289 ( .A(n3186), .B(n4721), .Y(n422) );
  INVX1 U2290 ( .A(n422), .Y(n2502) );
  INVX1 U2291 ( .A(n2505), .Y(n2503) );
  INVX1 U2292 ( .A(n2503), .Y(n2504) );
  AND2X1 U2293 ( .A(n3189), .B(n4721), .Y(n421) );
  INVX1 U2294 ( .A(n421), .Y(n2505) );
  INVX1 U2295 ( .A(n2508), .Y(n2506) );
  INVX1 U2296 ( .A(n2506), .Y(n2507) );
  AND2X1 U2297 ( .A(n3192), .B(n4721), .Y(n420) );
  INVX1 U2298 ( .A(n420), .Y(n2508) );
  INVX1 U2299 ( .A(n2511), .Y(n2509) );
  INVX1 U2300 ( .A(n2509), .Y(n2510) );
  AND2X1 U2301 ( .A(n3195), .B(n4721), .Y(n419) );
  INVX1 U2302 ( .A(n419), .Y(n2511) );
  INVX1 U2303 ( .A(n2514), .Y(n2512) );
  INVX1 U2304 ( .A(n2512), .Y(n2513) );
  AND2X1 U2305 ( .A(n3198), .B(n4721), .Y(n418) );
  INVX1 U2306 ( .A(n418), .Y(n2514) );
  INVX1 U2307 ( .A(n2517), .Y(n2515) );
  INVX1 U2308 ( .A(n2515), .Y(n2516) );
  AND2X1 U2309 ( .A(n3201), .B(n4721), .Y(n417) );
  INVX1 U2310 ( .A(n417), .Y(n2517) );
  INVX1 U2311 ( .A(n2520), .Y(n2518) );
  INVX1 U2312 ( .A(n2518), .Y(n2519) );
  AND2X1 U2313 ( .A(n3204), .B(n4721), .Y(n416) );
  INVX1 U2314 ( .A(n416), .Y(n2520) );
  INVX1 U2315 ( .A(n2523), .Y(n2521) );
  INVX1 U2316 ( .A(n2521), .Y(n2522) );
  AND2X1 U2317 ( .A(n4167), .B(n4724), .Y(n414) );
  INVX1 U2318 ( .A(n414), .Y(n2523) );
  INVX1 U2319 ( .A(n2526), .Y(n2524) );
  INVX1 U2320 ( .A(n2524), .Y(n2525) );
  AND2X1 U2321 ( .A(n4170), .B(n4724), .Y(n413) );
  INVX1 U2322 ( .A(n413), .Y(n2526) );
  INVX1 U2323 ( .A(n2529), .Y(n2527) );
  INVX1 U2324 ( .A(n2527), .Y(n2528) );
  AND2X1 U2325 ( .A(n4173), .B(n4724), .Y(n412) );
  INVX1 U2326 ( .A(n412), .Y(n2529) );
  INVX1 U2327 ( .A(n2532), .Y(n2530) );
  INVX1 U2328 ( .A(n2530), .Y(n2531) );
  AND2X1 U2329 ( .A(n4176), .B(n4724), .Y(n411) );
  INVX1 U2330 ( .A(n411), .Y(n2532) );
  INVX1 U2331 ( .A(n2535), .Y(n2533) );
  INVX1 U2332 ( .A(n2533), .Y(n2534) );
  AND2X1 U2333 ( .A(n4179), .B(n4724), .Y(n410) );
  INVX1 U2334 ( .A(n410), .Y(n2535) );
  INVX1 U2335 ( .A(n2538), .Y(n2536) );
  INVX1 U2336 ( .A(n2536), .Y(n2537) );
  AND2X1 U2337 ( .A(n4182), .B(n4724), .Y(n409) );
  INVX1 U2338 ( .A(n409), .Y(n2538) );
  INVX1 U2339 ( .A(n2541), .Y(n2539) );
  INVX1 U2340 ( .A(n2539), .Y(n2540) );
  AND2X1 U2341 ( .A(n4185), .B(n4724), .Y(n408) );
  INVX1 U2342 ( .A(n408), .Y(n2541) );
  INVX1 U2343 ( .A(n2544), .Y(n2542) );
  INVX1 U2344 ( .A(n2542), .Y(n2543) );
  AND2X1 U2345 ( .A(n4188), .B(n4724), .Y(n407) );
  INVX1 U2346 ( .A(n407), .Y(n2544) );
  INVX1 U2347 ( .A(n2547), .Y(n2545) );
  INVX1 U2348 ( .A(n2545), .Y(n2546) );
  AND2X1 U2349 ( .A(n4191), .B(n4724), .Y(n406) );
  INVX1 U2350 ( .A(n406), .Y(n2547) );
  INVX1 U2351 ( .A(n2550), .Y(n2548) );
  INVX1 U2352 ( .A(n2548), .Y(n2549) );
  AND2X1 U2353 ( .A(n4194), .B(n4724), .Y(n405) );
  INVX1 U2354 ( .A(n405), .Y(n2550) );
  INVX1 U2355 ( .A(n2553), .Y(n2551) );
  INVX1 U2356 ( .A(n2551), .Y(n2552) );
  AND2X1 U2357 ( .A(n4197), .B(n4724), .Y(n404) );
  INVX1 U2358 ( .A(n404), .Y(n2553) );
  INVX1 U2359 ( .A(n2556), .Y(n2554) );
  INVX1 U2360 ( .A(n2554), .Y(n2555) );
  AND2X1 U2361 ( .A(n4200), .B(n4724), .Y(n403) );
  INVX1 U2362 ( .A(n403), .Y(n2556) );
  INVX1 U2363 ( .A(n2559), .Y(n2557) );
  INVX1 U2364 ( .A(n2557), .Y(n2558) );
  AND2X1 U2365 ( .A(n4203), .B(n4724), .Y(n402) );
  INVX1 U2366 ( .A(n402), .Y(n2559) );
  INVX1 U2367 ( .A(n2562), .Y(n2560) );
  INVX1 U2368 ( .A(n2560), .Y(n2561) );
  AND2X1 U2369 ( .A(n4206), .B(n4724), .Y(n401) );
  INVX1 U2370 ( .A(n401), .Y(n2562) );
  INVX1 U2371 ( .A(n2565), .Y(n2563) );
  INVX1 U2372 ( .A(n2563), .Y(n2564) );
  AND2X1 U2373 ( .A(n4209), .B(n4724), .Y(n400) );
  INVX1 U2374 ( .A(n400), .Y(n2565) );
  INVX1 U2375 ( .A(n2568), .Y(n2566) );
  INVX1 U2376 ( .A(n2566), .Y(n2567) );
  AND2X1 U2377 ( .A(n4212), .B(n4724), .Y(n399) );
  INVX1 U2378 ( .A(n399), .Y(n2568) );
  INVX1 U2379 ( .A(n2571), .Y(n2569) );
  INVX1 U2380 ( .A(n2569), .Y(n2570) );
  AND2X1 U2381 ( .A(n3399), .B(n4727), .Y(n396) );
  INVX1 U2382 ( .A(n396), .Y(n2571) );
  INVX1 U2383 ( .A(n2574), .Y(n2572) );
  INVX1 U2384 ( .A(n2572), .Y(n2573) );
  AND2X1 U2385 ( .A(n3402), .B(n4727), .Y(n395) );
  INVX1 U2386 ( .A(n395), .Y(n2574) );
  INVX1 U2387 ( .A(n2577), .Y(n2575) );
  INVX1 U2388 ( .A(n2575), .Y(n2576) );
  AND2X1 U2389 ( .A(n3405), .B(n4727), .Y(n394) );
  INVX1 U2390 ( .A(n394), .Y(n2577) );
  INVX1 U2391 ( .A(n2580), .Y(n2578) );
  INVX1 U2392 ( .A(n2578), .Y(n2579) );
  AND2X1 U2393 ( .A(n3408), .B(n4727), .Y(n393) );
  INVX1 U2394 ( .A(n393), .Y(n2580) );
  INVX1 U2395 ( .A(n2583), .Y(n2581) );
  INVX1 U2396 ( .A(n2581), .Y(n2582) );
  AND2X1 U2397 ( .A(n3411), .B(n4727), .Y(n392) );
  INVX1 U2398 ( .A(n392), .Y(n2583) );
  INVX1 U2399 ( .A(n2586), .Y(n2584) );
  INVX1 U2400 ( .A(n2584), .Y(n2585) );
  AND2X1 U2401 ( .A(n3414), .B(n4727), .Y(n391) );
  INVX1 U2402 ( .A(n391), .Y(n2586) );
  INVX1 U2403 ( .A(n2589), .Y(n2587) );
  INVX1 U2404 ( .A(n2587), .Y(n2588) );
  AND2X1 U2405 ( .A(n3417), .B(n4727), .Y(n390) );
  INVX1 U2406 ( .A(n390), .Y(n2589) );
  INVX1 U2407 ( .A(n2592), .Y(n2590) );
  INVX1 U2408 ( .A(n2590), .Y(n2591) );
  AND2X1 U2409 ( .A(n3420), .B(n4727), .Y(n389) );
  INVX1 U2410 ( .A(n389), .Y(n2592) );
  INVX1 U2411 ( .A(n2595), .Y(n2593) );
  INVX1 U2412 ( .A(n2593), .Y(n2594) );
  AND2X1 U2413 ( .A(n3423), .B(n4727), .Y(n388) );
  INVX1 U2414 ( .A(n388), .Y(n2595) );
  INVX1 U2415 ( .A(n2598), .Y(n2596) );
  INVX1 U2416 ( .A(n2596), .Y(n2597) );
  AND2X1 U2417 ( .A(n3426), .B(n4727), .Y(n387) );
  INVX1 U2418 ( .A(n387), .Y(n2598) );
  INVX1 U2419 ( .A(n2601), .Y(n2599) );
  INVX1 U2420 ( .A(n2599), .Y(n2600) );
  AND2X1 U2421 ( .A(n3429), .B(n4727), .Y(n386) );
  INVX1 U2422 ( .A(n386), .Y(n2601) );
  INVX1 U2423 ( .A(n2604), .Y(n2602) );
  INVX1 U2424 ( .A(n2602), .Y(n2603) );
  AND2X1 U2425 ( .A(n3432), .B(n4727), .Y(n385) );
  INVX1 U2426 ( .A(n385), .Y(n2604) );
  INVX1 U2427 ( .A(n2607), .Y(n2605) );
  INVX1 U2428 ( .A(n2605), .Y(n2606) );
  AND2X1 U2429 ( .A(n3435), .B(n4727), .Y(n384) );
  INVX1 U2430 ( .A(n384), .Y(n2607) );
  INVX1 U2431 ( .A(n2610), .Y(n2608) );
  INVX1 U2432 ( .A(n2608), .Y(n2609) );
  AND2X1 U2433 ( .A(n3438), .B(n4727), .Y(n383) );
  INVX1 U2434 ( .A(n383), .Y(n2610) );
  INVX1 U2435 ( .A(n2613), .Y(n2611) );
  INVX1 U2436 ( .A(n2611), .Y(n2612) );
  AND2X1 U2437 ( .A(n3441), .B(n4727), .Y(n382) );
  INVX1 U2438 ( .A(n382), .Y(n2613) );
  INVX1 U2439 ( .A(n2616), .Y(n2614) );
  INVX1 U2440 ( .A(n2614), .Y(n2615) );
  AND2X1 U2441 ( .A(n3444), .B(n4727), .Y(n381) );
  INVX1 U2442 ( .A(n381), .Y(n2616) );
  INVX1 U2443 ( .A(n2619), .Y(n2617) );
  INVX1 U2444 ( .A(n2617), .Y(n2618) );
  AND2X1 U2445 ( .A(n4551), .B(n4730), .Y(n377) );
  INVX1 U2446 ( .A(n377), .Y(n2619) );
  INVX1 U2447 ( .A(n2622), .Y(n2620) );
  INVX1 U2448 ( .A(n2620), .Y(n2621) );
  AND2X1 U2449 ( .A(n4554), .B(n4730), .Y(n376) );
  INVX1 U2450 ( .A(n376), .Y(n2622) );
  INVX1 U2451 ( .A(n2625), .Y(n2623) );
  INVX1 U2452 ( .A(n2623), .Y(n2624) );
  AND2X1 U2453 ( .A(n4557), .B(n4730), .Y(n375) );
  INVX1 U2454 ( .A(n375), .Y(n2625) );
  INVX1 U2455 ( .A(n2628), .Y(n2626) );
  INVX1 U2456 ( .A(n2626), .Y(n2627) );
  AND2X1 U2457 ( .A(n4560), .B(n4730), .Y(n374) );
  INVX1 U2458 ( .A(n374), .Y(n2628) );
  INVX1 U2459 ( .A(n2631), .Y(n2629) );
  INVX1 U2460 ( .A(n2629), .Y(n2630) );
  AND2X1 U2461 ( .A(n4563), .B(n4730), .Y(n373) );
  INVX1 U2462 ( .A(n373), .Y(n2631) );
  INVX1 U2463 ( .A(n2634), .Y(n2632) );
  INVX1 U2464 ( .A(n2632), .Y(n2633) );
  AND2X1 U2465 ( .A(n4566), .B(n4730), .Y(n372) );
  INVX1 U2466 ( .A(n372), .Y(n2634) );
  INVX1 U2467 ( .A(n2637), .Y(n2635) );
  INVX1 U2468 ( .A(n2635), .Y(n2636) );
  AND2X1 U2469 ( .A(n4569), .B(n4730), .Y(n371) );
  INVX1 U2470 ( .A(n371), .Y(n2637) );
  INVX1 U2471 ( .A(n2640), .Y(n2638) );
  INVX1 U2472 ( .A(n2638), .Y(n2639) );
  AND2X1 U2473 ( .A(n4572), .B(n4730), .Y(n370) );
  INVX1 U2474 ( .A(n370), .Y(n2640) );
  INVX1 U2475 ( .A(n2643), .Y(n2641) );
  INVX1 U2476 ( .A(n2641), .Y(n2642) );
  AND2X1 U2477 ( .A(n4575), .B(n4730), .Y(n369) );
  INVX1 U2478 ( .A(n369), .Y(n2643) );
  INVX1 U2479 ( .A(n2646), .Y(n2644) );
  INVX1 U2480 ( .A(n2644), .Y(n2645) );
  AND2X1 U2481 ( .A(n4578), .B(n4730), .Y(n368) );
  INVX1 U2482 ( .A(n368), .Y(n2646) );
  INVX1 U2483 ( .A(n2649), .Y(n2647) );
  INVX1 U2484 ( .A(n2647), .Y(n2648) );
  AND2X1 U2485 ( .A(n4581), .B(n4730), .Y(n367) );
  INVX1 U2486 ( .A(n367), .Y(n2649) );
  INVX1 U2487 ( .A(n2652), .Y(n2650) );
  INVX1 U2488 ( .A(n2650), .Y(n2651) );
  AND2X1 U2489 ( .A(n4584), .B(n4730), .Y(n366) );
  INVX1 U2490 ( .A(n366), .Y(n2652) );
  INVX1 U2491 ( .A(n2655), .Y(n2653) );
  INVX1 U2492 ( .A(n2653), .Y(n2654) );
  AND2X1 U2493 ( .A(n4587), .B(n4730), .Y(n365) );
  INVX1 U2494 ( .A(n365), .Y(n2655) );
  INVX1 U2495 ( .A(n2658), .Y(n2656) );
  INVX1 U2496 ( .A(n2656), .Y(n2657) );
  AND2X1 U2497 ( .A(n4590), .B(n4730), .Y(n364) );
  INVX1 U2498 ( .A(n364), .Y(n2658) );
  INVX1 U2499 ( .A(n2661), .Y(n2659) );
  INVX1 U2500 ( .A(n2659), .Y(n2660) );
  AND2X1 U2501 ( .A(n4593), .B(n4730), .Y(n363) );
  INVX1 U2502 ( .A(n363), .Y(n2661) );
  INVX1 U2503 ( .A(n2664), .Y(n2662) );
  INVX1 U2504 ( .A(n2662), .Y(n2663) );
  AND2X1 U2505 ( .A(n4596), .B(n4730), .Y(n362) );
  INVX1 U2506 ( .A(n362), .Y(n2664) );
  INVX1 U2507 ( .A(n2667), .Y(n2665) );
  INVX1 U2508 ( .A(n2665), .Y(n2666) );
  AND2X1 U2509 ( .A(n3735), .B(n4733), .Y(n359) );
  INVX1 U2510 ( .A(n359), .Y(n2667) );
  INVX1 U2511 ( .A(n2670), .Y(n2668) );
  INVX1 U2512 ( .A(n2668), .Y(n2669) );
  AND2X1 U2513 ( .A(n3738), .B(n4733), .Y(n358) );
  INVX1 U2514 ( .A(n358), .Y(n2670) );
  INVX1 U2515 ( .A(n2673), .Y(n2671) );
  INVX1 U2516 ( .A(n2671), .Y(n2672) );
  AND2X1 U2517 ( .A(n3741), .B(n4733), .Y(n357) );
  INVX1 U2518 ( .A(n357), .Y(n2673) );
  INVX1 U2519 ( .A(n2676), .Y(n2674) );
  INVX1 U2520 ( .A(n2674), .Y(n2675) );
  AND2X1 U2521 ( .A(n3744), .B(n4733), .Y(n356) );
  INVX1 U2522 ( .A(n356), .Y(n2676) );
  INVX1 U2523 ( .A(n2679), .Y(n2677) );
  INVX1 U2524 ( .A(n2677), .Y(n2678) );
  AND2X1 U2525 ( .A(n3747), .B(n4733), .Y(n355) );
  INVX1 U2526 ( .A(n355), .Y(n2679) );
  INVX1 U2527 ( .A(n2682), .Y(n2680) );
  INVX1 U2528 ( .A(n2680), .Y(n2681) );
  AND2X1 U2529 ( .A(n3750), .B(n4733), .Y(n354) );
  INVX1 U2530 ( .A(n354), .Y(n2682) );
  INVX1 U2531 ( .A(n2685), .Y(n2683) );
  INVX1 U2532 ( .A(n2683), .Y(n2684) );
  AND2X1 U2533 ( .A(n3753), .B(n4733), .Y(n353) );
  INVX1 U2534 ( .A(n353), .Y(n2685) );
  INVX1 U2535 ( .A(n2688), .Y(n2686) );
  INVX1 U2536 ( .A(n2686), .Y(n2687) );
  AND2X1 U2537 ( .A(n3756), .B(n4733), .Y(n352) );
  INVX1 U2538 ( .A(n352), .Y(n2688) );
  INVX1 U2539 ( .A(n2691), .Y(n2689) );
  INVX1 U2540 ( .A(n2689), .Y(n2690) );
  AND2X1 U2541 ( .A(n3759), .B(n4733), .Y(n351) );
  INVX1 U2542 ( .A(n351), .Y(n2691) );
  INVX1 U2543 ( .A(n2694), .Y(n2692) );
  INVX1 U2544 ( .A(n2692), .Y(n2693) );
  AND2X1 U2545 ( .A(n3762), .B(n4733), .Y(n350) );
  INVX1 U2546 ( .A(n350), .Y(n2694) );
  INVX1 U2547 ( .A(n2697), .Y(n2695) );
  INVX1 U2548 ( .A(n2695), .Y(n2696) );
  AND2X1 U2549 ( .A(n3765), .B(n4733), .Y(n349) );
  INVX1 U2550 ( .A(n349), .Y(n2697) );
  INVX1 U2551 ( .A(n2700), .Y(n2698) );
  INVX1 U2552 ( .A(n2698), .Y(n2699) );
  AND2X1 U2553 ( .A(n3768), .B(n4733), .Y(n348) );
  INVX1 U2554 ( .A(n348), .Y(n2700) );
  INVX1 U2555 ( .A(n2703), .Y(n2701) );
  INVX1 U2556 ( .A(n2701), .Y(n2702) );
  AND2X1 U2557 ( .A(n3771), .B(n4733), .Y(n347) );
  INVX1 U2558 ( .A(n347), .Y(n2703) );
  INVX1 U2559 ( .A(n2706), .Y(n2704) );
  INVX1 U2560 ( .A(n2704), .Y(n2705) );
  AND2X1 U2561 ( .A(n3774), .B(n4733), .Y(n346) );
  INVX1 U2562 ( .A(n346), .Y(n2706) );
  INVX1 U2563 ( .A(n2709), .Y(n2707) );
  INVX1 U2564 ( .A(n2707), .Y(n2708) );
  AND2X1 U2565 ( .A(n3777), .B(n4733), .Y(n345) );
  INVX1 U2566 ( .A(n345), .Y(n2709) );
  INVX1 U2567 ( .A(n2712), .Y(n2710) );
  INVX1 U2568 ( .A(n2710), .Y(n2711) );
  AND2X1 U2569 ( .A(n3780), .B(n4733), .Y(n344) );
  INVX1 U2570 ( .A(n344), .Y(n2712) );
  INVX1 U2571 ( .A(n2715), .Y(n2713) );
  INVX1 U2572 ( .A(n2713), .Y(n2714) );
  AND2X1 U2573 ( .A(n4503), .B(n4736), .Y(n341) );
  INVX1 U2574 ( .A(n341), .Y(n2715) );
  INVX1 U2575 ( .A(n2718), .Y(n2716) );
  INVX1 U2576 ( .A(n2716), .Y(n2717) );
  AND2X1 U2577 ( .A(n4506), .B(n4736), .Y(n340) );
  INVX1 U2578 ( .A(n340), .Y(n2718) );
  INVX1 U2579 ( .A(n2721), .Y(n2719) );
  INVX1 U2580 ( .A(n2719), .Y(n2720) );
  AND2X1 U2581 ( .A(n4509), .B(n4736), .Y(n339) );
  INVX1 U2582 ( .A(n339), .Y(n2721) );
  INVX1 U2583 ( .A(n2724), .Y(n2722) );
  INVX1 U2584 ( .A(n2722), .Y(n2723) );
  AND2X1 U2585 ( .A(n4512), .B(n4736), .Y(n338) );
  INVX1 U2586 ( .A(n338), .Y(n2724) );
  INVX1 U2587 ( .A(n2727), .Y(n2725) );
  INVX1 U2588 ( .A(n2725), .Y(n2726) );
  AND2X1 U2589 ( .A(n4515), .B(n4736), .Y(n337) );
  INVX1 U2590 ( .A(n337), .Y(n2727) );
  INVX1 U2591 ( .A(n2730), .Y(n2728) );
  INVX1 U2592 ( .A(n2728), .Y(n2729) );
  AND2X1 U2593 ( .A(n4518), .B(n4736), .Y(n336) );
  INVX1 U2594 ( .A(n336), .Y(n2730) );
  INVX1 U2595 ( .A(n2733), .Y(n2731) );
  INVX1 U2596 ( .A(n2731), .Y(n2732) );
  AND2X1 U2597 ( .A(n4521), .B(n4736), .Y(n335) );
  INVX1 U2598 ( .A(n335), .Y(n2733) );
  INVX1 U2599 ( .A(n2736), .Y(n2734) );
  INVX1 U2600 ( .A(n2734), .Y(n2735) );
  AND2X1 U2601 ( .A(n4524), .B(n4736), .Y(n334) );
  INVX1 U2602 ( .A(n334), .Y(n2736) );
  INVX1 U2603 ( .A(n2739), .Y(n2737) );
  INVX1 U2604 ( .A(n2737), .Y(n2738) );
  AND2X1 U2605 ( .A(n4527), .B(n4736), .Y(n333) );
  INVX1 U2606 ( .A(n333), .Y(n2739) );
  INVX1 U2607 ( .A(n2742), .Y(n2740) );
  INVX1 U2608 ( .A(n2740), .Y(n2741) );
  AND2X1 U2609 ( .A(n4530), .B(n4736), .Y(n332) );
  INVX1 U2610 ( .A(n332), .Y(n2742) );
  INVX1 U2611 ( .A(n2745), .Y(n2743) );
  INVX1 U2612 ( .A(n2743), .Y(n2744) );
  AND2X1 U2613 ( .A(n4533), .B(n4736), .Y(n331) );
  INVX1 U2614 ( .A(n331), .Y(n2745) );
  INVX1 U2615 ( .A(n2748), .Y(n2746) );
  INVX1 U2616 ( .A(n2746), .Y(n2747) );
  AND2X1 U2617 ( .A(n4536), .B(n4736), .Y(n330) );
  INVX1 U2618 ( .A(n330), .Y(n2748) );
  INVX1 U2619 ( .A(n2751), .Y(n2749) );
  INVX1 U2620 ( .A(n2749), .Y(n2750) );
  AND2X1 U2621 ( .A(n4539), .B(n4736), .Y(n329) );
  INVX1 U2622 ( .A(n329), .Y(n2751) );
  INVX1 U2623 ( .A(n2754), .Y(n2752) );
  INVX1 U2624 ( .A(n2752), .Y(n2753) );
  AND2X1 U2625 ( .A(n4542), .B(n4736), .Y(n328) );
  INVX1 U2626 ( .A(n328), .Y(n2754) );
  INVX1 U2627 ( .A(n2757), .Y(n2755) );
  INVX1 U2628 ( .A(n2755), .Y(n2756) );
  AND2X1 U2629 ( .A(n4545), .B(n4736), .Y(n327) );
  INVX1 U2630 ( .A(n327), .Y(n2757) );
  INVX1 U2631 ( .A(n2760), .Y(n2758) );
  INVX1 U2632 ( .A(n2758), .Y(n2759) );
  AND2X1 U2633 ( .A(n4548), .B(n4736), .Y(n326) );
  INVX1 U2634 ( .A(n326), .Y(n2760) );
  INVX1 U2635 ( .A(n2763), .Y(n2761) );
  INVX1 U2636 ( .A(n2761), .Y(n2762) );
  AND2X1 U2637 ( .A(n3687), .B(n4739), .Y(n323) );
  INVX1 U2638 ( .A(n323), .Y(n2763) );
  INVX1 U2639 ( .A(n2766), .Y(n2764) );
  INVX1 U2640 ( .A(n2764), .Y(n2765) );
  AND2X1 U2641 ( .A(n3690), .B(n4739), .Y(n322) );
  INVX1 U2642 ( .A(n322), .Y(n2766) );
  INVX1 U2643 ( .A(n2769), .Y(n2767) );
  INVX1 U2644 ( .A(n2767), .Y(n2768) );
  AND2X1 U2645 ( .A(n3693), .B(n4739), .Y(n321) );
  INVX1 U2646 ( .A(n321), .Y(n2769) );
  INVX1 U2647 ( .A(n2772), .Y(n2770) );
  INVX1 U2648 ( .A(n2770), .Y(n2771) );
  AND2X1 U2649 ( .A(n3696), .B(n4739), .Y(n320) );
  INVX1 U2650 ( .A(n320), .Y(n2772) );
  INVX1 U2651 ( .A(n2775), .Y(n2773) );
  INVX1 U2652 ( .A(n2773), .Y(n2774) );
  AND2X1 U2653 ( .A(n3699), .B(n4739), .Y(n319) );
  INVX1 U2654 ( .A(n319), .Y(n2775) );
  INVX1 U2655 ( .A(n2778), .Y(n2776) );
  INVX1 U2656 ( .A(n2776), .Y(n2777) );
  AND2X1 U2657 ( .A(n3702), .B(n4739), .Y(n318) );
  INVX1 U2658 ( .A(n318), .Y(n2778) );
  INVX1 U2659 ( .A(n2781), .Y(n2779) );
  INVX1 U2660 ( .A(n2779), .Y(n2780) );
  AND2X1 U2661 ( .A(n3705), .B(n4739), .Y(n317) );
  INVX1 U2662 ( .A(n317), .Y(n2781) );
  INVX1 U2663 ( .A(n2784), .Y(n2782) );
  INVX1 U2664 ( .A(n2782), .Y(n2783) );
  AND2X1 U2665 ( .A(n3708), .B(n4739), .Y(n316) );
  INVX1 U2666 ( .A(n316), .Y(n2784) );
  INVX1 U2667 ( .A(n2787), .Y(n2785) );
  INVX1 U2668 ( .A(n2785), .Y(n2786) );
  AND2X1 U2669 ( .A(n3711), .B(n4739), .Y(n315) );
  INVX1 U2670 ( .A(n315), .Y(n2787) );
  INVX1 U2671 ( .A(n2790), .Y(n2788) );
  INVX1 U2672 ( .A(n2788), .Y(n2789) );
  AND2X1 U2673 ( .A(n3714), .B(n4739), .Y(n314) );
  INVX1 U2674 ( .A(n314), .Y(n2790) );
  INVX1 U2675 ( .A(n2793), .Y(n2791) );
  INVX1 U2676 ( .A(n2791), .Y(n2792) );
  AND2X1 U2677 ( .A(n3717), .B(n4739), .Y(n313) );
  INVX1 U2678 ( .A(n313), .Y(n2793) );
  INVX1 U2679 ( .A(n2796), .Y(n2794) );
  INVX1 U2680 ( .A(n2794), .Y(n2795) );
  AND2X1 U2681 ( .A(n3720), .B(n4739), .Y(n312) );
  INVX1 U2682 ( .A(n312), .Y(n2796) );
  INVX1 U2683 ( .A(n2799), .Y(n2797) );
  INVX1 U2684 ( .A(n2797), .Y(n2798) );
  AND2X1 U2685 ( .A(n3723), .B(n4739), .Y(n311) );
  INVX1 U2686 ( .A(n311), .Y(n2799) );
  INVX1 U2687 ( .A(n2802), .Y(n2800) );
  INVX1 U2688 ( .A(n2800), .Y(n2801) );
  AND2X1 U2689 ( .A(n3726), .B(n4739), .Y(n310) );
  INVX1 U2690 ( .A(n310), .Y(n2802) );
  INVX1 U2691 ( .A(n2805), .Y(n2803) );
  INVX1 U2692 ( .A(n2803), .Y(n2804) );
  AND2X1 U2693 ( .A(n3729), .B(n4739), .Y(n309) );
  INVX1 U2694 ( .A(n309), .Y(n2805) );
  INVX1 U2695 ( .A(n2808), .Y(n2806) );
  INVX1 U2696 ( .A(n2806), .Y(n2807) );
  AND2X1 U2697 ( .A(n3732), .B(n4739), .Y(n308) );
  INVX1 U2698 ( .A(n308), .Y(n2808) );
  INVX1 U2699 ( .A(n2811), .Y(n2809) );
  INVX1 U2700 ( .A(n2809), .Y(n2810) );
  AND2X1 U2701 ( .A(n4455), .B(n4742), .Y(n305) );
  INVX1 U2702 ( .A(n305), .Y(n2811) );
  INVX1 U2703 ( .A(n2814), .Y(n2812) );
  INVX1 U2704 ( .A(n2812), .Y(n2813) );
  AND2X1 U2705 ( .A(n4458), .B(n4742), .Y(n304) );
  INVX1 U2706 ( .A(n304), .Y(n2814) );
  INVX1 U2707 ( .A(n2817), .Y(n2815) );
  INVX1 U2708 ( .A(n2815), .Y(n2816) );
  AND2X1 U2709 ( .A(n4461), .B(n4742), .Y(n303) );
  INVX1 U2710 ( .A(n303), .Y(n2817) );
  INVX1 U2711 ( .A(n2820), .Y(n2818) );
  INVX1 U2712 ( .A(n2818), .Y(n2819) );
  AND2X1 U2713 ( .A(n4464), .B(n4742), .Y(n302) );
  INVX1 U2714 ( .A(n302), .Y(n2820) );
  INVX1 U2715 ( .A(n2823), .Y(n2821) );
  INVX1 U2716 ( .A(n2821), .Y(n2822) );
  AND2X1 U2717 ( .A(n4467), .B(n4742), .Y(n301) );
  INVX1 U2718 ( .A(n301), .Y(n2823) );
  INVX1 U2719 ( .A(n2826), .Y(n2824) );
  INVX1 U2720 ( .A(n2824), .Y(n2825) );
  AND2X1 U2721 ( .A(n4470), .B(n4742), .Y(n300) );
  INVX1 U2722 ( .A(n300), .Y(n2826) );
  INVX1 U2723 ( .A(n2829), .Y(n2827) );
  INVX1 U2724 ( .A(n2827), .Y(n2828) );
  AND2X1 U2725 ( .A(n4473), .B(n4742), .Y(n299) );
  INVX1 U2726 ( .A(n299), .Y(n2829) );
  INVX1 U2727 ( .A(n2832), .Y(n2830) );
  INVX1 U2728 ( .A(n2830), .Y(n2831) );
  AND2X1 U2729 ( .A(n4476), .B(n4742), .Y(n298) );
  INVX1 U2730 ( .A(n298), .Y(n2832) );
  INVX1 U2731 ( .A(n2835), .Y(n2833) );
  INVX1 U2732 ( .A(n2833), .Y(n2834) );
  AND2X1 U2733 ( .A(n4479), .B(n4742), .Y(n297) );
  INVX1 U2734 ( .A(n297), .Y(n2835) );
  INVX1 U2735 ( .A(n2838), .Y(n2836) );
  INVX1 U2736 ( .A(n2836), .Y(n2837) );
  AND2X1 U2737 ( .A(n4482), .B(n4742), .Y(n296) );
  INVX1 U2738 ( .A(n296), .Y(n2838) );
  INVX1 U2739 ( .A(n2841), .Y(n2839) );
  INVX1 U2740 ( .A(n2839), .Y(n2840) );
  AND2X1 U2741 ( .A(n4485), .B(n4742), .Y(n295) );
  INVX1 U2742 ( .A(n295), .Y(n2841) );
  INVX1 U2743 ( .A(n2844), .Y(n2842) );
  INVX1 U2744 ( .A(n2842), .Y(n2843) );
  AND2X1 U2745 ( .A(n4488), .B(n4742), .Y(n294) );
  INVX1 U2746 ( .A(n294), .Y(n2844) );
  INVX1 U2747 ( .A(n2847), .Y(n2845) );
  INVX1 U2748 ( .A(n2845), .Y(n2846) );
  AND2X1 U2749 ( .A(n4491), .B(n4742), .Y(n293) );
  INVX1 U2750 ( .A(n293), .Y(n2847) );
  INVX1 U2751 ( .A(n2850), .Y(n2848) );
  INVX1 U2752 ( .A(n2848), .Y(n2849) );
  AND2X1 U2753 ( .A(n4494), .B(n4742), .Y(n292) );
  INVX1 U2754 ( .A(n292), .Y(n2850) );
  INVX1 U2755 ( .A(n2853), .Y(n2851) );
  INVX1 U2756 ( .A(n2851), .Y(n2852) );
  AND2X1 U2757 ( .A(n4497), .B(n4742), .Y(n291) );
  INVX1 U2758 ( .A(n291), .Y(n2853) );
  INVX1 U2759 ( .A(n2856), .Y(n2854) );
  INVX1 U2760 ( .A(n2854), .Y(n2855) );
  AND2X1 U2761 ( .A(n4500), .B(n4742), .Y(n290) );
  INVX1 U2762 ( .A(n290), .Y(n2856) );
  INVX1 U2763 ( .A(n2859), .Y(n2857) );
  INVX1 U2764 ( .A(n2857), .Y(n2858) );
  AND2X1 U2765 ( .A(n3639), .B(n4745), .Y(n287) );
  INVX1 U2766 ( .A(n287), .Y(n2859) );
  INVX1 U2767 ( .A(n2862), .Y(n2860) );
  INVX1 U2768 ( .A(n2860), .Y(n2861) );
  AND2X1 U2769 ( .A(n3642), .B(n4745), .Y(n286) );
  INVX1 U2770 ( .A(n286), .Y(n2862) );
  INVX1 U2771 ( .A(n2865), .Y(n2863) );
  INVX1 U2772 ( .A(n2863), .Y(n2864) );
  AND2X1 U2773 ( .A(n3645), .B(n4745), .Y(n285) );
  INVX1 U2774 ( .A(n285), .Y(n2865) );
  INVX1 U2775 ( .A(n2868), .Y(n2866) );
  INVX1 U2776 ( .A(n2866), .Y(n2867) );
  AND2X1 U2777 ( .A(n3648), .B(n4745), .Y(n284) );
  INVX1 U2778 ( .A(n284), .Y(n2868) );
  INVX1 U2779 ( .A(n2871), .Y(n2869) );
  INVX1 U2780 ( .A(n2869), .Y(n2870) );
  AND2X1 U2781 ( .A(n3651), .B(n4745), .Y(n283) );
  INVX1 U2782 ( .A(n283), .Y(n2871) );
  INVX1 U2783 ( .A(n2874), .Y(n2872) );
  INVX1 U2784 ( .A(n2872), .Y(n2873) );
  AND2X1 U2785 ( .A(n3654), .B(n4745), .Y(n282) );
  INVX1 U2786 ( .A(n282), .Y(n2874) );
  INVX1 U2787 ( .A(n2877), .Y(n2875) );
  INVX1 U2788 ( .A(n2875), .Y(n2876) );
  AND2X1 U2789 ( .A(n3657), .B(n4745), .Y(n281) );
  INVX1 U2790 ( .A(n281), .Y(n2877) );
  INVX1 U2791 ( .A(n2880), .Y(n2878) );
  INVX1 U2792 ( .A(n2878), .Y(n2879) );
  AND2X1 U2793 ( .A(n3660), .B(n4745), .Y(n280) );
  INVX1 U2794 ( .A(n280), .Y(n2880) );
  INVX1 U2795 ( .A(n2883), .Y(n2881) );
  INVX1 U2796 ( .A(n2881), .Y(n2882) );
  AND2X1 U2797 ( .A(n3663), .B(n4745), .Y(n279) );
  INVX1 U2798 ( .A(n279), .Y(n2883) );
  INVX1 U2799 ( .A(n2886), .Y(n2884) );
  INVX1 U2800 ( .A(n2884), .Y(n2885) );
  AND2X1 U2801 ( .A(n3666), .B(n4745), .Y(n278) );
  INVX1 U2802 ( .A(n278), .Y(n2886) );
  INVX1 U2803 ( .A(n2889), .Y(n2887) );
  INVX1 U2804 ( .A(n2887), .Y(n2888) );
  AND2X1 U2805 ( .A(n3669), .B(n4745), .Y(n277) );
  INVX1 U2806 ( .A(n277), .Y(n2889) );
  INVX1 U2807 ( .A(n2892), .Y(n2890) );
  INVX1 U2808 ( .A(n2890), .Y(n2891) );
  AND2X1 U2809 ( .A(n3672), .B(n4745), .Y(n276) );
  INVX1 U2810 ( .A(n276), .Y(n2892) );
  INVX1 U2811 ( .A(n2895), .Y(n2893) );
  INVX1 U2812 ( .A(n2893), .Y(n2894) );
  AND2X1 U2813 ( .A(n3675), .B(n4745), .Y(n275) );
  INVX1 U2814 ( .A(n275), .Y(n2895) );
  INVX1 U2815 ( .A(n2898), .Y(n2896) );
  INVX1 U2816 ( .A(n2896), .Y(n2897) );
  AND2X1 U2817 ( .A(n3678), .B(n4745), .Y(n274) );
  INVX1 U2818 ( .A(n274), .Y(n2898) );
  INVX1 U2819 ( .A(n2901), .Y(n2899) );
  INVX1 U2820 ( .A(n2899), .Y(n2900) );
  AND2X1 U2821 ( .A(n3681), .B(n4745), .Y(n273) );
  INVX1 U2822 ( .A(n273), .Y(n2901) );
  INVX1 U2823 ( .A(n2904), .Y(n2902) );
  INVX1 U2824 ( .A(n2902), .Y(n2903) );
  AND2X1 U2825 ( .A(n3684), .B(n4745), .Y(n272) );
  INVX1 U2826 ( .A(n272), .Y(n2904) );
  INVX1 U2827 ( .A(n2907), .Y(n2905) );
  INVX1 U2828 ( .A(n2905), .Y(n2906) );
  AND2X1 U2829 ( .A(n4407), .B(n4748), .Y(n269) );
  INVX1 U2830 ( .A(n269), .Y(n2907) );
  INVX1 U2831 ( .A(n2910), .Y(n2908) );
  INVX1 U2832 ( .A(n2908), .Y(n2909) );
  AND2X1 U2833 ( .A(n4410), .B(n4748), .Y(n268) );
  INVX1 U2834 ( .A(n268), .Y(n2910) );
  INVX1 U2835 ( .A(n2913), .Y(n2911) );
  INVX1 U2836 ( .A(n2911), .Y(n2912) );
  AND2X1 U2837 ( .A(n4413), .B(n4748), .Y(n267) );
  INVX1 U2838 ( .A(n267), .Y(n2913) );
  INVX1 U2839 ( .A(n2916), .Y(n2914) );
  INVX1 U2840 ( .A(n2914), .Y(n2915) );
  AND2X1 U2841 ( .A(n4416), .B(n4748), .Y(n266) );
  INVX1 U2842 ( .A(n266), .Y(n2916) );
  INVX1 U2843 ( .A(n2919), .Y(n2917) );
  INVX1 U2844 ( .A(n2917), .Y(n2918) );
  AND2X1 U2845 ( .A(n4419), .B(n4748), .Y(n265) );
  INVX1 U2846 ( .A(n265), .Y(n2919) );
  INVX1 U2847 ( .A(n2922), .Y(n2920) );
  INVX1 U2848 ( .A(n2920), .Y(n2921) );
  AND2X1 U2849 ( .A(n4422), .B(n4748), .Y(n264) );
  INVX1 U2850 ( .A(n264), .Y(n2922) );
  INVX1 U2851 ( .A(n2925), .Y(n2923) );
  INVX1 U2852 ( .A(n2923), .Y(n2924) );
  AND2X1 U2853 ( .A(n4425), .B(n4748), .Y(n263) );
  INVX1 U2854 ( .A(n263), .Y(n2925) );
  INVX1 U2855 ( .A(n2928), .Y(n2926) );
  INVX1 U2856 ( .A(n2926), .Y(n2927) );
  AND2X1 U2857 ( .A(n4428), .B(n4748), .Y(n262) );
  INVX1 U2858 ( .A(n262), .Y(n2928) );
  INVX1 U2859 ( .A(n2931), .Y(n2929) );
  INVX1 U2860 ( .A(n2929), .Y(n2930) );
  AND2X1 U2861 ( .A(n4431), .B(n4748), .Y(n261) );
  INVX1 U2862 ( .A(n261), .Y(n2931) );
  INVX1 U2863 ( .A(n2934), .Y(n2932) );
  INVX1 U2864 ( .A(n2932), .Y(n2933) );
  AND2X1 U2865 ( .A(n4434), .B(n4748), .Y(n260) );
  INVX1 U2866 ( .A(n260), .Y(n2934) );
  INVX1 U2867 ( .A(n2937), .Y(n2935) );
  INVX1 U2868 ( .A(n2935), .Y(n2936) );
  AND2X1 U2869 ( .A(n4437), .B(n4748), .Y(n259) );
  INVX1 U2870 ( .A(n259), .Y(n2937) );
  INVX1 U2871 ( .A(n2940), .Y(n2938) );
  INVX1 U2872 ( .A(n2938), .Y(n2939) );
  AND2X1 U2873 ( .A(n4440), .B(n4748), .Y(n258) );
  INVX1 U2874 ( .A(n258), .Y(n2940) );
  INVX1 U2875 ( .A(n2943), .Y(n2941) );
  INVX1 U2876 ( .A(n2941), .Y(n2942) );
  AND2X1 U2877 ( .A(n4443), .B(n4748), .Y(n257) );
  INVX1 U2878 ( .A(n257), .Y(n2943) );
  INVX1 U2879 ( .A(n2946), .Y(n2944) );
  INVX1 U2880 ( .A(n2944), .Y(n2945) );
  AND2X1 U2881 ( .A(n4446), .B(n4748), .Y(n256) );
  INVX1 U2882 ( .A(n256), .Y(n2946) );
  INVX1 U2883 ( .A(n2949), .Y(n2947) );
  INVX1 U2884 ( .A(n2947), .Y(n2948) );
  AND2X1 U2885 ( .A(n4449), .B(n4748), .Y(n255) );
  INVX1 U2886 ( .A(n255), .Y(n2949) );
  INVX1 U2887 ( .A(n2952), .Y(n2950) );
  INVX1 U2888 ( .A(n2950), .Y(n2951) );
  AND2X1 U2889 ( .A(n4452), .B(n4748), .Y(n254) );
  INVX1 U2890 ( .A(n254), .Y(n2952) );
  INVX1 U2891 ( .A(n2955), .Y(n2953) );
  INVX1 U2892 ( .A(n2953), .Y(n2954) );
  AND2X1 U2893 ( .A(n3783), .B(n4655), .Y(n250) );
  INVX1 U2894 ( .A(n250), .Y(n2955) );
  INVX1 U2895 ( .A(n2958), .Y(n2956) );
  INVX1 U2896 ( .A(n2956), .Y(n2957) );
  AND2X1 U2897 ( .A(n3786), .B(n4655), .Y(n248) );
  INVX1 U2898 ( .A(n248), .Y(n2958) );
  INVX1 U2899 ( .A(n2961), .Y(n2959) );
  INVX1 U2900 ( .A(n2959), .Y(n2960) );
  AND2X1 U2901 ( .A(n3789), .B(n4655), .Y(n246) );
  INVX1 U2902 ( .A(n246), .Y(n2961) );
  INVX1 U2903 ( .A(n2964), .Y(n2962) );
  INVX1 U2904 ( .A(n2962), .Y(n2963) );
  AND2X1 U2905 ( .A(n3792), .B(n4655), .Y(n244) );
  INVX1 U2906 ( .A(n244), .Y(n2964) );
  INVX1 U2907 ( .A(n2967), .Y(n2965) );
  INVX1 U2908 ( .A(n2965), .Y(n2966) );
  AND2X1 U2909 ( .A(n3795), .B(n4655), .Y(n242) );
  INVX1 U2910 ( .A(n242), .Y(n2967) );
  INVX1 U2911 ( .A(n2970), .Y(n2968) );
  INVX1 U2912 ( .A(n2968), .Y(n2969) );
  AND2X1 U2913 ( .A(n3798), .B(n4655), .Y(n240) );
  INVX1 U2914 ( .A(n240), .Y(n2970) );
  INVX1 U2915 ( .A(n2973), .Y(n2971) );
  INVX1 U2916 ( .A(n2971), .Y(n2972) );
  AND2X1 U2917 ( .A(n3801), .B(n4655), .Y(n238) );
  INVX1 U2918 ( .A(n238), .Y(n2973) );
  INVX1 U2919 ( .A(n2976), .Y(n2974) );
  INVX1 U2920 ( .A(n2974), .Y(n2975) );
  AND2X1 U2921 ( .A(n3804), .B(n4655), .Y(n236) );
  INVX1 U2922 ( .A(n236), .Y(n2976) );
  INVX1 U2923 ( .A(n2979), .Y(n2977) );
  INVX1 U2924 ( .A(n2977), .Y(n2978) );
  AND2X1 U2925 ( .A(n3807), .B(n4655), .Y(n234) );
  INVX1 U2926 ( .A(n234), .Y(n2979) );
  INVX1 U2927 ( .A(n2982), .Y(n2980) );
  INVX1 U2928 ( .A(n2980), .Y(n2981) );
  AND2X1 U2929 ( .A(n3810), .B(n4655), .Y(n232) );
  INVX1 U2930 ( .A(n232), .Y(n2982) );
  INVX1 U2931 ( .A(n2985), .Y(n2983) );
  INVX1 U2932 ( .A(n2983), .Y(n2984) );
  AND2X1 U2933 ( .A(n3813), .B(n4655), .Y(n230) );
  INVX1 U2934 ( .A(n230), .Y(n2985) );
  INVX1 U2935 ( .A(n2988), .Y(n2986) );
  INVX1 U2936 ( .A(n2986), .Y(n2987) );
  AND2X1 U2937 ( .A(n3816), .B(n4655), .Y(n228) );
  INVX1 U2938 ( .A(n228), .Y(n2988) );
  INVX1 U2939 ( .A(n2991), .Y(n2989) );
  INVX1 U2940 ( .A(n2989), .Y(n2990) );
  AND2X1 U2941 ( .A(n3819), .B(n4655), .Y(n226) );
  INVX1 U2942 ( .A(n226), .Y(n2991) );
  INVX1 U2943 ( .A(n2994), .Y(n2992) );
  INVX1 U2944 ( .A(n2992), .Y(n2993) );
  AND2X1 U2945 ( .A(n3822), .B(n4655), .Y(n224) );
  INVX1 U2946 ( .A(n224), .Y(n2994) );
  INVX1 U2947 ( .A(n2997), .Y(n2995) );
  INVX1 U2948 ( .A(n2995), .Y(n2996) );
  AND2X1 U2949 ( .A(n3825), .B(n4655), .Y(n222) );
  INVX1 U2950 ( .A(n222), .Y(n2997) );
  INVX1 U2951 ( .A(n3000), .Y(n2998) );
  INVX1 U2952 ( .A(n2998), .Y(n2999) );
  AND2X1 U2953 ( .A(n3828), .B(n4655), .Y(n220) );
  INVX1 U2954 ( .A(n220), .Y(n3000) );
  INVX1 U2955 ( .A(n3003), .Y(n3001) );
  INVX1 U2956 ( .A(n3001), .Y(n3002) );
  AND2X1 U2957 ( .A(n5315), .B(n175), .Y(n217) );
  INVX1 U2958 ( .A(n217), .Y(n3003) );
  INVX1 U2959 ( .A(n3006), .Y(n3004) );
  INVX1 U2960 ( .A(n3004), .Y(n3005) );
  AND2X1 U2961 ( .A(n92), .B(n175), .Y(n215) );
  INVX1 U2962 ( .A(n215), .Y(n3006) );
  INVX1 U2963 ( .A(n3009), .Y(n3007) );
  INVX1 U2964 ( .A(n3007), .Y(n3008) );
  AND2X1 U2965 ( .A(n38), .B(n201), .Y(n213) );
  INVX1 U2966 ( .A(n213), .Y(n3009) );
  INVX1 U2967 ( .A(n3012), .Y(n3010) );
  INVX1 U2968 ( .A(n3010), .Y(n3011) );
  AND2X1 U2969 ( .A(n33), .B(n201), .Y(n211) );
  INVX1 U2970 ( .A(n211), .Y(n3012) );
  INVX1 U2971 ( .A(n3015), .Y(n3013) );
  INVX1 U2972 ( .A(n3013), .Y(n3014) );
  AND2X1 U2973 ( .A(n34), .B(n201), .Y(n209) );
  INVX1 U2974 ( .A(n209), .Y(n3015) );
  INVX1 U2975 ( .A(n3018), .Y(n3016) );
  INVX1 U2976 ( .A(n3016), .Y(n3017) );
  AND2X1 U2977 ( .A(n35), .B(n201), .Y(n207) );
  INVX1 U2978 ( .A(n207), .Y(n3018) );
  INVX1 U2979 ( .A(n3021), .Y(n3019) );
  INVX1 U2980 ( .A(n3019), .Y(n3020) );
  AND2X1 U2981 ( .A(n36), .B(n201), .Y(n205) );
  INVX1 U2982 ( .A(n205), .Y(n3021) );
  AND2X1 U2983 ( .A(n37), .B(n201), .Y(n203) );
  INVX1 U2984 ( .A(n203), .Y(n3022) );
  AND2X2 U2985 ( .A(we), .B(full_bar), .Y(n201) );
  INVX1 U2986 ( .A(n3025), .Y(n3023) );
  INVX1 U2987 ( .A(n3023), .Y(n3024) );
  AND2X1 U2988 ( .A(n88), .B(n175), .Y(n183) );
  INVX1 U2989 ( .A(n183), .Y(n3025) );
  INVX1 U2990 ( .A(n3028), .Y(n3026) );
  INVX1 U2991 ( .A(n3026), .Y(n3027) );
  AND2X1 U2992 ( .A(n89), .B(n175), .Y(n181) );
  INVX1 U2993 ( .A(n181), .Y(n3028) );
  INVX1 U2994 ( .A(n3031), .Y(n3029) );
  INVX1 U2995 ( .A(n3029), .Y(n3030) );
  AND2X1 U2996 ( .A(n90), .B(n175), .Y(n179) );
  INVX1 U2997 ( .A(n179), .Y(n3031) );
  INVX1 U2998 ( .A(n3034), .Y(n3032) );
  INVX1 U2999 ( .A(n3032), .Y(n3033) );
  AND2X1 U3000 ( .A(n91), .B(n175), .Y(n177) );
  INVX1 U3001 ( .A(n177), .Y(n3034) );
  INVX1 U3002 ( .A(n3037), .Y(n3035) );
  INVX1 U3003 ( .A(n3035), .Y(n3036) );
  OR2X1 U3004 ( .A(fillcount[1]), .B(fillcount[0]), .Y(n796) );
  INVX1 U3005 ( .A(n796), .Y(n3037) );
  INVX1 U3006 ( .A(n3040), .Y(n3038) );
  INVX1 U3007 ( .A(n3038), .Y(n3039) );
  BUFX2 U3008 ( .A(n808), .Y(n3040) );
  INVX1 U3009 ( .A(n3043), .Y(n3041) );
  INVX1 U3010 ( .A(n3041), .Y(n3042) );
  OR2X1 U3011 ( .A(n801), .B(n802), .Y(n800) );
  INVX1 U3012 ( .A(n800), .Y(n3043) );
  INVX1 U3013 ( .A(n3046), .Y(n3044) );
  INVX1 U3014 ( .A(n3044), .Y(n3045) );
  BUFX2 U3015 ( .A(rd_ptr_gray_ss[0]), .Y(n3046) );
  INVX1 U3016 ( .A(n3049), .Y(n3047) );
  INVX1 U3017 ( .A(n3047), .Y(n3048) );
  BUFX2 U3018 ( .A(wr_ptr_gray_ss[2]), .Y(n3049) );
  INVX1 U3019 ( .A(n3052), .Y(n3050) );
  INVX1 U3020 ( .A(n3050), .Y(n3051) );
  BUFX2 U3021 ( .A(rd_ptr_gray_ss[3]), .Y(n3052) );
  INVX1 U3022 ( .A(n3055), .Y(n3053) );
  INVX1 U3023 ( .A(n3053), .Y(n3054) );
  BUFX2 U3024 ( .A(wr_ptr_gray_ss[4]), .Y(n3055) );
  INVX1 U3025 ( .A(n3058), .Y(n3056) );
  INVX1 U3026 ( .A(n3056), .Y(n3057) );
  BUFX2 U3027 ( .A(wr_ptr_gray_ss[3]), .Y(n3058) );
  INVX1 U3028 ( .A(n3061), .Y(n3059) );
  INVX1 U3029 ( .A(n3059), .Y(n3060) );
  BUFX2 U3030 ( .A(wr_ptr_gray_ss[0]), .Y(n3061) );
  INVX1 U3031 ( .A(n3064), .Y(n3062) );
  INVX1 U3032 ( .A(n3062), .Y(n3063) );
  BUFX2 U3033 ( .A(fifo[208]), .Y(n3064) );
  INVX1 U3034 ( .A(n3067), .Y(n3065) );
  INVX1 U3035 ( .A(n3065), .Y(n3066) );
  BUFX2 U3036 ( .A(fifo[209]), .Y(n3067) );
  INVX1 U3037 ( .A(n3070), .Y(n3068) );
  INVX1 U3038 ( .A(n3068), .Y(n3069) );
  BUFX2 U3039 ( .A(fifo[210]), .Y(n3070) );
  INVX1 U3040 ( .A(n3073), .Y(n3071) );
  INVX1 U3041 ( .A(n3071), .Y(n3072) );
  BUFX2 U3042 ( .A(fifo[211]), .Y(n3073) );
  INVX1 U3043 ( .A(n3076), .Y(n3074) );
  INVX1 U3044 ( .A(n3074), .Y(n3075) );
  BUFX2 U3045 ( .A(fifo[212]), .Y(n3076) );
  INVX1 U3046 ( .A(n3079), .Y(n3077) );
  INVX1 U3047 ( .A(n3077), .Y(n3078) );
  BUFX2 U3048 ( .A(fifo[213]), .Y(n3079) );
  INVX1 U3049 ( .A(n3082), .Y(n3080) );
  INVX1 U3050 ( .A(n3080), .Y(n3081) );
  BUFX2 U3051 ( .A(fifo[214]), .Y(n3082) );
  INVX1 U3052 ( .A(n3085), .Y(n3083) );
  INVX1 U3053 ( .A(n3083), .Y(n3084) );
  BUFX2 U3054 ( .A(fifo[215]), .Y(n3085) );
  INVX1 U3055 ( .A(n3088), .Y(n3086) );
  INVX1 U3056 ( .A(n3086), .Y(n3087) );
  BUFX2 U3057 ( .A(fifo[216]), .Y(n3088) );
  INVX1 U3058 ( .A(n3091), .Y(n3089) );
  INVX1 U3059 ( .A(n3089), .Y(n3090) );
  BUFX2 U3060 ( .A(fifo[217]), .Y(n3091) );
  INVX1 U3061 ( .A(n3094), .Y(n3092) );
  INVX1 U3062 ( .A(n3092), .Y(n3093) );
  BUFX2 U3063 ( .A(fifo[218]), .Y(n3094) );
  INVX1 U3064 ( .A(n3097), .Y(n3095) );
  INVX1 U3065 ( .A(n3095), .Y(n3096) );
  BUFX2 U3066 ( .A(fifo[219]), .Y(n3097) );
  INVX1 U3067 ( .A(n3100), .Y(n3098) );
  INVX1 U3068 ( .A(n3098), .Y(n3099) );
  BUFX2 U3069 ( .A(fifo[220]), .Y(n3100) );
  INVX1 U3070 ( .A(n3103), .Y(n3101) );
  INVX1 U3071 ( .A(n3101), .Y(n3102) );
  BUFX2 U3072 ( .A(fifo[221]), .Y(n3103) );
  INVX1 U3073 ( .A(n3106), .Y(n3104) );
  INVX1 U3074 ( .A(n3104), .Y(n3105) );
  BUFX2 U3075 ( .A(fifo[222]), .Y(n3106) );
  INVX1 U3076 ( .A(n3109), .Y(n3107) );
  INVX1 U3077 ( .A(n3107), .Y(n3108) );
  BUFX2 U3078 ( .A(fifo[223]), .Y(n3109) );
  INVX1 U3079 ( .A(n3112), .Y(n3110) );
  INVX1 U3080 ( .A(n3110), .Y(n3111) );
  BUFX2 U3081 ( .A(fifo[176]), .Y(n3112) );
  INVX1 U3082 ( .A(n3115), .Y(n3113) );
  INVX1 U3083 ( .A(n3113), .Y(n3114) );
  BUFX2 U3084 ( .A(fifo[177]), .Y(n3115) );
  INVX1 U3085 ( .A(n3118), .Y(n3116) );
  INVX1 U3086 ( .A(n3116), .Y(n3117) );
  BUFX2 U3087 ( .A(fifo[178]), .Y(n3118) );
  INVX1 U3088 ( .A(n3121), .Y(n3119) );
  INVX1 U3089 ( .A(n3119), .Y(n3120) );
  BUFX2 U3090 ( .A(fifo[179]), .Y(n3121) );
  INVX1 U3091 ( .A(n3124), .Y(n3122) );
  INVX1 U3092 ( .A(n3122), .Y(n3123) );
  BUFX2 U3093 ( .A(fifo[180]), .Y(n3124) );
  INVX1 U3094 ( .A(n3127), .Y(n3125) );
  INVX1 U3095 ( .A(n3125), .Y(n3126) );
  BUFX2 U3096 ( .A(fifo[181]), .Y(n3127) );
  INVX1 U3097 ( .A(n3130), .Y(n3128) );
  INVX1 U3098 ( .A(n3128), .Y(n3129) );
  BUFX2 U3099 ( .A(fifo[182]), .Y(n3130) );
  INVX1 U3100 ( .A(n3133), .Y(n3131) );
  INVX1 U3101 ( .A(n3131), .Y(n3132) );
  BUFX2 U3102 ( .A(fifo[183]), .Y(n3133) );
  INVX1 U3103 ( .A(n3136), .Y(n3134) );
  INVX1 U3104 ( .A(n3134), .Y(n3135) );
  BUFX2 U3105 ( .A(fifo[184]), .Y(n3136) );
  INVX1 U3106 ( .A(n3139), .Y(n3137) );
  INVX1 U3107 ( .A(n3137), .Y(n3138) );
  BUFX2 U3108 ( .A(fifo[185]), .Y(n3139) );
  INVX1 U3109 ( .A(n3142), .Y(n3140) );
  INVX1 U3110 ( .A(n3140), .Y(n3141) );
  BUFX2 U3111 ( .A(fifo[186]), .Y(n3142) );
  INVX1 U3112 ( .A(n3145), .Y(n3143) );
  INVX1 U3113 ( .A(n3143), .Y(n3144) );
  BUFX2 U3114 ( .A(fifo[187]), .Y(n3145) );
  INVX1 U3115 ( .A(n3148), .Y(n3146) );
  INVX1 U3116 ( .A(n3146), .Y(n3147) );
  BUFX2 U3117 ( .A(fifo[188]), .Y(n3148) );
  INVX1 U3118 ( .A(n3151), .Y(n3149) );
  INVX1 U3119 ( .A(n3149), .Y(n3150) );
  BUFX2 U3120 ( .A(fifo[189]), .Y(n3151) );
  INVX1 U3121 ( .A(n3154), .Y(n3152) );
  INVX1 U3122 ( .A(n3152), .Y(n3153) );
  BUFX2 U3123 ( .A(fifo[190]), .Y(n3154) );
  INVX1 U3124 ( .A(n3157), .Y(n3155) );
  INVX1 U3125 ( .A(n3155), .Y(n3156) );
  BUFX2 U3126 ( .A(fifo[191]), .Y(n3157) );
  INVX1 U3127 ( .A(n3160), .Y(n3158) );
  INVX1 U3128 ( .A(n3158), .Y(n3159) );
  BUFX2 U3129 ( .A(fifo[336]), .Y(n3160) );
  INVX1 U3130 ( .A(n3163), .Y(n3161) );
  INVX1 U3131 ( .A(n3161), .Y(n3162) );
  BUFX2 U3132 ( .A(fifo[337]), .Y(n3163) );
  INVX1 U3133 ( .A(n3166), .Y(n3164) );
  INVX1 U3134 ( .A(n3164), .Y(n3165) );
  BUFX2 U3135 ( .A(fifo[338]), .Y(n3166) );
  INVX1 U3136 ( .A(n3169), .Y(n3167) );
  INVX1 U3137 ( .A(n3167), .Y(n3168) );
  BUFX2 U3138 ( .A(fifo[339]), .Y(n3169) );
  INVX1 U3139 ( .A(n3172), .Y(n3170) );
  INVX1 U3140 ( .A(n3170), .Y(n3171) );
  BUFX2 U3141 ( .A(fifo[340]), .Y(n3172) );
  INVX1 U3142 ( .A(n3175), .Y(n3173) );
  INVX1 U3143 ( .A(n3173), .Y(n3174) );
  BUFX2 U3144 ( .A(fifo[341]), .Y(n3175) );
  INVX1 U3145 ( .A(n3178), .Y(n3176) );
  INVX1 U3146 ( .A(n3176), .Y(n3177) );
  BUFX2 U3147 ( .A(fifo[342]), .Y(n3178) );
  INVX1 U3148 ( .A(n3181), .Y(n3179) );
  INVX1 U3149 ( .A(n3179), .Y(n3180) );
  BUFX2 U3150 ( .A(fifo[343]), .Y(n3181) );
  INVX1 U3151 ( .A(n3184), .Y(n3182) );
  INVX1 U3152 ( .A(n3182), .Y(n3183) );
  BUFX2 U3153 ( .A(fifo[344]), .Y(n3184) );
  INVX1 U3154 ( .A(n3187), .Y(n3185) );
  INVX1 U3155 ( .A(n3185), .Y(n3186) );
  BUFX2 U3156 ( .A(fifo[345]), .Y(n3187) );
  INVX1 U3157 ( .A(n3190), .Y(n3188) );
  INVX1 U3158 ( .A(n3188), .Y(n3189) );
  BUFX2 U3159 ( .A(fifo[346]), .Y(n3190) );
  INVX1 U3160 ( .A(n3193), .Y(n3191) );
  INVX1 U3161 ( .A(n3191), .Y(n3192) );
  BUFX2 U3162 ( .A(fifo[347]), .Y(n3193) );
  INVX1 U3163 ( .A(n3196), .Y(n3194) );
  INVX1 U3164 ( .A(n3194), .Y(n3195) );
  BUFX2 U3165 ( .A(fifo[348]), .Y(n3196) );
  INVX1 U3166 ( .A(n3199), .Y(n3197) );
  INVX1 U3167 ( .A(n3197), .Y(n3198) );
  BUFX2 U3168 ( .A(fifo[349]), .Y(n3199) );
  INVX1 U3169 ( .A(n3202), .Y(n3200) );
  INVX1 U3170 ( .A(n3200), .Y(n3201) );
  BUFX2 U3171 ( .A(fifo[350]), .Y(n3202) );
  INVX1 U3172 ( .A(n3205), .Y(n3203) );
  INVX1 U3173 ( .A(n3203), .Y(n3204) );
  BUFX2 U3174 ( .A(fifo[351]), .Y(n3205) );
  INVX1 U3175 ( .A(n3208), .Y(n3206) );
  INVX1 U3176 ( .A(n3206), .Y(n3207) );
  BUFX2 U3177 ( .A(fifo[304]), .Y(n3208) );
  INVX1 U3178 ( .A(n3211), .Y(n3209) );
  INVX1 U3179 ( .A(n3209), .Y(n3210) );
  BUFX2 U3180 ( .A(fifo[305]), .Y(n3211) );
  INVX1 U3181 ( .A(n3214), .Y(n3212) );
  INVX1 U3182 ( .A(n3212), .Y(n3213) );
  BUFX2 U3183 ( .A(fifo[306]), .Y(n3214) );
  INVX1 U3184 ( .A(n3217), .Y(n3215) );
  INVX1 U3185 ( .A(n3215), .Y(n3216) );
  BUFX2 U3186 ( .A(fifo[307]), .Y(n3217) );
  INVX1 U3187 ( .A(n3220), .Y(n3218) );
  INVX1 U3188 ( .A(n3218), .Y(n3219) );
  BUFX2 U3189 ( .A(fifo[308]), .Y(n3220) );
  INVX1 U3190 ( .A(n3223), .Y(n3221) );
  INVX1 U3191 ( .A(n3221), .Y(n3222) );
  BUFX2 U3192 ( .A(fifo[309]), .Y(n3223) );
  INVX1 U3193 ( .A(n3226), .Y(n3224) );
  INVX1 U3194 ( .A(n3224), .Y(n3225) );
  BUFX2 U3195 ( .A(fifo[310]), .Y(n3226) );
  INVX1 U3196 ( .A(n3229), .Y(n3227) );
  INVX1 U3197 ( .A(n3227), .Y(n3228) );
  BUFX2 U3198 ( .A(fifo[311]), .Y(n3229) );
  INVX1 U3199 ( .A(n3232), .Y(n3230) );
  INVX1 U3200 ( .A(n3230), .Y(n3231) );
  BUFX2 U3201 ( .A(fifo[312]), .Y(n3232) );
  INVX1 U3202 ( .A(n3235), .Y(n3233) );
  INVX1 U3203 ( .A(n3233), .Y(n3234) );
  BUFX2 U3204 ( .A(fifo[313]), .Y(n3235) );
  INVX1 U3205 ( .A(n3238), .Y(n3236) );
  INVX1 U3206 ( .A(n3236), .Y(n3237) );
  BUFX2 U3207 ( .A(fifo[314]), .Y(n3238) );
  INVX1 U3208 ( .A(n3241), .Y(n3239) );
  INVX1 U3209 ( .A(n3239), .Y(n3240) );
  BUFX2 U3210 ( .A(fifo[315]), .Y(n3241) );
  INVX1 U3211 ( .A(n3244), .Y(n3242) );
  INVX1 U3212 ( .A(n3242), .Y(n3243) );
  BUFX2 U3213 ( .A(fifo[316]), .Y(n3244) );
  INVX1 U3214 ( .A(n3247), .Y(n3245) );
  INVX1 U3215 ( .A(n3245), .Y(n3246) );
  BUFX2 U3216 ( .A(fifo[317]), .Y(n3247) );
  INVX1 U3217 ( .A(n3250), .Y(n3248) );
  INVX1 U3218 ( .A(n3248), .Y(n3249) );
  BUFX2 U3219 ( .A(fifo[318]), .Y(n3250) );
  INVX1 U3220 ( .A(n3253), .Y(n3251) );
  INVX1 U3221 ( .A(n3251), .Y(n3252) );
  BUFX2 U3222 ( .A(fifo[319]), .Y(n3253) );
  INVX1 U3223 ( .A(n3256), .Y(n3254) );
  INVX1 U3224 ( .A(n3254), .Y(n3255) );
  BUFX2 U3225 ( .A(fifo[144]), .Y(n3256) );
  INVX1 U3226 ( .A(n3259), .Y(n3257) );
  INVX1 U3227 ( .A(n3257), .Y(n3258) );
  BUFX2 U3228 ( .A(fifo[145]), .Y(n3259) );
  INVX1 U3229 ( .A(n3262), .Y(n3260) );
  INVX1 U3230 ( .A(n3260), .Y(n3261) );
  BUFX2 U3231 ( .A(fifo[146]), .Y(n3262) );
  INVX1 U3232 ( .A(n3265), .Y(n3263) );
  INVX1 U3233 ( .A(n3263), .Y(n3264) );
  BUFX2 U3234 ( .A(fifo[147]), .Y(n3265) );
  INVX1 U3235 ( .A(n3268), .Y(n3266) );
  INVX1 U3236 ( .A(n3266), .Y(n3267) );
  BUFX2 U3237 ( .A(fifo[148]), .Y(n3268) );
  INVX1 U3238 ( .A(n3271), .Y(n3269) );
  INVX1 U3239 ( .A(n3269), .Y(n3270) );
  BUFX2 U3240 ( .A(fifo[149]), .Y(n3271) );
  INVX1 U3241 ( .A(n3274), .Y(n3272) );
  INVX1 U3242 ( .A(n3272), .Y(n3273) );
  BUFX2 U3243 ( .A(fifo[150]), .Y(n3274) );
  INVX1 U3244 ( .A(n3277), .Y(n3275) );
  INVX1 U3245 ( .A(n3275), .Y(n3276) );
  BUFX2 U3246 ( .A(fifo[151]), .Y(n3277) );
  INVX1 U3247 ( .A(n3280), .Y(n3278) );
  INVX1 U3248 ( .A(n3278), .Y(n3279) );
  BUFX2 U3249 ( .A(fifo[152]), .Y(n3280) );
  INVX1 U3250 ( .A(n3283), .Y(n3281) );
  INVX1 U3251 ( .A(n3281), .Y(n3282) );
  BUFX2 U3252 ( .A(fifo[153]), .Y(n3283) );
  INVX1 U3253 ( .A(n3286), .Y(n3284) );
  INVX1 U3254 ( .A(n3284), .Y(n3285) );
  BUFX2 U3255 ( .A(fifo[154]), .Y(n3286) );
  INVX1 U3256 ( .A(n3289), .Y(n3287) );
  INVX1 U3257 ( .A(n3287), .Y(n3288) );
  BUFX2 U3258 ( .A(fifo[155]), .Y(n3289) );
  INVX1 U3259 ( .A(n3292), .Y(n3290) );
  INVX1 U3260 ( .A(n3290), .Y(n3291) );
  BUFX2 U3261 ( .A(fifo[156]), .Y(n3292) );
  INVX1 U3262 ( .A(n3295), .Y(n3293) );
  INVX1 U3263 ( .A(n3293), .Y(n3294) );
  BUFX2 U3264 ( .A(fifo[157]), .Y(n3295) );
  INVX1 U3265 ( .A(n3298), .Y(n3296) );
  INVX1 U3266 ( .A(n3296), .Y(n3297) );
  BUFX2 U3267 ( .A(fifo[158]), .Y(n3298) );
  INVX1 U3268 ( .A(n3301), .Y(n3299) );
  INVX1 U3269 ( .A(n3299), .Y(n3300) );
  BUFX2 U3270 ( .A(fifo[159]), .Y(n3301) );
  INVX1 U3271 ( .A(n3304), .Y(n3302) );
  INVX1 U3272 ( .A(n3302), .Y(n3303) );
  BUFX2 U3273 ( .A(fifo[272]), .Y(n3304) );
  INVX1 U3274 ( .A(n3307), .Y(n3305) );
  INVX1 U3275 ( .A(n3305), .Y(n3306) );
  BUFX2 U3276 ( .A(fifo[273]), .Y(n3307) );
  INVX1 U3277 ( .A(n3310), .Y(n3308) );
  INVX1 U3278 ( .A(n3308), .Y(n3309) );
  BUFX2 U3279 ( .A(fifo[274]), .Y(n3310) );
  INVX1 U3280 ( .A(n3313), .Y(n3311) );
  INVX1 U3281 ( .A(n3311), .Y(n3312) );
  BUFX2 U3282 ( .A(fifo[275]), .Y(n3313) );
  INVX1 U3283 ( .A(n3316), .Y(n3314) );
  INVX1 U3284 ( .A(n3314), .Y(n3315) );
  BUFX2 U3285 ( .A(fifo[276]), .Y(n3316) );
  INVX1 U3286 ( .A(n3319), .Y(n3317) );
  INVX1 U3287 ( .A(n3317), .Y(n3318) );
  BUFX2 U3288 ( .A(fifo[277]), .Y(n3319) );
  INVX1 U3289 ( .A(n3322), .Y(n3320) );
  INVX1 U3290 ( .A(n3320), .Y(n3321) );
  BUFX2 U3291 ( .A(fifo[278]), .Y(n3322) );
  INVX1 U3292 ( .A(n3325), .Y(n3323) );
  INVX1 U3293 ( .A(n3323), .Y(n3324) );
  BUFX2 U3294 ( .A(fifo[279]), .Y(n3325) );
  INVX1 U3295 ( .A(n3328), .Y(n3326) );
  INVX1 U3296 ( .A(n3326), .Y(n3327) );
  BUFX2 U3297 ( .A(fifo[280]), .Y(n3328) );
  INVX1 U3298 ( .A(n3331), .Y(n3329) );
  INVX1 U3299 ( .A(n3329), .Y(n3330) );
  BUFX2 U3300 ( .A(fifo[281]), .Y(n3331) );
  INVX1 U3301 ( .A(n3334), .Y(n3332) );
  INVX1 U3302 ( .A(n3332), .Y(n3333) );
  BUFX2 U3303 ( .A(fifo[282]), .Y(n3334) );
  INVX1 U3304 ( .A(n3337), .Y(n3335) );
  INVX1 U3305 ( .A(n3335), .Y(n3336) );
  BUFX2 U3306 ( .A(fifo[283]), .Y(n3337) );
  INVX1 U3307 ( .A(n3340), .Y(n3338) );
  INVX1 U3308 ( .A(n3338), .Y(n3339) );
  BUFX2 U3309 ( .A(fifo[284]), .Y(n3340) );
  INVX1 U3310 ( .A(n3343), .Y(n3341) );
  INVX1 U3311 ( .A(n3341), .Y(n3342) );
  BUFX2 U3312 ( .A(fifo[285]), .Y(n3343) );
  INVX1 U3313 ( .A(n3346), .Y(n3344) );
  INVX1 U3314 ( .A(n3344), .Y(n3345) );
  BUFX2 U3315 ( .A(fifo[286]), .Y(n3346) );
  INVX1 U3316 ( .A(n3349), .Y(n3347) );
  INVX1 U3317 ( .A(n3347), .Y(n3348) );
  BUFX2 U3318 ( .A(fifo[287]), .Y(n3349) );
  INVX1 U3319 ( .A(n3352), .Y(n3350) );
  INVX1 U3320 ( .A(n3350), .Y(n3351) );
  BUFX2 U3321 ( .A(fifo[240]), .Y(n3352) );
  INVX1 U3322 ( .A(n3355), .Y(n3353) );
  INVX1 U3323 ( .A(n3353), .Y(n3354) );
  BUFX2 U3324 ( .A(fifo[241]), .Y(n3355) );
  INVX1 U3325 ( .A(n3358), .Y(n3356) );
  INVX1 U3326 ( .A(n3356), .Y(n3357) );
  BUFX2 U3327 ( .A(fifo[242]), .Y(n3358) );
  INVX1 U3328 ( .A(n3361), .Y(n3359) );
  INVX1 U3329 ( .A(n3359), .Y(n3360) );
  BUFX2 U3330 ( .A(fifo[243]), .Y(n3361) );
  INVX1 U3331 ( .A(n3364), .Y(n3362) );
  INVX1 U3332 ( .A(n3362), .Y(n3363) );
  BUFX2 U3333 ( .A(fifo[244]), .Y(n3364) );
  INVX1 U3334 ( .A(n3367), .Y(n3365) );
  INVX1 U3335 ( .A(n3365), .Y(n3366) );
  BUFX2 U3336 ( .A(fifo[245]), .Y(n3367) );
  INVX1 U3337 ( .A(n3370), .Y(n3368) );
  INVX1 U3338 ( .A(n3368), .Y(n3369) );
  BUFX2 U3339 ( .A(fifo[246]), .Y(n3370) );
  INVX1 U3340 ( .A(n3373), .Y(n3371) );
  INVX1 U3341 ( .A(n3371), .Y(n3372) );
  BUFX2 U3342 ( .A(fifo[247]), .Y(n3373) );
  INVX1 U3343 ( .A(n3376), .Y(n3374) );
  INVX1 U3344 ( .A(n3374), .Y(n3375) );
  BUFX2 U3345 ( .A(fifo[248]), .Y(n3376) );
  INVX1 U3346 ( .A(n3379), .Y(n3377) );
  INVX1 U3347 ( .A(n3377), .Y(n3378) );
  BUFX2 U3348 ( .A(fifo[249]), .Y(n3379) );
  INVX1 U3349 ( .A(n3382), .Y(n3380) );
  INVX1 U3350 ( .A(n3380), .Y(n3381) );
  BUFX2 U3351 ( .A(fifo[250]), .Y(n3382) );
  INVX1 U3352 ( .A(n3385), .Y(n3383) );
  INVX1 U3353 ( .A(n3383), .Y(n3384) );
  BUFX2 U3354 ( .A(fifo[251]), .Y(n3385) );
  INVX1 U3355 ( .A(n3388), .Y(n3386) );
  INVX1 U3356 ( .A(n3386), .Y(n3387) );
  BUFX2 U3357 ( .A(fifo[252]), .Y(n3388) );
  INVX1 U3358 ( .A(n3391), .Y(n3389) );
  INVX1 U3359 ( .A(n3389), .Y(n3390) );
  BUFX2 U3360 ( .A(fifo[253]), .Y(n3391) );
  INVX1 U3361 ( .A(n3394), .Y(n3392) );
  INVX1 U3362 ( .A(n3392), .Y(n3393) );
  BUFX2 U3363 ( .A(fifo[254]), .Y(n3394) );
  INVX1 U3364 ( .A(n3397), .Y(n3395) );
  INVX1 U3365 ( .A(n3395), .Y(n3396) );
  BUFX2 U3366 ( .A(fifo[255]), .Y(n3397) );
  INVX1 U3367 ( .A(n3400), .Y(n3398) );
  INVX1 U3368 ( .A(n3398), .Y(n3399) );
  BUFX2 U3369 ( .A(fifo[368]), .Y(n3400) );
  INVX1 U3370 ( .A(n3403), .Y(n3401) );
  INVX1 U3371 ( .A(n3401), .Y(n3402) );
  BUFX2 U3372 ( .A(fifo[369]), .Y(n3403) );
  INVX1 U3373 ( .A(n3406), .Y(n3404) );
  INVX1 U3374 ( .A(n3404), .Y(n3405) );
  BUFX2 U3375 ( .A(fifo[370]), .Y(n3406) );
  INVX1 U3376 ( .A(n3409), .Y(n3407) );
  INVX1 U3377 ( .A(n3407), .Y(n3408) );
  BUFX2 U3378 ( .A(fifo[371]), .Y(n3409) );
  INVX1 U3379 ( .A(n3412), .Y(n3410) );
  INVX1 U3380 ( .A(n3410), .Y(n3411) );
  BUFX2 U3381 ( .A(fifo[372]), .Y(n3412) );
  INVX1 U3382 ( .A(n3415), .Y(n3413) );
  INVX1 U3383 ( .A(n3413), .Y(n3414) );
  BUFX2 U3384 ( .A(fifo[373]), .Y(n3415) );
  INVX1 U3385 ( .A(n3418), .Y(n3416) );
  INVX1 U3386 ( .A(n3416), .Y(n3417) );
  BUFX2 U3387 ( .A(fifo[374]), .Y(n3418) );
  INVX1 U3388 ( .A(n3421), .Y(n3419) );
  INVX1 U3389 ( .A(n3419), .Y(n3420) );
  BUFX2 U3390 ( .A(fifo[375]), .Y(n3421) );
  INVX1 U3391 ( .A(n3424), .Y(n3422) );
  INVX1 U3392 ( .A(n3422), .Y(n3423) );
  BUFX2 U3393 ( .A(fifo[376]), .Y(n3424) );
  INVX1 U3394 ( .A(n3427), .Y(n3425) );
  INVX1 U3395 ( .A(n3425), .Y(n3426) );
  BUFX2 U3396 ( .A(fifo[377]), .Y(n3427) );
  INVX1 U3397 ( .A(n3430), .Y(n3428) );
  INVX1 U3398 ( .A(n3428), .Y(n3429) );
  BUFX2 U3399 ( .A(fifo[378]), .Y(n3430) );
  INVX1 U3400 ( .A(n3433), .Y(n3431) );
  INVX1 U3401 ( .A(n3431), .Y(n3432) );
  BUFX2 U3402 ( .A(fifo[379]), .Y(n3433) );
  INVX1 U3403 ( .A(n3436), .Y(n3434) );
  INVX1 U3404 ( .A(n3434), .Y(n3435) );
  BUFX2 U3405 ( .A(fifo[380]), .Y(n3436) );
  INVX1 U3406 ( .A(n3439), .Y(n3437) );
  INVX1 U3407 ( .A(n3437), .Y(n3438) );
  BUFX2 U3408 ( .A(fifo[381]), .Y(n3439) );
  INVX1 U3409 ( .A(n3442), .Y(n3440) );
  INVX1 U3410 ( .A(n3440), .Y(n3441) );
  BUFX2 U3411 ( .A(fifo[382]), .Y(n3442) );
  INVX1 U3412 ( .A(n3445), .Y(n3443) );
  INVX1 U3413 ( .A(n3443), .Y(n3444) );
  BUFX2 U3414 ( .A(fifo[383]), .Y(n3445) );
  INVX1 U3415 ( .A(n3448), .Y(n3446) );
  INVX1 U3416 ( .A(n3446), .Y(n3447) );
  BUFX2 U3417 ( .A(fifo[80]), .Y(n3448) );
  INVX1 U3418 ( .A(n3451), .Y(n3449) );
  INVX1 U3419 ( .A(n3449), .Y(n3450) );
  BUFX2 U3420 ( .A(fifo[81]), .Y(n3451) );
  INVX1 U3421 ( .A(n3454), .Y(n3452) );
  INVX1 U3422 ( .A(n3452), .Y(n3453) );
  BUFX2 U3423 ( .A(fifo[82]), .Y(n3454) );
  INVX1 U3424 ( .A(n3457), .Y(n3455) );
  INVX1 U3425 ( .A(n3455), .Y(n3456) );
  BUFX2 U3426 ( .A(fifo[83]), .Y(n3457) );
  INVX1 U3427 ( .A(n3460), .Y(n3458) );
  INVX1 U3428 ( .A(n3458), .Y(n3459) );
  BUFX2 U3429 ( .A(fifo[84]), .Y(n3460) );
  INVX1 U3430 ( .A(n3463), .Y(n3461) );
  INVX1 U3431 ( .A(n3461), .Y(n3462) );
  BUFX2 U3432 ( .A(fifo[85]), .Y(n3463) );
  INVX1 U3433 ( .A(n3466), .Y(n3464) );
  INVX1 U3434 ( .A(n3464), .Y(n3465) );
  BUFX2 U3435 ( .A(fifo[86]), .Y(n3466) );
  INVX1 U3436 ( .A(n3469), .Y(n3467) );
  INVX1 U3437 ( .A(n3467), .Y(n3468) );
  BUFX2 U3438 ( .A(fifo[87]), .Y(n3469) );
  INVX1 U3439 ( .A(n3472), .Y(n3470) );
  INVX1 U3440 ( .A(n3470), .Y(n3471) );
  BUFX2 U3441 ( .A(fifo[88]), .Y(n3472) );
  INVX1 U3442 ( .A(n3475), .Y(n3473) );
  INVX1 U3443 ( .A(n3473), .Y(n3474) );
  BUFX2 U3444 ( .A(fifo[89]), .Y(n3475) );
  INVX1 U3445 ( .A(n3478), .Y(n3476) );
  INVX1 U3446 ( .A(n3476), .Y(n3477) );
  BUFX2 U3447 ( .A(fifo[90]), .Y(n3478) );
  INVX1 U3448 ( .A(n3481), .Y(n3479) );
  INVX1 U3449 ( .A(n3479), .Y(n3480) );
  BUFX2 U3450 ( .A(fifo[91]), .Y(n3481) );
  INVX1 U3451 ( .A(n3484), .Y(n3482) );
  INVX1 U3452 ( .A(n3482), .Y(n3483) );
  BUFX2 U3453 ( .A(fifo[92]), .Y(n3484) );
  INVX1 U3454 ( .A(n3487), .Y(n3485) );
  INVX1 U3455 ( .A(n3485), .Y(n3486) );
  BUFX2 U3456 ( .A(fifo[93]), .Y(n3487) );
  INVX1 U3457 ( .A(n3490), .Y(n3488) );
  INVX1 U3458 ( .A(n3488), .Y(n3489) );
  BUFX2 U3459 ( .A(fifo[94]), .Y(n3490) );
  INVX1 U3460 ( .A(n3493), .Y(n3491) );
  INVX1 U3461 ( .A(n3491), .Y(n3492) );
  BUFX2 U3462 ( .A(fifo[95]), .Y(n3493) );
  INVX1 U3463 ( .A(n3496), .Y(n3494) );
  INVX1 U3464 ( .A(n3494), .Y(n3495) );
  BUFX2 U3465 ( .A(fifo[48]), .Y(n3496) );
  INVX1 U3466 ( .A(n3499), .Y(n3497) );
  INVX1 U3467 ( .A(n3497), .Y(n3498) );
  BUFX2 U3468 ( .A(fifo[49]), .Y(n3499) );
  INVX1 U3469 ( .A(n3502), .Y(n3500) );
  INVX1 U3470 ( .A(n3500), .Y(n3501) );
  BUFX2 U3471 ( .A(fifo[50]), .Y(n3502) );
  INVX1 U3472 ( .A(n3505), .Y(n3503) );
  INVX1 U3473 ( .A(n3503), .Y(n3504) );
  BUFX2 U3474 ( .A(fifo[51]), .Y(n3505) );
  INVX1 U3475 ( .A(n3508), .Y(n3506) );
  INVX1 U3476 ( .A(n3506), .Y(n3507) );
  BUFX2 U3477 ( .A(fifo[52]), .Y(n3508) );
  INVX1 U3478 ( .A(n3511), .Y(n3509) );
  INVX1 U3479 ( .A(n3509), .Y(n3510) );
  BUFX2 U3480 ( .A(fifo[53]), .Y(n3511) );
  INVX1 U3481 ( .A(n3514), .Y(n3512) );
  INVX1 U3482 ( .A(n3512), .Y(n3513) );
  BUFX2 U3483 ( .A(fifo[54]), .Y(n3514) );
  INVX1 U3484 ( .A(n3517), .Y(n3515) );
  INVX1 U3485 ( .A(n3515), .Y(n3516) );
  BUFX2 U3486 ( .A(fifo[55]), .Y(n3517) );
  INVX1 U3487 ( .A(n3520), .Y(n3518) );
  INVX1 U3488 ( .A(n3518), .Y(n3519) );
  BUFX2 U3489 ( .A(fifo[56]), .Y(n3520) );
  INVX1 U3490 ( .A(n3523), .Y(n3521) );
  INVX1 U3491 ( .A(n3521), .Y(n3522) );
  BUFX2 U3492 ( .A(fifo[57]), .Y(n3523) );
  INVX1 U3493 ( .A(n3526), .Y(n3524) );
  INVX1 U3494 ( .A(n3524), .Y(n3525) );
  BUFX2 U3495 ( .A(fifo[58]), .Y(n3526) );
  INVX1 U3496 ( .A(n3529), .Y(n3527) );
  INVX1 U3497 ( .A(n3527), .Y(n3528) );
  BUFX2 U3498 ( .A(fifo[59]), .Y(n3529) );
  INVX1 U3499 ( .A(n3532), .Y(n3530) );
  INVX1 U3500 ( .A(n3530), .Y(n3531) );
  BUFX2 U3501 ( .A(fifo[60]), .Y(n3532) );
  INVX1 U3502 ( .A(n3535), .Y(n3533) );
  INVX1 U3503 ( .A(n3533), .Y(n3534) );
  BUFX2 U3504 ( .A(fifo[61]), .Y(n3535) );
  INVX1 U3505 ( .A(n3538), .Y(n3536) );
  INVX1 U3506 ( .A(n3536), .Y(n3537) );
  BUFX2 U3507 ( .A(fifo[62]), .Y(n3538) );
  INVX1 U3508 ( .A(n3541), .Y(n3539) );
  INVX1 U3509 ( .A(n3539), .Y(n3540) );
  BUFX2 U3510 ( .A(fifo[63]), .Y(n3541) );
  INVX1 U3511 ( .A(n3544), .Y(n3542) );
  INVX1 U3512 ( .A(n3542), .Y(n3543) );
  BUFX2 U3513 ( .A(fifo[16]), .Y(n3544) );
  INVX1 U3514 ( .A(n3547), .Y(n3545) );
  INVX1 U3515 ( .A(n3545), .Y(n3546) );
  BUFX2 U3516 ( .A(fifo[17]), .Y(n3547) );
  INVX1 U3517 ( .A(n3550), .Y(n3548) );
  INVX1 U3518 ( .A(n3548), .Y(n3549) );
  BUFX2 U3519 ( .A(fifo[18]), .Y(n3550) );
  INVX1 U3520 ( .A(n3553), .Y(n3551) );
  INVX1 U3521 ( .A(n3551), .Y(n3552) );
  BUFX2 U3522 ( .A(fifo[19]), .Y(n3553) );
  INVX1 U3523 ( .A(n3556), .Y(n3554) );
  INVX1 U3524 ( .A(n3554), .Y(n3555) );
  BUFX2 U3525 ( .A(fifo[20]), .Y(n3556) );
  INVX1 U3526 ( .A(n3559), .Y(n3557) );
  INVX1 U3527 ( .A(n3557), .Y(n3558) );
  BUFX2 U3528 ( .A(fifo[21]), .Y(n3559) );
  INVX1 U3529 ( .A(n3562), .Y(n3560) );
  INVX1 U3530 ( .A(n3560), .Y(n3561) );
  BUFX2 U3531 ( .A(fifo[22]), .Y(n3562) );
  INVX1 U3532 ( .A(n3565), .Y(n3563) );
  INVX1 U3533 ( .A(n3563), .Y(n3564) );
  BUFX2 U3534 ( .A(fifo[23]), .Y(n3565) );
  INVX1 U3535 ( .A(n3568), .Y(n3566) );
  INVX1 U3536 ( .A(n3566), .Y(n3567) );
  BUFX2 U3537 ( .A(fifo[24]), .Y(n3568) );
  INVX1 U3538 ( .A(n3571), .Y(n3569) );
  INVX1 U3539 ( .A(n3569), .Y(n3570) );
  BUFX2 U3540 ( .A(fifo[25]), .Y(n3571) );
  INVX1 U3541 ( .A(n3574), .Y(n3572) );
  INVX1 U3542 ( .A(n3572), .Y(n3573) );
  BUFX2 U3543 ( .A(fifo[26]), .Y(n3574) );
  INVX1 U3544 ( .A(n3577), .Y(n3575) );
  INVX1 U3545 ( .A(n3575), .Y(n3576) );
  BUFX2 U3546 ( .A(fifo[27]), .Y(n3577) );
  INVX1 U3547 ( .A(n3580), .Y(n3578) );
  INVX1 U3548 ( .A(n3578), .Y(n3579) );
  BUFX2 U3549 ( .A(fifo[28]), .Y(n3580) );
  INVX1 U3550 ( .A(n3583), .Y(n3581) );
  INVX1 U3551 ( .A(n3581), .Y(n3582) );
  BUFX2 U3552 ( .A(fifo[29]), .Y(n3583) );
  INVX1 U3553 ( .A(n3586), .Y(n3584) );
  INVX1 U3554 ( .A(n3584), .Y(n3585) );
  BUFX2 U3555 ( .A(fifo[30]), .Y(n3586) );
  INVX1 U3556 ( .A(n3589), .Y(n3587) );
  INVX1 U3557 ( .A(n3587), .Y(n3588) );
  BUFX2 U3558 ( .A(fifo[31]), .Y(n3589) );
  INVX1 U3559 ( .A(n3592), .Y(n3590) );
  INVX1 U3560 ( .A(n3590), .Y(n3591) );
  BUFX2 U3561 ( .A(fifo[112]), .Y(n3592) );
  INVX1 U3562 ( .A(n3595), .Y(n3593) );
  INVX1 U3563 ( .A(n3593), .Y(n3594) );
  BUFX2 U3564 ( .A(fifo[113]), .Y(n3595) );
  INVX1 U3565 ( .A(n3598), .Y(n3596) );
  INVX1 U3566 ( .A(n3596), .Y(n3597) );
  BUFX2 U3567 ( .A(fifo[114]), .Y(n3598) );
  INVX1 U3568 ( .A(n3601), .Y(n3599) );
  INVX1 U3569 ( .A(n3599), .Y(n3600) );
  BUFX2 U3570 ( .A(fifo[115]), .Y(n3601) );
  INVX1 U3571 ( .A(n3604), .Y(n3602) );
  INVX1 U3572 ( .A(n3602), .Y(n3603) );
  BUFX2 U3573 ( .A(fifo[116]), .Y(n3604) );
  INVX1 U3574 ( .A(n3607), .Y(n3605) );
  INVX1 U3575 ( .A(n3605), .Y(n3606) );
  BUFX2 U3576 ( .A(fifo[117]), .Y(n3607) );
  INVX1 U3577 ( .A(n3610), .Y(n3608) );
  INVX1 U3578 ( .A(n3608), .Y(n3609) );
  BUFX2 U3579 ( .A(fifo[118]), .Y(n3610) );
  INVX1 U3580 ( .A(n3613), .Y(n3611) );
  INVX1 U3581 ( .A(n3611), .Y(n3612) );
  BUFX2 U3582 ( .A(fifo[119]), .Y(n3613) );
  INVX1 U3583 ( .A(n3616), .Y(n3614) );
  INVX1 U3584 ( .A(n3614), .Y(n3615) );
  BUFX2 U3585 ( .A(fifo[120]), .Y(n3616) );
  INVX1 U3586 ( .A(n3619), .Y(n3617) );
  INVX1 U3587 ( .A(n3617), .Y(n3618) );
  BUFX2 U3588 ( .A(fifo[121]), .Y(n3619) );
  INVX1 U3589 ( .A(n3622), .Y(n3620) );
  INVX1 U3590 ( .A(n3620), .Y(n3621) );
  BUFX2 U3591 ( .A(fifo[122]), .Y(n3622) );
  INVX1 U3592 ( .A(n3625), .Y(n3623) );
  INVX1 U3593 ( .A(n3623), .Y(n3624) );
  BUFX2 U3594 ( .A(fifo[123]), .Y(n3625) );
  INVX1 U3595 ( .A(n3628), .Y(n3626) );
  INVX1 U3596 ( .A(n3626), .Y(n3627) );
  BUFX2 U3597 ( .A(fifo[124]), .Y(n3628) );
  INVX1 U3598 ( .A(n3631), .Y(n3629) );
  INVX1 U3599 ( .A(n3629), .Y(n3630) );
  BUFX2 U3600 ( .A(fifo[125]), .Y(n3631) );
  INVX1 U3601 ( .A(n3634), .Y(n3632) );
  INVX1 U3602 ( .A(n3632), .Y(n3633) );
  BUFX2 U3603 ( .A(fifo[126]), .Y(n3634) );
  INVX1 U3604 ( .A(n3637), .Y(n3635) );
  INVX1 U3605 ( .A(n3635), .Y(n3636) );
  BUFX2 U3606 ( .A(fifo[127]), .Y(n3637) );
  INVX1 U3607 ( .A(n3640), .Y(n3638) );
  INVX1 U3608 ( .A(n3638), .Y(n3639) );
  BUFX2 U3609 ( .A(fifo[464]), .Y(n3640) );
  INVX1 U3610 ( .A(n3643), .Y(n3641) );
  INVX1 U3611 ( .A(n3641), .Y(n3642) );
  BUFX2 U3612 ( .A(fifo[465]), .Y(n3643) );
  INVX1 U3613 ( .A(n3646), .Y(n3644) );
  INVX1 U3614 ( .A(n3644), .Y(n3645) );
  BUFX2 U3615 ( .A(fifo[466]), .Y(n3646) );
  INVX1 U3616 ( .A(n3649), .Y(n3647) );
  INVX1 U3617 ( .A(n3647), .Y(n3648) );
  BUFX2 U3618 ( .A(fifo[467]), .Y(n3649) );
  INVX1 U3619 ( .A(n3652), .Y(n3650) );
  INVX1 U3620 ( .A(n3650), .Y(n3651) );
  BUFX2 U3621 ( .A(fifo[468]), .Y(n3652) );
  INVX1 U3622 ( .A(n3655), .Y(n3653) );
  INVX1 U3623 ( .A(n3653), .Y(n3654) );
  BUFX2 U3624 ( .A(fifo[469]), .Y(n3655) );
  INVX1 U3625 ( .A(n3658), .Y(n3656) );
  INVX1 U3626 ( .A(n3656), .Y(n3657) );
  BUFX2 U3627 ( .A(fifo[470]), .Y(n3658) );
  INVX1 U3628 ( .A(n3661), .Y(n3659) );
  INVX1 U3629 ( .A(n3659), .Y(n3660) );
  BUFX2 U3630 ( .A(fifo[471]), .Y(n3661) );
  INVX1 U3631 ( .A(n3664), .Y(n3662) );
  INVX1 U3632 ( .A(n3662), .Y(n3663) );
  BUFX2 U3633 ( .A(fifo[472]), .Y(n3664) );
  INVX1 U3634 ( .A(n3667), .Y(n3665) );
  INVX1 U3635 ( .A(n3665), .Y(n3666) );
  BUFX2 U3636 ( .A(fifo[473]), .Y(n3667) );
  INVX1 U3637 ( .A(n3670), .Y(n3668) );
  INVX1 U3638 ( .A(n3668), .Y(n3669) );
  BUFX2 U3639 ( .A(fifo[474]), .Y(n3670) );
  INVX1 U3640 ( .A(n3673), .Y(n3671) );
  INVX1 U3641 ( .A(n3671), .Y(n3672) );
  BUFX2 U3642 ( .A(fifo[475]), .Y(n3673) );
  INVX1 U3643 ( .A(n3676), .Y(n3674) );
  INVX1 U3644 ( .A(n3674), .Y(n3675) );
  BUFX2 U3645 ( .A(fifo[476]), .Y(n3676) );
  INVX1 U3646 ( .A(n3679), .Y(n3677) );
  INVX1 U3647 ( .A(n3677), .Y(n3678) );
  BUFX2 U3648 ( .A(fifo[477]), .Y(n3679) );
  INVX1 U3649 ( .A(n3682), .Y(n3680) );
  INVX1 U3650 ( .A(n3680), .Y(n3681) );
  BUFX2 U3651 ( .A(fifo[478]), .Y(n3682) );
  INVX1 U3652 ( .A(n3685), .Y(n3683) );
  INVX1 U3653 ( .A(n3683), .Y(n3684) );
  BUFX2 U3654 ( .A(fifo[479]), .Y(n3685) );
  INVX1 U3655 ( .A(n3688), .Y(n3686) );
  INVX1 U3656 ( .A(n3686), .Y(n3687) );
  BUFX2 U3657 ( .A(fifo[432]), .Y(n3688) );
  INVX1 U3658 ( .A(n3691), .Y(n3689) );
  INVX1 U3659 ( .A(n3689), .Y(n3690) );
  BUFX2 U3660 ( .A(fifo[433]), .Y(n3691) );
  INVX1 U3661 ( .A(n3694), .Y(n3692) );
  INVX1 U3662 ( .A(n3692), .Y(n3693) );
  BUFX2 U3663 ( .A(fifo[434]), .Y(n3694) );
  INVX1 U3664 ( .A(n3697), .Y(n3695) );
  INVX1 U3665 ( .A(n3695), .Y(n3696) );
  BUFX2 U3666 ( .A(fifo[435]), .Y(n3697) );
  INVX1 U3667 ( .A(n3700), .Y(n3698) );
  INVX1 U3668 ( .A(n3698), .Y(n3699) );
  BUFX2 U3669 ( .A(fifo[436]), .Y(n3700) );
  INVX1 U3670 ( .A(n3703), .Y(n3701) );
  INVX1 U3671 ( .A(n3701), .Y(n3702) );
  BUFX2 U3672 ( .A(fifo[437]), .Y(n3703) );
  INVX1 U3673 ( .A(n3706), .Y(n3704) );
  INVX1 U3674 ( .A(n3704), .Y(n3705) );
  BUFX2 U3675 ( .A(fifo[438]), .Y(n3706) );
  INVX1 U3676 ( .A(n3709), .Y(n3707) );
  INVX1 U3677 ( .A(n3707), .Y(n3708) );
  BUFX2 U3678 ( .A(fifo[439]), .Y(n3709) );
  INVX1 U3679 ( .A(n3712), .Y(n3710) );
  INVX1 U3680 ( .A(n3710), .Y(n3711) );
  BUFX2 U3681 ( .A(fifo[440]), .Y(n3712) );
  INVX1 U3682 ( .A(n3715), .Y(n3713) );
  INVX1 U3683 ( .A(n3713), .Y(n3714) );
  BUFX2 U3684 ( .A(fifo[441]), .Y(n3715) );
  INVX1 U3685 ( .A(n3718), .Y(n3716) );
  INVX1 U3686 ( .A(n3716), .Y(n3717) );
  BUFX2 U3687 ( .A(fifo[442]), .Y(n3718) );
  INVX1 U3688 ( .A(n3721), .Y(n3719) );
  INVX1 U3689 ( .A(n3719), .Y(n3720) );
  BUFX2 U3690 ( .A(fifo[443]), .Y(n3721) );
  INVX1 U3691 ( .A(n3724), .Y(n3722) );
  INVX1 U3692 ( .A(n3722), .Y(n3723) );
  BUFX2 U3693 ( .A(fifo[444]), .Y(n3724) );
  INVX1 U3694 ( .A(n3727), .Y(n3725) );
  INVX1 U3695 ( .A(n3725), .Y(n3726) );
  BUFX2 U3696 ( .A(fifo[445]), .Y(n3727) );
  INVX1 U3697 ( .A(n3730), .Y(n3728) );
  INVX1 U3698 ( .A(n3728), .Y(n3729) );
  BUFX2 U3699 ( .A(fifo[446]), .Y(n3730) );
  INVX1 U3700 ( .A(n3733), .Y(n3731) );
  INVX1 U3701 ( .A(n3731), .Y(n3732) );
  BUFX2 U3702 ( .A(fifo[447]), .Y(n3733) );
  INVX1 U3703 ( .A(n3736), .Y(n3734) );
  INVX1 U3704 ( .A(n3734), .Y(n3735) );
  BUFX2 U3705 ( .A(fifo[400]), .Y(n3736) );
  INVX1 U3706 ( .A(n3739), .Y(n3737) );
  INVX1 U3707 ( .A(n3737), .Y(n3738) );
  BUFX2 U3708 ( .A(fifo[401]), .Y(n3739) );
  INVX1 U3709 ( .A(n3742), .Y(n3740) );
  INVX1 U3710 ( .A(n3740), .Y(n3741) );
  BUFX2 U3711 ( .A(fifo[402]), .Y(n3742) );
  INVX1 U3712 ( .A(n3745), .Y(n3743) );
  INVX1 U3713 ( .A(n3743), .Y(n3744) );
  BUFX2 U3714 ( .A(fifo[403]), .Y(n3745) );
  INVX1 U3715 ( .A(n3748), .Y(n3746) );
  INVX1 U3716 ( .A(n3746), .Y(n3747) );
  BUFX2 U3717 ( .A(fifo[404]), .Y(n3748) );
  INVX1 U3718 ( .A(n3751), .Y(n3749) );
  INVX1 U3719 ( .A(n3749), .Y(n3750) );
  BUFX2 U3720 ( .A(fifo[405]), .Y(n3751) );
  INVX1 U3721 ( .A(n3754), .Y(n3752) );
  INVX1 U3722 ( .A(n3752), .Y(n3753) );
  BUFX2 U3723 ( .A(fifo[406]), .Y(n3754) );
  INVX1 U3724 ( .A(n3757), .Y(n3755) );
  INVX1 U3725 ( .A(n3755), .Y(n3756) );
  BUFX2 U3726 ( .A(fifo[407]), .Y(n3757) );
  INVX1 U3727 ( .A(n3760), .Y(n3758) );
  INVX1 U3728 ( .A(n3758), .Y(n3759) );
  BUFX2 U3729 ( .A(fifo[408]), .Y(n3760) );
  INVX1 U3730 ( .A(n3763), .Y(n3761) );
  INVX1 U3731 ( .A(n3761), .Y(n3762) );
  BUFX2 U3732 ( .A(fifo[409]), .Y(n3763) );
  INVX1 U3733 ( .A(n3766), .Y(n3764) );
  INVX1 U3734 ( .A(n3764), .Y(n3765) );
  BUFX2 U3735 ( .A(fifo[410]), .Y(n3766) );
  INVX1 U3736 ( .A(n3769), .Y(n3767) );
  INVX1 U3737 ( .A(n3767), .Y(n3768) );
  BUFX2 U3738 ( .A(fifo[411]), .Y(n3769) );
  INVX1 U3739 ( .A(n3772), .Y(n3770) );
  INVX1 U3740 ( .A(n3770), .Y(n3771) );
  BUFX2 U3741 ( .A(fifo[412]), .Y(n3772) );
  INVX1 U3742 ( .A(n3775), .Y(n3773) );
  INVX1 U3743 ( .A(n3773), .Y(n3774) );
  BUFX2 U3744 ( .A(fifo[413]), .Y(n3775) );
  INVX1 U3745 ( .A(n3778), .Y(n3776) );
  INVX1 U3746 ( .A(n3776), .Y(n3777) );
  BUFX2 U3747 ( .A(fifo[414]), .Y(n3778) );
  INVX1 U3748 ( .A(n3781), .Y(n3779) );
  INVX1 U3749 ( .A(n3779), .Y(n3780) );
  BUFX2 U3750 ( .A(fifo[415]), .Y(n3781) );
  INVX1 U3751 ( .A(n3784), .Y(n3782) );
  INVX1 U3752 ( .A(n3782), .Y(n3783) );
  BUFX2 U3753 ( .A(fifo[496]), .Y(n3784) );
  INVX1 U3754 ( .A(n3787), .Y(n3785) );
  INVX1 U3755 ( .A(n3785), .Y(n3786) );
  BUFX2 U3756 ( .A(fifo[497]), .Y(n3787) );
  INVX1 U3757 ( .A(n3790), .Y(n3788) );
  INVX1 U3758 ( .A(n3788), .Y(n3789) );
  BUFX2 U3759 ( .A(fifo[498]), .Y(n3790) );
  INVX1 U3760 ( .A(n3793), .Y(n3791) );
  INVX1 U3761 ( .A(n3791), .Y(n3792) );
  BUFX2 U3762 ( .A(fifo[499]), .Y(n3793) );
  INVX1 U3763 ( .A(n3796), .Y(n3794) );
  INVX1 U3764 ( .A(n3794), .Y(n3795) );
  BUFX2 U3765 ( .A(fifo[500]), .Y(n3796) );
  INVX1 U3766 ( .A(n3799), .Y(n3797) );
  INVX1 U3767 ( .A(n3797), .Y(n3798) );
  BUFX2 U3768 ( .A(fifo[501]), .Y(n3799) );
  INVX1 U3769 ( .A(n3802), .Y(n3800) );
  INVX1 U3770 ( .A(n3800), .Y(n3801) );
  BUFX2 U3771 ( .A(fifo[502]), .Y(n3802) );
  INVX1 U3772 ( .A(n3805), .Y(n3803) );
  INVX1 U3773 ( .A(n3803), .Y(n3804) );
  BUFX2 U3774 ( .A(fifo[503]), .Y(n3805) );
  INVX1 U3775 ( .A(n3808), .Y(n3806) );
  INVX1 U3776 ( .A(n3806), .Y(n3807) );
  BUFX2 U3777 ( .A(fifo[504]), .Y(n3808) );
  INVX1 U3778 ( .A(n3811), .Y(n3809) );
  INVX1 U3779 ( .A(n3809), .Y(n3810) );
  BUFX2 U3780 ( .A(fifo[505]), .Y(n3811) );
  INVX1 U3781 ( .A(n3814), .Y(n3812) );
  INVX1 U3782 ( .A(n3812), .Y(n3813) );
  BUFX2 U3783 ( .A(fifo[506]), .Y(n3814) );
  INVX1 U3784 ( .A(n3817), .Y(n3815) );
  INVX1 U3785 ( .A(n3815), .Y(n3816) );
  BUFX2 U3786 ( .A(fifo[507]), .Y(n3817) );
  INVX1 U3787 ( .A(n3820), .Y(n3818) );
  INVX1 U3788 ( .A(n3818), .Y(n3819) );
  BUFX2 U3789 ( .A(fifo[508]), .Y(n3820) );
  INVX1 U3790 ( .A(n3823), .Y(n3821) );
  INVX1 U3791 ( .A(n3821), .Y(n3822) );
  BUFX2 U3792 ( .A(fifo[509]), .Y(n3823) );
  INVX1 U3793 ( .A(n3826), .Y(n3824) );
  INVX1 U3794 ( .A(n3824), .Y(n3825) );
  BUFX2 U3795 ( .A(fifo[510]), .Y(n3826) );
  INVX1 U3796 ( .A(n3829), .Y(n3827) );
  INVX1 U3797 ( .A(n3827), .Y(n3828) );
  BUFX2 U3798 ( .A(fifo[511]), .Y(n3829) );
  INVX1 U3799 ( .A(n3832), .Y(n3830) );
  INVX1 U3800 ( .A(n3830), .Y(n3831) );
  BUFX2 U3801 ( .A(fifo[192]), .Y(n3832) );
  INVX1 U3802 ( .A(n3835), .Y(n3833) );
  INVX1 U3803 ( .A(n3833), .Y(n3834) );
  BUFX2 U3804 ( .A(fifo[193]), .Y(n3835) );
  INVX1 U3805 ( .A(n3838), .Y(n3836) );
  INVX1 U3806 ( .A(n3836), .Y(n3837) );
  BUFX2 U3807 ( .A(fifo[194]), .Y(n3838) );
  INVX1 U3808 ( .A(n3841), .Y(n3839) );
  INVX1 U3809 ( .A(n3839), .Y(n3840) );
  BUFX2 U3810 ( .A(fifo[195]), .Y(n3841) );
  INVX1 U3811 ( .A(n3844), .Y(n3842) );
  INVX1 U3812 ( .A(n3842), .Y(n3843) );
  BUFX2 U3813 ( .A(fifo[196]), .Y(n3844) );
  INVX1 U3814 ( .A(n3847), .Y(n3845) );
  INVX1 U3815 ( .A(n3845), .Y(n3846) );
  BUFX2 U3816 ( .A(fifo[197]), .Y(n3847) );
  INVX1 U3817 ( .A(n3850), .Y(n3848) );
  INVX1 U3818 ( .A(n3848), .Y(n3849) );
  BUFX2 U3819 ( .A(fifo[198]), .Y(n3850) );
  INVX1 U3820 ( .A(n3853), .Y(n3851) );
  INVX1 U3821 ( .A(n3851), .Y(n3852) );
  BUFX2 U3822 ( .A(fifo[199]), .Y(n3853) );
  INVX1 U3823 ( .A(n3856), .Y(n3854) );
  INVX1 U3824 ( .A(n3854), .Y(n3855) );
  BUFX2 U3825 ( .A(fifo[200]), .Y(n3856) );
  INVX1 U3826 ( .A(n3859), .Y(n3857) );
  INVX1 U3827 ( .A(n3857), .Y(n3858) );
  BUFX2 U3828 ( .A(fifo[201]), .Y(n3859) );
  INVX1 U3829 ( .A(n3862), .Y(n3860) );
  INVX1 U3830 ( .A(n3860), .Y(n3861) );
  BUFX2 U3831 ( .A(fifo[202]), .Y(n3862) );
  INVX1 U3832 ( .A(n3865), .Y(n3863) );
  INVX1 U3833 ( .A(n3863), .Y(n3864) );
  BUFX2 U3834 ( .A(fifo[203]), .Y(n3865) );
  INVX1 U3835 ( .A(n3868), .Y(n3866) );
  INVX1 U3836 ( .A(n3866), .Y(n3867) );
  BUFX2 U3837 ( .A(fifo[204]), .Y(n3868) );
  INVX1 U3838 ( .A(n3871), .Y(n3869) );
  INVX1 U3839 ( .A(n3869), .Y(n3870) );
  BUFX2 U3840 ( .A(fifo[205]), .Y(n3871) );
  INVX1 U3841 ( .A(n3874), .Y(n3872) );
  INVX1 U3842 ( .A(n3872), .Y(n3873) );
  BUFX2 U3843 ( .A(fifo[206]), .Y(n3874) );
  INVX1 U3844 ( .A(n3877), .Y(n3875) );
  INVX1 U3845 ( .A(n3875), .Y(n3876) );
  BUFX2 U3846 ( .A(fifo[207]), .Y(n3877) );
  INVX1 U3847 ( .A(n3880), .Y(n3878) );
  INVX1 U3848 ( .A(n3878), .Y(n3879) );
  BUFX2 U3849 ( .A(fifo[160]), .Y(n3880) );
  INVX1 U3850 ( .A(n3883), .Y(n3881) );
  INVX1 U3851 ( .A(n3881), .Y(n3882) );
  BUFX2 U3852 ( .A(fifo[161]), .Y(n3883) );
  INVX1 U3853 ( .A(n3886), .Y(n3884) );
  INVX1 U3854 ( .A(n3884), .Y(n3885) );
  BUFX2 U3855 ( .A(fifo[162]), .Y(n3886) );
  INVX1 U3856 ( .A(n3889), .Y(n3887) );
  INVX1 U3857 ( .A(n3887), .Y(n3888) );
  BUFX2 U3858 ( .A(fifo[163]), .Y(n3889) );
  INVX1 U3859 ( .A(n3892), .Y(n3890) );
  INVX1 U3860 ( .A(n3890), .Y(n3891) );
  BUFX2 U3861 ( .A(fifo[164]), .Y(n3892) );
  INVX1 U3862 ( .A(n3895), .Y(n3893) );
  INVX1 U3863 ( .A(n3893), .Y(n3894) );
  BUFX2 U3864 ( .A(fifo[165]), .Y(n3895) );
  INVX1 U3865 ( .A(n3898), .Y(n3896) );
  INVX1 U3866 ( .A(n3896), .Y(n3897) );
  BUFX2 U3867 ( .A(fifo[166]), .Y(n3898) );
  INVX1 U3868 ( .A(n3901), .Y(n3899) );
  INVX1 U3869 ( .A(n3899), .Y(n3900) );
  BUFX2 U3870 ( .A(fifo[167]), .Y(n3901) );
  INVX1 U3871 ( .A(n3904), .Y(n3902) );
  INVX1 U3872 ( .A(n3902), .Y(n3903) );
  BUFX2 U3873 ( .A(fifo[168]), .Y(n3904) );
  INVX1 U3874 ( .A(n3907), .Y(n3905) );
  INVX1 U3875 ( .A(n3905), .Y(n3906) );
  BUFX2 U3876 ( .A(fifo[169]), .Y(n3907) );
  INVX1 U3877 ( .A(n3910), .Y(n3908) );
  INVX1 U3878 ( .A(n3908), .Y(n3909) );
  BUFX2 U3879 ( .A(fifo[170]), .Y(n3910) );
  INVX1 U3880 ( .A(n3913), .Y(n3911) );
  INVX1 U3881 ( .A(n3911), .Y(n3912) );
  BUFX2 U3882 ( .A(fifo[171]), .Y(n3913) );
  INVX1 U3883 ( .A(n3916), .Y(n3914) );
  INVX1 U3884 ( .A(n3914), .Y(n3915) );
  BUFX2 U3885 ( .A(fifo[172]), .Y(n3916) );
  INVX1 U3886 ( .A(n3919), .Y(n3917) );
  INVX1 U3887 ( .A(n3917), .Y(n3918) );
  BUFX2 U3888 ( .A(fifo[173]), .Y(n3919) );
  INVX1 U3889 ( .A(n3922), .Y(n3920) );
  INVX1 U3890 ( .A(n3920), .Y(n3921) );
  BUFX2 U3891 ( .A(fifo[174]), .Y(n3922) );
  INVX1 U3892 ( .A(n3925), .Y(n3923) );
  INVX1 U3893 ( .A(n3923), .Y(n3924) );
  BUFX2 U3894 ( .A(fifo[175]), .Y(n3925) );
  INVX1 U3895 ( .A(n3928), .Y(n3926) );
  INVX1 U3896 ( .A(n3926), .Y(n3927) );
  BUFX2 U3897 ( .A(fifo[320]), .Y(n3928) );
  INVX1 U3898 ( .A(n3931), .Y(n3929) );
  INVX1 U3899 ( .A(n3929), .Y(n3930) );
  BUFX2 U3900 ( .A(fifo[321]), .Y(n3931) );
  INVX1 U3901 ( .A(n3934), .Y(n3932) );
  INVX1 U3902 ( .A(n3932), .Y(n3933) );
  BUFX2 U3903 ( .A(fifo[322]), .Y(n3934) );
  INVX1 U3904 ( .A(n3937), .Y(n3935) );
  INVX1 U3905 ( .A(n3935), .Y(n3936) );
  BUFX2 U3906 ( .A(fifo[323]), .Y(n3937) );
  INVX1 U3907 ( .A(n3940), .Y(n3938) );
  INVX1 U3908 ( .A(n3938), .Y(n3939) );
  BUFX2 U3909 ( .A(fifo[324]), .Y(n3940) );
  INVX1 U3910 ( .A(n3943), .Y(n3941) );
  INVX1 U3911 ( .A(n3941), .Y(n3942) );
  BUFX2 U3912 ( .A(fifo[325]), .Y(n3943) );
  INVX1 U3913 ( .A(n3946), .Y(n3944) );
  INVX1 U3914 ( .A(n3944), .Y(n3945) );
  BUFX2 U3915 ( .A(fifo[326]), .Y(n3946) );
  INVX1 U3916 ( .A(n3949), .Y(n3947) );
  INVX1 U3917 ( .A(n3947), .Y(n3948) );
  BUFX2 U3918 ( .A(fifo[327]), .Y(n3949) );
  INVX1 U3919 ( .A(n3952), .Y(n3950) );
  INVX1 U3920 ( .A(n3950), .Y(n3951) );
  BUFX2 U3921 ( .A(fifo[328]), .Y(n3952) );
  INVX1 U3922 ( .A(n3955), .Y(n3953) );
  INVX1 U3923 ( .A(n3953), .Y(n3954) );
  BUFX2 U3924 ( .A(fifo[329]), .Y(n3955) );
  INVX1 U3925 ( .A(n3958), .Y(n3956) );
  INVX1 U3926 ( .A(n3956), .Y(n3957) );
  BUFX2 U3927 ( .A(fifo[330]), .Y(n3958) );
  INVX1 U3928 ( .A(n3961), .Y(n3959) );
  INVX1 U3929 ( .A(n3959), .Y(n3960) );
  BUFX2 U3930 ( .A(fifo[331]), .Y(n3961) );
  INVX1 U3931 ( .A(n3964), .Y(n3962) );
  INVX1 U3932 ( .A(n3962), .Y(n3963) );
  BUFX2 U3933 ( .A(fifo[332]), .Y(n3964) );
  INVX1 U3934 ( .A(n3967), .Y(n3965) );
  INVX1 U3935 ( .A(n3965), .Y(n3966) );
  BUFX2 U3936 ( .A(fifo[333]), .Y(n3967) );
  INVX1 U3937 ( .A(n3970), .Y(n3968) );
  INVX1 U3938 ( .A(n3968), .Y(n3969) );
  BUFX2 U3939 ( .A(fifo[334]), .Y(n3970) );
  INVX1 U3940 ( .A(n3973), .Y(n3971) );
  INVX1 U3941 ( .A(n3971), .Y(n3972) );
  BUFX2 U3942 ( .A(fifo[335]), .Y(n3973) );
  INVX1 U3943 ( .A(n3976), .Y(n3974) );
  INVX1 U3944 ( .A(n3974), .Y(n3975) );
  BUFX2 U3945 ( .A(fifo[288]), .Y(n3976) );
  INVX1 U3946 ( .A(n3979), .Y(n3977) );
  INVX1 U3947 ( .A(n3977), .Y(n3978) );
  BUFX2 U3948 ( .A(fifo[289]), .Y(n3979) );
  INVX1 U3949 ( .A(n3982), .Y(n3980) );
  INVX1 U3950 ( .A(n3980), .Y(n3981) );
  BUFX2 U3951 ( .A(fifo[290]), .Y(n3982) );
  INVX1 U3952 ( .A(n3985), .Y(n3983) );
  INVX1 U3953 ( .A(n3983), .Y(n3984) );
  BUFX2 U3954 ( .A(fifo[291]), .Y(n3985) );
  INVX1 U3955 ( .A(n3988), .Y(n3986) );
  INVX1 U3956 ( .A(n3986), .Y(n3987) );
  BUFX2 U3957 ( .A(fifo[292]), .Y(n3988) );
  INVX1 U3958 ( .A(n3991), .Y(n3989) );
  INVX1 U3959 ( .A(n3989), .Y(n3990) );
  BUFX2 U3960 ( .A(fifo[293]), .Y(n3991) );
  INVX1 U3961 ( .A(n3994), .Y(n3992) );
  INVX1 U3962 ( .A(n3992), .Y(n3993) );
  BUFX2 U3963 ( .A(fifo[294]), .Y(n3994) );
  INVX1 U3964 ( .A(n3997), .Y(n3995) );
  INVX1 U3965 ( .A(n3995), .Y(n3996) );
  BUFX2 U3966 ( .A(fifo[295]), .Y(n3997) );
  INVX1 U3967 ( .A(n4000), .Y(n3998) );
  INVX1 U3968 ( .A(n3998), .Y(n3999) );
  BUFX2 U3969 ( .A(fifo[296]), .Y(n4000) );
  INVX1 U3970 ( .A(n4003), .Y(n4001) );
  INVX1 U3971 ( .A(n4001), .Y(n4002) );
  BUFX2 U3972 ( .A(fifo[297]), .Y(n4003) );
  INVX1 U3973 ( .A(n4006), .Y(n4004) );
  INVX1 U3974 ( .A(n4004), .Y(n4005) );
  BUFX2 U3975 ( .A(fifo[298]), .Y(n4006) );
  INVX1 U3976 ( .A(n4009), .Y(n4007) );
  INVX1 U3977 ( .A(n4007), .Y(n4008) );
  BUFX2 U3978 ( .A(fifo[299]), .Y(n4009) );
  INVX1 U3979 ( .A(n4012), .Y(n4010) );
  INVX1 U3980 ( .A(n4010), .Y(n4011) );
  BUFX2 U3981 ( .A(fifo[300]), .Y(n4012) );
  INVX1 U3982 ( .A(n4015), .Y(n4013) );
  INVX1 U3983 ( .A(n4013), .Y(n4014) );
  BUFX2 U3984 ( .A(fifo[301]), .Y(n4015) );
  INVX1 U3985 ( .A(n4018), .Y(n4016) );
  INVX1 U3986 ( .A(n4016), .Y(n4017) );
  BUFX2 U3987 ( .A(fifo[302]), .Y(n4018) );
  INVX1 U3988 ( .A(n4021), .Y(n4019) );
  INVX1 U3989 ( .A(n4019), .Y(n4020) );
  BUFX2 U3990 ( .A(fifo[303]), .Y(n4021) );
  INVX1 U3991 ( .A(n4024), .Y(n4022) );
  INVX1 U3992 ( .A(n4022), .Y(n4023) );
  BUFX2 U3993 ( .A(fifo[128]), .Y(n4024) );
  INVX1 U3994 ( .A(n4027), .Y(n4025) );
  INVX1 U3995 ( .A(n4025), .Y(n4026) );
  BUFX2 U3996 ( .A(fifo[129]), .Y(n4027) );
  INVX1 U3997 ( .A(n4030), .Y(n4028) );
  INVX1 U3998 ( .A(n4028), .Y(n4029) );
  BUFX2 U3999 ( .A(fifo[130]), .Y(n4030) );
  INVX1 U4000 ( .A(n4033), .Y(n4031) );
  INVX1 U4001 ( .A(n4031), .Y(n4032) );
  BUFX2 U4002 ( .A(fifo[131]), .Y(n4033) );
  INVX1 U4003 ( .A(n4036), .Y(n4034) );
  INVX1 U4004 ( .A(n4034), .Y(n4035) );
  BUFX2 U4005 ( .A(fifo[132]), .Y(n4036) );
  INVX1 U4006 ( .A(n4039), .Y(n4037) );
  INVX1 U4007 ( .A(n4037), .Y(n4038) );
  BUFX2 U4008 ( .A(fifo[133]), .Y(n4039) );
  INVX1 U4009 ( .A(n4042), .Y(n4040) );
  INVX1 U4010 ( .A(n4040), .Y(n4041) );
  BUFX2 U4011 ( .A(fifo[134]), .Y(n4042) );
  INVX1 U4012 ( .A(n4045), .Y(n4043) );
  INVX1 U4013 ( .A(n4043), .Y(n4044) );
  BUFX2 U4014 ( .A(fifo[135]), .Y(n4045) );
  INVX1 U4015 ( .A(n4048), .Y(n4046) );
  INVX1 U4016 ( .A(n4046), .Y(n4047) );
  BUFX2 U4017 ( .A(fifo[136]), .Y(n4048) );
  INVX1 U4018 ( .A(n4051), .Y(n4049) );
  INVX1 U4019 ( .A(n4049), .Y(n4050) );
  BUFX2 U4020 ( .A(fifo[137]), .Y(n4051) );
  INVX1 U4021 ( .A(n4054), .Y(n4052) );
  INVX1 U4022 ( .A(n4052), .Y(n4053) );
  BUFX2 U4023 ( .A(fifo[138]), .Y(n4054) );
  INVX1 U4024 ( .A(n4057), .Y(n4055) );
  INVX1 U4025 ( .A(n4055), .Y(n4056) );
  BUFX2 U4026 ( .A(fifo[139]), .Y(n4057) );
  INVX1 U4027 ( .A(n4060), .Y(n4058) );
  INVX1 U4028 ( .A(n4058), .Y(n4059) );
  BUFX2 U4029 ( .A(fifo[140]), .Y(n4060) );
  INVX1 U4030 ( .A(n4063), .Y(n4061) );
  INVX1 U4031 ( .A(n4061), .Y(n4062) );
  BUFX2 U4032 ( .A(fifo[141]), .Y(n4063) );
  INVX1 U4033 ( .A(n4066), .Y(n4064) );
  INVX1 U4034 ( .A(n4064), .Y(n4065) );
  BUFX2 U4035 ( .A(fifo[142]), .Y(n4066) );
  INVX1 U4036 ( .A(n4069), .Y(n4067) );
  INVX1 U4037 ( .A(n4067), .Y(n4068) );
  BUFX2 U4038 ( .A(fifo[143]), .Y(n4069) );
  INVX1 U4039 ( .A(n4072), .Y(n4070) );
  INVX1 U4040 ( .A(n4070), .Y(n4071) );
  BUFX2 U4041 ( .A(fifo[256]), .Y(n4072) );
  INVX1 U4042 ( .A(n4075), .Y(n4073) );
  INVX1 U4043 ( .A(n4073), .Y(n4074) );
  BUFX2 U4044 ( .A(fifo[257]), .Y(n4075) );
  INVX1 U4045 ( .A(n4078), .Y(n4076) );
  INVX1 U4046 ( .A(n4076), .Y(n4077) );
  BUFX2 U4047 ( .A(fifo[258]), .Y(n4078) );
  INVX1 U4048 ( .A(n4081), .Y(n4079) );
  INVX1 U4049 ( .A(n4079), .Y(n4080) );
  BUFX2 U4050 ( .A(fifo[259]), .Y(n4081) );
  INVX1 U4051 ( .A(n4084), .Y(n4082) );
  INVX1 U4052 ( .A(n4082), .Y(n4083) );
  BUFX2 U4053 ( .A(fifo[260]), .Y(n4084) );
  INVX1 U4054 ( .A(n4087), .Y(n4085) );
  INVX1 U4055 ( .A(n4085), .Y(n4086) );
  BUFX2 U4056 ( .A(fifo[261]), .Y(n4087) );
  INVX1 U4057 ( .A(n4090), .Y(n4088) );
  INVX1 U4058 ( .A(n4088), .Y(n4089) );
  BUFX2 U4059 ( .A(fifo[262]), .Y(n4090) );
  INVX1 U4060 ( .A(n4093), .Y(n4091) );
  INVX1 U4061 ( .A(n4091), .Y(n4092) );
  BUFX2 U4062 ( .A(fifo[263]), .Y(n4093) );
  INVX1 U4063 ( .A(n4096), .Y(n4094) );
  INVX1 U4064 ( .A(n4094), .Y(n4095) );
  BUFX2 U4065 ( .A(fifo[264]), .Y(n4096) );
  INVX1 U4066 ( .A(n4099), .Y(n4097) );
  INVX1 U4067 ( .A(n4097), .Y(n4098) );
  BUFX2 U4068 ( .A(fifo[265]), .Y(n4099) );
  INVX1 U4069 ( .A(n4102), .Y(n4100) );
  INVX1 U4070 ( .A(n4100), .Y(n4101) );
  BUFX2 U4071 ( .A(fifo[266]), .Y(n4102) );
  INVX1 U4072 ( .A(n4105), .Y(n4103) );
  INVX1 U4073 ( .A(n4103), .Y(n4104) );
  BUFX2 U4074 ( .A(fifo[267]), .Y(n4105) );
  INVX1 U4075 ( .A(n4108), .Y(n4106) );
  INVX1 U4076 ( .A(n4106), .Y(n4107) );
  BUFX2 U4077 ( .A(fifo[268]), .Y(n4108) );
  INVX1 U4078 ( .A(n4111), .Y(n4109) );
  INVX1 U4079 ( .A(n4109), .Y(n4110) );
  BUFX2 U4080 ( .A(fifo[269]), .Y(n4111) );
  INVX1 U4081 ( .A(n4114), .Y(n4112) );
  INVX1 U4082 ( .A(n4112), .Y(n4113) );
  BUFX2 U4083 ( .A(fifo[270]), .Y(n4114) );
  INVX1 U4084 ( .A(n4117), .Y(n4115) );
  INVX1 U4085 ( .A(n4115), .Y(n4116) );
  BUFX2 U4086 ( .A(fifo[271]), .Y(n4117) );
  INVX1 U4087 ( .A(n4120), .Y(n4118) );
  INVX1 U4088 ( .A(n4118), .Y(n4119) );
  BUFX2 U4089 ( .A(fifo[224]), .Y(n4120) );
  INVX1 U4090 ( .A(n4123), .Y(n4121) );
  INVX1 U4091 ( .A(n4121), .Y(n4122) );
  BUFX2 U4092 ( .A(fifo[225]), .Y(n4123) );
  INVX1 U4093 ( .A(n4126), .Y(n4124) );
  INVX1 U4094 ( .A(n4124), .Y(n4125) );
  BUFX2 U4095 ( .A(fifo[226]), .Y(n4126) );
  INVX1 U4096 ( .A(n4129), .Y(n4127) );
  INVX1 U4097 ( .A(n4127), .Y(n4128) );
  BUFX2 U4098 ( .A(fifo[227]), .Y(n4129) );
  INVX1 U4099 ( .A(n4132), .Y(n4130) );
  INVX1 U4100 ( .A(n4130), .Y(n4131) );
  BUFX2 U4101 ( .A(fifo[228]), .Y(n4132) );
  INVX1 U4102 ( .A(n4135), .Y(n4133) );
  INVX1 U4103 ( .A(n4133), .Y(n4134) );
  BUFX2 U4104 ( .A(fifo[229]), .Y(n4135) );
  INVX1 U4105 ( .A(n4138), .Y(n4136) );
  INVX1 U4106 ( .A(n4136), .Y(n4137) );
  BUFX2 U4107 ( .A(fifo[230]), .Y(n4138) );
  INVX1 U4108 ( .A(n4141), .Y(n4139) );
  INVX1 U4109 ( .A(n4139), .Y(n4140) );
  BUFX2 U4110 ( .A(fifo[231]), .Y(n4141) );
  INVX1 U4111 ( .A(n4144), .Y(n4142) );
  INVX1 U4112 ( .A(n4142), .Y(n4143) );
  BUFX2 U4113 ( .A(fifo[232]), .Y(n4144) );
  INVX1 U4114 ( .A(n4147), .Y(n4145) );
  INVX1 U4115 ( .A(n4145), .Y(n4146) );
  BUFX2 U4116 ( .A(fifo[233]), .Y(n4147) );
  INVX1 U4117 ( .A(n4150), .Y(n4148) );
  INVX1 U4118 ( .A(n4148), .Y(n4149) );
  BUFX2 U4119 ( .A(fifo[234]), .Y(n4150) );
  INVX1 U4120 ( .A(n4153), .Y(n4151) );
  INVX1 U4121 ( .A(n4151), .Y(n4152) );
  BUFX2 U4122 ( .A(fifo[235]), .Y(n4153) );
  INVX1 U4123 ( .A(n4156), .Y(n4154) );
  INVX1 U4124 ( .A(n4154), .Y(n4155) );
  BUFX2 U4125 ( .A(fifo[236]), .Y(n4156) );
  INVX1 U4126 ( .A(n4159), .Y(n4157) );
  INVX1 U4127 ( .A(n4157), .Y(n4158) );
  BUFX2 U4128 ( .A(fifo[237]), .Y(n4159) );
  INVX1 U4129 ( .A(n4162), .Y(n4160) );
  INVX1 U4130 ( .A(n4160), .Y(n4161) );
  BUFX2 U4131 ( .A(fifo[238]), .Y(n4162) );
  INVX1 U4132 ( .A(n4165), .Y(n4163) );
  INVX1 U4133 ( .A(n4163), .Y(n4164) );
  BUFX2 U4134 ( .A(fifo[239]), .Y(n4165) );
  INVX1 U4135 ( .A(n4168), .Y(n4166) );
  INVX1 U4136 ( .A(n4166), .Y(n4167) );
  BUFX2 U4137 ( .A(fifo[352]), .Y(n4168) );
  INVX1 U4138 ( .A(n4171), .Y(n4169) );
  INVX1 U4139 ( .A(n4169), .Y(n4170) );
  BUFX2 U4140 ( .A(fifo[353]), .Y(n4171) );
  INVX1 U4141 ( .A(n4174), .Y(n4172) );
  INVX1 U4142 ( .A(n4172), .Y(n4173) );
  BUFX2 U4143 ( .A(fifo[354]), .Y(n4174) );
  INVX1 U4144 ( .A(n4177), .Y(n4175) );
  INVX1 U4145 ( .A(n4175), .Y(n4176) );
  BUFX2 U4146 ( .A(fifo[355]), .Y(n4177) );
  INVX1 U4147 ( .A(n4180), .Y(n4178) );
  INVX1 U4148 ( .A(n4178), .Y(n4179) );
  BUFX2 U4149 ( .A(fifo[356]), .Y(n4180) );
  INVX1 U4150 ( .A(n4183), .Y(n4181) );
  INVX1 U4151 ( .A(n4181), .Y(n4182) );
  BUFX2 U4152 ( .A(fifo[357]), .Y(n4183) );
  INVX1 U4153 ( .A(n4186), .Y(n4184) );
  INVX1 U4154 ( .A(n4184), .Y(n4185) );
  BUFX2 U4155 ( .A(fifo[358]), .Y(n4186) );
  INVX1 U4156 ( .A(n4189), .Y(n4187) );
  INVX1 U4157 ( .A(n4187), .Y(n4188) );
  BUFX2 U4158 ( .A(fifo[359]), .Y(n4189) );
  INVX1 U4159 ( .A(n4192), .Y(n4190) );
  INVX1 U4160 ( .A(n4190), .Y(n4191) );
  BUFX2 U4161 ( .A(fifo[360]), .Y(n4192) );
  INVX1 U4162 ( .A(n4195), .Y(n4193) );
  INVX1 U4163 ( .A(n4193), .Y(n4194) );
  BUFX2 U4164 ( .A(fifo[361]), .Y(n4195) );
  INVX1 U4165 ( .A(n4198), .Y(n4196) );
  INVX1 U4166 ( .A(n4196), .Y(n4197) );
  BUFX2 U4167 ( .A(fifo[362]), .Y(n4198) );
  INVX1 U4168 ( .A(n4201), .Y(n4199) );
  INVX1 U4169 ( .A(n4199), .Y(n4200) );
  BUFX2 U4170 ( .A(fifo[363]), .Y(n4201) );
  INVX1 U4171 ( .A(n4204), .Y(n4202) );
  INVX1 U4172 ( .A(n4202), .Y(n4203) );
  BUFX2 U4173 ( .A(fifo[364]), .Y(n4204) );
  INVX1 U4174 ( .A(n4207), .Y(n4205) );
  INVX1 U4175 ( .A(n4205), .Y(n4206) );
  BUFX2 U4176 ( .A(fifo[365]), .Y(n4207) );
  INVX1 U4177 ( .A(n4210), .Y(n4208) );
  INVX1 U4178 ( .A(n4208), .Y(n4209) );
  BUFX2 U4179 ( .A(fifo[366]), .Y(n4210) );
  INVX1 U4180 ( .A(n4213), .Y(n4211) );
  INVX1 U4181 ( .A(n4211), .Y(n4212) );
  BUFX2 U4182 ( .A(fifo[367]), .Y(n4213) );
  INVX1 U4183 ( .A(n4216), .Y(n4214) );
  INVX1 U4184 ( .A(n4214), .Y(n4215) );
  BUFX2 U4185 ( .A(fifo[64]), .Y(n4216) );
  INVX1 U4186 ( .A(n4219), .Y(n4217) );
  INVX1 U4187 ( .A(n4217), .Y(n4218) );
  BUFX2 U4188 ( .A(fifo[65]), .Y(n4219) );
  INVX1 U4189 ( .A(n4222), .Y(n4220) );
  INVX1 U4190 ( .A(n4220), .Y(n4221) );
  BUFX2 U4191 ( .A(fifo[66]), .Y(n4222) );
  INVX1 U4192 ( .A(n4225), .Y(n4223) );
  INVX1 U4193 ( .A(n4223), .Y(n4224) );
  BUFX2 U4194 ( .A(fifo[67]), .Y(n4225) );
  INVX1 U4195 ( .A(n4228), .Y(n4226) );
  INVX1 U4196 ( .A(n4226), .Y(n4227) );
  BUFX2 U4197 ( .A(fifo[68]), .Y(n4228) );
  INVX1 U4198 ( .A(n4231), .Y(n4229) );
  INVX1 U4199 ( .A(n4229), .Y(n4230) );
  BUFX2 U4200 ( .A(fifo[69]), .Y(n4231) );
  INVX1 U4201 ( .A(n4234), .Y(n4232) );
  INVX1 U4202 ( .A(n4232), .Y(n4233) );
  BUFX2 U4203 ( .A(fifo[70]), .Y(n4234) );
  INVX1 U4204 ( .A(n4237), .Y(n4235) );
  INVX1 U4205 ( .A(n4235), .Y(n4236) );
  BUFX2 U4206 ( .A(fifo[71]), .Y(n4237) );
  INVX1 U4207 ( .A(n4240), .Y(n4238) );
  INVX1 U4208 ( .A(n4238), .Y(n4239) );
  BUFX2 U4209 ( .A(fifo[72]), .Y(n4240) );
  INVX1 U4210 ( .A(n4243), .Y(n4241) );
  INVX1 U4211 ( .A(n4241), .Y(n4242) );
  BUFX2 U4212 ( .A(fifo[73]), .Y(n4243) );
  INVX1 U4213 ( .A(n4246), .Y(n4244) );
  INVX1 U4214 ( .A(n4244), .Y(n4245) );
  BUFX2 U4215 ( .A(fifo[74]), .Y(n4246) );
  INVX1 U4216 ( .A(n4249), .Y(n4247) );
  INVX1 U4217 ( .A(n4247), .Y(n4248) );
  BUFX2 U4218 ( .A(fifo[75]), .Y(n4249) );
  INVX1 U4219 ( .A(n4252), .Y(n4250) );
  INVX1 U4220 ( .A(n4250), .Y(n4251) );
  BUFX2 U4221 ( .A(fifo[76]), .Y(n4252) );
  INVX1 U4222 ( .A(n4255), .Y(n4253) );
  INVX1 U4223 ( .A(n4253), .Y(n4254) );
  BUFX2 U4224 ( .A(fifo[77]), .Y(n4255) );
  INVX1 U4225 ( .A(n4258), .Y(n4256) );
  INVX1 U4226 ( .A(n4256), .Y(n4257) );
  BUFX2 U4227 ( .A(fifo[78]), .Y(n4258) );
  INVX1 U4228 ( .A(n4261), .Y(n4259) );
  INVX1 U4229 ( .A(n4259), .Y(n4260) );
  BUFX2 U4230 ( .A(fifo[79]), .Y(n4261) );
  INVX1 U4231 ( .A(n4264), .Y(n4262) );
  INVX1 U4232 ( .A(n4262), .Y(n4263) );
  BUFX2 U4233 ( .A(fifo[32]), .Y(n4264) );
  INVX1 U4234 ( .A(n4267), .Y(n4265) );
  INVX1 U4235 ( .A(n4265), .Y(n4266) );
  BUFX2 U4236 ( .A(fifo[33]), .Y(n4267) );
  INVX1 U4237 ( .A(n4270), .Y(n4268) );
  INVX1 U4238 ( .A(n4268), .Y(n4269) );
  BUFX2 U4239 ( .A(fifo[34]), .Y(n4270) );
  INVX1 U4240 ( .A(n4273), .Y(n4271) );
  INVX1 U4241 ( .A(n4271), .Y(n4272) );
  BUFX2 U4242 ( .A(fifo[35]), .Y(n4273) );
  INVX1 U4243 ( .A(n4276), .Y(n4274) );
  INVX1 U4244 ( .A(n4274), .Y(n4275) );
  BUFX2 U4245 ( .A(fifo[36]), .Y(n4276) );
  INVX1 U4246 ( .A(n4279), .Y(n4277) );
  INVX1 U4247 ( .A(n4277), .Y(n4278) );
  BUFX2 U4248 ( .A(fifo[37]), .Y(n4279) );
  INVX1 U4249 ( .A(n4282), .Y(n4280) );
  INVX1 U4250 ( .A(n4280), .Y(n4281) );
  BUFX2 U4251 ( .A(fifo[38]), .Y(n4282) );
  INVX1 U4252 ( .A(n4285), .Y(n4283) );
  INVX1 U4253 ( .A(n4283), .Y(n4284) );
  BUFX2 U4254 ( .A(fifo[39]), .Y(n4285) );
  INVX1 U4255 ( .A(n4288), .Y(n4286) );
  INVX1 U4256 ( .A(n4286), .Y(n4287) );
  BUFX2 U4257 ( .A(fifo[40]), .Y(n4288) );
  INVX1 U4258 ( .A(n4291), .Y(n4289) );
  INVX1 U4259 ( .A(n4289), .Y(n4290) );
  BUFX2 U4260 ( .A(fifo[41]), .Y(n4291) );
  INVX1 U4261 ( .A(n4294), .Y(n4292) );
  INVX1 U4262 ( .A(n4292), .Y(n4293) );
  BUFX2 U4263 ( .A(fifo[42]), .Y(n4294) );
  INVX1 U4264 ( .A(n4297), .Y(n4295) );
  INVX1 U4265 ( .A(n4295), .Y(n4296) );
  BUFX2 U4266 ( .A(fifo[43]), .Y(n4297) );
  INVX1 U4267 ( .A(n4300), .Y(n4298) );
  INVX1 U4268 ( .A(n4298), .Y(n4299) );
  BUFX2 U4269 ( .A(fifo[44]), .Y(n4300) );
  INVX1 U4270 ( .A(n4303), .Y(n4301) );
  INVX1 U4271 ( .A(n4301), .Y(n4302) );
  BUFX2 U4272 ( .A(fifo[45]), .Y(n4303) );
  INVX1 U4273 ( .A(n4306), .Y(n4304) );
  INVX1 U4274 ( .A(n4304), .Y(n4305) );
  BUFX2 U4275 ( .A(fifo[46]), .Y(n4306) );
  INVX1 U4276 ( .A(n4309), .Y(n4307) );
  INVX1 U4277 ( .A(n4307), .Y(n4308) );
  BUFX2 U4278 ( .A(fifo[47]), .Y(n4309) );
  INVX1 U4279 ( .A(n4312), .Y(n4310) );
  INVX1 U4280 ( .A(n4310), .Y(n4311) );
  BUFX2 U4281 ( .A(fifo[0]), .Y(n4312) );
  INVX1 U4282 ( .A(n4315), .Y(n4313) );
  INVX1 U4283 ( .A(n4313), .Y(n4314) );
  BUFX2 U4284 ( .A(fifo[1]), .Y(n4315) );
  INVX1 U4285 ( .A(n4318), .Y(n4316) );
  INVX1 U4286 ( .A(n4316), .Y(n4317) );
  BUFX2 U4287 ( .A(fifo[2]), .Y(n4318) );
  INVX1 U4288 ( .A(n4321), .Y(n4319) );
  INVX1 U4289 ( .A(n4319), .Y(n4320) );
  BUFX2 U4290 ( .A(fifo[3]), .Y(n4321) );
  INVX1 U4291 ( .A(n4324), .Y(n4322) );
  INVX1 U4292 ( .A(n4322), .Y(n4323) );
  BUFX2 U4293 ( .A(fifo[4]), .Y(n4324) );
  INVX1 U4294 ( .A(n4327), .Y(n4325) );
  INVX1 U4295 ( .A(n4325), .Y(n4326) );
  BUFX2 U4296 ( .A(fifo[5]), .Y(n4327) );
  INVX1 U4297 ( .A(n4330), .Y(n4328) );
  INVX1 U4298 ( .A(n4328), .Y(n4329) );
  BUFX2 U4299 ( .A(fifo[6]), .Y(n4330) );
  INVX1 U4300 ( .A(n4333), .Y(n4331) );
  INVX1 U4301 ( .A(n4331), .Y(n4332) );
  BUFX2 U4302 ( .A(fifo[7]), .Y(n4333) );
  INVX1 U4303 ( .A(n4336), .Y(n4334) );
  INVX1 U4304 ( .A(n4334), .Y(n4335) );
  BUFX2 U4305 ( .A(fifo[8]), .Y(n4336) );
  INVX1 U4306 ( .A(n4339), .Y(n4337) );
  INVX1 U4307 ( .A(n4337), .Y(n4338) );
  BUFX2 U4308 ( .A(fifo[9]), .Y(n4339) );
  INVX1 U4309 ( .A(n4342), .Y(n4340) );
  INVX1 U4310 ( .A(n4340), .Y(n4341) );
  BUFX2 U4311 ( .A(fifo[10]), .Y(n4342) );
  INVX1 U4312 ( .A(n4345), .Y(n4343) );
  INVX1 U4313 ( .A(n4343), .Y(n4344) );
  BUFX2 U4314 ( .A(fifo[11]), .Y(n4345) );
  INVX1 U4315 ( .A(n4348), .Y(n4346) );
  INVX1 U4316 ( .A(n4346), .Y(n4347) );
  BUFX2 U4317 ( .A(fifo[12]), .Y(n4348) );
  INVX1 U4318 ( .A(n4351), .Y(n4349) );
  INVX1 U4319 ( .A(n4349), .Y(n4350) );
  BUFX2 U4320 ( .A(fifo[13]), .Y(n4351) );
  INVX1 U4321 ( .A(n4354), .Y(n4352) );
  INVX1 U4322 ( .A(n4352), .Y(n4353) );
  BUFX2 U4323 ( .A(fifo[14]), .Y(n4354) );
  INVX1 U4324 ( .A(n4357), .Y(n4355) );
  INVX1 U4325 ( .A(n4355), .Y(n4356) );
  BUFX2 U4326 ( .A(fifo[15]), .Y(n4357) );
  INVX1 U4327 ( .A(n4360), .Y(n4358) );
  INVX1 U4328 ( .A(n4358), .Y(n4359) );
  BUFX2 U4329 ( .A(fifo[96]), .Y(n4360) );
  INVX1 U4330 ( .A(n4363), .Y(n4361) );
  INVX1 U4331 ( .A(n4361), .Y(n4362) );
  BUFX2 U4332 ( .A(fifo[97]), .Y(n4363) );
  INVX1 U4333 ( .A(n4366), .Y(n4364) );
  INVX1 U4334 ( .A(n4364), .Y(n4365) );
  BUFX2 U4335 ( .A(fifo[98]), .Y(n4366) );
  INVX1 U4336 ( .A(n4369), .Y(n4367) );
  INVX1 U4337 ( .A(n4367), .Y(n4368) );
  BUFX2 U4338 ( .A(fifo[99]), .Y(n4369) );
  INVX1 U4339 ( .A(n4372), .Y(n4370) );
  INVX1 U4340 ( .A(n4370), .Y(n4371) );
  BUFX2 U4341 ( .A(fifo[100]), .Y(n4372) );
  INVX1 U4342 ( .A(n4375), .Y(n4373) );
  INVX1 U4343 ( .A(n4373), .Y(n4374) );
  BUFX2 U4344 ( .A(fifo[101]), .Y(n4375) );
  INVX1 U4345 ( .A(n4378), .Y(n4376) );
  INVX1 U4346 ( .A(n4376), .Y(n4377) );
  BUFX2 U4347 ( .A(fifo[102]), .Y(n4378) );
  INVX1 U4348 ( .A(n4381), .Y(n4379) );
  INVX1 U4349 ( .A(n4379), .Y(n4380) );
  BUFX2 U4350 ( .A(fifo[103]), .Y(n4381) );
  INVX1 U4351 ( .A(n4384), .Y(n4382) );
  INVX1 U4352 ( .A(n4382), .Y(n4383) );
  BUFX2 U4353 ( .A(fifo[104]), .Y(n4384) );
  INVX1 U4354 ( .A(n4387), .Y(n4385) );
  INVX1 U4355 ( .A(n4385), .Y(n4386) );
  BUFX2 U4356 ( .A(fifo[105]), .Y(n4387) );
  INVX1 U4357 ( .A(n4390), .Y(n4388) );
  INVX1 U4358 ( .A(n4388), .Y(n4389) );
  BUFX2 U4359 ( .A(fifo[106]), .Y(n4390) );
  INVX1 U4360 ( .A(n4393), .Y(n4391) );
  INVX1 U4361 ( .A(n4391), .Y(n4392) );
  BUFX2 U4362 ( .A(fifo[107]), .Y(n4393) );
  INVX1 U4363 ( .A(n4396), .Y(n4394) );
  INVX1 U4364 ( .A(n4394), .Y(n4395) );
  BUFX2 U4365 ( .A(fifo[108]), .Y(n4396) );
  INVX1 U4366 ( .A(n4399), .Y(n4397) );
  INVX1 U4367 ( .A(n4397), .Y(n4398) );
  BUFX2 U4368 ( .A(fifo[109]), .Y(n4399) );
  INVX1 U4369 ( .A(n4402), .Y(n4400) );
  INVX1 U4370 ( .A(n4400), .Y(n4401) );
  BUFX2 U4371 ( .A(fifo[110]), .Y(n4402) );
  INVX1 U4372 ( .A(n4405), .Y(n4403) );
  INVX1 U4373 ( .A(n4403), .Y(n4404) );
  BUFX2 U4374 ( .A(fifo[111]), .Y(n4405) );
  INVX1 U4375 ( .A(n4408), .Y(n4406) );
  INVX1 U4376 ( .A(n4406), .Y(n4407) );
  BUFX2 U4377 ( .A(fifo[480]), .Y(n4408) );
  INVX1 U4378 ( .A(n4411), .Y(n4409) );
  INVX1 U4379 ( .A(n4409), .Y(n4410) );
  BUFX2 U4380 ( .A(fifo[481]), .Y(n4411) );
  INVX1 U4381 ( .A(n4414), .Y(n4412) );
  INVX1 U4382 ( .A(n4412), .Y(n4413) );
  BUFX2 U4383 ( .A(fifo[482]), .Y(n4414) );
  INVX1 U4384 ( .A(n4417), .Y(n4415) );
  INVX1 U4385 ( .A(n4415), .Y(n4416) );
  BUFX2 U4386 ( .A(fifo[483]), .Y(n4417) );
  INVX1 U4387 ( .A(n4420), .Y(n4418) );
  INVX1 U4388 ( .A(n4418), .Y(n4419) );
  BUFX2 U4389 ( .A(fifo[484]), .Y(n4420) );
  INVX1 U4390 ( .A(n4423), .Y(n4421) );
  INVX1 U4391 ( .A(n4421), .Y(n4422) );
  BUFX2 U4392 ( .A(fifo[485]), .Y(n4423) );
  INVX1 U4393 ( .A(n4426), .Y(n4424) );
  INVX1 U4394 ( .A(n4424), .Y(n4425) );
  BUFX2 U4395 ( .A(fifo[486]), .Y(n4426) );
  INVX1 U4396 ( .A(n4429), .Y(n4427) );
  INVX1 U4397 ( .A(n4427), .Y(n4428) );
  BUFX2 U4398 ( .A(fifo[487]), .Y(n4429) );
  INVX1 U4399 ( .A(n4432), .Y(n4430) );
  INVX1 U4400 ( .A(n4430), .Y(n4431) );
  BUFX2 U4401 ( .A(fifo[488]), .Y(n4432) );
  INVX1 U4402 ( .A(n4435), .Y(n4433) );
  INVX1 U4403 ( .A(n4433), .Y(n4434) );
  BUFX2 U4404 ( .A(fifo[489]), .Y(n4435) );
  INVX1 U4405 ( .A(n4438), .Y(n4436) );
  INVX1 U4406 ( .A(n4436), .Y(n4437) );
  BUFX2 U4407 ( .A(fifo[490]), .Y(n4438) );
  INVX1 U4408 ( .A(n4441), .Y(n4439) );
  INVX1 U4409 ( .A(n4439), .Y(n4440) );
  BUFX2 U4410 ( .A(fifo[491]), .Y(n4441) );
  INVX1 U4411 ( .A(n4444), .Y(n4442) );
  INVX1 U4412 ( .A(n4442), .Y(n4443) );
  BUFX2 U4413 ( .A(fifo[492]), .Y(n4444) );
  INVX1 U4414 ( .A(n4447), .Y(n4445) );
  INVX1 U4415 ( .A(n4445), .Y(n4446) );
  BUFX2 U4416 ( .A(fifo[493]), .Y(n4447) );
  INVX1 U4417 ( .A(n4450), .Y(n4448) );
  INVX1 U4418 ( .A(n4448), .Y(n4449) );
  BUFX2 U4419 ( .A(fifo[494]), .Y(n4450) );
  INVX1 U4420 ( .A(n4453), .Y(n4451) );
  INVX1 U4421 ( .A(n4451), .Y(n4452) );
  BUFX2 U4422 ( .A(fifo[495]), .Y(n4453) );
  INVX1 U4423 ( .A(n4456), .Y(n4454) );
  INVX1 U4424 ( .A(n4454), .Y(n4455) );
  BUFX2 U4425 ( .A(fifo[448]), .Y(n4456) );
  INVX1 U4426 ( .A(n4459), .Y(n4457) );
  INVX1 U4427 ( .A(n4457), .Y(n4458) );
  BUFX2 U4428 ( .A(fifo[449]), .Y(n4459) );
  INVX1 U4429 ( .A(n4462), .Y(n4460) );
  INVX1 U4430 ( .A(n4460), .Y(n4461) );
  BUFX2 U4431 ( .A(fifo[450]), .Y(n4462) );
  INVX1 U4432 ( .A(n4465), .Y(n4463) );
  INVX1 U4433 ( .A(n4463), .Y(n4464) );
  BUFX2 U4434 ( .A(fifo[451]), .Y(n4465) );
  INVX1 U4435 ( .A(n4468), .Y(n4466) );
  INVX1 U4436 ( .A(n4466), .Y(n4467) );
  BUFX2 U4437 ( .A(fifo[452]), .Y(n4468) );
  INVX1 U4438 ( .A(n4471), .Y(n4469) );
  INVX1 U4439 ( .A(n4469), .Y(n4470) );
  BUFX2 U4440 ( .A(fifo[453]), .Y(n4471) );
  INVX1 U4441 ( .A(n4474), .Y(n4472) );
  INVX1 U4442 ( .A(n4472), .Y(n4473) );
  BUFX2 U4443 ( .A(fifo[454]), .Y(n4474) );
  INVX1 U4444 ( .A(n4477), .Y(n4475) );
  INVX1 U4445 ( .A(n4475), .Y(n4476) );
  BUFX2 U4446 ( .A(fifo[455]), .Y(n4477) );
  INVX1 U4447 ( .A(n4480), .Y(n4478) );
  INVX1 U4448 ( .A(n4478), .Y(n4479) );
  BUFX2 U4449 ( .A(fifo[456]), .Y(n4480) );
  INVX1 U4450 ( .A(n4483), .Y(n4481) );
  INVX1 U4451 ( .A(n4481), .Y(n4482) );
  BUFX2 U4452 ( .A(fifo[457]), .Y(n4483) );
  INVX1 U4453 ( .A(n4486), .Y(n4484) );
  INVX1 U4454 ( .A(n4484), .Y(n4485) );
  BUFX2 U4455 ( .A(fifo[458]), .Y(n4486) );
  INVX1 U4456 ( .A(n4489), .Y(n4487) );
  INVX1 U4457 ( .A(n4487), .Y(n4488) );
  BUFX2 U4458 ( .A(fifo[459]), .Y(n4489) );
  INVX1 U4459 ( .A(n4492), .Y(n4490) );
  INVX1 U4460 ( .A(n4490), .Y(n4491) );
  BUFX2 U4461 ( .A(fifo[460]), .Y(n4492) );
  INVX1 U4462 ( .A(n4495), .Y(n4493) );
  INVX1 U4463 ( .A(n4493), .Y(n4494) );
  BUFX2 U4464 ( .A(fifo[461]), .Y(n4495) );
  INVX1 U4465 ( .A(n4498), .Y(n4496) );
  INVX1 U4466 ( .A(n4496), .Y(n4497) );
  BUFX2 U4467 ( .A(fifo[462]), .Y(n4498) );
  INVX1 U4468 ( .A(n4501), .Y(n4499) );
  INVX1 U4469 ( .A(n4499), .Y(n4500) );
  BUFX2 U4470 ( .A(fifo[463]), .Y(n4501) );
  INVX1 U4471 ( .A(n4504), .Y(n4502) );
  INVX1 U4472 ( .A(n4502), .Y(n4503) );
  BUFX2 U4473 ( .A(fifo[416]), .Y(n4504) );
  INVX1 U4474 ( .A(n4507), .Y(n4505) );
  INVX1 U4475 ( .A(n4505), .Y(n4506) );
  BUFX2 U4476 ( .A(fifo[417]), .Y(n4507) );
  INVX1 U4477 ( .A(n4510), .Y(n4508) );
  INVX1 U4478 ( .A(n4508), .Y(n4509) );
  BUFX2 U4479 ( .A(fifo[418]), .Y(n4510) );
  INVX1 U4480 ( .A(n4513), .Y(n4511) );
  INVX1 U4481 ( .A(n4511), .Y(n4512) );
  BUFX2 U4482 ( .A(fifo[419]), .Y(n4513) );
  INVX1 U4483 ( .A(n4516), .Y(n4514) );
  INVX1 U4484 ( .A(n4514), .Y(n4515) );
  BUFX2 U4485 ( .A(fifo[420]), .Y(n4516) );
  INVX1 U4486 ( .A(n4519), .Y(n4517) );
  INVX1 U4487 ( .A(n4517), .Y(n4518) );
  BUFX2 U4488 ( .A(fifo[421]), .Y(n4519) );
  INVX1 U4489 ( .A(n4522), .Y(n4520) );
  INVX1 U4490 ( .A(n4520), .Y(n4521) );
  BUFX2 U4491 ( .A(fifo[422]), .Y(n4522) );
  INVX1 U4492 ( .A(n4525), .Y(n4523) );
  INVX1 U4493 ( .A(n4523), .Y(n4524) );
  BUFX2 U4494 ( .A(fifo[423]), .Y(n4525) );
  INVX1 U4495 ( .A(n4528), .Y(n4526) );
  INVX1 U4496 ( .A(n4526), .Y(n4527) );
  BUFX2 U4497 ( .A(fifo[424]), .Y(n4528) );
  INVX1 U4498 ( .A(n4531), .Y(n4529) );
  INVX1 U4499 ( .A(n4529), .Y(n4530) );
  BUFX2 U4500 ( .A(fifo[425]), .Y(n4531) );
  INVX1 U4501 ( .A(n4534), .Y(n4532) );
  INVX1 U4502 ( .A(n4532), .Y(n4533) );
  BUFX2 U4503 ( .A(fifo[426]), .Y(n4534) );
  INVX1 U4504 ( .A(n4537), .Y(n4535) );
  INVX1 U4505 ( .A(n4535), .Y(n4536) );
  BUFX2 U4506 ( .A(fifo[427]), .Y(n4537) );
  INVX1 U4507 ( .A(n4540), .Y(n4538) );
  INVX1 U4508 ( .A(n4538), .Y(n4539) );
  BUFX2 U4509 ( .A(fifo[428]), .Y(n4540) );
  INVX1 U4510 ( .A(n4543), .Y(n4541) );
  INVX1 U4511 ( .A(n4541), .Y(n4542) );
  BUFX2 U4512 ( .A(fifo[429]), .Y(n4543) );
  INVX1 U4513 ( .A(n4546), .Y(n4544) );
  INVX1 U4514 ( .A(n4544), .Y(n4545) );
  BUFX2 U4515 ( .A(fifo[430]), .Y(n4546) );
  INVX1 U4516 ( .A(n4549), .Y(n4547) );
  INVX1 U4517 ( .A(n4547), .Y(n4548) );
  BUFX2 U4518 ( .A(fifo[431]), .Y(n4549) );
  INVX1 U4519 ( .A(n4552), .Y(n4550) );
  INVX1 U4520 ( .A(n4550), .Y(n4551) );
  BUFX2 U4521 ( .A(fifo[384]), .Y(n4552) );
  INVX1 U4522 ( .A(n4555), .Y(n4553) );
  INVX1 U4523 ( .A(n4553), .Y(n4554) );
  BUFX2 U4524 ( .A(fifo[385]), .Y(n4555) );
  INVX1 U4525 ( .A(n4558), .Y(n4556) );
  INVX1 U4526 ( .A(n4556), .Y(n4557) );
  BUFX2 U4527 ( .A(fifo[386]), .Y(n4558) );
  INVX1 U4528 ( .A(n4561), .Y(n4559) );
  INVX1 U4529 ( .A(n4559), .Y(n4560) );
  BUFX2 U4530 ( .A(fifo[387]), .Y(n4561) );
  INVX1 U4531 ( .A(n4564), .Y(n4562) );
  INVX1 U4532 ( .A(n4562), .Y(n4563) );
  BUFX2 U4533 ( .A(fifo[388]), .Y(n4564) );
  INVX1 U4534 ( .A(n4567), .Y(n4565) );
  INVX1 U4535 ( .A(n4565), .Y(n4566) );
  BUFX2 U4536 ( .A(fifo[389]), .Y(n4567) );
  INVX1 U4537 ( .A(n4570), .Y(n4568) );
  INVX1 U4538 ( .A(n4568), .Y(n4569) );
  BUFX2 U4539 ( .A(fifo[390]), .Y(n4570) );
  INVX1 U4540 ( .A(n4573), .Y(n4571) );
  INVX1 U4541 ( .A(n4571), .Y(n4572) );
  BUFX2 U4542 ( .A(fifo[391]), .Y(n4573) );
  INVX1 U4543 ( .A(n4576), .Y(n4574) );
  INVX1 U4544 ( .A(n4574), .Y(n4575) );
  BUFX2 U4545 ( .A(fifo[392]), .Y(n4576) );
  INVX1 U4546 ( .A(n4579), .Y(n4577) );
  INVX1 U4547 ( .A(n4577), .Y(n4578) );
  BUFX2 U4548 ( .A(fifo[393]), .Y(n4579) );
  INVX1 U4549 ( .A(n4582), .Y(n4580) );
  INVX1 U4550 ( .A(n4580), .Y(n4581) );
  BUFX2 U4551 ( .A(fifo[394]), .Y(n4582) );
  INVX1 U4552 ( .A(n4585), .Y(n4583) );
  INVX1 U4553 ( .A(n4583), .Y(n4584) );
  BUFX2 U4554 ( .A(fifo[395]), .Y(n4585) );
  INVX1 U4555 ( .A(n4588), .Y(n4586) );
  INVX1 U4556 ( .A(n4586), .Y(n4587) );
  BUFX2 U4557 ( .A(fifo[396]), .Y(n4588) );
  INVX1 U4558 ( .A(n4591), .Y(n4589) );
  INVX1 U4559 ( .A(n4589), .Y(n4590) );
  BUFX2 U4560 ( .A(fifo[397]), .Y(n4591) );
  INVX1 U4561 ( .A(n4594), .Y(n4592) );
  INVX1 U4562 ( .A(n4592), .Y(n4593) );
  BUFX2 U4563 ( .A(fifo[398]), .Y(n4594) );
  INVX1 U4564 ( .A(n4597), .Y(n4595) );
  INVX1 U4565 ( .A(n4595), .Y(n4596) );
  BUFX2 U4566 ( .A(fifo[399]), .Y(n4597) );
  INVX1 U4567 ( .A(rd_ptr_gray_ss[2]), .Y(n5272) );
  INVX1 U4568 ( .A(rd_ptr_gray_ss[1]), .Y(n5273) );
  BUFX2 U4569 ( .A(n11), .Y(n4598) );
  INVX1 U4570 ( .A(n4598), .Y(n5297) );
  BUFX2 U4571 ( .A(n10), .Y(n4599) );
  INVX1 U4572 ( .A(n4599), .Y(n5322) );
  INVX1 U4573 ( .A(rd_ptr_gray_ss[5]), .Y(n4600) );
  INVX1 U4574 ( .A(n4600), .Y(n4601) );
  INVX1 U4575 ( .A(n4604), .Y(n4602) );
  INVX1 U4576 ( .A(n4602), .Y(n4603) );
  AND2X2 U4577 ( .A(n4633), .B(n206), .Y(n708) );
  INVX1 U4578 ( .A(n708), .Y(n4604) );
  INVX1 U4579 ( .A(n4607), .Y(n4605) );
  INVX1 U4580 ( .A(n4605), .Y(n4606) );
  AND2X1 U4581 ( .A(n4636), .B(n208), .Y(n743) );
  INVX1 U4582 ( .A(n743), .Y(n4607) );
  INVX1 U4583 ( .A(n4610), .Y(n4608) );
  INVX1 U4584 ( .A(n4608), .Y(n4609) );
  BUFX2 U4585 ( .A(wr_ptr_gray_ss[5]), .Y(n4610) );
  INVX1 U4586 ( .A(n4613), .Y(n4611) );
  INVX1 U4587 ( .A(n4611), .Y(n4612) );
  OR2X2 U4588 ( .A(n4606), .B(n210), .Y(n342) );
  INVX1 U4589 ( .A(n342), .Y(n4613) );
  INVX1 U4590 ( .A(n4616), .Y(n4614) );
  INVX1 U4591 ( .A(n4614), .Y(n4615) );
  OR2X2 U4592 ( .A(n4606), .B(n4645), .Y(n324) );
  INVX1 U4593 ( .A(n324), .Y(n4616) );
  INVX1 U4594 ( .A(n4619), .Y(n4617) );
  INVX1 U4595 ( .A(n4617), .Y(n4618) );
  OR2X2 U4596 ( .A(n4603), .B(n210), .Y(n306) );
  INVX1 U4597 ( .A(n306), .Y(n4619) );
  INVX1 U4598 ( .A(n4622), .Y(n4620) );
  INVX1 U4599 ( .A(n4620), .Y(n4621) );
  OR2X2 U4600 ( .A(n4603), .B(n4646), .Y(n288) );
  INVX1 U4601 ( .A(n288), .Y(n4622) );
  INVX1 U4602 ( .A(n4625), .Y(n4623) );
  INVX1 U4603 ( .A(n4623), .Y(n4624) );
  BUFX2 U4604 ( .A(wr_ptr_gray_ss[1]), .Y(n4625) );
  INVX1 U4605 ( .A(n4628), .Y(n4626) );
  INVX1 U4606 ( .A(n4626), .Y(n4627) );
  BUFX2 U4607 ( .A(rd_ptr_bin_5_), .Y(n4628) );
  INVX1 U4608 ( .A(n4631), .Y(n4629) );
  INVX1 U4609 ( .A(n4629), .Y(n4630) );
  BUFX2 U4610 ( .A(wr_ptr_bin[5]), .Y(n4631) );
  INVX1 U4611 ( .A(n4634), .Y(n4632) );
  INVX2 U4612 ( .A(n4632), .Y(n4633) );
  BUFX2 U4613 ( .A(wr_ptr_bin[1]), .Y(n4634) );
  INVX1 U4614 ( .A(n4637), .Y(n4635) );
  INVX1 U4615 ( .A(n4635), .Y(n4636) );
  BUFX2 U4616 ( .A(wr_ptr_bin[2]), .Y(n4637) );
  INVX1 U4617 ( .A(n4640), .Y(n4638) );
  INVX1 U4618 ( .A(n4638), .Y(n4639) );
  BUFX2 U4619 ( .A(wr_ptr_bin[4]), .Y(n4640) );
  INVX1 U4620 ( .A(n4643), .Y(n4641) );
  INVX1 U4621 ( .A(n4641), .Y(n4642) );
  BUFX2 U4622 ( .A(wr_ptr_bin[3]), .Y(n4643) );
  INVX1 U4623 ( .A(n4647), .Y(n4644) );
  INVX1 U4624 ( .A(n4644), .Y(n4645) );
  INVX1 U4625 ( .A(n4644), .Y(n4646) );
  BUFX2 U4626 ( .A(wr_ptr_bin[0]), .Y(n4647) );
  INVX1 U4627 ( .A(n4650), .Y(n4648) );
  INVX1 U4628 ( .A(n4648), .Y(n4649) );
  AND2X2 U4629 ( .A(re), .B(empty_bar), .Y(n185) );
  INVX1 U4630 ( .A(n185), .Y(n4650) );
  INVX1 U4631 ( .A(n4653), .Y(n4651) );
  INVX1 U4632 ( .A(n4651), .Y(n4652) );
  BUFX2 U4633 ( .A(n14), .Y(n4653) );
  INVX1 U4634 ( .A(n4656), .Y(n4654) );
  INVX2 U4635 ( .A(n4654), .Y(n4655) );
  AND2X1 U4636 ( .A(n251), .B(n252), .Y(n218) );
  INVX1 U4637 ( .A(n218), .Y(n4656) );
  INVX1 U4638 ( .A(n4659), .Y(n4657) );
  INVX2 U4639 ( .A(n4657), .Y(n4658) );
  AND2X1 U4640 ( .A(n673), .B(n378), .Y(n778) );
  INVX1 U4641 ( .A(n778), .Y(n4659) );
  INVX1 U4642 ( .A(n4662), .Y(n4660) );
  INVX2 U4643 ( .A(n4660), .Y(n4661) );
  INVX1 U4644 ( .A(n761), .Y(n4662) );
  INVX1 U4645 ( .A(n4665), .Y(n4663) );
  INVX2 U4646 ( .A(n4663), .Y(n4664) );
  INVX1 U4647 ( .A(n744), .Y(n4665) );
  INVX1 U4648 ( .A(n4668), .Y(n4666) );
  INVX2 U4649 ( .A(n4666), .Y(n4667) );
  INVX1 U4650 ( .A(n726), .Y(n4668) );
  INVX1 U4651 ( .A(n4671), .Y(n4669) );
  INVX2 U4652 ( .A(n4669), .Y(n4670) );
  INVX1 U4653 ( .A(n709), .Y(n4671) );
  INVX1 U4654 ( .A(n4674), .Y(n4672) );
  INVX2 U4655 ( .A(n4672), .Y(n4673) );
  INVX1 U4656 ( .A(n691), .Y(n4674) );
  INVX1 U4657 ( .A(n4677), .Y(n4675) );
  INVX2 U4658 ( .A(n4675), .Y(n4676) );
  INVX1 U4659 ( .A(n674), .Y(n4677) );
  INVX1 U4660 ( .A(n4680), .Y(n4678) );
  INVX2 U4661 ( .A(n4678), .Y(n4679) );
  INVX1 U4662 ( .A(n656), .Y(n4680) );
  INVX1 U4663 ( .A(n4683), .Y(n4681) );
  INVX2 U4664 ( .A(n4681), .Y(n4682) );
  AND2X1 U4665 ( .A(n535), .B(n378), .Y(n638) );
  INVX1 U4666 ( .A(n638), .Y(n4683) );
  INVX1 U4667 ( .A(n4686), .Y(n4684) );
  INVX2 U4668 ( .A(n4684), .Y(n4685) );
  INVX1 U4669 ( .A(n621), .Y(n4686) );
  INVX1 U4670 ( .A(n4689), .Y(n4687) );
  INVX2 U4671 ( .A(n4687), .Y(n4688) );
  INVX1 U4672 ( .A(n604), .Y(n4689) );
  INVX1 U4673 ( .A(n4692), .Y(n4690) );
  INVX2 U4674 ( .A(n4690), .Y(n4691) );
  INVX1 U4675 ( .A(n587), .Y(n4692) );
  INVX1 U4676 ( .A(n4695), .Y(n4693) );
  INVX2 U4677 ( .A(n4693), .Y(n4694) );
  INVX1 U4678 ( .A(n570), .Y(n4695) );
  INVX1 U4679 ( .A(n4698), .Y(n4696) );
  INVX2 U4680 ( .A(n4696), .Y(n4697) );
  INVX1 U4681 ( .A(n553), .Y(n4698) );
  INVX1 U4682 ( .A(n4701), .Y(n4699) );
  INVX2 U4683 ( .A(n4699), .Y(n4700) );
  INVX1 U4684 ( .A(n536), .Y(n4701) );
  INVX1 U4685 ( .A(n4704), .Y(n4702) );
  INVX2 U4686 ( .A(n4702), .Y(n4703) );
  INVX1 U4687 ( .A(n518), .Y(n4704) );
  INVX1 U4688 ( .A(n4707), .Y(n4705) );
  INVX2 U4689 ( .A(n4705), .Y(n4706) );
  AND2X1 U4690 ( .A(n397), .B(n378), .Y(n500) );
  INVX1 U4691 ( .A(n500), .Y(n4707) );
  INVX1 U4692 ( .A(n4710), .Y(n4708) );
  INVX2 U4693 ( .A(n4708), .Y(n4709) );
  INVX1 U4694 ( .A(n483), .Y(n4710) );
  INVX1 U4695 ( .A(n4713), .Y(n4711) );
  INVX2 U4696 ( .A(n4711), .Y(n4712) );
  INVX1 U4697 ( .A(n466), .Y(n4713) );
  INVX1 U4698 ( .A(n4716), .Y(n4714) );
  INVX2 U4699 ( .A(n4714), .Y(n4715) );
  INVX1 U4700 ( .A(n449), .Y(n4716) );
  INVX1 U4701 ( .A(n4719), .Y(n4717) );
  INVX2 U4702 ( .A(n4717), .Y(n4718) );
  INVX1 U4703 ( .A(n432), .Y(n4719) );
  INVX1 U4704 ( .A(n4722), .Y(n4720) );
  INVX2 U4705 ( .A(n4720), .Y(n4721) );
  INVX1 U4706 ( .A(n415), .Y(n4722) );
  INVX1 U4707 ( .A(n4725), .Y(n4723) );
  INVX2 U4708 ( .A(n4723), .Y(n4724) );
  INVX1 U4709 ( .A(n398), .Y(n4725) );
  INVX1 U4710 ( .A(n4728), .Y(n4726) );
  INVX2 U4711 ( .A(n4726), .Y(n4727) );
  INVX1 U4712 ( .A(n380), .Y(n4728) );
  INVX1 U4713 ( .A(n4731), .Y(n4729) );
  INVX2 U4714 ( .A(n4729), .Y(n4730) );
  AND2X1 U4715 ( .A(n378), .B(n252), .Y(n361) );
  INVX1 U4716 ( .A(n361), .Y(n4731) );
  INVX1 U4717 ( .A(n4734), .Y(n4732) );
  INVX2 U4718 ( .A(n4732), .Y(n4733) );
  INVX1 U4719 ( .A(n343), .Y(n4734) );
  INVX1 U4720 ( .A(n4737), .Y(n4735) );
  INVX2 U4721 ( .A(n4735), .Y(n4736) );
  INVX1 U4722 ( .A(n325), .Y(n4737) );
  INVX1 U4723 ( .A(n4740), .Y(n4738) );
  INVX2 U4724 ( .A(n4738), .Y(n4739) );
  INVX1 U4725 ( .A(n307), .Y(n4740) );
  INVX1 U4726 ( .A(n4743), .Y(n4741) );
  INVX2 U4727 ( .A(n4741), .Y(n4742) );
  INVX1 U4728 ( .A(n289), .Y(n4743) );
  INVX1 U4729 ( .A(n4746), .Y(n4744) );
  INVX2 U4730 ( .A(n4744), .Y(n4745) );
  INVX1 U4731 ( .A(n271), .Y(n4746) );
  INVX1 U4732 ( .A(n4749), .Y(n4747) );
  INVX2 U4733 ( .A(n4747), .Y(n4748) );
  INVX1 U4734 ( .A(n253), .Y(n4749) );
  INVX1 U4735 ( .A(n4752), .Y(n4750) );
  INVX1 U4736 ( .A(n4750), .Y(n4751) );
  BUFX2 U4737 ( .A(n13), .Y(n4752) );
  INVX1 U4738 ( .A(n1416), .Y(n4753) );
  INVX8 U4739 ( .A(n4753), .Y(n4754) );
  INVX8 U4740 ( .A(n4753), .Y(n4755) );
  XNOR2X1 U5256 ( .A(n3045), .B(rd_ptr_bin_ss[1]), .Y(n5271) );
  INVX1 U5257 ( .A(n5271), .Y(rd_ptr_bin_ss[0]) );
  XNOR2X1 U5258 ( .A(rd_ptr_bin_ss[3]), .B(n5272), .Y(rd_ptr_bin_ss[2]) );
  XNOR2X1 U5259 ( .A(rd_ptr_bin_ss[2]), .B(n5273), .Y(rd_ptr_bin_ss[1]) );
  INVX1 U5260 ( .A(n12), .Y(n5274) );
  INVX8 U5261 ( .A(n5274), .Y(n5275) );
  INVX8 U5262 ( .A(n5284), .Y(n5276) );
  INVX8 U5263 ( .A(n5284), .Y(n5277) );
  INVX8 U5264 ( .A(n5284), .Y(n5278) );
  INVX8 U5265 ( .A(n5283), .Y(n5279) );
  INVX8 U5266 ( .A(n5282), .Y(n5280) );
  INVX8 U5267 ( .A(n5282), .Y(n5281) );
  INVX8 U5268 ( .A(n4754), .Y(n5282) );
  INVX8 U5269 ( .A(n4755), .Y(n5283) );
  INVX8 U5270 ( .A(n4754), .Y(n5284) );
  INVX8 U5271 ( .A(n5295), .Y(n5285) );
  INVX8 U5272 ( .A(n5295), .Y(n5286) );
  INVX8 U5273 ( .A(n5294), .Y(n5287) );
  INVX8 U5274 ( .A(n5294), .Y(n5288) );
  INVX8 U5275 ( .A(n5294), .Y(n5289) );
  INVX8 U5276 ( .A(n5293), .Y(n5290) );
  INVX8 U5277 ( .A(n5293), .Y(n5291) );
  INVX8 U5278 ( .A(n5293), .Y(n5292) );
  INVX8 U5279 ( .A(n5296), .Y(n5293) );
  INVX8 U5280 ( .A(n5296), .Y(n5294) );
  INVX8 U5281 ( .A(n5296), .Y(n5295) );
  INVX8 U5282 ( .A(n5297), .Y(n5296) );
  INVX8 U5283 ( .A(n5314), .Y(n5298) );
  INVX8 U5284 ( .A(n5314), .Y(n5299) );
  INVX8 U5285 ( .A(n5314), .Y(n5300) );
  INVX8 U5286 ( .A(n5315), .Y(n5301) );
  INVX8 U5287 ( .A(n5315), .Y(n5302) );
  INVX8 U5288 ( .A(n5315), .Y(n5303) );
  INVX8 U5289 ( .A(n5316), .Y(n5304) );
  INVX8 U5290 ( .A(n5316), .Y(n5305) );
  INVX8 U5291 ( .A(n5317), .Y(n5306) );
  INVX8 U5292 ( .A(n5317), .Y(n5307) );
  INVX8 U5293 ( .A(n5317), .Y(n5308) );
  INVX8 U5294 ( .A(n5318), .Y(n5309) );
  INVX8 U5295 ( .A(n5318), .Y(n5310) );
  INVX8 U5296 ( .A(n5318), .Y(n5311) );
  INVX8 U5297 ( .A(n5319), .Y(n5312) );
  INVX8 U5298 ( .A(n5316), .Y(n5313) );
  INVX8 U5299 ( .A(n5321), .Y(n5314) );
  INVX8 U5300 ( .A(n5321), .Y(n5315) );
  INVX8 U5301 ( .A(n5321), .Y(n5316) );
  INVX8 U5302 ( .A(n5320), .Y(n5317) );
  INVX8 U5303 ( .A(n5320), .Y(n5318) );
  INVX8 U5304 ( .A(n5320), .Y(n5319) );
  INVX8 U5305 ( .A(n5322), .Y(n5320) );
  INVX8 U5306 ( .A(n5322), .Y(n5321) );
  MUX2X1 U5307 ( .B(n5324), .A(n5325), .S(n5292), .Y(n5323) );
  MUX2X1 U5308 ( .B(n5327), .A(n5328), .S(n5292), .Y(n5326) );
  MUX2X1 U5309 ( .B(n5330), .A(n5331), .S(n5292), .Y(n5329) );
  MUX2X1 U5310 ( .B(n5333), .A(n5334), .S(n5292), .Y(n5332) );
  MUX2X1 U5311 ( .B(n5336), .A(n5337), .S(n4751), .Y(n5335) );
  MUX2X1 U5312 ( .B(n5339), .A(n5340), .S(n5292), .Y(n5338) );
  MUX2X1 U5313 ( .B(n5342), .A(n5343), .S(n5292), .Y(n5341) );
  MUX2X1 U5314 ( .B(n5345), .A(n5346), .S(n5292), .Y(n5344) );
  MUX2X1 U5315 ( .B(n5348), .A(n5349), .S(n5292), .Y(n5347) );
  MUX2X1 U5316 ( .B(n5351), .A(n5352), .S(n4751), .Y(n5350) );
  MUX2X1 U5317 ( .B(n5354), .A(n5355), .S(n5292), .Y(n5353) );
  MUX2X1 U5318 ( .B(n5357), .A(n5358), .S(n5292), .Y(n5356) );
  MUX2X1 U5319 ( .B(n5360), .A(n5361), .S(n5292), .Y(n5359) );
  MUX2X1 U5320 ( .B(n5363), .A(n5364), .S(n5292), .Y(n5362) );
  MUX2X1 U5321 ( .B(n5366), .A(n5367), .S(n4751), .Y(n5365) );
  MUX2X1 U5322 ( .B(n5369), .A(n5370), .S(n5292), .Y(n5368) );
  MUX2X1 U5323 ( .B(n5372), .A(n5373), .S(n5292), .Y(n5371) );
  MUX2X1 U5324 ( .B(n5375), .A(n5376), .S(n5291), .Y(n5374) );
  MUX2X1 U5325 ( .B(n5378), .A(n5379), .S(n5291), .Y(n5377) );
  MUX2X1 U5326 ( .B(n5381), .A(n5382), .S(n4751), .Y(n5380) );
  MUX2X1 U5327 ( .B(n5384), .A(n5385), .S(n5291), .Y(n5383) );
  MUX2X1 U5328 ( .B(n5387), .A(n5388), .S(n5291), .Y(n5386) );
  MUX2X1 U5329 ( .B(n5390), .A(n5391), .S(n5291), .Y(n5389) );
  MUX2X1 U5330 ( .B(n5393), .A(n5394), .S(n5291), .Y(n5392) );
  MUX2X1 U5331 ( .B(n5396), .A(n5397), .S(n4751), .Y(n5395) );
  MUX2X1 U5332 ( .B(n5399), .A(n5400), .S(n5291), .Y(n5398) );
  MUX2X1 U5333 ( .B(n5402), .A(n5403), .S(n5291), .Y(n5401) );
  MUX2X1 U5334 ( .B(n5405), .A(n5406), .S(n5291), .Y(n5404) );
  MUX2X1 U5335 ( .B(n5408), .A(n5409), .S(n5291), .Y(n5407) );
  MUX2X1 U5336 ( .B(n5411), .A(n5412), .S(n4751), .Y(n5410) );
  MUX2X1 U5337 ( .B(n5414), .A(n5415), .S(n5291), .Y(n5413) );
  MUX2X1 U5338 ( .B(n5417), .A(n5418), .S(n5291), .Y(n5416) );
  MUX2X1 U5339 ( .B(n5420), .A(n5421), .S(n5291), .Y(n5419) );
  MUX2X1 U5340 ( .B(n5423), .A(n5424), .S(n5291), .Y(n5422) );
  MUX2X1 U5341 ( .B(n5426), .A(n5427), .S(n4751), .Y(n5425) );
  MUX2X1 U5342 ( .B(n5429), .A(n5430), .S(n5291), .Y(n5428) );
  MUX2X1 U5343 ( .B(n5432), .A(n5433), .S(n5291), .Y(n5431) );
  MUX2X1 U5344 ( .B(n5435), .A(n5436), .S(n5291), .Y(n5434) );
  MUX2X1 U5345 ( .B(n5438), .A(n5439), .S(n5290), .Y(n5437) );
  MUX2X1 U5346 ( .B(n5441), .A(n5442), .S(n4751), .Y(n5440) );
  MUX2X1 U5347 ( .B(n5444), .A(n5445), .S(n5290), .Y(n5443) );
  MUX2X1 U5348 ( .B(n5447), .A(n5448), .S(n5290), .Y(n5446) );
  MUX2X1 U5349 ( .B(n5450), .A(n5451), .S(n5290), .Y(n5449) );
  MUX2X1 U5350 ( .B(n5453), .A(n5454), .S(n5290), .Y(n5452) );
  MUX2X1 U5351 ( .B(n5456), .A(n5457), .S(n4751), .Y(n5455) );
  MUX2X1 U5352 ( .B(n5459), .A(n5460), .S(n5290), .Y(n5458) );
  MUX2X1 U5353 ( .B(n5462), .A(n5463), .S(n5290), .Y(n5461) );
  MUX2X1 U5354 ( .B(n5465), .A(n5466), .S(n5290), .Y(n5464) );
  MUX2X1 U5355 ( .B(n5468), .A(n5469), .S(n5290), .Y(n5467) );
  MUX2X1 U5356 ( .B(n5471), .A(n5472), .S(n4751), .Y(n5470) );
  MUX2X1 U5357 ( .B(n5474), .A(n5475), .S(n5290), .Y(n5473) );
  MUX2X1 U5358 ( .B(n5477), .A(n5478), .S(n5290), .Y(n5476) );
  MUX2X1 U5359 ( .B(n5480), .A(n5481), .S(n5290), .Y(n5479) );
  MUX2X1 U5360 ( .B(n5483), .A(n5484), .S(n5290), .Y(n5482) );
  MUX2X1 U5361 ( .B(n5486), .A(n5487), .S(n4751), .Y(n5485) );
  MUX2X1 U5362 ( .B(n5489), .A(n5490), .S(n5290), .Y(n5488) );
  MUX2X1 U5363 ( .B(n5492), .A(n5493), .S(n5290), .Y(n5491) );
  MUX2X1 U5364 ( .B(n5495), .A(n5496), .S(n5290), .Y(n5494) );
  MUX2X1 U5365 ( .B(n5498), .A(n5499), .S(n5290), .Y(n5497) );
  MUX2X1 U5366 ( .B(n5501), .A(n5502), .S(n4751), .Y(n5500) );
  MUX2X1 U5367 ( .B(n5504), .A(n5505), .S(n5289), .Y(n5503) );
  MUX2X1 U5368 ( .B(n5507), .A(n5508), .S(n5289), .Y(n5506) );
  MUX2X1 U5369 ( .B(n5510), .A(n5511), .S(n5289), .Y(n5509) );
  MUX2X1 U5370 ( .B(n5513), .A(n5514), .S(n5289), .Y(n5512) );
  MUX2X1 U5371 ( .B(n5516), .A(n5517), .S(n4751), .Y(n5515) );
  MUX2X1 U5372 ( .B(n5519), .A(n5520), .S(n5289), .Y(n5518) );
  MUX2X1 U5373 ( .B(n5522), .A(n5523), .S(n5289), .Y(n5521) );
  MUX2X1 U5374 ( .B(n5525), .A(n5526), .S(n5289), .Y(n5524) );
  MUX2X1 U5375 ( .B(n5528), .A(n5529), .S(n5289), .Y(n5527) );
  MUX2X1 U5376 ( .B(n5531), .A(n5532), .S(n4751), .Y(n5530) );
  MUX2X1 U5377 ( .B(n5534), .A(n5535), .S(n5289), .Y(n5533) );
  MUX2X1 U5378 ( .B(n5537), .A(n5538), .S(n5289), .Y(n5536) );
  MUX2X1 U5379 ( .B(n5540), .A(n5541), .S(n5289), .Y(n5539) );
  MUX2X1 U5380 ( .B(n5543), .A(n5544), .S(n5289), .Y(n5542) );
  MUX2X1 U5381 ( .B(n5546), .A(n5547), .S(n4751), .Y(n5545) );
  MUX2X1 U5382 ( .B(n5549), .A(n5550), .S(n5289), .Y(n5548) );
  MUX2X1 U5383 ( .B(n5552), .A(n5553), .S(n5289), .Y(n5551) );
  MUX2X1 U5384 ( .B(n5555), .A(n5556), .S(n5289), .Y(n5554) );
  MUX2X1 U5385 ( .B(n5558), .A(n5559), .S(n5289), .Y(n5557) );
  MUX2X1 U5386 ( .B(n5561), .A(n5562), .S(n4751), .Y(n5560) );
  MUX2X1 U5387 ( .B(n5564), .A(n5565), .S(n5289), .Y(n5563) );
  MUX2X1 U5388 ( .B(n5567), .A(n5568), .S(n5288), .Y(n5566) );
  MUX2X1 U5389 ( .B(n5570), .A(n5571), .S(n5288), .Y(n5569) );
  MUX2X1 U5390 ( .B(n5573), .A(n5574), .S(n5288), .Y(n5572) );
  MUX2X1 U5391 ( .B(n5576), .A(n5577), .S(n4751), .Y(n5575) );
  MUX2X1 U5392 ( .B(n5579), .A(n5580), .S(n5288), .Y(n5578) );
  MUX2X1 U5393 ( .B(n5582), .A(n5583), .S(n5288), .Y(n5581) );
  MUX2X1 U5394 ( .B(n5585), .A(n5586), .S(n5288), .Y(n5584) );
  MUX2X1 U5395 ( .B(n5588), .A(n5589), .S(n5288), .Y(n5587) );
  MUX2X1 U5396 ( .B(n5591), .A(n5592), .S(n4751), .Y(n5590) );
  MUX2X1 U5397 ( .B(n5594), .A(n5595), .S(n5288), .Y(n5593) );
  MUX2X1 U5398 ( .B(n5597), .A(n5598), .S(n5288), .Y(n5596) );
  MUX2X1 U5399 ( .B(n5600), .A(n5601), .S(n5288), .Y(n5599) );
  MUX2X1 U5400 ( .B(n5603), .A(n5604), .S(n5288), .Y(n5602) );
  MUX2X1 U5401 ( .B(n5606), .A(n5607), .S(n4751), .Y(n5605) );
  MUX2X1 U5402 ( .B(n5609), .A(n5610), .S(n5288), .Y(n5608) );
  MUX2X1 U5403 ( .B(n5612), .A(n5613), .S(n5288), .Y(n5611) );
  MUX2X1 U5404 ( .B(n5615), .A(n5616), .S(n5288), .Y(n5614) );
  MUX2X1 U5405 ( .B(n5618), .A(n5619), .S(n5288), .Y(n5617) );
  MUX2X1 U5406 ( .B(n5621), .A(n5622), .S(n4751), .Y(n5620) );
  MUX2X1 U5407 ( .B(n5624), .A(n5625), .S(n5288), .Y(n5623) );
  MUX2X1 U5408 ( .B(n5627), .A(n5628), .S(n5288), .Y(n5626) );
  MUX2X1 U5409 ( .B(n5630), .A(n5631), .S(n5287), .Y(n5629) );
  MUX2X1 U5410 ( .B(n5633), .A(n5634), .S(n5287), .Y(n5632) );
  MUX2X1 U5411 ( .B(n5636), .A(n5637), .S(n4751), .Y(n5635) );
  MUX2X1 U5412 ( .B(n5639), .A(n5640), .S(n5287), .Y(n5638) );
  MUX2X1 U5413 ( .B(n5642), .A(n5643), .S(n5287), .Y(n5641) );
  MUX2X1 U5414 ( .B(n5645), .A(n5646), .S(n5287), .Y(n5644) );
  MUX2X1 U5415 ( .B(n5648), .A(n5649), .S(n5287), .Y(n5647) );
  MUX2X1 U5416 ( .B(n5651), .A(n5652), .S(n4751), .Y(n5650) );
  MUX2X1 U5417 ( .B(n5654), .A(n5655), .S(n5287), .Y(n5653) );
  MUX2X1 U5418 ( .B(n5657), .A(n5658), .S(n5287), .Y(n5656) );
  MUX2X1 U5419 ( .B(n5660), .A(n5661), .S(n5287), .Y(n5659) );
  MUX2X1 U5420 ( .B(n5663), .A(n5664), .S(n5287), .Y(n5662) );
  MUX2X1 U5421 ( .B(n5666), .A(n5667), .S(n4751), .Y(n5665) );
  MUX2X1 U5422 ( .B(n5669), .A(n5670), .S(n5287), .Y(n5668) );
  MUX2X1 U5423 ( .B(n5672), .A(n5673), .S(n5287), .Y(n5671) );
  MUX2X1 U5424 ( .B(n5675), .A(n5676), .S(n5287), .Y(n5674) );
  MUX2X1 U5425 ( .B(n5678), .A(n5679), .S(n5287), .Y(n5677) );
  MUX2X1 U5426 ( .B(n5681), .A(n5682), .S(n4751), .Y(n5680) );
  MUX2X1 U5427 ( .B(n5684), .A(n5685), .S(n5287), .Y(n5683) );
  MUX2X1 U5428 ( .B(n5687), .A(n5688), .S(n5287), .Y(n5686) );
  MUX2X1 U5429 ( .B(n5690), .A(n5691), .S(n5287), .Y(n5689) );
  MUX2X1 U5430 ( .B(n5693), .A(n5694), .S(n5286), .Y(n5692) );
  MUX2X1 U5431 ( .B(n5696), .A(n5697), .S(n4751), .Y(n5695) );
  MUX2X1 U5432 ( .B(n5699), .A(n5700), .S(n5286), .Y(n5698) );
  MUX2X1 U5433 ( .B(n5702), .A(n5703), .S(n5286), .Y(n5701) );
  MUX2X1 U5434 ( .B(n5705), .A(n5706), .S(n5286), .Y(n5704) );
  MUX2X1 U5435 ( .B(n5708), .A(n5709), .S(n5286), .Y(n5707) );
  MUX2X1 U5436 ( .B(n5711), .A(n5712), .S(n4751), .Y(n5710) );
  MUX2X1 U5437 ( .B(n5714), .A(n5715), .S(n5286), .Y(n5713) );
  MUX2X1 U5438 ( .B(n5717), .A(n5718), .S(n5286), .Y(n5716) );
  MUX2X1 U5439 ( .B(n5720), .A(n5721), .S(n5286), .Y(n5719) );
  MUX2X1 U5440 ( .B(n5723), .A(n5724), .S(n5286), .Y(n5722) );
  MUX2X1 U5441 ( .B(n5726), .A(n5727), .S(n4751), .Y(n5725) );
  MUX2X1 U5442 ( .B(n5729), .A(n5730), .S(n5286), .Y(n5728) );
  MUX2X1 U5443 ( .B(n5732), .A(n5733), .S(n5286), .Y(n5731) );
  MUX2X1 U5444 ( .B(n5735), .A(n5736), .S(n5286), .Y(n5734) );
  MUX2X1 U5445 ( .B(n5738), .A(n5739), .S(n5286), .Y(n5737) );
  MUX2X1 U5446 ( .B(n5741), .A(n5742), .S(n4751), .Y(n5740) );
  MUX2X1 U5447 ( .B(n5744), .A(n5745), .S(n5286), .Y(n5743) );
  MUX2X1 U5448 ( .B(n5747), .A(n5748), .S(n5286), .Y(n5746) );
  MUX2X1 U5449 ( .B(n5750), .A(n5751), .S(n5286), .Y(n5749) );
  MUX2X1 U5450 ( .B(n5753), .A(n5754), .S(n5286), .Y(n5752) );
  MUX2X1 U5451 ( .B(n5756), .A(n5757), .S(n4751), .Y(n5755) );
  MUX2X1 U5452 ( .B(n5759), .A(n5760), .S(n5285), .Y(n5758) );
  MUX2X1 U5453 ( .B(n5762), .A(n5763), .S(n5285), .Y(n5761) );
  MUX2X1 U5454 ( .B(n5765), .A(n5766), .S(n5285), .Y(n5764) );
  MUX2X1 U5455 ( .B(n5768), .A(n5769), .S(n5285), .Y(n5767) );
  MUX2X1 U5456 ( .B(n5771), .A(n5772), .S(n4751), .Y(n5770) );
  MUX2X1 U5457 ( .B(n5774), .A(n5775), .S(n5285), .Y(n5773) );
  MUX2X1 U5458 ( .B(n5777), .A(n5778), .S(n5285), .Y(n5776) );
  MUX2X1 U5459 ( .B(n5780), .A(n5781), .S(n5285), .Y(n5779) );
  MUX2X1 U5460 ( .B(n5783), .A(n5784), .S(n5285), .Y(n5782) );
  MUX2X1 U5461 ( .B(n5786), .A(n5787), .S(n4751), .Y(n5785) );
  MUX2X1 U5462 ( .B(n5789), .A(n5790), .S(n5285), .Y(n5788) );
  MUX2X1 U5463 ( .B(n5792), .A(n5793), .S(n5285), .Y(n5791) );
  MUX2X1 U5464 ( .B(n5795), .A(n5796), .S(n5285), .Y(n5794) );
  MUX2X1 U5465 ( .B(n5798), .A(n5799), .S(n5285), .Y(n5797) );
  MUX2X1 U5466 ( .B(n5801), .A(n5802), .S(n4751), .Y(n5800) );
  MUX2X1 U5467 ( .B(n3543), .A(n4311), .S(n5298), .Y(n5325) );
  MUX2X1 U5468 ( .B(n3495), .A(n4263), .S(n5309), .Y(n5324) );
  MUX2X1 U5469 ( .B(n3447), .A(n4215), .S(n5305), .Y(n5328) );
  MUX2X1 U5470 ( .B(n3591), .A(n4359), .S(n5305), .Y(n5327) );
  MUX2X1 U5471 ( .B(n5326), .A(n5323), .S(n5275), .Y(n5337) );
  MUX2X1 U5472 ( .B(n3255), .A(n4023), .S(n5305), .Y(n5331) );
  MUX2X1 U5473 ( .B(n3111), .A(n3879), .S(n5305), .Y(n5330) );
  MUX2X1 U5474 ( .B(n3063), .A(n3831), .S(n5305), .Y(n5334) );
  MUX2X1 U5475 ( .B(n3351), .A(n4119), .S(n5306), .Y(n5333) );
  MUX2X1 U5476 ( .B(n5332), .A(n5329), .S(n5275), .Y(n5336) );
  MUX2X1 U5477 ( .B(n3303), .A(n4071), .S(n5306), .Y(n5340) );
  MUX2X1 U5478 ( .B(n3207), .A(n3975), .S(n5306), .Y(n5339) );
  MUX2X1 U5479 ( .B(n3159), .A(n3927), .S(n5306), .Y(n5343) );
  MUX2X1 U5480 ( .B(n3399), .A(n4167), .S(n5306), .Y(n5342) );
  MUX2X1 U5481 ( .B(n5341), .A(n5338), .S(n5275), .Y(n5352) );
  MUX2X1 U5482 ( .B(n3735), .A(n4551), .S(n5306), .Y(n5346) );
  MUX2X1 U5483 ( .B(n3687), .A(n4503), .S(n5306), .Y(n5345) );
  MUX2X1 U5484 ( .B(n3639), .A(n4455), .S(n5306), .Y(n5349) );
  MUX2X1 U5485 ( .B(n3783), .A(n4407), .S(n5306), .Y(n5348) );
  MUX2X1 U5486 ( .B(n5347), .A(n5344), .S(n5275), .Y(n5351) );
  MUX2X1 U5487 ( .B(n5350), .A(n5335), .S(n4652), .Y(n5803) );
  INVX2 U5488 ( .A(n5803), .Y(n86) );
  MUX2X1 U5489 ( .B(n3546), .A(n4314), .S(n5306), .Y(n5355) );
  MUX2X1 U5490 ( .B(n3498), .A(n4266), .S(n5306), .Y(n5354) );
  MUX2X1 U5491 ( .B(n3450), .A(n4218), .S(n5306), .Y(n5358) );
  MUX2X1 U5492 ( .B(n3594), .A(n4362), .S(n5306), .Y(n5357) );
  MUX2X1 U5493 ( .B(n5356), .A(n5353), .S(n5275), .Y(n5367) );
  MUX2X1 U5494 ( .B(n3258), .A(n4026), .S(n5306), .Y(n5361) );
  MUX2X1 U5495 ( .B(n3114), .A(n3882), .S(n5306), .Y(n5360) );
  MUX2X1 U5496 ( .B(n3066), .A(n3834), .S(n5306), .Y(n5364) );
  MUX2X1 U5497 ( .B(n3354), .A(n4122), .S(n5306), .Y(n5363) );
  MUX2X1 U5498 ( .B(n5362), .A(n5359), .S(n5275), .Y(n5366) );
  MUX2X1 U5499 ( .B(n3306), .A(n4074), .S(n5307), .Y(n5370) );
  MUX2X1 U5500 ( .B(n3210), .A(n3978), .S(n5307), .Y(n5369) );
  MUX2X1 U5501 ( .B(n3162), .A(n3930), .S(n5307), .Y(n5373) );
  MUX2X1 U5502 ( .B(n3402), .A(n4170), .S(n5307), .Y(n5372) );
  MUX2X1 U5503 ( .B(n5371), .A(n5368), .S(n5275), .Y(n5382) );
  MUX2X1 U5504 ( .B(n3738), .A(n4554), .S(n5307), .Y(n5376) );
  MUX2X1 U5505 ( .B(n3690), .A(n4506), .S(n5307), .Y(n5375) );
  MUX2X1 U5506 ( .B(n3642), .A(n4458), .S(n5307), .Y(n5379) );
  MUX2X1 U5507 ( .B(n3786), .A(n4410), .S(n5307), .Y(n5378) );
  MUX2X1 U5508 ( .B(n5377), .A(n5374), .S(n5275), .Y(n5381) );
  MUX2X1 U5509 ( .B(n5380), .A(n5365), .S(n4652), .Y(n5804) );
  MUX2X1 U5510 ( .B(n3549), .A(n4317), .S(n5307), .Y(n5385) );
  MUX2X1 U5511 ( .B(n3501), .A(n4269), .S(n5307), .Y(n5384) );
  MUX2X1 U5512 ( .B(n3453), .A(n4221), .S(n5307), .Y(n5388) );
  MUX2X1 U5513 ( .B(n3597), .A(n4365), .S(n5307), .Y(n5387) );
  MUX2X1 U5514 ( .B(n5386), .A(n5383), .S(n5275), .Y(n5397) );
  MUX2X1 U5515 ( .B(n3261), .A(n4029), .S(n5307), .Y(n5391) );
  MUX2X1 U5516 ( .B(n3117), .A(n3885), .S(n5307), .Y(n5390) );
  MUX2X1 U5517 ( .B(n3069), .A(n3837), .S(n5307), .Y(n5394) );
  MUX2X1 U5518 ( .B(n3357), .A(n4125), .S(n5307), .Y(n5393) );
  MUX2X1 U5519 ( .B(n5392), .A(n5389), .S(n5275), .Y(n5396) );
  MUX2X1 U5520 ( .B(n3309), .A(n4077), .S(n5307), .Y(n5400) );
  MUX2X1 U5521 ( .B(n3213), .A(n3981), .S(n5308), .Y(n5399) );
  MUX2X1 U5522 ( .B(n3165), .A(n3933), .S(n5308), .Y(n5403) );
  MUX2X1 U5523 ( .B(n3405), .A(n4173), .S(n5308), .Y(n5402) );
  MUX2X1 U5524 ( .B(n5401), .A(n5398), .S(n5275), .Y(n5412) );
  MUX2X1 U5525 ( .B(n3741), .A(n4557), .S(n5308), .Y(n5406) );
  MUX2X1 U5526 ( .B(n3693), .A(n4509), .S(n5308), .Y(n5405) );
  MUX2X1 U5527 ( .B(n3645), .A(n4461), .S(n5308), .Y(n5409) );
  MUX2X1 U5528 ( .B(n3789), .A(n4413), .S(n5308), .Y(n5408) );
  MUX2X1 U5529 ( .B(n5407), .A(n5404), .S(n5275), .Y(n5411) );
  MUX2X1 U5530 ( .B(n5410), .A(n5395), .S(n4652), .Y(n5805) );
  INVX2 U5531 ( .A(n5805), .Y(n84) );
  MUX2X1 U5532 ( .B(n3552), .A(n4320), .S(n5308), .Y(n5415) );
  MUX2X1 U5533 ( .B(n3504), .A(n4272), .S(n5308), .Y(n5414) );
  MUX2X1 U5534 ( .B(n3456), .A(n4224), .S(n5308), .Y(n5418) );
  MUX2X1 U5535 ( .B(n3600), .A(n4368), .S(n5308), .Y(n5417) );
  MUX2X1 U5536 ( .B(n5416), .A(n5413), .S(n5275), .Y(n5427) );
  MUX2X1 U5537 ( .B(n3264), .A(n4032), .S(n5308), .Y(n5421) );
  MUX2X1 U5538 ( .B(n3120), .A(n3888), .S(n5308), .Y(n5420) );
  MUX2X1 U5539 ( .B(n3072), .A(n3840), .S(n5308), .Y(n5424) );
  MUX2X1 U5540 ( .B(n3360), .A(n4128), .S(n5308), .Y(n5423) );
  MUX2X1 U5541 ( .B(n5422), .A(n5419), .S(n5275), .Y(n5426) );
  MUX2X1 U5542 ( .B(n3312), .A(n4080), .S(n5308), .Y(n5430) );
  MUX2X1 U5543 ( .B(n3216), .A(n3984), .S(n5308), .Y(n5429) );
  MUX2X1 U5544 ( .B(n3168), .A(n3936), .S(n5309), .Y(n5433) );
  MUX2X1 U5545 ( .B(n3408), .A(n4176), .S(n5309), .Y(n5432) );
  MUX2X1 U5546 ( .B(n5431), .A(n5428), .S(n5275), .Y(n5442) );
  MUX2X1 U5547 ( .B(n3744), .A(n4560), .S(n5309), .Y(n5436) );
  MUX2X1 U5548 ( .B(n3696), .A(n4512), .S(n5309), .Y(n5435) );
  MUX2X1 U5549 ( .B(n3648), .A(n4464), .S(n5309), .Y(n5439) );
  MUX2X1 U5550 ( .B(n3792), .A(n4416), .S(n5309), .Y(n5438) );
  MUX2X1 U5551 ( .B(n5437), .A(n5434), .S(n5275), .Y(n5441) );
  MUX2X1 U5552 ( .B(n5440), .A(n5425), .S(n4652), .Y(n5806) );
  INVX2 U5553 ( .A(n5806), .Y(n83) );
  MUX2X1 U5554 ( .B(n3555), .A(n4323), .S(n5309), .Y(n5445) );
  MUX2X1 U5555 ( .B(n3507), .A(n4275), .S(n5309), .Y(n5444) );
  MUX2X1 U5556 ( .B(n3459), .A(n4227), .S(n5309), .Y(n5448) );
  MUX2X1 U5557 ( .B(n3603), .A(n4371), .S(n5309), .Y(n5447) );
  MUX2X1 U5558 ( .B(n5446), .A(n5443), .S(n5275), .Y(n5457) );
  MUX2X1 U5559 ( .B(n3267), .A(n4035), .S(n5309), .Y(n5451) );
  MUX2X1 U5560 ( .B(n3123), .A(n3891), .S(n5309), .Y(n5450) );
  MUX2X1 U5561 ( .B(n3075), .A(n3843), .S(n5309), .Y(n5454) );
  MUX2X1 U5562 ( .B(n3363), .A(n4131), .S(n5309), .Y(n5453) );
  MUX2X1 U5563 ( .B(n5452), .A(n5449), .S(n5275), .Y(n5456) );
  MUX2X1 U5564 ( .B(n3315), .A(n4083), .S(n5309), .Y(n5460) );
  MUX2X1 U5565 ( .B(n3219), .A(n3987), .S(n5309), .Y(n5459) );
  MUX2X1 U5566 ( .B(n3171), .A(n3939), .S(n5310), .Y(n5463) );
  MUX2X1 U5567 ( .B(n3411), .A(n4179), .S(n5310), .Y(n5462) );
  MUX2X1 U5568 ( .B(n5461), .A(n5458), .S(n5275), .Y(n5472) );
  MUX2X1 U5569 ( .B(n3747), .A(n4563), .S(n5310), .Y(n5466) );
  MUX2X1 U5570 ( .B(n3699), .A(n4515), .S(n5310), .Y(n5465) );
  MUX2X1 U5571 ( .B(n3651), .A(n4467), .S(n5310), .Y(n5469) );
  MUX2X1 U5572 ( .B(n3795), .A(n4419), .S(n5310), .Y(n5468) );
  MUX2X1 U5573 ( .B(n5467), .A(n5464), .S(n5275), .Y(n5471) );
  MUX2X1 U5574 ( .B(n5470), .A(n5455), .S(n4652), .Y(n5807) );
  MUX2X1 U5575 ( .B(n3558), .A(n4326), .S(n5310), .Y(n5475) );
  MUX2X1 U5576 ( .B(n3510), .A(n4278), .S(n5310), .Y(n5474) );
  MUX2X1 U5577 ( .B(n3462), .A(n4230), .S(n5310), .Y(n5478) );
  MUX2X1 U5578 ( .B(n3606), .A(n4374), .S(n5310), .Y(n5477) );
  MUX2X1 U5579 ( .B(n5476), .A(n5473), .S(n5275), .Y(n5487) );
  MUX2X1 U5580 ( .B(n3270), .A(n4038), .S(n5310), .Y(n5481) );
  MUX2X1 U5581 ( .B(n3126), .A(n3894), .S(n5310), .Y(n5480) );
  MUX2X1 U5582 ( .B(n3078), .A(n3846), .S(n5310), .Y(n5484) );
  MUX2X1 U5583 ( .B(n3366), .A(n4134), .S(n5310), .Y(n5483) );
  MUX2X1 U5584 ( .B(n5482), .A(n5479), .S(n5275), .Y(n5486) );
  MUX2X1 U5585 ( .B(n3318), .A(n4086), .S(n5310), .Y(n5490) );
  MUX2X1 U5586 ( .B(n3222), .A(n3990), .S(n5310), .Y(n5489) );
  MUX2X1 U5587 ( .B(n3174), .A(n3942), .S(n5310), .Y(n5493) );
  MUX2X1 U5588 ( .B(n3414), .A(n4182), .S(n5311), .Y(n5492) );
  MUX2X1 U5589 ( .B(n5491), .A(n5488), .S(n5275), .Y(n5502) );
  MUX2X1 U5590 ( .B(n3750), .A(n4566), .S(n5311), .Y(n5496) );
  MUX2X1 U5591 ( .B(n3702), .A(n4518), .S(n5311), .Y(n5495) );
  MUX2X1 U5592 ( .B(n3654), .A(n4470), .S(n5311), .Y(n5499) );
  MUX2X1 U5593 ( .B(n3798), .A(n4422), .S(n5311), .Y(n5498) );
  MUX2X1 U5594 ( .B(n5497), .A(n5494), .S(n5275), .Y(n5501) );
  MUX2X1 U5595 ( .B(n5500), .A(n5485), .S(n4652), .Y(n5808) );
  INVX2 U5596 ( .A(n5808), .Y(n81) );
  MUX2X1 U5597 ( .B(n3561), .A(n4329), .S(n5311), .Y(n5505) );
  MUX2X1 U5598 ( .B(n3513), .A(n4281), .S(n5311), .Y(n5504) );
  MUX2X1 U5599 ( .B(n3465), .A(n4233), .S(n5311), .Y(n5508) );
  MUX2X1 U5600 ( .B(n3609), .A(n4377), .S(n5311), .Y(n5507) );
  MUX2X1 U5601 ( .B(n5506), .A(n5503), .S(n5275), .Y(n5517) );
  MUX2X1 U5602 ( .B(n3273), .A(n4041), .S(n5311), .Y(n5511) );
  MUX2X1 U5603 ( .B(n3129), .A(n3897), .S(n5311), .Y(n5510) );
  MUX2X1 U5604 ( .B(n3081), .A(n3849), .S(n5311), .Y(n5514) );
  MUX2X1 U5605 ( .B(n3369), .A(n4137), .S(n5311), .Y(n5513) );
  MUX2X1 U5606 ( .B(n5512), .A(n5509), .S(n5275), .Y(n5516) );
  MUX2X1 U5607 ( .B(n3321), .A(n4089), .S(n5311), .Y(n5520) );
  MUX2X1 U5608 ( .B(n3225), .A(n3993), .S(n5311), .Y(n5519) );
  MUX2X1 U5609 ( .B(n3177), .A(n3945), .S(n5311), .Y(n5523) );
  MUX2X1 U5610 ( .B(n3417), .A(n4185), .S(n5311), .Y(n5522) );
  MUX2X1 U5611 ( .B(n5521), .A(n5518), .S(n5275), .Y(n5532) );
  MUX2X1 U5612 ( .B(n3753), .A(n4569), .S(n5312), .Y(n5526) );
  MUX2X1 U5613 ( .B(n3705), .A(n4521), .S(n5312), .Y(n5525) );
  MUX2X1 U5614 ( .B(n3657), .A(n4473), .S(n5312), .Y(n5529) );
  MUX2X1 U5615 ( .B(n3801), .A(n4425), .S(n5312), .Y(n5528) );
  MUX2X1 U5616 ( .B(n5527), .A(n5524), .S(n5275), .Y(n5531) );
  MUX2X1 U5617 ( .B(n5530), .A(n5515), .S(n4652), .Y(n5809) );
  INVX2 U5618 ( .A(n5809), .Y(n80) );
  MUX2X1 U5619 ( .B(n3564), .A(n4332), .S(n5312), .Y(n5535) );
  MUX2X1 U5620 ( .B(n3516), .A(n4284), .S(n5312), .Y(n5534) );
  MUX2X1 U5621 ( .B(n3468), .A(n4236), .S(n5312), .Y(n5538) );
  MUX2X1 U5622 ( .B(n3612), .A(n4380), .S(n5312), .Y(n5537) );
  MUX2X1 U5623 ( .B(n5536), .A(n5533), .S(n5275), .Y(n5547) );
  MUX2X1 U5624 ( .B(n3276), .A(n4044), .S(n5312), .Y(n5541) );
  MUX2X1 U5625 ( .B(n3132), .A(n3900), .S(n5312), .Y(n5540) );
  MUX2X1 U5626 ( .B(n3084), .A(n3852), .S(n5312), .Y(n5544) );
  MUX2X1 U5627 ( .B(n3372), .A(n4140), .S(n5312), .Y(n5543) );
  MUX2X1 U5628 ( .B(n5542), .A(n5539), .S(n5275), .Y(n5546) );
  MUX2X1 U5629 ( .B(n3324), .A(n4092), .S(n5312), .Y(n5550) );
  MUX2X1 U5630 ( .B(n3228), .A(n3996), .S(n5312), .Y(n5549) );
  MUX2X1 U5631 ( .B(n3180), .A(n3948), .S(n5312), .Y(n5553) );
  MUX2X1 U5632 ( .B(n3420), .A(n4188), .S(n5312), .Y(n5552) );
  MUX2X1 U5633 ( .B(n5551), .A(n5548), .S(n5275), .Y(n5562) );
  MUX2X1 U5634 ( .B(n3756), .A(n4572), .S(n5312), .Y(n5556) );
  MUX2X1 U5635 ( .B(n3708), .A(n4524), .S(n5313), .Y(n5555) );
  MUX2X1 U5636 ( .B(n3660), .A(n4476), .S(n5313), .Y(n5559) );
  MUX2X1 U5637 ( .B(n3804), .A(n4428), .S(n5313), .Y(n5558) );
  MUX2X1 U5638 ( .B(n5557), .A(n5554), .S(n5275), .Y(n5561) );
  MUX2X1 U5639 ( .B(n5560), .A(n5545), .S(n4652), .Y(n5810) );
  MUX2X1 U5640 ( .B(n3567), .A(n4335), .S(n5313), .Y(n5565) );
  MUX2X1 U5641 ( .B(n3519), .A(n4287), .S(n5301), .Y(n5564) );
  MUX2X1 U5642 ( .B(n3471), .A(n4239), .S(n5298), .Y(n5568) );
  MUX2X1 U5643 ( .B(n3615), .A(n4383), .S(n5298), .Y(n5567) );
  MUX2X1 U5644 ( .B(n5566), .A(n5563), .S(n5275), .Y(n5577) );
  MUX2X1 U5645 ( .B(n3279), .A(n4047), .S(n5298), .Y(n5571) );
  MUX2X1 U5646 ( .B(n3135), .A(n3903), .S(n5298), .Y(n5570) );
  MUX2X1 U5647 ( .B(n3087), .A(n3855), .S(n5298), .Y(n5574) );
  MUX2X1 U5648 ( .B(n3375), .A(n4143), .S(n5298), .Y(n5573) );
  MUX2X1 U5649 ( .B(n5572), .A(n5569), .S(n5275), .Y(n5576) );
  MUX2X1 U5650 ( .B(n3327), .A(n4095), .S(n5298), .Y(n5580) );
  MUX2X1 U5651 ( .B(n3231), .A(n3999), .S(n5298), .Y(n5579) );
  MUX2X1 U5652 ( .B(n3183), .A(n3951), .S(n5298), .Y(n5583) );
  MUX2X1 U5653 ( .B(n3423), .A(n4191), .S(n5298), .Y(n5582) );
  MUX2X1 U5654 ( .B(n5581), .A(n5578), .S(n5275), .Y(n5592) );
  MUX2X1 U5655 ( .B(n3759), .A(n4575), .S(n5298), .Y(n5586) );
  MUX2X1 U5656 ( .B(n3711), .A(n4527), .S(n5298), .Y(n5585) );
  MUX2X1 U5657 ( .B(n3663), .A(n4479), .S(n5298), .Y(n5589) );
  MUX2X1 U5658 ( .B(n3807), .A(n4431), .S(n5299), .Y(n5588) );
  MUX2X1 U5659 ( .B(n5587), .A(n5584), .S(n5275), .Y(n5591) );
  MUX2X1 U5660 ( .B(n5590), .A(n5575), .S(n4652), .Y(n5811) );
  INVX2 U5661 ( .A(n5811), .Y(n78) );
  MUX2X1 U5662 ( .B(n3570), .A(n4338), .S(n5299), .Y(n5595) );
  MUX2X1 U5663 ( .B(n3522), .A(n4290), .S(n5299), .Y(n5594) );
  MUX2X1 U5664 ( .B(n3474), .A(n4242), .S(n5299), .Y(n5598) );
  MUX2X1 U5665 ( .B(n3618), .A(n4386), .S(n5299), .Y(n5597) );
  MUX2X1 U5666 ( .B(n5596), .A(n5593), .S(n5275), .Y(n5607) );
  MUX2X1 U5667 ( .B(n3282), .A(n4050), .S(n5299), .Y(n5601) );
  MUX2X1 U5668 ( .B(n3138), .A(n3906), .S(n5299), .Y(n5600) );
  MUX2X1 U5669 ( .B(n3090), .A(n3858), .S(n5299), .Y(n5604) );
  MUX2X1 U5670 ( .B(n3378), .A(n4146), .S(n5299), .Y(n5603) );
  MUX2X1 U5671 ( .B(n5602), .A(n5599), .S(n5275), .Y(n5606) );
  MUX2X1 U5672 ( .B(n3330), .A(n4098), .S(n5299), .Y(n5610) );
  MUX2X1 U5673 ( .B(n3234), .A(n4002), .S(n5299), .Y(n5609) );
  MUX2X1 U5674 ( .B(n3186), .A(n3954), .S(n5299), .Y(n5613) );
  MUX2X1 U5675 ( .B(n3426), .A(n4194), .S(n5299), .Y(n5612) );
  MUX2X1 U5676 ( .B(n5611), .A(n5608), .S(n5275), .Y(n5622) );
  MUX2X1 U5677 ( .B(n3762), .A(n4578), .S(n5299), .Y(n5616) );
  MUX2X1 U5678 ( .B(n3714), .A(n4530), .S(n5299), .Y(n5615) );
  MUX2X1 U5679 ( .B(n3666), .A(n4482), .S(n5299), .Y(n5619) );
  MUX2X1 U5680 ( .B(n3810), .A(n4434), .S(n5299), .Y(n5618) );
  MUX2X1 U5681 ( .B(n5617), .A(n5614), .S(n5275), .Y(n5621) );
  MUX2X1 U5682 ( .B(n5620), .A(n5605), .S(n4652), .Y(n5812) );
  INVX2 U5683 ( .A(n5812), .Y(n77) );
  MUX2X1 U5684 ( .B(n3573), .A(n4341), .S(n5300), .Y(n5625) );
  MUX2X1 U5685 ( .B(n3525), .A(n4293), .S(n5300), .Y(n5624) );
  MUX2X1 U5686 ( .B(n3477), .A(n4245), .S(n5300), .Y(n5628) );
  MUX2X1 U5687 ( .B(n3621), .A(n4389), .S(n5300), .Y(n5627) );
  MUX2X1 U5688 ( .B(n5626), .A(n5623), .S(n5275), .Y(n5637) );
  MUX2X1 U5689 ( .B(n3285), .A(n4053), .S(n5300), .Y(n5631) );
  MUX2X1 U5690 ( .B(n3141), .A(n3909), .S(n5300), .Y(n5630) );
  MUX2X1 U5691 ( .B(n3093), .A(n3861), .S(n5300), .Y(n5634) );
  MUX2X1 U5692 ( .B(n3381), .A(n4149), .S(n5300), .Y(n5633) );
  MUX2X1 U5693 ( .B(n5632), .A(n5629), .S(n5275), .Y(n5636) );
  MUX2X1 U5694 ( .B(n3333), .A(n4101), .S(n5300), .Y(n5640) );
  MUX2X1 U5695 ( .B(n3237), .A(n4005), .S(n5300), .Y(n5639) );
  MUX2X1 U5696 ( .B(n3189), .A(n3957), .S(n5300), .Y(n5643) );
  MUX2X1 U5697 ( .B(n3429), .A(n4197), .S(n5300), .Y(n5642) );
  MUX2X1 U5698 ( .B(n5641), .A(n5638), .S(n5275), .Y(n5652) );
  MUX2X1 U5699 ( .B(n3765), .A(n4581), .S(n5300), .Y(n5646) );
  MUX2X1 U5700 ( .B(n3717), .A(n4533), .S(n5300), .Y(n5645) );
  MUX2X1 U5701 ( .B(n3669), .A(n4485), .S(n5300), .Y(n5649) );
  MUX2X1 U5702 ( .B(n3813), .A(n4437), .S(n5300), .Y(n5648) );
  MUX2X1 U5703 ( .B(n5647), .A(n5644), .S(n5275), .Y(n5651) );
  MUX2X1 U5704 ( .B(n5650), .A(n5635), .S(n4652), .Y(n5813) );
  MUX2X1 U5705 ( .B(n3576), .A(n4344), .S(n5300), .Y(n5655) );
  MUX2X1 U5706 ( .B(n3528), .A(n4296), .S(n5301), .Y(n5654) );
  MUX2X1 U5707 ( .B(n3480), .A(n4248), .S(n5301), .Y(n5658) );
  MUX2X1 U5708 ( .B(n3624), .A(n4392), .S(n5301), .Y(n5657) );
  MUX2X1 U5709 ( .B(n5656), .A(n5653), .S(n5275), .Y(n5667) );
  MUX2X1 U5710 ( .B(n3288), .A(n4056), .S(n5301), .Y(n5661) );
  MUX2X1 U5711 ( .B(n3144), .A(n3912), .S(n5301), .Y(n5660) );
  MUX2X1 U5712 ( .B(n3096), .A(n3864), .S(n5301), .Y(n5664) );
  MUX2X1 U5713 ( .B(n3384), .A(n4152), .S(n5301), .Y(n5663) );
  MUX2X1 U5714 ( .B(n5662), .A(n5659), .S(n5275), .Y(n5666) );
  MUX2X1 U5715 ( .B(n3336), .A(n4104), .S(n5301), .Y(n5670) );
  MUX2X1 U5716 ( .B(n3240), .A(n4008), .S(n5301), .Y(n5669) );
  MUX2X1 U5717 ( .B(n3192), .A(n3960), .S(n5301), .Y(n5673) );
  MUX2X1 U5718 ( .B(n3432), .A(n4200), .S(n5301), .Y(n5672) );
  MUX2X1 U5719 ( .B(n5671), .A(n5668), .S(n5275), .Y(n5682) );
  MUX2X1 U5720 ( .B(n3768), .A(n4584), .S(n5301), .Y(n5676) );
  MUX2X1 U5721 ( .B(n3720), .A(n4536), .S(n5301), .Y(n5675) );
  MUX2X1 U5722 ( .B(n3672), .A(n4488), .S(n5301), .Y(n5679) );
  MUX2X1 U5723 ( .B(n3816), .A(n4440), .S(n5301), .Y(n5678) );
  MUX2X1 U5724 ( .B(n5677), .A(n5674), .S(n5275), .Y(n5681) );
  MUX2X1 U5725 ( .B(n5680), .A(n5665), .S(n4652), .Y(n5814) );
  INVX2 U5726 ( .A(n5814), .Y(n75) );
  MUX2X1 U5727 ( .B(n3579), .A(n4347), .S(n5301), .Y(n5685) );
  MUX2X1 U5728 ( .B(n3531), .A(n4299), .S(n5302), .Y(n5684) );
  MUX2X1 U5729 ( .B(n3483), .A(n4251), .S(n5305), .Y(n5688) );
  MUX2X1 U5730 ( .B(n3627), .A(n4395), .S(n5302), .Y(n5687) );
  MUX2X1 U5731 ( .B(n5686), .A(n5683), .S(n5275), .Y(n5697) );
  MUX2X1 U5732 ( .B(n3291), .A(n4059), .S(n5302), .Y(n5691) );
  MUX2X1 U5733 ( .B(n3147), .A(n3915), .S(n5302), .Y(n5690) );
  MUX2X1 U5734 ( .B(n3099), .A(n3867), .S(n5302), .Y(n5694) );
  MUX2X1 U5735 ( .B(n3387), .A(n4155), .S(n5302), .Y(n5693) );
  MUX2X1 U5736 ( .B(n5692), .A(n5689), .S(n5275), .Y(n5696) );
  MUX2X1 U5737 ( .B(n3339), .A(n4107), .S(n5302), .Y(n5700) );
  MUX2X1 U5738 ( .B(n3243), .A(n4011), .S(n5302), .Y(n5699) );
  MUX2X1 U5739 ( .B(n3195), .A(n3963), .S(n5302), .Y(n5703) );
  MUX2X1 U5740 ( .B(n3435), .A(n4203), .S(n5302), .Y(n5702) );
  MUX2X1 U5741 ( .B(n5701), .A(n5698), .S(n5275), .Y(n5712) );
  MUX2X1 U5742 ( .B(n3771), .A(n4587), .S(n5302), .Y(n5706) );
  MUX2X1 U5743 ( .B(n3723), .A(n4539), .S(n5302), .Y(n5705) );
  MUX2X1 U5744 ( .B(n3675), .A(n4491), .S(n5302), .Y(n5709) );
  MUX2X1 U5745 ( .B(n3819), .A(n4443), .S(n5302), .Y(n5708) );
  MUX2X1 U5746 ( .B(n5707), .A(n5704), .S(n5275), .Y(n5711) );
  MUX2X1 U5747 ( .B(n5710), .A(n5695), .S(n4652), .Y(n5815) );
  INVX2 U5748 ( .A(n5815), .Y(n74) );
  MUX2X1 U5749 ( .B(n3582), .A(n4350), .S(n5302), .Y(n5715) );
  MUX2X1 U5750 ( .B(n3534), .A(n4302), .S(n5302), .Y(n5714) );
  MUX2X1 U5751 ( .B(n3486), .A(n4254), .S(n5302), .Y(n5718) );
  MUX2X1 U5752 ( .B(n3630), .A(n4398), .S(n5303), .Y(n5717) );
  MUX2X1 U5753 ( .B(n5716), .A(n5713), .S(n5275), .Y(n5727) );
  MUX2X1 U5754 ( .B(n3294), .A(n4062), .S(n5303), .Y(n5721) );
  MUX2X1 U5755 ( .B(n3150), .A(n3918), .S(n5303), .Y(n5720) );
  MUX2X1 U5756 ( .B(n3102), .A(n3870), .S(n5303), .Y(n5724) );
  MUX2X1 U5757 ( .B(n3390), .A(n4158), .S(n5303), .Y(n5723) );
  MUX2X1 U5758 ( .B(n5722), .A(n5719), .S(n5275), .Y(n5726) );
  MUX2X1 U5759 ( .B(n3342), .A(n4110), .S(n5303), .Y(n5730) );
  MUX2X1 U5760 ( .B(n3246), .A(n4014), .S(n5303), .Y(n5729) );
  MUX2X1 U5761 ( .B(n3198), .A(n3966), .S(n5303), .Y(n5733) );
  MUX2X1 U5762 ( .B(n3438), .A(n4206), .S(n5303), .Y(n5732) );
  MUX2X1 U5763 ( .B(n5731), .A(n5728), .S(n5275), .Y(n5742) );
  MUX2X1 U5764 ( .B(n3774), .A(n4590), .S(n5303), .Y(n5736) );
  MUX2X1 U5765 ( .B(n3726), .A(n4542), .S(n5303), .Y(n5735) );
  MUX2X1 U5766 ( .B(n3678), .A(n4494), .S(n5303), .Y(n5739) );
  MUX2X1 U5767 ( .B(n3822), .A(n4446), .S(n5303), .Y(n5738) );
  MUX2X1 U5768 ( .B(n5737), .A(n5734), .S(n5275), .Y(n5741) );
  MUX2X1 U5769 ( .B(n5740), .A(n5725), .S(n4652), .Y(n5816) );
  MUX2X1 U5770 ( .B(n3585), .A(n4353), .S(n5303), .Y(n5745) );
  MUX2X1 U5771 ( .B(n3537), .A(n4305), .S(n5303), .Y(n5744) );
  MUX2X1 U5772 ( .B(n3489), .A(n4257), .S(n5303), .Y(n5748) );
  MUX2X1 U5773 ( .B(n3633), .A(n4401), .S(n5303), .Y(n5747) );
  MUX2X1 U5774 ( .B(n5746), .A(n5743), .S(n5275), .Y(n5757) );
  MUX2X1 U5775 ( .B(n3297), .A(n4065), .S(n5304), .Y(n5751) );
  MUX2X1 U5776 ( .B(n3153), .A(n3921), .S(n5304), .Y(n5750) );
  MUX2X1 U5777 ( .B(n3105), .A(n3873), .S(n5304), .Y(n5754) );
  MUX2X1 U5778 ( .B(n3393), .A(n4161), .S(n5304), .Y(n5753) );
  MUX2X1 U5779 ( .B(n5752), .A(n5749), .S(n5275), .Y(n5756) );
  MUX2X1 U5780 ( .B(n3345), .A(n4113), .S(n5304), .Y(n5760) );
  MUX2X1 U5781 ( .B(n3249), .A(n4017), .S(n5304), .Y(n5759) );
  MUX2X1 U5782 ( .B(n3201), .A(n3969), .S(n5304), .Y(n5763) );
  MUX2X1 U5783 ( .B(n3441), .A(n4209), .S(n5304), .Y(n5762) );
  MUX2X1 U5784 ( .B(n5761), .A(n5758), .S(n5275), .Y(n5772) );
  MUX2X1 U5785 ( .B(n3777), .A(n4593), .S(n5304), .Y(n5766) );
  MUX2X1 U5786 ( .B(n3729), .A(n4545), .S(n5304), .Y(n5765) );
  MUX2X1 U5787 ( .B(n3681), .A(n4497), .S(n5304), .Y(n5769) );
  MUX2X1 U5788 ( .B(n3825), .A(n4449), .S(n5304), .Y(n5768) );
  MUX2X1 U5789 ( .B(n5767), .A(n5764), .S(n5275), .Y(n5771) );
  MUX2X1 U5790 ( .B(n5770), .A(n5755), .S(n4652), .Y(n5817) );
  INVX2 U5791 ( .A(n5817), .Y(n72) );
  MUX2X1 U5792 ( .B(n3588), .A(n4356), .S(n5304), .Y(n5775) );
  MUX2X1 U5793 ( .B(n3540), .A(n4308), .S(n5304), .Y(n5774) );
  MUX2X1 U5794 ( .B(n3492), .A(n4260), .S(n5304), .Y(n5778) );
  MUX2X1 U5795 ( .B(n3636), .A(n4404), .S(n5304), .Y(n5777) );
  MUX2X1 U5796 ( .B(n5776), .A(n5773), .S(n5275), .Y(n5787) );
  MUX2X1 U5797 ( .B(n3300), .A(n4068), .S(n5304), .Y(n5781) );
  MUX2X1 U5798 ( .B(n3156), .A(n3924), .S(n5305), .Y(n5780) );
  MUX2X1 U5799 ( .B(n3108), .A(n3876), .S(n5305), .Y(n5784) );
  MUX2X1 U5800 ( .B(n3396), .A(n4164), .S(n5305), .Y(n5783) );
  MUX2X1 U5801 ( .B(n5782), .A(n5779), .S(n5275), .Y(n5786) );
  MUX2X1 U5802 ( .B(n3348), .A(n4116), .S(n5305), .Y(n5790) );
  MUX2X1 U5803 ( .B(n3252), .A(n4020), .S(n5305), .Y(n5789) );
  MUX2X1 U5804 ( .B(n3204), .A(n3972), .S(n5305), .Y(n5793) );
  MUX2X1 U5805 ( .B(n3444), .A(n4212), .S(n5305), .Y(n5792) );
  MUX2X1 U5806 ( .B(n5791), .A(n5788), .S(n5275), .Y(n5802) );
  MUX2X1 U5807 ( .B(n3780), .A(n4596), .S(n5305), .Y(n5796) );
  MUX2X1 U5808 ( .B(n3732), .A(n4548), .S(n5305), .Y(n5795) );
  MUX2X1 U5809 ( .B(n3684), .A(n4500), .S(n5305), .Y(n5799) );
  MUX2X1 U5810 ( .B(n3828), .A(n4452), .S(n5305), .Y(n5798) );
  MUX2X1 U5811 ( .B(n5797), .A(n5794), .S(n5275), .Y(n5801) );
  MUX2X1 U5812 ( .B(n5800), .A(n5785), .S(n4652), .Y(n5818) );
  INVX1 U5813 ( .A(rd_ptr_bin_ss[0]), .Y(r301_B_not_0_) );
  INVX1 U5814 ( .A(rd_ptr_bin_ss[1]), .Y(r301_B_not_1_) );
  INVX1 U5815 ( .A(rd_ptr_bin_ss[2]), .Y(r301_B_not_2_) );
  INVX1 U5816 ( .A(rd_ptr_bin_ss[3]), .Y(r301_B_not_3_) );
  INVX1 U5817 ( .A(rd_ptr_bin_ss[4]), .Y(r301_B_not_4_) );
  INVX1 U5818 ( .A(n4601), .Y(r301_B_not_5_) );
  XNOR2X1 U5819 ( .A(r301_B_not_0_), .B(n4646), .Y(fillcount[0]) );
  INVX2 U5820 ( .A(n1), .Y(r301_carry[1]) );
  INVX1 U5821 ( .A(n4646), .Y(n33) );
  XOR2X1 U5822 ( .A(add_158_carry[5]), .B(n4630), .Y(n38) );
  XOR2X1 U5823 ( .A(add_176_carry[5]), .B(n4627), .Y(n92) );
endmodule


module FIFO_2clk_DATA_WIDTH34_FIFO_DEPTH32_PTR_WIDTH6 ( rclk, wclk, reset, we, 
        re, data_in, empty_bar, full_bar, data_out, fillcount );
  input [33:0] data_in;
  output [33:0] data_out;
  output [5:0] fillcount;
  input rclk, wclk, reset, we, re;
  output empty_bar, full_bar;
  wire   n10, n11, n12, n13, n14, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, rd_ptr_bin_5_, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n33, n34, n35, n36, n37,
         n38, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n106, n107, n108, n109, n110,
         n193, n194, n195, n196, n197, n199, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n2536, n2541, n2546, n2551, n2553, n2555, n2557, n2559,
         n2561, n2563, n2565, n2567, n2569, n2571, n2573, n2575, n2577, n2579,
         n2581, n2583, n2585, n2587, n2589, n2591, n2593, n2595, n2597, n2599,
         n2601, n2603, n2605, n2607, n2609, n2611, n2613, n2615, n2617, n2619,
         n2627, n2632, n2637, n2642, n2644, n2649, n2657, n2658, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, r301_B_not_0_,
         r301_B_not_1_, r301_B_not_2_, r301_B_not_3_, r301_B_not_4_,
         r301_B_not_5_, n1, n2, n3, n4, n5, n6, n7, n8, n25, n26, n27, n28,
         n29, n30, n31, n32, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n105, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n155, n156, n158, n159, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n198, n200,
         n252, n1141, n1431, n1432, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2535, n2540, n2545, n2550, n2552, n2558, n2560, n2562, n2564, n2566,
         n2568, n2570, n2572, n2574, n2576, n2578, n2580, n2582, n2584, n2586,
         n2588, n2590, n2592, n2594, n2596, n2598, n2600, n2602, n2604, n2606,
         n2608, n2610, n2612, n2614, n2616, n2618, n2620, n2645, n2656, n2659,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
         n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9969,
         n9970, n9972, n9973, n9975, n9976, n9978, n9979, n9981, n9982, n9984,
         n9985, n9987, n9988, n9990, n9991, n9993, n9994, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10005, n10006, n10008, n10009,
         n10011, n10012, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10029, n10030, n10031, n10032, n10033, n10035, n10036, n10038,
         n10039, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10051, n10052, n10054, n10056, n10058, n10059,
         n10061, n10062, n10064, n10065, n10067, n10068, n10070, n10071,
         n10073, n10074, n10076, n10077, n10079, n10080, n10081, n10082,
         n10083, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10485, n10486,
         n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494,
         n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
         n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510,
         n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518,
         n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526,
         n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534,
         n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542,
         n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550,
         n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558,
         n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
         n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574,
         n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582,
         n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590,
         n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598,
         n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606,
         n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614,
         n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
         n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630,
         n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638,
         n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646,
         n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654,
         n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662,
         n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670,
         n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678,
         n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686,
         n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694,
         n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702,
         n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710,
         n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718,
         n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726,
         n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734,
         n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742,
         n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750,
         n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758,
         n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766,
         n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774,
         n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782,
         n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790,
         n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798,
         n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806,
         n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814,
         n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822,
         n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830,
         n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838,
         n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846,
         n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854,
         n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862,
         n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870,
         n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878,
         n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886,
         n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894,
         n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902,
         n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910,
         n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
         n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926,
         n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
         n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942,
         n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950,
         n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958,
         n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
         n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974,
         n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982,
         n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990,
         n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
         n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
         n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
         n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022,
         n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030,
         n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
         n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046,
         n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054,
         n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
         n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
         n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
         n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
         n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094,
         n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
         n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
         n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
         n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126,
         n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134,
         n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
         n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
         n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158,
         n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
         n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174,
         n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182,
         n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190,
         n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198,
         n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206,
         n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214,
         n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222,
         n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230,
         n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238,
         n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246,
         n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254,
         n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262,
         n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270,
         n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278,
         n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286,
         n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294,
         n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302,
         n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310,
         n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318,
         n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326,
         n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334,
         n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
         n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
         n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
         n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
         n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374,
         n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382,
         n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390,
         n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398,
         n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406,
         n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414,
         n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422,
         n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430,
         n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438,
         n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446,
         n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454,
         n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462,
         n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470,
         n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478,
         n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486,
         n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494,
         n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502,
         n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510,
         n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518,
         n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526,
         n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534,
         n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542,
         n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550,
         n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558,
         n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566,
         n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
         n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582,
         n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590,
         n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598,
         n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606,
         n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614,
         n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622,
         n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630,
         n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638,
         n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
         n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654,
         n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662,
         n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670,
         n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678,
         n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686,
         n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694,
         n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702,
         n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710,
         n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718,
         n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726,
         n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734,
         n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742,
         n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750,
         n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758,
         n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766,
         n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774,
         n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782,
         n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790,
         n11791, n11792, n11793, n11794, n11795;
  wire   [5:0] wr_ptr_gray;
  wire   [5:0] wr_ptr_gray_ss;
  wire   [5:0] wr_ptr_gray_s;
  wire   [5:0] rd_ptr_gray;
  wire   [5:0] rd_ptr_gray_ss;
  wire   [5:0] rd_ptr_gray_s;
  wire   [4:0] rd_ptr_bin_ss;
  wire   [5:0] wr_ptr_bin;
  wire   [1087:0] fifo;
  wire   [5:2] add_176_carry;
  wire   [5:2] add_158_carry;
  wire   [4:2] r301_carry;

  DFFSR rd_ptr_gray_reg_5_ ( .D(n10047), .CLK(rclk), .R(n10539), .S(1'b1), .Q(
        rd_ptr_gray[5]) );
  DFFSR rd_ptr_gray_s_reg_5_ ( .D(n149), .CLK(wclk), .R(n10539), .S(1'b1), .Q(
        rd_ptr_gray_s[5]) );
  DFFSR rd_ptr_gray_ss_reg_5_ ( .D(n146), .CLK(wclk), .R(n10539), .S(1'b1), 
        .Q(rd_ptr_gray_ss[5]) );
  DFFSR rd_ptr_gray_reg_4_ ( .D(n15), .CLK(rclk), .R(n10539), .S(1'b1), .Q(
        rd_ptr_gray[4]) );
  DFFSR rd_ptr_gray_s_reg_4_ ( .D(n143), .CLK(wclk), .R(n10538), .S(1'b1), .Q(
        rd_ptr_gray_s[4]) );
  DFFSR rd_ptr_gray_ss_reg_4_ ( .D(n140), .CLK(wclk), .R(n10538), .S(1'b1), 
        .Q(rd_ptr_gray_ss[4]) );
  DFFSR wr_ptr_bin_reg_5_ ( .D(n2649), .CLK(wclk), .R(n10607), .S(1'b1), .Q(
        wr_ptr_bin[5]) );
  DFFSR wr_ptr_gray_reg_5_ ( .D(n10081), .CLK(wclk), .R(n10607), .S(1'b1), .Q(
        wr_ptr_gray[5]) );
  DFFSR wr_ptr_gray_s_reg_5_ ( .D(n137), .CLK(rclk), .R(n10607), .S(1'b1), .Q(
        wr_ptr_gray_s[5]) );
  DFFSR wr_ptr_bin_reg_0_ ( .D(n2644), .CLK(wclk), .R(n10608), .S(1'b1), .Q(
        wr_ptr_bin[0]) );
  DFFSR wr_ptr_bin_reg_1_ ( .D(n2642), .CLK(wclk), .R(n10608), .S(1'b1), .Q(
        wr_ptr_bin[1]) );
  DFFSR wr_ptr_gray_reg_0_ ( .D(n24), .CLK(wclk), .R(n10608), .S(1'b1), .Q(
        wr_ptr_gray[0]) );
  DFFSR wr_ptr_gray_s_reg_0_ ( .D(n131), .CLK(rclk), .R(n10608), .S(1'b1), .Q(
        wr_ptr_gray_s[0]) );
  DFFSR wr_ptr_gray_ss_reg_0_ ( .D(n128), .CLK(rclk), .R(n10608), .S(1'b1), 
        .Q(wr_ptr_gray_ss[0]) );
  DFFSR wr_ptr_bin_reg_2_ ( .D(n2637), .CLK(wclk), .R(n10608), .S(1'b1), .Q(
        wr_ptr_bin[2]) );
  DFFSR wr_ptr_gray_reg_1_ ( .D(n174), .CLK(wclk), .R(n10607), .S(1'b1), .Q(
        wr_ptr_gray[1]) );
  DFFSR wr_ptr_gray_s_reg_1_ ( .D(n125), .CLK(rclk), .R(n10607), .S(1'b1), .Q(
        wr_ptr_gray_s[1]) );
  DFFSR wr_ptr_gray_ss_reg_1_ ( .D(n122), .CLK(rclk), .R(n10607), .S(1'b1), 
        .Q(wr_ptr_gray_ss[1]) );
  DFFSR wr_ptr_bin_reg_3_ ( .D(n2632), .CLK(wclk), .R(n10607), .S(1'b1), .Q(
        wr_ptr_bin[3]) );
  DFFSR wr_ptr_gray_reg_2_ ( .D(n22), .CLK(wclk), .R(n10607), .S(1'b1), .Q(
        wr_ptr_gray[2]) );
  DFFSR wr_ptr_gray_s_reg_2_ ( .D(n119), .CLK(rclk), .R(n10607), .S(1'b1), .Q(
        wr_ptr_gray_s[2]) );
  DFFSR wr_ptr_gray_ss_reg_2_ ( .D(n116), .CLK(rclk), .R(n10607), .S(1'b1), 
        .Q(wr_ptr_gray_ss[2]) );
  DFFSR wr_ptr_bin_reg_4_ ( .D(n2627), .CLK(wclk), .R(n10607), .S(1'b1), .Q(
        wr_ptr_bin[4]) );
  DFFSR wr_ptr_gray_reg_3_ ( .D(n21), .CLK(wclk), .R(n10541), .S(1'b1), .Q(
        wr_ptr_gray[3]) );
  DFFSR wr_ptr_gray_s_reg_3_ ( .D(n113), .CLK(rclk), .R(n10541), .S(1'b1), .Q(
        wr_ptr_gray_s[3]) );
  DFFSR wr_ptr_gray_ss_reg_3_ ( .D(n105), .CLK(rclk), .R(n10541), .S(1'b1), 
        .Q(wr_ptr_gray_ss[3]) );
  DFFSR wr_ptr_gray_reg_4_ ( .D(n20), .CLK(wclk), .R(n10541), .S(1'b1), .Q(
        wr_ptr_gray[4]) );
  DFFSR wr_ptr_gray_s_reg_4_ ( .D(n68), .CLK(rclk), .R(n10540), .S(1'b1), .Q(
        wr_ptr_gray_s[4]) );
  DFFSR data_out_reg_31_ ( .D(n2557), .CLK(rclk), .R(n10537), .S(1'b1), .Q(
        n11799) );
  DFFSR data_out_reg_32_ ( .D(n2555), .CLK(rclk), .R(n10537), .S(1'b1), .Q(
        n11798) );
  DFFSR rd_ptr_gray_reg_0_ ( .D(n19), .CLK(rclk), .R(n10540), .S(1'b1), .Q(
        rd_ptr_gray[0]) );
  DFFSR rd_ptr_gray_s_reg_0_ ( .D(n62), .CLK(wclk), .R(n10540), .S(1'b1), .Q(
        rd_ptr_gray_s[0]) );
  DFFSR rd_ptr_gray_ss_reg_0_ ( .D(n59), .CLK(wclk), .R(n10540), .S(1'b1), .Q(
        rd_ptr_gray_ss[0]) );
  DFFSR rd_ptr_gray_reg_1_ ( .D(n18), .CLK(rclk), .R(n10540), .S(1'b1), .Q(
        rd_ptr_gray[1]) );
  DFFSR rd_ptr_gray_s_reg_1_ ( .D(n56), .CLK(wclk), .R(n10540), .S(1'b1), .Q(
        rd_ptr_gray_s[1]) );
  DFFSR rd_ptr_gray_ss_reg_1_ ( .D(n53), .CLK(wclk), .R(n10540), .S(1'b1), .Q(
        rd_ptr_gray_ss[1]) );
  DFFSR rd_ptr_gray_reg_2_ ( .D(n17), .CLK(rclk), .R(n10539), .S(1'b1), .Q(
        rd_ptr_gray[2]) );
  DFFSR rd_ptr_gray_s_reg_2_ ( .D(n50), .CLK(wclk), .R(n10539), .S(1'b1), .Q(
        rd_ptr_gray_s[2]) );
  DFFSR rd_ptr_gray_ss_reg_2_ ( .D(n47), .CLK(wclk), .R(n10539), .S(1'b1), .Q(
        rd_ptr_gray_ss[2]) );
  DFFSR rd_ptr_gray_reg_3_ ( .D(n16), .CLK(rclk), .R(n10539), .S(1'b1), .Q(
        rd_ptr_gray[3]) );
  DFFSR rd_ptr_gray_s_reg_3_ ( .D(n44), .CLK(wclk), .R(n10539), .S(1'b1), .Q(
        rd_ptr_gray_s[3]) );
  DFFSR rd_ptr_gray_ss_reg_3_ ( .D(n41), .CLK(wclk), .R(n10539), .S(1'b1), .Q(
        rd_ptr_gray_ss[3]) );
  DFFSR fifo_reg_1__33_ ( .D(n2695), .CLK(wclk), .R(n10564), .S(1'b1), .Q(
        fifo[1053]) );
  DFFSR fifo_reg_1__32_ ( .D(n2696), .CLK(wclk), .R(n10564), .S(1'b1), .Q(
        fifo[1052]) );
  DFFSR fifo_reg_1__31_ ( .D(n2697), .CLK(wclk), .R(n10564), .S(1'b1), .Q(
        fifo[1051]) );
  DFFSR fifo_reg_1__30_ ( .D(n2698), .CLK(wclk), .R(n10564), .S(1'b1), .Q(
        fifo[1050]) );
  DFFSR fifo_reg_1__29_ ( .D(n2699), .CLK(wclk), .R(n10564), .S(1'b1), .Q(
        fifo[1049]) );
  DFFSR fifo_reg_1__28_ ( .D(n2700), .CLK(wclk), .R(n10564), .S(1'b1), .Q(
        fifo[1048]) );
  DFFSR fifo_reg_1__27_ ( .D(n2701), .CLK(wclk), .R(n10565), .S(1'b1), .Q(
        fifo[1047]) );
  DFFSR fifo_reg_1__26_ ( .D(n2702), .CLK(wclk), .R(n10565), .S(1'b1), .Q(
        fifo[1046]) );
  DFFSR fifo_reg_1__25_ ( .D(n2703), .CLK(wclk), .R(n10565), .S(1'b1), .Q(
        fifo[1045]) );
  DFFSR fifo_reg_1__24_ ( .D(n2704), .CLK(wclk), .R(n10565), .S(1'b1), .Q(
        fifo[1044]) );
  DFFSR fifo_reg_1__23_ ( .D(n2705), .CLK(wclk), .R(n10565), .S(1'b1), .Q(
        fifo[1043]) );
  DFFSR fifo_reg_1__22_ ( .D(n2706), .CLK(wclk), .R(n10565), .S(1'b1), .Q(
        fifo[1042]) );
  DFFSR fifo_reg_1__21_ ( .D(n2707), .CLK(wclk), .R(n10565), .S(1'b1), .Q(
        fifo[1041]) );
  DFFSR fifo_reg_1__20_ ( .D(n2708), .CLK(wclk), .R(n10565), .S(1'b1), .Q(
        fifo[1040]) );
  DFFSR fifo_reg_1__19_ ( .D(n2709), .CLK(wclk), .R(n10565), .S(1'b1), .Q(
        fifo[1039]) );
  DFFSR fifo_reg_1__18_ ( .D(n2710), .CLK(wclk), .R(n10565), .S(1'b1), .Q(
        fifo[1038]) );
  DFFSR fifo_reg_1__17_ ( .D(n2711), .CLK(wclk), .R(n10565), .S(1'b1), .Q(
        fifo[1037]) );
  DFFSR fifo_reg_1__16_ ( .D(n2712), .CLK(wclk), .R(n10565), .S(1'b1), .Q(
        fifo[1036]) );
  DFFSR fifo_reg_1__15_ ( .D(n2713), .CLK(wclk), .R(n10566), .S(1'b1), .Q(
        fifo[1035]) );
  DFFSR fifo_reg_1__14_ ( .D(n2714), .CLK(wclk), .R(n10566), .S(1'b1), .Q(
        fifo[1034]) );
  DFFSR fifo_reg_1__13_ ( .D(n2715), .CLK(wclk), .R(n10566), .S(1'b1), .Q(
        fifo[1033]) );
  DFFSR fifo_reg_1__12_ ( .D(n2716), .CLK(wclk), .R(n10566), .S(1'b1), .Q(
        fifo[1032]) );
  DFFSR fifo_reg_1__11_ ( .D(n2717), .CLK(wclk), .R(n10566), .S(1'b1), .Q(
        fifo[1031]) );
  DFFSR fifo_reg_1__10_ ( .D(n2718), .CLK(wclk), .R(n10566), .S(1'b1), .Q(
        fifo[1030]) );
  DFFSR fifo_reg_1__9_ ( .D(n2719), .CLK(wclk), .R(n10566), .S(1'b1), .Q(
        fifo[1029]) );
  DFFSR fifo_reg_1__8_ ( .D(n2720), .CLK(wclk), .R(n10566), .S(1'b1), .Q(
        fifo[1028]) );
  DFFSR fifo_reg_1__7_ ( .D(n2721), .CLK(wclk), .R(n10566), .S(1'b1), .Q(
        fifo[1027]) );
  DFFSR fifo_reg_1__6_ ( .D(n2722), .CLK(wclk), .R(n10566), .S(1'b1), .Q(
        fifo[1026]) );
  DFFSR fifo_reg_1__5_ ( .D(n2723), .CLK(wclk), .R(n10566), .S(1'b1), .Q(
        fifo[1025]) );
  DFFSR fifo_reg_1__4_ ( .D(n2724), .CLK(wclk), .R(n10566), .S(1'b1), .Q(
        fifo[1024]) );
  DFFSR fifo_reg_1__3_ ( .D(n2725), .CLK(wclk), .R(n10567), .S(1'b1), .Q(
        fifo[1023]) );
  DFFSR fifo_reg_1__2_ ( .D(n2726), .CLK(wclk), .R(n10567), .S(1'b1), .Q(
        fifo[1022]) );
  DFFSR fifo_reg_1__1_ ( .D(n2727), .CLK(wclk), .R(n10567), .S(1'b1), .Q(
        fifo[1021]) );
  DFFSR fifo_reg_1__0_ ( .D(n2728), .CLK(wclk), .R(n10567), .S(1'b1), .Q(
        fifo[1020]) );
  DFFSR fifo_reg_2__33_ ( .D(n2729), .CLK(wclk), .R(n10567), .S(1'b1), .Q(
        fifo[1019]) );
  DFFSR fifo_reg_2__32_ ( .D(n2730), .CLK(wclk), .R(n10567), .S(1'b1), .Q(
        fifo[1018]) );
  DFFSR fifo_reg_2__31_ ( .D(n2731), .CLK(wclk), .R(n10567), .S(1'b1), .Q(
        fifo[1017]) );
  DFFSR fifo_reg_2__30_ ( .D(n2732), .CLK(wclk), .R(n10567), .S(1'b1), .Q(
        fifo[1016]) );
  DFFSR fifo_reg_2__29_ ( .D(n2733), .CLK(wclk), .R(n10567), .S(1'b1), .Q(
        fifo[1015]) );
  DFFSR fifo_reg_2__28_ ( .D(n2734), .CLK(wclk), .R(n10567), .S(1'b1), .Q(
        fifo[1014]) );
  DFFSR fifo_reg_2__27_ ( .D(n2735), .CLK(wclk), .R(n10567), .S(1'b1), .Q(
        fifo[1013]) );
  DFFSR fifo_reg_2__26_ ( .D(n2736), .CLK(wclk), .R(n10567), .S(1'b1), .Q(
        fifo[1012]) );
  DFFSR fifo_reg_2__25_ ( .D(n2737), .CLK(wclk), .R(n10568), .S(1'b1), .Q(
        fifo[1011]) );
  DFFSR fifo_reg_2__24_ ( .D(n2738), .CLK(wclk), .R(n10568), .S(1'b1), .Q(
        fifo[1010]) );
  DFFSR fifo_reg_2__23_ ( .D(n2739), .CLK(wclk), .R(n10568), .S(1'b1), .Q(
        fifo[1009]) );
  DFFSR fifo_reg_2__22_ ( .D(n2740), .CLK(wclk), .R(n10568), .S(1'b1), .Q(
        fifo[1008]) );
  DFFSR fifo_reg_2__21_ ( .D(n2741), .CLK(wclk), .R(n10568), .S(1'b1), .Q(
        fifo[1007]) );
  DFFSR fifo_reg_2__20_ ( .D(n2742), .CLK(wclk), .R(n10568), .S(1'b1), .Q(
        fifo[1006]) );
  DFFSR fifo_reg_2__19_ ( .D(n2743), .CLK(wclk), .R(n10568), .S(1'b1), .Q(
        fifo[1005]) );
  DFFSR fifo_reg_2__18_ ( .D(n2744), .CLK(wclk), .R(n10568), .S(1'b1), .Q(
        fifo[1004]) );
  DFFSR fifo_reg_2__17_ ( .D(n2745), .CLK(wclk), .R(n10568), .S(1'b1), .Q(
        fifo[1003]) );
  DFFSR fifo_reg_2__16_ ( .D(n2746), .CLK(wclk), .R(n10568), .S(1'b1), .Q(
        fifo[1002]) );
  DFFSR fifo_reg_2__15_ ( .D(n2747), .CLK(wclk), .R(n10568), .S(1'b1), .Q(
        fifo[1001]) );
  DFFSR fifo_reg_2__14_ ( .D(n2748), .CLK(wclk), .R(n10568), .S(1'b1), .Q(
        fifo[1000]) );
  DFFSR fifo_reg_2__13_ ( .D(n2749), .CLK(wclk), .R(n10569), .S(1'b1), .Q(
        fifo[999]) );
  DFFSR fifo_reg_2__12_ ( .D(n2750), .CLK(wclk), .R(n10569), .S(1'b1), .Q(
        fifo[998]) );
  DFFSR fifo_reg_2__11_ ( .D(n2751), .CLK(wclk), .R(n10569), .S(1'b1), .Q(
        fifo[997]) );
  DFFSR fifo_reg_2__10_ ( .D(n2752), .CLK(wclk), .R(n10569), .S(1'b1), .Q(
        fifo[996]) );
  DFFSR fifo_reg_2__9_ ( .D(n2753), .CLK(wclk), .R(n10569), .S(1'b1), .Q(
        fifo[995]) );
  DFFSR fifo_reg_2__8_ ( .D(n2754), .CLK(wclk), .R(n10569), .S(1'b1), .Q(
        fifo[994]) );
  DFFSR fifo_reg_2__7_ ( .D(n2755), .CLK(wclk), .R(n10569), .S(1'b1), .Q(
        fifo[993]) );
  DFFSR fifo_reg_2__6_ ( .D(n2756), .CLK(wclk), .R(n10569), .S(1'b1), .Q(
        fifo[992]) );
  DFFSR fifo_reg_2__5_ ( .D(n2757), .CLK(wclk), .R(n10569), .S(1'b1), .Q(
        fifo[991]) );
  DFFSR fifo_reg_2__4_ ( .D(n2758), .CLK(wclk), .R(n10569), .S(1'b1), .Q(
        fifo[990]) );
  DFFSR fifo_reg_2__3_ ( .D(n2759), .CLK(wclk), .R(n10569), .S(1'b1), .Q(
        fifo[989]) );
  DFFSR fifo_reg_2__2_ ( .D(n2760), .CLK(wclk), .R(n10569), .S(1'b1), .Q(
        fifo[988]) );
  DFFSR fifo_reg_2__1_ ( .D(n2761), .CLK(wclk), .R(n10570), .S(1'b1), .Q(
        fifo[987]) );
  DFFSR fifo_reg_2__0_ ( .D(n2762), .CLK(wclk), .R(n10570), .S(1'b1), .Q(
        fifo[986]) );
  DFFSR fifo_reg_3__33_ ( .D(n2763), .CLK(wclk), .R(n10570), .S(1'b1), .Q(
        fifo[985]) );
  DFFSR fifo_reg_3__32_ ( .D(n2764), .CLK(wclk), .R(n10570), .S(1'b1), .Q(
        fifo[984]) );
  DFFSR fifo_reg_3__31_ ( .D(n2765), .CLK(wclk), .R(n10570), .S(1'b1), .Q(
        fifo[983]) );
  DFFSR fifo_reg_3__30_ ( .D(n2766), .CLK(wclk), .R(n10570), .S(1'b1), .Q(
        fifo[982]) );
  DFFSR fifo_reg_3__29_ ( .D(n2767), .CLK(wclk), .R(n10570), .S(1'b1), .Q(
        fifo[981]) );
  DFFSR fifo_reg_3__28_ ( .D(n2768), .CLK(wclk), .R(n10570), .S(1'b1), .Q(
        fifo[980]) );
  DFFSR fifo_reg_3__27_ ( .D(n2769), .CLK(wclk), .R(n10570), .S(1'b1), .Q(
        fifo[979]) );
  DFFSR fifo_reg_3__26_ ( .D(n2770), .CLK(wclk), .R(n10570), .S(1'b1), .Q(
        fifo[978]) );
  DFFSR fifo_reg_3__25_ ( .D(n2771), .CLK(wclk), .R(n10570), .S(1'b1), .Q(
        fifo[977]) );
  DFFSR fifo_reg_3__24_ ( .D(n2772), .CLK(wclk), .R(n10570), .S(1'b1), .Q(
        fifo[976]) );
  DFFSR fifo_reg_3__23_ ( .D(n2773), .CLK(wclk), .R(n10571), .S(1'b1), .Q(
        fifo[975]) );
  DFFSR fifo_reg_3__22_ ( .D(n2774), .CLK(wclk), .R(n10571), .S(1'b1), .Q(
        fifo[974]) );
  DFFSR fifo_reg_3__21_ ( .D(n2775), .CLK(wclk), .R(n10571), .S(1'b1), .Q(
        fifo[973]) );
  DFFSR fifo_reg_3__20_ ( .D(n2776), .CLK(wclk), .R(n10571), .S(1'b1), .Q(
        fifo[972]) );
  DFFSR fifo_reg_3__19_ ( .D(n2777), .CLK(wclk), .R(n10571), .S(1'b1), .Q(
        fifo[971]) );
  DFFSR fifo_reg_3__18_ ( .D(n2778), .CLK(wclk), .R(n10571), .S(1'b1), .Q(
        fifo[970]) );
  DFFSR fifo_reg_3__17_ ( .D(n2779), .CLK(wclk), .R(n10571), .S(1'b1), .Q(
        fifo[969]) );
  DFFSR fifo_reg_3__16_ ( .D(n2780), .CLK(wclk), .R(n10571), .S(1'b1), .Q(
        fifo[968]) );
  DFFSR fifo_reg_3__15_ ( .D(n2781), .CLK(wclk), .R(n10571), .S(1'b1), .Q(
        fifo[967]) );
  DFFSR fifo_reg_3__14_ ( .D(n2782), .CLK(wclk), .R(n10571), .S(1'b1), .Q(
        fifo[966]) );
  DFFSR fifo_reg_3__13_ ( .D(n2783), .CLK(wclk), .R(n10571), .S(1'b1), .Q(
        fifo[965]) );
  DFFSR fifo_reg_3__12_ ( .D(n2784), .CLK(wclk), .R(n10571), .S(1'b1), .Q(
        fifo[964]) );
  DFFSR fifo_reg_3__11_ ( .D(n2785), .CLK(wclk), .R(n10572), .S(1'b1), .Q(
        fifo[963]) );
  DFFSR fifo_reg_3__10_ ( .D(n2786), .CLK(wclk), .R(n10572), .S(1'b1), .Q(
        fifo[962]) );
  DFFSR fifo_reg_3__9_ ( .D(n2787), .CLK(wclk), .R(n10572), .S(1'b1), .Q(
        fifo[961]) );
  DFFSR fifo_reg_3__8_ ( .D(n2788), .CLK(wclk), .R(n10572), .S(1'b1), .Q(
        fifo[960]) );
  DFFSR fifo_reg_3__7_ ( .D(n2789), .CLK(wclk), .R(n10572), .S(1'b1), .Q(
        fifo[959]) );
  DFFSR fifo_reg_3__6_ ( .D(n2790), .CLK(wclk), .R(n10572), .S(1'b1), .Q(
        fifo[958]) );
  DFFSR fifo_reg_3__5_ ( .D(n2791), .CLK(wclk), .R(n10572), .S(1'b1), .Q(
        fifo[957]) );
  DFFSR fifo_reg_3__4_ ( .D(n2792), .CLK(wclk), .R(n10572), .S(1'b1), .Q(
        fifo[956]) );
  DFFSR fifo_reg_3__3_ ( .D(n2793), .CLK(wclk), .R(n10572), .S(1'b1), .Q(
        fifo[955]) );
  DFFSR fifo_reg_3__2_ ( .D(n2794), .CLK(wclk), .R(n10572), .S(1'b1), .Q(
        fifo[954]) );
  DFFSR fifo_reg_3__1_ ( .D(n2795), .CLK(wclk), .R(n10572), .S(1'b1), .Q(
        fifo[953]) );
  DFFSR fifo_reg_3__0_ ( .D(n2796), .CLK(wclk), .R(n10572), .S(1'b1), .Q(
        fifo[952]) );
  DFFSR fifo_reg_4__33_ ( .D(n2797), .CLK(wclk), .R(n10573), .S(1'b1), .Q(
        fifo[951]) );
  DFFSR fifo_reg_4__32_ ( .D(n2798), .CLK(wclk), .R(n10573), .S(1'b1), .Q(
        fifo[950]) );
  DFFSR fifo_reg_4__31_ ( .D(n2799), .CLK(wclk), .R(n10573), .S(1'b1), .Q(
        fifo[949]) );
  DFFSR fifo_reg_4__30_ ( .D(n2800), .CLK(wclk), .R(n10573), .S(1'b1), .Q(
        fifo[948]) );
  DFFSR fifo_reg_4__29_ ( .D(n2801), .CLK(wclk), .R(n10573), .S(1'b1), .Q(
        fifo[947]) );
  DFFSR fifo_reg_4__28_ ( .D(n2802), .CLK(wclk), .R(n10573), .S(1'b1), .Q(
        fifo[946]) );
  DFFSR fifo_reg_4__27_ ( .D(n2803), .CLK(wclk), .R(n10573), .S(1'b1), .Q(
        fifo[945]) );
  DFFSR fifo_reg_4__26_ ( .D(n2804), .CLK(wclk), .R(n10573), .S(1'b1), .Q(
        fifo[944]) );
  DFFSR fifo_reg_4__25_ ( .D(n2805), .CLK(wclk), .R(n10573), .S(1'b1), .Q(
        fifo[943]) );
  DFFSR fifo_reg_4__24_ ( .D(n2806), .CLK(wclk), .R(n10573), .S(1'b1), .Q(
        fifo[942]) );
  DFFSR fifo_reg_4__23_ ( .D(n2807), .CLK(wclk), .R(n10573), .S(1'b1), .Q(
        fifo[941]) );
  DFFSR fifo_reg_4__22_ ( .D(n2808), .CLK(wclk), .R(n10573), .S(1'b1), .Q(
        fifo[940]) );
  DFFSR fifo_reg_4__21_ ( .D(n2809), .CLK(wclk), .R(n10574), .S(1'b1), .Q(
        fifo[939]) );
  DFFSR fifo_reg_4__20_ ( .D(n2810), .CLK(wclk), .R(n10574), .S(1'b1), .Q(
        fifo[938]) );
  DFFSR fifo_reg_4__19_ ( .D(n2811), .CLK(wclk), .R(n10574), .S(1'b1), .Q(
        fifo[937]) );
  DFFSR fifo_reg_4__18_ ( .D(n2812), .CLK(wclk), .R(n10574), .S(1'b1), .Q(
        fifo[936]) );
  DFFSR fifo_reg_4__17_ ( .D(n2813), .CLK(wclk), .R(n10574), .S(1'b1), .Q(
        fifo[935]) );
  DFFSR fifo_reg_4__16_ ( .D(n2814), .CLK(wclk), .R(n10574), .S(1'b1), .Q(
        fifo[934]) );
  DFFSR fifo_reg_4__15_ ( .D(n2815), .CLK(wclk), .R(n10574), .S(1'b1), .Q(
        fifo[933]) );
  DFFSR fifo_reg_4__14_ ( .D(n2816), .CLK(wclk), .R(n10574), .S(1'b1), .Q(
        fifo[932]) );
  DFFSR fifo_reg_4__13_ ( .D(n2817), .CLK(wclk), .R(n10574), .S(1'b1), .Q(
        fifo[931]) );
  DFFSR fifo_reg_4__12_ ( .D(n2818), .CLK(wclk), .R(n10574), .S(1'b1), .Q(
        fifo[930]) );
  DFFSR fifo_reg_4__11_ ( .D(n2819), .CLK(wclk), .R(n10574), .S(1'b1), .Q(
        fifo[929]) );
  DFFSR fifo_reg_4__10_ ( .D(n2820), .CLK(wclk), .R(n10574), .S(1'b1), .Q(
        fifo[928]) );
  DFFSR fifo_reg_4__9_ ( .D(n2821), .CLK(wclk), .R(n10575), .S(1'b1), .Q(
        fifo[927]) );
  DFFSR fifo_reg_4__8_ ( .D(n2822), .CLK(wclk), .R(n10575), .S(1'b1), .Q(
        fifo[926]) );
  DFFSR fifo_reg_4__7_ ( .D(n2823), .CLK(wclk), .R(n10575), .S(1'b1), .Q(
        fifo[925]) );
  DFFSR fifo_reg_4__6_ ( .D(n2824), .CLK(wclk), .R(n10575), .S(1'b1), .Q(
        fifo[924]) );
  DFFSR fifo_reg_4__5_ ( .D(n2825), .CLK(wclk), .R(n10575), .S(1'b1), .Q(
        fifo[923]) );
  DFFSR fifo_reg_4__4_ ( .D(n2826), .CLK(wclk), .R(n10575), .S(1'b1), .Q(
        fifo[922]) );
  DFFSR fifo_reg_4__3_ ( .D(n2827), .CLK(wclk), .R(n10575), .S(1'b1), .Q(
        fifo[921]) );
  DFFSR fifo_reg_4__2_ ( .D(n2828), .CLK(wclk), .R(n10575), .S(1'b1), .Q(
        fifo[920]) );
  DFFSR fifo_reg_4__1_ ( .D(n2829), .CLK(wclk), .R(n10575), .S(1'b1), .Q(
        fifo[919]) );
  DFFSR fifo_reg_4__0_ ( .D(n2830), .CLK(wclk), .R(n10575), .S(1'b1), .Q(
        fifo[918]) );
  DFFSR fifo_reg_5__33_ ( .D(n2831), .CLK(wclk), .R(n10575), .S(1'b1), .Q(
        fifo[917]) );
  DFFSR fifo_reg_5__32_ ( .D(n2832), .CLK(wclk), .R(n10575), .S(1'b1), .Q(
        fifo[916]) );
  DFFSR fifo_reg_5__31_ ( .D(n2833), .CLK(wclk), .R(n10576), .S(1'b1), .Q(
        fifo[915]) );
  DFFSR fifo_reg_5__30_ ( .D(n2834), .CLK(wclk), .R(n10576), .S(1'b1), .Q(
        fifo[914]) );
  DFFSR fifo_reg_5__29_ ( .D(n2835), .CLK(wclk), .R(n10576), .S(1'b1), .Q(
        fifo[913]) );
  DFFSR fifo_reg_5__28_ ( .D(n2836), .CLK(wclk), .R(n10576), .S(1'b1), .Q(
        fifo[912]) );
  DFFSR fifo_reg_5__27_ ( .D(n2837), .CLK(wclk), .R(n10576), .S(1'b1), .Q(
        fifo[911]) );
  DFFSR fifo_reg_5__26_ ( .D(n2838), .CLK(wclk), .R(n10576), .S(1'b1), .Q(
        fifo[910]) );
  DFFSR fifo_reg_5__25_ ( .D(n2839), .CLK(wclk), .R(n10576), .S(1'b1), .Q(
        fifo[909]) );
  DFFSR fifo_reg_5__24_ ( .D(n2840), .CLK(wclk), .R(n10576), .S(1'b1), .Q(
        fifo[908]) );
  DFFSR fifo_reg_5__23_ ( .D(n2841), .CLK(wclk), .R(n10576), .S(1'b1), .Q(
        fifo[907]) );
  DFFSR fifo_reg_5__22_ ( .D(n2842), .CLK(wclk), .R(n10576), .S(1'b1), .Q(
        fifo[906]) );
  DFFSR fifo_reg_5__21_ ( .D(n2843), .CLK(wclk), .R(n10576), .S(1'b1), .Q(
        fifo[905]) );
  DFFSR fifo_reg_5__20_ ( .D(n2844), .CLK(wclk), .R(n10576), .S(1'b1), .Q(
        fifo[904]) );
  DFFSR fifo_reg_5__19_ ( .D(n2845), .CLK(wclk), .R(n10577), .S(1'b1), .Q(
        fifo[903]) );
  DFFSR fifo_reg_5__18_ ( .D(n2846), .CLK(wclk), .R(n10577), .S(1'b1), .Q(
        fifo[902]) );
  DFFSR fifo_reg_5__17_ ( .D(n2847), .CLK(wclk), .R(n10577), .S(1'b1), .Q(
        fifo[901]) );
  DFFSR fifo_reg_5__16_ ( .D(n2848), .CLK(wclk), .R(n10577), .S(1'b1), .Q(
        fifo[900]) );
  DFFSR fifo_reg_5__15_ ( .D(n2849), .CLK(wclk), .R(n10577), .S(1'b1), .Q(
        fifo[899]) );
  DFFSR fifo_reg_5__14_ ( .D(n2850), .CLK(wclk), .R(n10577), .S(1'b1), .Q(
        fifo[898]) );
  DFFSR fifo_reg_5__13_ ( .D(n2851), .CLK(wclk), .R(n10577), .S(1'b1), .Q(
        fifo[897]) );
  DFFSR fifo_reg_5__12_ ( .D(n2852), .CLK(wclk), .R(n10577), .S(1'b1), .Q(
        fifo[896]) );
  DFFSR fifo_reg_5__11_ ( .D(n2853), .CLK(wclk), .R(n10577), .S(1'b1), .Q(
        fifo[895]) );
  DFFSR fifo_reg_5__10_ ( .D(n2854), .CLK(wclk), .R(n10577), .S(1'b1), .Q(
        fifo[894]) );
  DFFSR fifo_reg_5__9_ ( .D(n2855), .CLK(wclk), .R(n10577), .S(1'b1), .Q(
        fifo[893]) );
  DFFSR fifo_reg_5__8_ ( .D(n2856), .CLK(wclk), .R(n10577), .S(1'b1), .Q(
        fifo[892]) );
  DFFSR fifo_reg_5__7_ ( .D(n2857), .CLK(wclk), .R(n10578), .S(1'b1), .Q(
        fifo[891]) );
  DFFSR fifo_reg_5__6_ ( .D(n2858), .CLK(wclk), .R(n10578), .S(1'b1), .Q(
        fifo[890]) );
  DFFSR fifo_reg_5__5_ ( .D(n2859), .CLK(wclk), .R(n10578), .S(1'b1), .Q(
        fifo[889]) );
  DFFSR fifo_reg_5__4_ ( .D(n2860), .CLK(wclk), .R(n10578), .S(1'b1), .Q(
        fifo[888]) );
  DFFSR fifo_reg_5__3_ ( .D(n2861), .CLK(wclk), .R(n10578), .S(1'b1), .Q(
        fifo[887]) );
  DFFSR fifo_reg_5__2_ ( .D(n2862), .CLK(wclk), .R(n10578), .S(1'b1), .Q(
        fifo[886]) );
  DFFSR fifo_reg_5__1_ ( .D(n2863), .CLK(wclk), .R(n10578), .S(1'b1), .Q(
        fifo[885]) );
  DFFSR fifo_reg_5__0_ ( .D(n2864), .CLK(wclk), .R(n10578), .S(1'b1), .Q(
        fifo[884]) );
  DFFSR fifo_reg_6__33_ ( .D(n2865), .CLK(wclk), .R(n10578), .S(1'b1), .Q(
        fifo[883]) );
  DFFSR fifo_reg_6__32_ ( .D(n2866), .CLK(wclk), .R(n10578), .S(1'b1), .Q(
        fifo[882]) );
  DFFSR fifo_reg_6__31_ ( .D(n2867), .CLK(wclk), .R(n10578), .S(1'b1), .Q(
        fifo[881]) );
  DFFSR fifo_reg_6__30_ ( .D(n2868), .CLK(wclk), .R(n10578), .S(1'b1), .Q(
        fifo[880]) );
  DFFSR fifo_reg_6__29_ ( .D(n2869), .CLK(wclk), .R(n10579), .S(1'b1), .Q(
        fifo[879]) );
  DFFSR fifo_reg_6__28_ ( .D(n2870), .CLK(wclk), .R(n10579), .S(1'b1), .Q(
        fifo[878]) );
  DFFSR fifo_reg_6__27_ ( .D(n2871), .CLK(wclk), .R(n10579), .S(1'b1), .Q(
        fifo[877]) );
  DFFSR fifo_reg_6__26_ ( .D(n2872), .CLK(wclk), .R(n10579), .S(1'b1), .Q(
        fifo[876]) );
  DFFSR fifo_reg_6__25_ ( .D(n2873), .CLK(wclk), .R(n10579), .S(1'b1), .Q(
        fifo[875]) );
  DFFSR fifo_reg_6__24_ ( .D(n2874), .CLK(wclk), .R(n10579), .S(1'b1), .Q(
        fifo[874]) );
  DFFSR fifo_reg_6__23_ ( .D(n2875), .CLK(wclk), .R(n10579), .S(1'b1), .Q(
        fifo[873]) );
  DFFSR fifo_reg_6__22_ ( .D(n2876), .CLK(wclk), .R(n10579), .S(1'b1), .Q(
        fifo[872]) );
  DFFSR fifo_reg_6__21_ ( .D(n2877), .CLK(wclk), .R(n10579), .S(1'b1), .Q(
        fifo[871]) );
  DFFSR fifo_reg_6__20_ ( .D(n2878), .CLK(wclk), .R(n10579), .S(1'b1), .Q(
        fifo[870]) );
  DFFSR fifo_reg_6__19_ ( .D(n2879), .CLK(wclk), .R(n10579), .S(1'b1), .Q(
        fifo[869]) );
  DFFSR fifo_reg_6__18_ ( .D(n2880), .CLK(wclk), .R(n10579), .S(1'b1), .Q(
        fifo[868]) );
  DFFSR fifo_reg_6__17_ ( .D(n2881), .CLK(wclk), .R(n10580), .S(1'b1), .Q(
        fifo[867]) );
  DFFSR fifo_reg_6__16_ ( .D(n2882), .CLK(wclk), .R(n10580), .S(1'b1), .Q(
        fifo[866]) );
  DFFSR fifo_reg_6__15_ ( .D(n2883), .CLK(wclk), .R(n10580), .S(1'b1), .Q(
        fifo[865]) );
  DFFSR fifo_reg_6__14_ ( .D(n2884), .CLK(wclk), .R(n10580), .S(1'b1), .Q(
        fifo[864]) );
  DFFSR fifo_reg_6__13_ ( .D(n2885), .CLK(wclk), .R(n10580), .S(1'b1), .Q(
        fifo[863]) );
  DFFSR fifo_reg_6__12_ ( .D(n2886), .CLK(wclk), .R(n10580), .S(1'b1), .Q(
        fifo[862]) );
  DFFSR fifo_reg_6__11_ ( .D(n2887), .CLK(wclk), .R(n10580), .S(1'b1), .Q(
        fifo[861]) );
  DFFSR fifo_reg_6__10_ ( .D(n2888), .CLK(wclk), .R(n10580), .S(1'b1), .Q(
        fifo[860]) );
  DFFSR fifo_reg_6__9_ ( .D(n2889), .CLK(wclk), .R(n10580), .S(1'b1), .Q(
        fifo[859]) );
  DFFSR fifo_reg_6__8_ ( .D(n2890), .CLK(wclk), .R(n10580), .S(1'b1), .Q(
        fifo[858]) );
  DFFSR fifo_reg_6__7_ ( .D(n2891), .CLK(wclk), .R(n10580), .S(1'b1), .Q(
        fifo[857]) );
  DFFSR fifo_reg_6__6_ ( .D(n2892), .CLK(wclk), .R(n10580), .S(1'b1), .Q(
        fifo[856]) );
  DFFSR fifo_reg_6__5_ ( .D(n2893), .CLK(wclk), .R(n10581), .S(1'b1), .Q(
        fifo[855]) );
  DFFSR fifo_reg_6__4_ ( .D(n2894), .CLK(wclk), .R(n10581), .S(1'b1), .Q(
        fifo[854]) );
  DFFSR fifo_reg_6__3_ ( .D(n2895), .CLK(wclk), .R(n10581), .S(1'b1), .Q(
        fifo[853]) );
  DFFSR fifo_reg_6__2_ ( .D(n2896), .CLK(wclk), .R(n10581), .S(1'b1), .Q(
        fifo[852]) );
  DFFSR fifo_reg_6__1_ ( .D(n2897), .CLK(wclk), .R(n10581), .S(1'b1), .Q(
        fifo[851]) );
  DFFSR fifo_reg_6__0_ ( .D(n2898), .CLK(wclk), .R(n10581), .S(1'b1), .Q(
        fifo[850]) );
  DFFSR fifo_reg_7__33_ ( .D(n2899), .CLK(wclk), .R(n10581), .S(1'b1), .Q(
        fifo[849]) );
  DFFSR fifo_reg_7__32_ ( .D(n2900), .CLK(wclk), .R(n10581), .S(1'b1), .Q(
        fifo[848]) );
  DFFSR fifo_reg_7__31_ ( .D(n2901), .CLK(wclk), .R(n10581), .S(1'b1), .Q(
        fifo[847]) );
  DFFSR fifo_reg_7__30_ ( .D(n2902), .CLK(wclk), .R(n10581), .S(1'b1), .Q(
        fifo[846]) );
  DFFSR fifo_reg_7__29_ ( .D(n2903), .CLK(wclk), .R(n10581), .S(1'b1), .Q(
        fifo[845]) );
  DFFSR fifo_reg_7__28_ ( .D(n2904), .CLK(wclk), .R(n10581), .S(1'b1), .Q(
        fifo[844]) );
  DFFSR fifo_reg_7__27_ ( .D(n2905), .CLK(wclk), .R(n10582), .S(1'b1), .Q(
        fifo[843]) );
  DFFSR fifo_reg_7__26_ ( .D(n2906), .CLK(wclk), .R(n10582), .S(1'b1), .Q(
        fifo[842]) );
  DFFSR fifo_reg_7__25_ ( .D(n2907), .CLK(wclk), .R(n10582), .S(1'b1), .Q(
        fifo[841]) );
  DFFSR fifo_reg_7__24_ ( .D(n2908), .CLK(wclk), .R(n10582), .S(1'b1), .Q(
        fifo[840]) );
  DFFSR fifo_reg_7__23_ ( .D(n2909), .CLK(wclk), .R(n10582), .S(1'b1), .Q(
        fifo[839]) );
  DFFSR fifo_reg_7__22_ ( .D(n2910), .CLK(wclk), .R(n10582), .S(1'b1), .Q(
        fifo[838]) );
  DFFSR fifo_reg_7__21_ ( .D(n2911), .CLK(wclk), .R(n10582), .S(1'b1), .Q(
        fifo[837]) );
  DFFSR fifo_reg_7__20_ ( .D(n2912), .CLK(wclk), .R(n10582), .S(1'b1), .Q(
        fifo[836]) );
  DFFSR fifo_reg_7__19_ ( .D(n2913), .CLK(wclk), .R(n10582), .S(1'b1), .Q(
        fifo[835]) );
  DFFSR fifo_reg_7__18_ ( .D(n2914), .CLK(wclk), .R(n10582), .S(1'b1), .Q(
        fifo[834]) );
  DFFSR fifo_reg_7__17_ ( .D(n2915), .CLK(wclk), .R(n10582), .S(1'b1), .Q(
        fifo[833]) );
  DFFSR fifo_reg_7__16_ ( .D(n2916), .CLK(wclk), .R(n10582), .S(1'b1), .Q(
        fifo[832]) );
  DFFSR fifo_reg_7__15_ ( .D(n2917), .CLK(wclk), .R(n10583), .S(1'b1), .Q(
        fifo[831]) );
  DFFSR fifo_reg_7__14_ ( .D(n2918), .CLK(wclk), .R(n10583), .S(1'b1), .Q(
        fifo[830]) );
  DFFSR fifo_reg_7__13_ ( .D(n2919), .CLK(wclk), .R(n10583), .S(1'b1), .Q(
        fifo[829]) );
  DFFSR fifo_reg_7__12_ ( .D(n2920), .CLK(wclk), .R(n10583), .S(1'b1), .Q(
        fifo[828]) );
  DFFSR fifo_reg_7__11_ ( .D(n2921), .CLK(wclk), .R(n10583), .S(1'b1), .Q(
        fifo[827]) );
  DFFSR fifo_reg_7__10_ ( .D(n2922), .CLK(wclk), .R(n10583), .S(1'b1), .Q(
        fifo[826]) );
  DFFSR fifo_reg_7__9_ ( .D(n2923), .CLK(wclk), .R(n10583), .S(1'b1), .Q(
        fifo[825]) );
  DFFSR fifo_reg_7__8_ ( .D(n2924), .CLK(wclk), .R(n10583), .S(1'b1), .Q(
        fifo[824]) );
  DFFSR fifo_reg_7__7_ ( .D(n2925), .CLK(wclk), .R(n10583), .S(1'b1), .Q(
        fifo[823]) );
  DFFSR fifo_reg_7__6_ ( .D(n2926), .CLK(wclk), .R(n10583), .S(1'b1), .Q(
        fifo[822]) );
  DFFSR fifo_reg_7__5_ ( .D(n2927), .CLK(wclk), .R(n10583), .S(1'b1), .Q(
        fifo[821]) );
  DFFSR fifo_reg_7__4_ ( .D(n2928), .CLK(wclk), .R(n10583), .S(1'b1), .Q(
        fifo[820]) );
  DFFSR fifo_reg_7__3_ ( .D(n2929), .CLK(wclk), .R(n10584), .S(1'b1), .Q(
        fifo[819]) );
  DFFSR fifo_reg_7__2_ ( .D(n2930), .CLK(wclk), .R(n10584), .S(1'b1), .Q(
        fifo[818]) );
  DFFSR fifo_reg_7__1_ ( .D(n2931), .CLK(wclk), .R(n10584), .S(1'b1), .Q(
        fifo[817]) );
  DFFSR fifo_reg_7__0_ ( .D(n2932), .CLK(wclk), .R(n10584), .S(1'b1), .Q(
        fifo[816]) );
  DFFSR fifo_reg_8__33_ ( .D(n2933), .CLK(wclk), .R(n10584), .S(1'b1), .Q(
        fifo[815]) );
  DFFSR fifo_reg_8__32_ ( .D(n2934), .CLK(wclk), .R(n10584), .S(1'b1), .Q(
        fifo[814]) );
  DFFSR fifo_reg_8__31_ ( .D(n2935), .CLK(wclk), .R(n10584), .S(1'b1), .Q(
        fifo[813]) );
  DFFSR fifo_reg_8__30_ ( .D(n2936), .CLK(wclk), .R(n10584), .S(1'b1), .Q(
        fifo[812]) );
  DFFSR fifo_reg_8__29_ ( .D(n2937), .CLK(wclk), .R(n10584), .S(1'b1), .Q(
        fifo[811]) );
  DFFSR fifo_reg_8__28_ ( .D(n2938), .CLK(wclk), .R(n10584), .S(1'b1), .Q(
        fifo[810]) );
  DFFSR fifo_reg_8__27_ ( .D(n2939), .CLK(wclk), .R(n10584), .S(1'b1), .Q(
        fifo[809]) );
  DFFSR fifo_reg_8__26_ ( .D(n2940), .CLK(wclk), .R(n10584), .S(1'b1), .Q(
        fifo[808]) );
  DFFSR fifo_reg_8__25_ ( .D(n2941), .CLK(wclk), .R(n10585), .S(1'b1), .Q(
        fifo[807]) );
  DFFSR fifo_reg_8__24_ ( .D(n2942), .CLK(wclk), .R(n10585), .S(1'b1), .Q(
        fifo[806]) );
  DFFSR fifo_reg_8__23_ ( .D(n2943), .CLK(wclk), .R(n10585), .S(1'b1), .Q(
        fifo[805]) );
  DFFSR fifo_reg_8__22_ ( .D(n2944), .CLK(wclk), .R(n10585), .S(1'b1), .Q(
        fifo[804]) );
  DFFSR fifo_reg_8__21_ ( .D(n2945), .CLK(wclk), .R(n10585), .S(1'b1), .Q(
        fifo[803]) );
  DFFSR fifo_reg_8__20_ ( .D(n2946), .CLK(wclk), .R(n10585), .S(1'b1), .Q(
        fifo[802]) );
  DFFSR fifo_reg_8__19_ ( .D(n2947), .CLK(wclk), .R(n10585), .S(1'b1), .Q(
        fifo[801]) );
  DFFSR fifo_reg_8__18_ ( .D(n2948), .CLK(wclk), .R(n10585), .S(1'b1), .Q(
        fifo[800]) );
  DFFSR fifo_reg_8__17_ ( .D(n2949), .CLK(wclk), .R(n10585), .S(1'b1), .Q(
        fifo[799]) );
  DFFSR fifo_reg_8__16_ ( .D(n2950), .CLK(wclk), .R(n10585), .S(1'b1), .Q(
        fifo[798]) );
  DFFSR fifo_reg_8__15_ ( .D(n2951), .CLK(wclk), .R(n10585), .S(1'b1), .Q(
        fifo[797]) );
  DFFSR fifo_reg_8__14_ ( .D(n2952), .CLK(wclk), .R(n10585), .S(1'b1), .Q(
        fifo[796]) );
  DFFSR fifo_reg_8__13_ ( .D(n2953), .CLK(wclk), .R(n10586), .S(1'b1), .Q(
        fifo[795]) );
  DFFSR fifo_reg_8__12_ ( .D(n2954), .CLK(wclk), .R(n10586), .S(1'b1), .Q(
        fifo[794]) );
  DFFSR fifo_reg_8__11_ ( .D(n2955), .CLK(wclk), .R(n10586), .S(1'b1), .Q(
        fifo[793]) );
  DFFSR fifo_reg_8__10_ ( .D(n2956), .CLK(wclk), .R(n10586), .S(1'b1), .Q(
        fifo[792]) );
  DFFSR fifo_reg_8__9_ ( .D(n2957), .CLK(wclk), .R(n10586), .S(1'b1), .Q(
        fifo[791]) );
  DFFSR fifo_reg_8__8_ ( .D(n2958), .CLK(wclk), .R(n10586), .S(1'b1), .Q(
        fifo[790]) );
  DFFSR fifo_reg_8__7_ ( .D(n2959), .CLK(wclk), .R(n10586), .S(1'b1), .Q(
        fifo[789]) );
  DFFSR fifo_reg_8__6_ ( .D(n2960), .CLK(wclk), .R(n10586), .S(1'b1), .Q(
        fifo[788]) );
  DFFSR fifo_reg_8__5_ ( .D(n2961), .CLK(wclk), .R(n10586), .S(1'b1), .Q(
        fifo[787]) );
  DFFSR fifo_reg_8__4_ ( .D(n2962), .CLK(wclk), .R(n10586), .S(1'b1), .Q(
        fifo[786]) );
  DFFSR fifo_reg_8__3_ ( .D(n2963), .CLK(wclk), .R(n10586), .S(1'b1), .Q(
        fifo[785]) );
  DFFSR fifo_reg_8__2_ ( .D(n2964), .CLK(wclk), .R(n10586), .S(1'b1), .Q(
        fifo[784]) );
  DFFSR fifo_reg_8__1_ ( .D(n2965), .CLK(wclk), .R(n10587), .S(1'b1), .Q(
        fifo[783]) );
  DFFSR fifo_reg_8__0_ ( .D(n2966), .CLK(wclk), .R(n10587), .S(1'b1), .Q(
        fifo[782]) );
  DFFSR fifo_reg_9__33_ ( .D(n2967), .CLK(wclk), .R(n10587), .S(1'b1), .Q(
        fifo[781]) );
  DFFSR fifo_reg_9__32_ ( .D(n2968), .CLK(wclk), .R(n10587), .S(1'b1), .Q(
        fifo[780]) );
  DFFSR fifo_reg_9__31_ ( .D(n2969), .CLK(wclk), .R(n10587), .S(1'b1), .Q(
        fifo[779]) );
  DFFSR fifo_reg_9__30_ ( .D(n2970), .CLK(wclk), .R(n10587), .S(1'b1), .Q(
        fifo[778]) );
  DFFSR fifo_reg_9__29_ ( .D(n2971), .CLK(wclk), .R(n10587), .S(1'b1), .Q(
        fifo[777]) );
  DFFSR fifo_reg_9__28_ ( .D(n2972), .CLK(wclk), .R(n10587), .S(1'b1), .Q(
        fifo[776]) );
  DFFSR fifo_reg_9__27_ ( .D(n2973), .CLK(wclk), .R(n10587), .S(1'b1), .Q(
        fifo[775]) );
  DFFSR fifo_reg_9__26_ ( .D(n2974), .CLK(wclk), .R(n10587), .S(1'b1), .Q(
        fifo[774]) );
  DFFSR fifo_reg_9__25_ ( .D(n2975), .CLK(wclk), .R(n10587), .S(1'b1), .Q(
        fifo[773]) );
  DFFSR fifo_reg_9__24_ ( .D(n2976), .CLK(wclk), .R(n10587), .S(1'b1), .Q(
        fifo[772]) );
  DFFSR fifo_reg_9__23_ ( .D(n2977), .CLK(wclk), .R(n10588), .S(1'b1), .Q(
        fifo[771]) );
  DFFSR fifo_reg_9__22_ ( .D(n2978), .CLK(wclk), .R(n10588), .S(1'b1), .Q(
        fifo[770]) );
  DFFSR fifo_reg_9__21_ ( .D(n2979), .CLK(wclk), .R(n10588), .S(1'b1), .Q(
        fifo[769]) );
  DFFSR fifo_reg_9__20_ ( .D(n2980), .CLK(wclk), .R(n10588), .S(1'b1), .Q(
        fifo[768]) );
  DFFSR fifo_reg_9__19_ ( .D(n2981), .CLK(wclk), .R(n10588), .S(1'b1), .Q(
        fifo[767]) );
  DFFSR fifo_reg_9__18_ ( .D(n2982), .CLK(wclk), .R(n10588), .S(1'b1), .Q(
        fifo[766]) );
  DFFSR fifo_reg_9__17_ ( .D(n2983), .CLK(wclk), .R(n10588), .S(1'b1), .Q(
        fifo[765]) );
  DFFSR fifo_reg_9__16_ ( .D(n2984), .CLK(wclk), .R(n10588), .S(1'b1), .Q(
        fifo[764]) );
  DFFSR fifo_reg_9__15_ ( .D(n2985), .CLK(wclk), .R(n10588), .S(1'b1), .Q(
        fifo[763]) );
  DFFSR fifo_reg_9__14_ ( .D(n2986), .CLK(wclk), .R(n10588), .S(1'b1), .Q(
        fifo[762]) );
  DFFSR fifo_reg_9__13_ ( .D(n2987), .CLK(wclk), .R(n10588), .S(1'b1), .Q(
        fifo[761]) );
  DFFSR fifo_reg_9__12_ ( .D(n2988), .CLK(wclk), .R(n10588), .S(1'b1), .Q(
        fifo[760]) );
  DFFSR fifo_reg_9__11_ ( .D(n2989), .CLK(wclk), .R(n10589), .S(1'b1), .Q(
        fifo[759]) );
  DFFSR fifo_reg_9__10_ ( .D(n2990), .CLK(wclk), .R(n10589), .S(1'b1), .Q(
        fifo[758]) );
  DFFSR fifo_reg_9__9_ ( .D(n2991), .CLK(wclk), .R(n10589), .S(1'b1), .Q(
        fifo[757]) );
  DFFSR fifo_reg_9__8_ ( .D(n2992), .CLK(wclk), .R(n10589), .S(1'b1), .Q(
        fifo[756]) );
  DFFSR fifo_reg_9__7_ ( .D(n2993), .CLK(wclk), .R(n10589), .S(1'b1), .Q(
        fifo[755]) );
  DFFSR fifo_reg_9__6_ ( .D(n2994), .CLK(wclk), .R(n10589), .S(1'b1), .Q(
        fifo[754]) );
  DFFSR fifo_reg_9__5_ ( .D(n2995), .CLK(wclk), .R(n10589), .S(1'b1), .Q(
        fifo[753]) );
  DFFSR fifo_reg_9__4_ ( .D(n2996), .CLK(wclk), .R(n10589), .S(1'b1), .Q(
        fifo[752]) );
  DFFSR fifo_reg_9__3_ ( .D(n2997), .CLK(wclk), .R(n10589), .S(1'b1), .Q(
        fifo[751]) );
  DFFSR fifo_reg_9__2_ ( .D(n2998), .CLK(wclk), .R(n10589), .S(1'b1), .Q(
        fifo[750]) );
  DFFSR fifo_reg_9__1_ ( .D(n2999), .CLK(wclk), .R(n10589), .S(1'b1), .Q(
        fifo[749]) );
  DFFSR fifo_reg_9__0_ ( .D(n3000), .CLK(wclk), .R(n10589), .S(1'b1), .Q(
        fifo[748]) );
  DFFSR fifo_reg_10__33_ ( .D(n3001), .CLK(wclk), .R(n10590), .S(1'b1), .Q(
        fifo[747]) );
  DFFSR fifo_reg_10__32_ ( .D(n3002), .CLK(wclk), .R(n10590), .S(1'b1), .Q(
        fifo[746]) );
  DFFSR fifo_reg_10__31_ ( .D(n3003), .CLK(wclk), .R(n10590), .S(1'b1), .Q(
        fifo[745]) );
  DFFSR fifo_reg_10__30_ ( .D(n3004), .CLK(wclk), .R(n10590), .S(1'b1), .Q(
        fifo[744]) );
  DFFSR fifo_reg_10__29_ ( .D(n3005), .CLK(wclk), .R(n10590), .S(1'b1), .Q(
        fifo[743]) );
  DFFSR fifo_reg_10__28_ ( .D(n3006), .CLK(wclk), .R(n10590), .S(1'b1), .Q(
        fifo[742]) );
  DFFSR fifo_reg_10__27_ ( .D(n3007), .CLK(wclk), .R(n10590), .S(1'b1), .Q(
        fifo[741]) );
  DFFSR fifo_reg_10__26_ ( .D(n3008), .CLK(wclk), .R(n10590), .S(1'b1), .Q(
        fifo[740]) );
  DFFSR fifo_reg_10__25_ ( .D(n3009), .CLK(wclk), .R(n10590), .S(1'b1), .Q(
        fifo[739]) );
  DFFSR fifo_reg_10__24_ ( .D(n3010), .CLK(wclk), .R(n10590), .S(1'b1), .Q(
        fifo[738]) );
  DFFSR fifo_reg_10__23_ ( .D(n3011), .CLK(wclk), .R(n10590), .S(1'b1), .Q(
        fifo[737]) );
  DFFSR fifo_reg_10__22_ ( .D(n3012), .CLK(wclk), .R(n10590), .S(1'b1), .Q(
        fifo[736]) );
  DFFSR fifo_reg_10__21_ ( .D(n3013), .CLK(wclk), .R(n10591), .S(1'b1), .Q(
        fifo[735]) );
  DFFSR fifo_reg_10__20_ ( .D(n3014), .CLK(wclk), .R(n10591), .S(1'b1), .Q(
        fifo[734]) );
  DFFSR fifo_reg_10__19_ ( .D(n3015), .CLK(wclk), .R(n10591), .S(1'b1), .Q(
        fifo[733]) );
  DFFSR fifo_reg_10__18_ ( .D(n3016), .CLK(wclk), .R(n10591), .S(1'b1), .Q(
        fifo[732]) );
  DFFSR fifo_reg_10__17_ ( .D(n3017), .CLK(wclk), .R(n10591), .S(1'b1), .Q(
        fifo[731]) );
  DFFSR fifo_reg_10__16_ ( .D(n3018), .CLK(wclk), .R(n10591), .S(1'b1), .Q(
        fifo[730]) );
  DFFSR fifo_reg_10__15_ ( .D(n3019), .CLK(wclk), .R(n10591), .S(1'b1), .Q(
        fifo[729]) );
  DFFSR fifo_reg_10__14_ ( .D(n3020), .CLK(wclk), .R(n10591), .S(1'b1), .Q(
        fifo[728]) );
  DFFSR fifo_reg_10__13_ ( .D(n3021), .CLK(wclk), .R(n10591), .S(1'b1), .Q(
        fifo[727]) );
  DFFSR fifo_reg_10__12_ ( .D(n3022), .CLK(wclk), .R(n10591), .S(1'b1), .Q(
        fifo[726]) );
  DFFSR fifo_reg_10__11_ ( .D(n3023), .CLK(wclk), .R(n10591), .S(1'b1), .Q(
        fifo[725]) );
  DFFSR fifo_reg_10__10_ ( .D(n3024), .CLK(wclk), .R(n10591), .S(1'b1), .Q(
        fifo[724]) );
  DFFSR fifo_reg_10__9_ ( .D(n3025), .CLK(wclk), .R(n10592), .S(1'b1), .Q(
        fifo[723]) );
  DFFSR fifo_reg_10__8_ ( .D(n3026), .CLK(wclk), .R(n10592), .S(1'b1), .Q(
        fifo[722]) );
  DFFSR fifo_reg_10__7_ ( .D(n3027), .CLK(wclk), .R(n10592), .S(1'b1), .Q(
        fifo[721]) );
  DFFSR fifo_reg_10__6_ ( .D(n3028), .CLK(wclk), .R(n10592), .S(1'b1), .Q(
        fifo[720]) );
  DFFSR fifo_reg_10__5_ ( .D(n3029), .CLK(wclk), .R(n10592), .S(1'b1), .Q(
        fifo[719]) );
  DFFSR fifo_reg_10__4_ ( .D(n3030), .CLK(wclk), .R(n10592), .S(1'b1), .Q(
        fifo[718]) );
  DFFSR fifo_reg_10__3_ ( .D(n3031), .CLK(wclk), .R(n10592), .S(1'b1), .Q(
        fifo[717]) );
  DFFSR fifo_reg_10__2_ ( .D(n3032), .CLK(wclk), .R(n10592), .S(1'b1), .Q(
        fifo[716]) );
  DFFSR fifo_reg_10__1_ ( .D(n3033), .CLK(wclk), .R(n10592), .S(1'b1), .Q(
        fifo[715]) );
  DFFSR fifo_reg_10__0_ ( .D(n3034), .CLK(wclk), .R(n10592), .S(1'b1), .Q(
        fifo[714]) );
  DFFSR fifo_reg_11__33_ ( .D(n3035), .CLK(wclk), .R(n10592), .S(1'b1), .Q(
        fifo[713]) );
  DFFSR fifo_reg_11__32_ ( .D(n3036), .CLK(wclk), .R(n10592), .S(1'b1), .Q(
        fifo[712]) );
  DFFSR fifo_reg_11__31_ ( .D(n3037), .CLK(wclk), .R(n10593), .S(1'b1), .Q(
        fifo[711]) );
  DFFSR fifo_reg_11__30_ ( .D(n3038), .CLK(wclk), .R(n10593), .S(1'b1), .Q(
        fifo[710]) );
  DFFSR fifo_reg_11__29_ ( .D(n3039), .CLK(wclk), .R(n10593), .S(1'b1), .Q(
        fifo[709]) );
  DFFSR fifo_reg_11__28_ ( .D(n3040), .CLK(wclk), .R(n10593), .S(1'b1), .Q(
        fifo[708]) );
  DFFSR fifo_reg_11__27_ ( .D(n3041), .CLK(wclk), .R(n10593), .S(1'b1), .Q(
        fifo[707]) );
  DFFSR fifo_reg_11__26_ ( .D(n3042), .CLK(wclk), .R(n10593), .S(1'b1), .Q(
        fifo[706]) );
  DFFSR fifo_reg_11__25_ ( .D(n3043), .CLK(wclk), .R(n10593), .S(1'b1), .Q(
        fifo[705]) );
  DFFSR fifo_reg_11__24_ ( .D(n3044), .CLK(wclk), .R(n10593), .S(1'b1), .Q(
        fifo[704]) );
  DFFSR fifo_reg_11__23_ ( .D(n3045), .CLK(wclk), .R(n10593), .S(1'b1), .Q(
        fifo[703]) );
  DFFSR fifo_reg_11__22_ ( .D(n3046), .CLK(wclk), .R(n10593), .S(1'b1), .Q(
        fifo[702]) );
  DFFSR fifo_reg_11__21_ ( .D(n3047), .CLK(wclk), .R(n10593), .S(1'b1), .Q(
        fifo[701]) );
  DFFSR fifo_reg_11__20_ ( .D(n3048), .CLK(wclk), .R(n10593), .S(1'b1), .Q(
        fifo[700]) );
  DFFSR fifo_reg_11__19_ ( .D(n3049), .CLK(wclk), .R(n10594), .S(1'b1), .Q(
        fifo[699]) );
  DFFSR fifo_reg_11__18_ ( .D(n3050), .CLK(wclk), .R(n10594), .S(1'b1), .Q(
        fifo[698]) );
  DFFSR fifo_reg_11__17_ ( .D(n3051), .CLK(wclk), .R(n10594), .S(1'b1), .Q(
        fifo[697]) );
  DFFSR fifo_reg_11__16_ ( .D(n3052), .CLK(wclk), .R(n10594), .S(1'b1), .Q(
        fifo[696]) );
  DFFSR fifo_reg_11__15_ ( .D(n3053), .CLK(wclk), .R(n10594), .S(1'b1), .Q(
        fifo[695]) );
  DFFSR fifo_reg_11__14_ ( .D(n3054), .CLK(wclk), .R(n10594), .S(1'b1), .Q(
        fifo[694]) );
  DFFSR fifo_reg_11__13_ ( .D(n3055), .CLK(wclk), .R(n10594), .S(1'b1), .Q(
        fifo[693]) );
  DFFSR fifo_reg_11__12_ ( .D(n3056), .CLK(wclk), .R(n10594), .S(1'b1), .Q(
        fifo[692]) );
  DFFSR fifo_reg_11__11_ ( .D(n3057), .CLK(wclk), .R(n10594), .S(1'b1), .Q(
        fifo[691]) );
  DFFSR fifo_reg_11__10_ ( .D(n3058), .CLK(wclk), .R(n10594), .S(1'b1), .Q(
        fifo[690]) );
  DFFSR fifo_reg_11__9_ ( .D(n3059), .CLK(wclk), .R(n10594), .S(1'b1), .Q(
        fifo[689]) );
  DFFSR fifo_reg_11__8_ ( .D(n3060), .CLK(wclk), .R(n10594), .S(1'b1), .Q(
        fifo[688]) );
  DFFSR fifo_reg_11__7_ ( .D(n3061), .CLK(wclk), .R(n10595), .S(1'b1), .Q(
        fifo[687]) );
  DFFSR fifo_reg_11__6_ ( .D(n3062), .CLK(wclk), .R(n10595), .S(1'b1), .Q(
        fifo[686]) );
  DFFSR fifo_reg_11__5_ ( .D(n3063), .CLK(wclk), .R(n10595), .S(1'b1), .Q(
        fifo[685]) );
  DFFSR fifo_reg_11__4_ ( .D(n3064), .CLK(wclk), .R(n10595), .S(1'b1), .Q(
        fifo[684]) );
  DFFSR fifo_reg_11__3_ ( .D(n3065), .CLK(wclk), .R(n10595), .S(1'b1), .Q(
        fifo[683]) );
  DFFSR fifo_reg_11__2_ ( .D(n3066), .CLK(wclk), .R(n10595), .S(1'b1), .Q(
        fifo[682]) );
  DFFSR fifo_reg_11__1_ ( .D(n3067), .CLK(wclk), .R(n10595), .S(1'b1), .Q(
        fifo[681]) );
  DFFSR fifo_reg_11__0_ ( .D(n3068), .CLK(wclk), .R(n10595), .S(1'b1), .Q(
        fifo[680]) );
  DFFSR fifo_reg_12__33_ ( .D(n3069), .CLK(wclk), .R(n10595), .S(1'b1), .Q(
        fifo[679]) );
  DFFSR fifo_reg_12__32_ ( .D(n3070), .CLK(wclk), .R(n10595), .S(1'b1), .Q(
        fifo[678]) );
  DFFSR fifo_reg_12__31_ ( .D(n3071), .CLK(wclk), .R(n10595), .S(1'b1), .Q(
        fifo[677]) );
  DFFSR fifo_reg_12__30_ ( .D(n3072), .CLK(wclk), .R(n10595), .S(1'b1), .Q(
        fifo[676]) );
  DFFSR fifo_reg_12__29_ ( .D(n3073), .CLK(wclk), .R(n10596), .S(1'b1), .Q(
        fifo[675]) );
  DFFSR fifo_reg_12__28_ ( .D(n3074), .CLK(wclk), .R(n10596), .S(1'b1), .Q(
        fifo[674]) );
  DFFSR fifo_reg_12__27_ ( .D(n3075), .CLK(wclk), .R(n10596), .S(1'b1), .Q(
        fifo[673]) );
  DFFSR fifo_reg_12__26_ ( .D(n3076), .CLK(wclk), .R(n10596), .S(1'b1), .Q(
        fifo[672]) );
  DFFSR fifo_reg_12__25_ ( .D(n3077), .CLK(wclk), .R(n10596), .S(1'b1), .Q(
        fifo[671]) );
  DFFSR fifo_reg_12__24_ ( .D(n3078), .CLK(wclk), .R(n10596), .S(1'b1), .Q(
        fifo[670]) );
  DFFSR fifo_reg_12__23_ ( .D(n3079), .CLK(wclk), .R(n10596), .S(1'b1), .Q(
        fifo[669]) );
  DFFSR fifo_reg_12__22_ ( .D(n3080), .CLK(wclk), .R(n10596), .S(1'b1), .Q(
        fifo[668]) );
  DFFSR fifo_reg_12__21_ ( .D(n3081), .CLK(wclk), .R(n10596), .S(1'b1), .Q(
        fifo[667]) );
  DFFSR fifo_reg_12__20_ ( .D(n3082), .CLK(wclk), .R(n10596), .S(1'b1), .Q(
        fifo[666]) );
  DFFSR fifo_reg_12__19_ ( .D(n3083), .CLK(wclk), .R(n10596), .S(1'b1), .Q(
        fifo[665]) );
  DFFSR fifo_reg_12__18_ ( .D(n3084), .CLK(wclk), .R(n10596), .S(1'b1), .Q(
        fifo[664]) );
  DFFSR fifo_reg_12__17_ ( .D(n3085), .CLK(wclk), .R(n10597), .S(1'b1), .Q(
        fifo[663]) );
  DFFSR fifo_reg_12__16_ ( .D(n3086), .CLK(wclk), .R(n10597), .S(1'b1), .Q(
        fifo[662]) );
  DFFSR fifo_reg_12__15_ ( .D(n3087), .CLK(wclk), .R(n10597), .S(1'b1), .Q(
        fifo[661]) );
  DFFSR fifo_reg_12__14_ ( .D(n3088), .CLK(wclk), .R(n10597), .S(1'b1), .Q(
        fifo[660]) );
  DFFSR fifo_reg_12__13_ ( .D(n3089), .CLK(wclk), .R(n10597), .S(1'b1), .Q(
        fifo[659]) );
  DFFSR fifo_reg_12__12_ ( .D(n3090), .CLK(wclk), .R(n10597), .S(1'b1), .Q(
        fifo[658]) );
  DFFSR fifo_reg_12__11_ ( .D(n3091), .CLK(wclk), .R(n10597), .S(1'b1), .Q(
        fifo[657]) );
  DFFSR fifo_reg_12__10_ ( .D(n3092), .CLK(wclk), .R(n10597), .S(1'b1), .Q(
        fifo[656]) );
  DFFSR fifo_reg_12__9_ ( .D(n3093), .CLK(wclk), .R(n10597), .S(1'b1), .Q(
        fifo[655]) );
  DFFSR fifo_reg_12__8_ ( .D(n3094), .CLK(wclk), .R(n10597), .S(1'b1), .Q(
        fifo[654]) );
  DFFSR fifo_reg_12__7_ ( .D(n3095), .CLK(wclk), .R(n10597), .S(1'b1), .Q(
        fifo[653]) );
  DFFSR fifo_reg_12__6_ ( .D(n3096), .CLK(wclk), .R(n10597), .S(1'b1), .Q(
        fifo[652]) );
  DFFSR fifo_reg_12__5_ ( .D(n3097), .CLK(wclk), .R(n10598), .S(1'b1), .Q(
        fifo[651]) );
  DFFSR fifo_reg_12__4_ ( .D(n3098), .CLK(wclk), .R(n10598), .S(1'b1), .Q(
        fifo[650]) );
  DFFSR fifo_reg_12__3_ ( .D(n3099), .CLK(wclk), .R(n10598), .S(1'b1), .Q(
        fifo[649]) );
  DFFSR fifo_reg_12__2_ ( .D(n3100), .CLK(wclk), .R(n10598), .S(1'b1), .Q(
        fifo[648]) );
  DFFSR fifo_reg_12__1_ ( .D(n3101), .CLK(wclk), .R(n10598), .S(1'b1), .Q(
        fifo[647]) );
  DFFSR fifo_reg_12__0_ ( .D(n3102), .CLK(wclk), .R(n10598), .S(1'b1), .Q(
        fifo[646]) );
  DFFSR fifo_reg_13__33_ ( .D(n3103), .CLK(wclk), .R(n10598), .S(1'b1), .Q(
        fifo[645]) );
  DFFSR fifo_reg_13__32_ ( .D(n3104), .CLK(wclk), .R(n10598), .S(1'b1), .Q(
        fifo[644]) );
  DFFSR fifo_reg_13__31_ ( .D(n3105), .CLK(wclk), .R(n10598), .S(1'b1), .Q(
        fifo[643]) );
  DFFSR fifo_reg_13__30_ ( .D(n3106), .CLK(wclk), .R(n10598), .S(1'b1), .Q(
        fifo[642]) );
  DFFSR fifo_reg_13__29_ ( .D(n3107), .CLK(wclk), .R(n10598), .S(1'b1), .Q(
        fifo[641]) );
  DFFSR fifo_reg_13__28_ ( .D(n3108), .CLK(wclk), .R(n10598), .S(1'b1), .Q(
        fifo[640]) );
  DFFSR fifo_reg_13__27_ ( .D(n3109), .CLK(wclk), .R(n10599), .S(1'b1), .Q(
        fifo[639]) );
  DFFSR fifo_reg_13__26_ ( .D(n3110), .CLK(wclk), .R(n10599), .S(1'b1), .Q(
        fifo[638]) );
  DFFSR fifo_reg_13__25_ ( .D(n3111), .CLK(wclk), .R(n10599), .S(1'b1), .Q(
        fifo[637]) );
  DFFSR fifo_reg_13__24_ ( .D(n3112), .CLK(wclk), .R(n10599), .S(1'b1), .Q(
        fifo[636]) );
  DFFSR fifo_reg_13__23_ ( .D(n3113), .CLK(wclk), .R(n10599), .S(1'b1), .Q(
        fifo[635]) );
  DFFSR fifo_reg_13__22_ ( .D(n3114), .CLK(wclk), .R(n10599), .S(1'b1), .Q(
        fifo[634]) );
  DFFSR fifo_reg_13__21_ ( .D(n3115), .CLK(wclk), .R(n10599), .S(1'b1), .Q(
        fifo[633]) );
  DFFSR fifo_reg_13__20_ ( .D(n3116), .CLK(wclk), .R(n10599), .S(1'b1), .Q(
        fifo[632]) );
  DFFSR fifo_reg_13__19_ ( .D(n3117), .CLK(wclk), .R(n10599), .S(1'b1), .Q(
        fifo[631]) );
  DFFSR fifo_reg_13__18_ ( .D(n3118), .CLK(wclk), .R(n10599), .S(1'b1), .Q(
        fifo[630]) );
  DFFSR fifo_reg_13__17_ ( .D(n3119), .CLK(wclk), .R(n10599), .S(1'b1), .Q(
        fifo[629]) );
  DFFSR fifo_reg_13__16_ ( .D(n3120), .CLK(wclk), .R(n10599), .S(1'b1), .Q(
        fifo[628]) );
  DFFSR fifo_reg_13__15_ ( .D(n3121), .CLK(wclk), .R(n10600), .S(1'b1), .Q(
        fifo[627]) );
  DFFSR fifo_reg_13__14_ ( .D(n3122), .CLK(wclk), .R(n10600), .S(1'b1), .Q(
        fifo[626]) );
  DFFSR fifo_reg_13__13_ ( .D(n3123), .CLK(wclk), .R(n10600), .S(1'b1), .Q(
        fifo[625]) );
  DFFSR fifo_reg_13__12_ ( .D(n3124), .CLK(wclk), .R(n10600), .S(1'b1), .Q(
        fifo[624]) );
  DFFSR fifo_reg_13__11_ ( .D(n3125), .CLK(wclk), .R(n10600), .S(1'b1), .Q(
        fifo[623]) );
  DFFSR fifo_reg_13__10_ ( .D(n3126), .CLK(wclk), .R(n10600), .S(1'b1), .Q(
        fifo[622]) );
  DFFSR fifo_reg_13__9_ ( .D(n3127), .CLK(wclk), .R(n10600), .S(1'b1), .Q(
        fifo[621]) );
  DFFSR fifo_reg_13__8_ ( .D(n3128), .CLK(wclk), .R(n10600), .S(1'b1), .Q(
        fifo[620]) );
  DFFSR fifo_reg_13__7_ ( .D(n3129), .CLK(wclk), .R(n10600), .S(1'b1), .Q(
        fifo[619]) );
  DFFSR fifo_reg_13__6_ ( .D(n3130), .CLK(wclk), .R(n10600), .S(1'b1), .Q(
        fifo[618]) );
  DFFSR fifo_reg_13__5_ ( .D(n3131), .CLK(wclk), .R(n10600), .S(1'b1), .Q(
        fifo[617]) );
  DFFSR fifo_reg_13__4_ ( .D(n3132), .CLK(wclk), .R(n10600), .S(1'b1), .Q(
        fifo[616]) );
  DFFSR fifo_reg_13__3_ ( .D(n3133), .CLK(wclk), .R(n10601), .S(1'b1), .Q(
        fifo[615]) );
  DFFSR fifo_reg_13__2_ ( .D(n3134), .CLK(wclk), .R(n10601), .S(1'b1), .Q(
        fifo[614]) );
  DFFSR fifo_reg_13__1_ ( .D(n3135), .CLK(wclk), .R(n10601), .S(1'b1), .Q(
        fifo[613]) );
  DFFSR fifo_reg_13__0_ ( .D(n3136), .CLK(wclk), .R(n10601), .S(1'b1), .Q(
        fifo[612]) );
  DFFSR fifo_reg_14__33_ ( .D(n3137), .CLK(wclk), .R(n10601), .S(1'b1), .Q(
        fifo[611]) );
  DFFSR fifo_reg_14__32_ ( .D(n3138), .CLK(wclk), .R(n10601), .S(1'b1), .Q(
        fifo[610]) );
  DFFSR fifo_reg_14__31_ ( .D(n3139), .CLK(wclk), .R(n10601), .S(1'b1), .Q(
        fifo[609]) );
  DFFSR fifo_reg_14__30_ ( .D(n3140), .CLK(wclk), .R(n10601), .S(1'b1), .Q(
        fifo[608]) );
  DFFSR fifo_reg_14__29_ ( .D(n3141), .CLK(wclk), .R(n10601), .S(1'b1), .Q(
        fifo[607]) );
  DFFSR fifo_reg_14__28_ ( .D(n3142), .CLK(wclk), .R(n10601), .S(1'b1), .Q(
        fifo[606]) );
  DFFSR fifo_reg_14__27_ ( .D(n3143), .CLK(wclk), .R(n10601), .S(1'b1), .Q(
        fifo[605]) );
  DFFSR fifo_reg_14__26_ ( .D(n3144), .CLK(wclk), .R(n10601), .S(1'b1), .Q(
        fifo[604]) );
  DFFSR fifo_reg_14__25_ ( .D(n3145), .CLK(wclk), .R(n10602), .S(1'b1), .Q(
        fifo[603]) );
  DFFSR fifo_reg_14__24_ ( .D(n3146), .CLK(wclk), .R(n10602), .S(1'b1), .Q(
        fifo[602]) );
  DFFSR fifo_reg_14__23_ ( .D(n3147), .CLK(wclk), .R(n10602), .S(1'b1), .Q(
        fifo[601]) );
  DFFSR fifo_reg_14__22_ ( .D(n3148), .CLK(wclk), .R(n10602), .S(1'b1), .Q(
        fifo[600]) );
  DFFSR fifo_reg_14__21_ ( .D(n3149), .CLK(wclk), .R(n10602), .S(1'b1), .Q(
        fifo[599]) );
  DFFSR fifo_reg_14__20_ ( .D(n3150), .CLK(wclk), .R(n10602), .S(1'b1), .Q(
        fifo[598]) );
  DFFSR fifo_reg_14__19_ ( .D(n3151), .CLK(wclk), .R(n10602), .S(1'b1), .Q(
        fifo[597]) );
  DFFSR fifo_reg_14__18_ ( .D(n3152), .CLK(wclk), .R(n10602), .S(1'b1), .Q(
        fifo[596]) );
  DFFSR fifo_reg_14__17_ ( .D(n3153), .CLK(wclk), .R(n10602), .S(1'b1), .Q(
        fifo[595]) );
  DFFSR fifo_reg_14__16_ ( .D(n3154), .CLK(wclk), .R(n10602), .S(1'b1), .Q(
        fifo[594]) );
  DFFSR fifo_reg_14__15_ ( .D(n3155), .CLK(wclk), .R(n10602), .S(1'b1), .Q(
        fifo[593]) );
  DFFSR fifo_reg_14__14_ ( .D(n3156), .CLK(wclk), .R(n10602), .S(1'b1), .Q(
        fifo[592]) );
  DFFSR fifo_reg_14__13_ ( .D(n3157), .CLK(wclk), .R(n10603), .S(1'b1), .Q(
        fifo[591]) );
  DFFSR fifo_reg_14__12_ ( .D(n3158), .CLK(wclk), .R(n10603), .S(1'b1), .Q(
        fifo[590]) );
  DFFSR fifo_reg_14__11_ ( .D(n3159), .CLK(wclk), .R(n10603), .S(1'b1), .Q(
        fifo[589]) );
  DFFSR fifo_reg_14__10_ ( .D(n3160), .CLK(wclk), .R(n10603), .S(1'b1), .Q(
        fifo[588]) );
  DFFSR fifo_reg_14__9_ ( .D(n3161), .CLK(wclk), .R(n10603), .S(1'b1), .Q(
        fifo[587]) );
  DFFSR fifo_reg_14__8_ ( .D(n3162), .CLK(wclk), .R(n10603), .S(1'b1), .Q(
        fifo[586]) );
  DFFSR fifo_reg_14__7_ ( .D(n3163), .CLK(wclk), .R(n10603), .S(1'b1), .Q(
        fifo[585]) );
  DFFSR fifo_reg_14__6_ ( .D(n3164), .CLK(wclk), .R(n10603), .S(1'b1), .Q(
        fifo[584]) );
  DFFSR fifo_reg_14__5_ ( .D(n3165), .CLK(wclk), .R(n10603), .S(1'b1), .Q(
        fifo[583]) );
  DFFSR fifo_reg_14__4_ ( .D(n3166), .CLK(wclk), .R(n10603), .S(1'b1), .Q(
        fifo[582]) );
  DFFSR fifo_reg_14__3_ ( .D(n3167), .CLK(wclk), .R(n10603), .S(1'b1), .Q(
        fifo[581]) );
  DFFSR fifo_reg_14__2_ ( .D(n3168), .CLK(wclk), .R(n10603), .S(1'b1), .Q(
        fifo[580]) );
  DFFSR fifo_reg_14__1_ ( .D(n3169), .CLK(wclk), .R(n10604), .S(1'b1), .Q(
        fifo[579]) );
  DFFSR fifo_reg_14__0_ ( .D(n3170), .CLK(wclk), .R(n10604), .S(1'b1), .Q(
        fifo[578]) );
  DFFSR fifo_reg_15__33_ ( .D(n3171), .CLK(wclk), .R(n10604), .S(1'b1), .Q(
        fifo[577]) );
  DFFSR fifo_reg_15__32_ ( .D(n3172), .CLK(wclk), .R(n10604), .S(1'b1), .Q(
        fifo[576]) );
  DFFSR fifo_reg_15__31_ ( .D(n3173), .CLK(wclk), .R(n10604), .S(1'b1), .Q(
        fifo[575]) );
  DFFSR fifo_reg_15__30_ ( .D(n3174), .CLK(wclk), .R(n10604), .S(1'b1), .Q(
        fifo[574]) );
  DFFSR fifo_reg_15__29_ ( .D(n3175), .CLK(wclk), .R(n10604), .S(1'b1), .Q(
        fifo[573]) );
  DFFSR fifo_reg_15__28_ ( .D(n3176), .CLK(wclk), .R(n10604), .S(1'b1), .Q(
        fifo[572]) );
  DFFSR fifo_reg_15__27_ ( .D(n3177), .CLK(wclk), .R(n10604), .S(1'b1), .Q(
        fifo[571]) );
  DFFSR fifo_reg_15__26_ ( .D(n3178), .CLK(wclk), .R(n10604), .S(1'b1), .Q(
        fifo[570]) );
  DFFSR fifo_reg_15__25_ ( .D(n3179), .CLK(wclk), .R(n10604), .S(1'b1), .Q(
        fifo[569]) );
  DFFSR fifo_reg_15__24_ ( .D(n3180), .CLK(wclk), .R(n10604), .S(1'b1), .Q(
        fifo[568]) );
  DFFSR fifo_reg_15__23_ ( .D(n3181), .CLK(wclk), .R(n10605), .S(1'b1), .Q(
        fifo[567]) );
  DFFSR fifo_reg_15__22_ ( .D(n3182), .CLK(wclk), .R(n10605), .S(1'b1), .Q(
        fifo[566]) );
  DFFSR fifo_reg_15__21_ ( .D(n3183), .CLK(wclk), .R(n10605), .S(1'b1), .Q(
        fifo[565]) );
  DFFSR fifo_reg_15__20_ ( .D(n3184), .CLK(wclk), .R(n10605), .S(1'b1), .Q(
        fifo[564]) );
  DFFSR fifo_reg_15__19_ ( .D(n3185), .CLK(wclk), .R(n10605), .S(1'b1), .Q(
        fifo[563]) );
  DFFSR fifo_reg_15__18_ ( .D(n3186), .CLK(wclk), .R(n10605), .S(1'b1), .Q(
        fifo[562]) );
  DFFSR fifo_reg_15__17_ ( .D(n3187), .CLK(wclk), .R(n10605), .S(1'b1), .Q(
        fifo[561]) );
  DFFSR fifo_reg_15__16_ ( .D(n3188), .CLK(wclk), .R(n10605), .S(1'b1), .Q(
        fifo[560]) );
  DFFSR fifo_reg_15__15_ ( .D(n3189), .CLK(wclk), .R(n10605), .S(1'b1), .Q(
        fifo[559]) );
  DFFSR fifo_reg_15__14_ ( .D(n3190), .CLK(wclk), .R(n10605), .S(1'b1), .Q(
        fifo[558]) );
  DFFSR fifo_reg_15__13_ ( .D(n3191), .CLK(wclk), .R(n10605), .S(1'b1), .Q(
        fifo[557]) );
  DFFSR fifo_reg_15__12_ ( .D(n3192), .CLK(wclk), .R(n10605), .S(1'b1), .Q(
        fifo[556]) );
  DFFSR fifo_reg_15__11_ ( .D(n3193), .CLK(wclk), .R(n10606), .S(1'b1), .Q(
        fifo[555]) );
  DFFSR fifo_reg_15__10_ ( .D(n3194), .CLK(wclk), .R(n10606), .S(1'b1), .Q(
        fifo[554]) );
  DFFSR fifo_reg_15__9_ ( .D(n3195), .CLK(wclk), .R(n10606), .S(1'b1), .Q(
        fifo[553]) );
  DFFSR fifo_reg_15__8_ ( .D(n3196), .CLK(wclk), .R(n10606), .S(1'b1), .Q(
        fifo[552]) );
  DFFSR fifo_reg_15__7_ ( .D(n3197), .CLK(wclk), .R(n10606), .S(1'b1), .Q(
        fifo[551]) );
  DFFSR fifo_reg_15__6_ ( .D(n3198), .CLK(wclk), .R(n10606), .S(1'b1), .Q(
        fifo[550]) );
  DFFSR fifo_reg_15__5_ ( .D(n3199), .CLK(wclk), .R(n10606), .S(1'b1), .Q(
        fifo[549]) );
  DFFSR fifo_reg_15__4_ ( .D(n3200), .CLK(wclk), .R(n10606), .S(1'b1), .Q(
        fifo[548]) );
  DFFSR fifo_reg_15__3_ ( .D(n3201), .CLK(wclk), .R(n10606), .S(1'b1), .Q(
        fifo[547]) );
  DFFSR fifo_reg_15__2_ ( .D(n3202), .CLK(wclk), .R(n10606), .S(1'b1), .Q(
        fifo[546]) );
  DFFSR fifo_reg_15__1_ ( .D(n3203), .CLK(wclk), .R(n10606), .S(1'b1), .Q(
        fifo[545]) );
  DFFSR fifo_reg_15__0_ ( .D(n3204), .CLK(wclk), .R(n10606), .S(1'b1), .Q(
        fifo[544]) );
  DFFSR fifo_reg_24__33_ ( .D(n3477), .CLK(wclk), .R(n10541), .S(1'b1), .Q(
        fifo[271]) );
  DFFSR fifo_reg_24__32_ ( .D(n3478), .CLK(wclk), .R(n10541), .S(1'b1), .Q(
        fifo[270]) );
  DFFSR fifo_reg_24__31_ ( .D(n3479), .CLK(wclk), .R(n10541), .S(1'b1), .Q(
        fifo[269]) );
  DFFSR fifo_reg_24__30_ ( .D(n3480), .CLK(wclk), .R(n10541), .S(1'b1), .Q(
        fifo[268]) );
  DFFSR fifo_reg_24__29_ ( .D(n3481), .CLK(wclk), .R(n10541), .S(1'b1), .Q(
        fifo[267]) );
  DFFSR fifo_reg_24__28_ ( .D(n3482), .CLK(wclk), .R(n10541), .S(1'b1), .Q(
        fifo[266]) );
  DFFSR fifo_reg_24__27_ ( .D(n3483), .CLK(wclk), .R(n10541), .S(1'b1), .Q(
        fifo[265]) );
  DFFSR fifo_reg_24__26_ ( .D(n3484), .CLK(wclk), .R(n10541), .S(1'b1), .Q(
        fifo[264]) );
  DFFSR fifo_reg_24__25_ ( .D(n3485), .CLK(wclk), .R(n10542), .S(1'b1), .Q(
        fifo[263]) );
  DFFSR fifo_reg_24__24_ ( .D(n3486), .CLK(wclk), .R(n10542), .S(1'b1), .Q(
        fifo[262]) );
  DFFSR fifo_reg_24__23_ ( .D(n3487), .CLK(wclk), .R(n10542), .S(1'b1), .Q(
        fifo[261]) );
  DFFSR fifo_reg_24__22_ ( .D(n3488), .CLK(wclk), .R(n10542), .S(1'b1), .Q(
        fifo[260]) );
  DFFSR fifo_reg_24__21_ ( .D(n3489), .CLK(wclk), .R(n10542), .S(1'b1), .Q(
        fifo[259]) );
  DFFSR fifo_reg_24__20_ ( .D(n3490), .CLK(wclk), .R(n10542), .S(1'b1), .Q(
        fifo[258]) );
  DFFSR fifo_reg_24__19_ ( .D(n3491), .CLK(wclk), .R(n10542), .S(1'b1), .Q(
        fifo[257]) );
  DFFSR fifo_reg_24__18_ ( .D(n3492), .CLK(wclk), .R(n10542), .S(1'b1), .Q(
        fifo[256]) );
  DFFSR fifo_reg_24__17_ ( .D(n3493), .CLK(wclk), .R(n10542), .S(1'b1), .Q(
        fifo[255]) );
  DFFSR fifo_reg_24__16_ ( .D(n3494), .CLK(wclk), .R(n10542), .S(1'b1), .Q(
        fifo[254]) );
  DFFSR fifo_reg_24__15_ ( .D(n3495), .CLK(wclk), .R(n10542), .S(1'b1), .Q(
        fifo[253]) );
  DFFSR fifo_reg_24__14_ ( .D(n3496), .CLK(wclk), .R(n10542), .S(1'b1), .Q(
        fifo[252]) );
  DFFSR fifo_reg_24__13_ ( .D(n3497), .CLK(wclk), .R(n10543), .S(1'b1), .Q(
        fifo[251]) );
  DFFSR fifo_reg_24__12_ ( .D(n3498), .CLK(wclk), .R(n10543), .S(1'b1), .Q(
        fifo[250]) );
  DFFSR fifo_reg_24__11_ ( .D(n3499), .CLK(wclk), .R(n10543), .S(1'b1), .Q(
        fifo[249]) );
  DFFSR fifo_reg_24__10_ ( .D(n3500), .CLK(wclk), .R(n10543), .S(1'b1), .Q(
        fifo[248]) );
  DFFSR fifo_reg_24__9_ ( .D(n3501), .CLK(wclk), .R(n10543), .S(1'b1), .Q(
        fifo[247]) );
  DFFSR fifo_reg_24__8_ ( .D(n3502), .CLK(wclk), .R(n10543), .S(1'b1), .Q(
        fifo[246]) );
  DFFSR fifo_reg_24__7_ ( .D(n3503), .CLK(wclk), .R(n10543), .S(1'b1), .Q(
        fifo[245]) );
  DFFSR fifo_reg_24__6_ ( .D(n3504), .CLK(wclk), .R(n10543), .S(1'b1), .Q(
        fifo[244]) );
  DFFSR fifo_reg_24__5_ ( .D(n3505), .CLK(wclk), .R(n10543), .S(1'b1), .Q(
        fifo[243]) );
  DFFSR fifo_reg_24__4_ ( .D(n3506), .CLK(wclk), .R(n10543), .S(1'b1), .Q(
        fifo[242]) );
  DFFSR fifo_reg_24__3_ ( .D(n3507), .CLK(wclk), .R(n10543), .S(1'b1), .Q(
        fifo[241]) );
  DFFSR fifo_reg_24__2_ ( .D(n3508), .CLK(wclk), .R(n10543), .S(1'b1), .Q(
        fifo[240]) );
  DFFSR fifo_reg_24__1_ ( .D(n3509), .CLK(wclk), .R(n10544), .S(1'b1), .Q(
        fifo[239]) );
  DFFSR fifo_reg_24__0_ ( .D(n3510), .CLK(wclk), .R(n10544), .S(1'b1), .Q(
        fifo[238]) );
  DFFSR fifo_reg_25__33_ ( .D(n3511), .CLK(wclk), .R(n10544), .S(1'b1), .Q(
        fifo[237]) );
  DFFSR fifo_reg_25__32_ ( .D(n3512), .CLK(wclk), .R(n10544), .S(1'b1), .Q(
        fifo[236]) );
  DFFSR fifo_reg_25__31_ ( .D(n3513), .CLK(wclk), .R(n10544), .S(1'b1), .Q(
        fifo[235]) );
  DFFSR fifo_reg_25__30_ ( .D(n3514), .CLK(wclk), .R(n10544), .S(1'b1), .Q(
        fifo[234]) );
  DFFSR fifo_reg_25__29_ ( .D(n3515), .CLK(wclk), .R(n10544), .S(1'b1), .Q(
        fifo[233]) );
  DFFSR fifo_reg_25__28_ ( .D(n3516), .CLK(wclk), .R(n10544), .S(1'b1), .Q(
        fifo[232]) );
  DFFSR fifo_reg_25__27_ ( .D(n3517), .CLK(wclk), .R(n10544), .S(1'b1), .Q(
        fifo[231]) );
  DFFSR fifo_reg_25__26_ ( .D(n3518), .CLK(wclk), .R(n10544), .S(1'b1), .Q(
        fifo[230]) );
  DFFSR fifo_reg_25__25_ ( .D(n3519), .CLK(wclk), .R(n10544), .S(1'b1), .Q(
        fifo[229]) );
  DFFSR fifo_reg_25__24_ ( .D(n3520), .CLK(wclk), .R(n10544), .S(1'b1), .Q(
        fifo[228]) );
  DFFSR fifo_reg_25__23_ ( .D(n3521), .CLK(wclk), .R(n10545), .S(1'b1), .Q(
        fifo[227]) );
  DFFSR fifo_reg_25__22_ ( .D(n3522), .CLK(wclk), .R(n10545), .S(1'b1), .Q(
        fifo[226]) );
  DFFSR fifo_reg_25__21_ ( .D(n3523), .CLK(wclk), .R(n10545), .S(1'b1), .Q(
        fifo[225]) );
  DFFSR fifo_reg_25__20_ ( .D(n3524), .CLK(wclk), .R(n10545), .S(1'b1), .Q(
        fifo[224]) );
  DFFSR fifo_reg_25__19_ ( .D(n3525), .CLK(wclk), .R(n10545), .S(1'b1), .Q(
        fifo[223]) );
  DFFSR fifo_reg_25__18_ ( .D(n3526), .CLK(wclk), .R(n10545), .S(1'b1), .Q(
        fifo[222]) );
  DFFSR fifo_reg_25__17_ ( .D(n3527), .CLK(wclk), .R(n10545), .S(1'b1), .Q(
        fifo[221]) );
  DFFSR fifo_reg_25__16_ ( .D(n3528), .CLK(wclk), .R(n10545), .S(1'b1), .Q(
        fifo[220]) );
  DFFSR fifo_reg_25__15_ ( .D(n3529), .CLK(wclk), .R(n10545), .S(1'b1), .Q(
        fifo[219]) );
  DFFSR fifo_reg_25__14_ ( .D(n3530), .CLK(wclk), .R(n10545), .S(1'b1), .Q(
        fifo[218]) );
  DFFSR fifo_reg_25__13_ ( .D(n3531), .CLK(wclk), .R(n10545), .S(1'b1), .Q(
        fifo[217]) );
  DFFSR fifo_reg_25__12_ ( .D(n3532), .CLK(wclk), .R(n10545), .S(1'b1), .Q(
        fifo[216]) );
  DFFSR fifo_reg_25__11_ ( .D(n3533), .CLK(wclk), .R(n10546), .S(1'b1), .Q(
        fifo[215]) );
  DFFSR fifo_reg_25__10_ ( .D(n3534), .CLK(wclk), .R(n10546), .S(1'b1), .Q(
        fifo[214]) );
  DFFSR fifo_reg_25__9_ ( .D(n3535), .CLK(wclk), .R(n10546), .S(1'b1), .Q(
        fifo[213]) );
  DFFSR fifo_reg_25__8_ ( .D(n3536), .CLK(wclk), .R(n10546), .S(1'b1), .Q(
        fifo[212]) );
  DFFSR fifo_reg_25__7_ ( .D(n3537), .CLK(wclk), .R(n10546), .S(1'b1), .Q(
        fifo[211]) );
  DFFSR fifo_reg_25__6_ ( .D(n3538), .CLK(wclk), .R(n10546), .S(1'b1), .Q(
        fifo[210]) );
  DFFSR fifo_reg_25__5_ ( .D(n3539), .CLK(wclk), .R(n10546), .S(1'b1), .Q(
        fifo[209]) );
  DFFSR fifo_reg_25__4_ ( .D(n3540), .CLK(wclk), .R(n10546), .S(1'b1), .Q(
        fifo[208]) );
  DFFSR fifo_reg_25__3_ ( .D(n3541), .CLK(wclk), .R(n10546), .S(1'b1), .Q(
        fifo[207]) );
  DFFSR fifo_reg_25__2_ ( .D(n3542), .CLK(wclk), .R(n10546), .S(1'b1), .Q(
        fifo[206]) );
  DFFSR fifo_reg_25__1_ ( .D(n3543), .CLK(wclk), .R(n10546), .S(1'b1), .Q(
        fifo[205]) );
  DFFSR fifo_reg_25__0_ ( .D(n3544), .CLK(wclk), .R(n10546), .S(1'b1), .Q(
        fifo[204]) );
  DFFSR fifo_reg_26__33_ ( .D(n3545), .CLK(wclk), .R(n10547), .S(1'b1), .Q(
        fifo[203]) );
  DFFSR fifo_reg_26__32_ ( .D(n3546), .CLK(wclk), .R(n10547), .S(1'b1), .Q(
        fifo[202]) );
  DFFSR fifo_reg_26__31_ ( .D(n3547), .CLK(wclk), .R(n10547), .S(1'b1), .Q(
        fifo[201]) );
  DFFSR fifo_reg_26__30_ ( .D(n3548), .CLK(wclk), .R(n10547), .S(1'b1), .Q(
        fifo[200]) );
  DFFSR fifo_reg_26__29_ ( .D(n3549), .CLK(wclk), .R(n10547), .S(1'b1), .Q(
        fifo[199]) );
  DFFSR fifo_reg_26__28_ ( .D(n3550), .CLK(wclk), .R(n10547), .S(1'b1), .Q(
        fifo[198]) );
  DFFSR fifo_reg_26__27_ ( .D(n3551), .CLK(wclk), .R(n10547), .S(1'b1), .Q(
        fifo[197]) );
  DFFSR fifo_reg_26__26_ ( .D(n3552), .CLK(wclk), .R(n10547), .S(1'b1), .Q(
        fifo[196]) );
  DFFSR fifo_reg_26__25_ ( .D(n3553), .CLK(wclk), .R(n10547), .S(1'b1), .Q(
        fifo[195]) );
  DFFSR fifo_reg_26__24_ ( .D(n3554), .CLK(wclk), .R(n10547), .S(1'b1), .Q(
        fifo[194]) );
  DFFSR fifo_reg_26__23_ ( .D(n3555), .CLK(wclk), .R(n10547), .S(1'b1), .Q(
        fifo[193]) );
  DFFSR fifo_reg_26__22_ ( .D(n3556), .CLK(wclk), .R(n10547), .S(1'b1), .Q(
        fifo[192]) );
  DFFSR fifo_reg_26__21_ ( .D(n3557), .CLK(wclk), .R(n10548), .S(1'b1), .Q(
        fifo[191]) );
  DFFSR fifo_reg_26__20_ ( .D(n3558), .CLK(wclk), .R(n10548), .S(1'b1), .Q(
        fifo[190]) );
  DFFSR fifo_reg_26__19_ ( .D(n3559), .CLK(wclk), .R(n10548), .S(1'b1), .Q(
        fifo[189]) );
  DFFSR fifo_reg_26__18_ ( .D(n3560), .CLK(wclk), .R(n10548), .S(1'b1), .Q(
        fifo[188]) );
  DFFSR fifo_reg_26__17_ ( .D(n3561), .CLK(wclk), .R(n10548), .S(1'b1), .Q(
        fifo[187]) );
  DFFSR fifo_reg_26__16_ ( .D(n3562), .CLK(wclk), .R(n10548), .S(1'b1), .Q(
        fifo[186]) );
  DFFSR fifo_reg_26__15_ ( .D(n3563), .CLK(wclk), .R(n10548), .S(1'b1), .Q(
        fifo[185]) );
  DFFSR fifo_reg_26__14_ ( .D(n3564), .CLK(wclk), .R(n10548), .S(1'b1), .Q(
        fifo[184]) );
  DFFSR fifo_reg_26__13_ ( .D(n3565), .CLK(wclk), .R(n10548), .S(1'b1), .Q(
        fifo[183]) );
  DFFSR fifo_reg_26__12_ ( .D(n3566), .CLK(wclk), .R(n10548), .S(1'b1), .Q(
        fifo[182]) );
  DFFSR fifo_reg_26__11_ ( .D(n3567), .CLK(wclk), .R(n10548), .S(1'b1), .Q(
        fifo[181]) );
  DFFSR fifo_reg_26__10_ ( .D(n3568), .CLK(wclk), .R(n10548), .S(1'b1), .Q(
        fifo[180]) );
  DFFSR fifo_reg_26__9_ ( .D(n3569), .CLK(wclk), .R(n10549), .S(1'b1), .Q(
        fifo[179]) );
  DFFSR fifo_reg_26__8_ ( .D(n3570), .CLK(wclk), .R(n10549), .S(1'b1), .Q(
        fifo[178]) );
  DFFSR fifo_reg_26__7_ ( .D(n3571), .CLK(wclk), .R(n10549), .S(1'b1), .Q(
        fifo[177]) );
  DFFSR fifo_reg_26__6_ ( .D(n3572), .CLK(wclk), .R(n10549), .S(1'b1), .Q(
        fifo[176]) );
  DFFSR fifo_reg_26__5_ ( .D(n3573), .CLK(wclk), .R(n10549), .S(1'b1), .Q(
        fifo[175]) );
  DFFSR fifo_reg_26__4_ ( .D(n3574), .CLK(wclk), .R(n10549), .S(1'b1), .Q(
        fifo[174]) );
  DFFSR fifo_reg_26__3_ ( .D(n3575), .CLK(wclk), .R(n10549), .S(1'b1), .Q(
        fifo[173]) );
  DFFSR fifo_reg_26__2_ ( .D(n3576), .CLK(wclk), .R(n10549), .S(1'b1), .Q(
        fifo[172]) );
  DFFSR fifo_reg_26__1_ ( .D(n3577), .CLK(wclk), .R(n10549), .S(1'b1), .Q(
        fifo[171]) );
  DFFSR fifo_reg_26__0_ ( .D(n3578), .CLK(wclk), .R(n10549), .S(1'b1), .Q(
        fifo[170]) );
  DFFSR fifo_reg_27__33_ ( .D(n3579), .CLK(wclk), .R(n10549), .S(1'b1), .Q(
        fifo[169]) );
  DFFSR fifo_reg_27__32_ ( .D(n3580), .CLK(wclk), .R(n10549), .S(1'b1), .Q(
        fifo[168]) );
  DFFSR fifo_reg_27__31_ ( .D(n3581), .CLK(wclk), .R(n10550), .S(1'b1), .Q(
        fifo[167]) );
  DFFSR fifo_reg_27__30_ ( .D(n3582), .CLK(wclk), .R(n10550), .S(1'b1), .Q(
        fifo[166]) );
  DFFSR fifo_reg_27__29_ ( .D(n3583), .CLK(wclk), .R(n10550), .S(1'b1), .Q(
        fifo[165]) );
  DFFSR fifo_reg_27__28_ ( .D(n3584), .CLK(wclk), .R(n10550), .S(1'b1), .Q(
        fifo[164]) );
  DFFSR fifo_reg_27__27_ ( .D(n3585), .CLK(wclk), .R(n10550), .S(1'b1), .Q(
        fifo[163]) );
  DFFSR fifo_reg_27__26_ ( .D(n3586), .CLK(wclk), .R(n10550), .S(1'b1), .Q(
        fifo[162]) );
  DFFSR fifo_reg_27__25_ ( .D(n3587), .CLK(wclk), .R(n10550), .S(1'b1), .Q(
        fifo[161]) );
  DFFSR fifo_reg_27__24_ ( .D(n3588), .CLK(wclk), .R(n10550), .S(1'b1), .Q(
        fifo[160]) );
  DFFSR fifo_reg_27__23_ ( .D(n3589), .CLK(wclk), .R(n10550), .S(1'b1), .Q(
        fifo[159]) );
  DFFSR fifo_reg_27__22_ ( .D(n3590), .CLK(wclk), .R(n10550), .S(1'b1), .Q(
        fifo[158]) );
  DFFSR fifo_reg_27__21_ ( .D(n3591), .CLK(wclk), .R(n10550), .S(1'b1), .Q(
        fifo[157]) );
  DFFSR fifo_reg_27__20_ ( .D(n3592), .CLK(wclk), .R(n10550), .S(1'b1), .Q(
        fifo[156]) );
  DFFSR fifo_reg_27__19_ ( .D(n3593), .CLK(wclk), .R(n10551), .S(1'b1), .Q(
        fifo[155]) );
  DFFSR fifo_reg_27__18_ ( .D(n3594), .CLK(wclk), .R(n10551), .S(1'b1), .Q(
        fifo[154]) );
  DFFSR fifo_reg_27__17_ ( .D(n3595), .CLK(wclk), .R(n10551), .S(1'b1), .Q(
        fifo[153]) );
  DFFSR fifo_reg_27__16_ ( .D(n3596), .CLK(wclk), .R(n10551), .S(1'b1), .Q(
        fifo[152]) );
  DFFSR fifo_reg_27__15_ ( .D(n3597), .CLK(wclk), .R(n10551), .S(1'b1), .Q(
        fifo[151]) );
  DFFSR fifo_reg_27__14_ ( .D(n3598), .CLK(wclk), .R(n10551), .S(1'b1), .Q(
        fifo[150]) );
  DFFSR fifo_reg_27__13_ ( .D(n3599), .CLK(wclk), .R(n10551), .S(1'b1), .Q(
        fifo[149]) );
  DFFSR fifo_reg_27__12_ ( .D(n3600), .CLK(wclk), .R(n10551), .S(1'b1), .Q(
        fifo[148]) );
  DFFSR fifo_reg_27__11_ ( .D(n3601), .CLK(wclk), .R(n10551), .S(1'b1), .Q(
        fifo[147]) );
  DFFSR fifo_reg_27__10_ ( .D(n3602), .CLK(wclk), .R(n10551), .S(1'b1), .Q(
        fifo[146]) );
  DFFSR fifo_reg_27__9_ ( .D(n3603), .CLK(wclk), .R(n10551), .S(1'b1), .Q(
        fifo[145]) );
  DFFSR fifo_reg_27__8_ ( .D(n3604), .CLK(wclk), .R(n10551), .S(1'b1), .Q(
        fifo[144]) );
  DFFSR fifo_reg_27__7_ ( .D(n3605), .CLK(wclk), .R(n10552), .S(1'b1), .Q(
        fifo[143]) );
  DFFSR fifo_reg_27__6_ ( .D(n3606), .CLK(wclk), .R(n10552), .S(1'b1), .Q(
        fifo[142]) );
  DFFSR fifo_reg_27__5_ ( .D(n3607), .CLK(wclk), .R(n10552), .S(1'b1), .Q(
        fifo[141]) );
  DFFSR fifo_reg_27__4_ ( .D(n3608), .CLK(wclk), .R(n10552), .S(1'b1), .Q(
        fifo[140]) );
  DFFSR fifo_reg_27__3_ ( .D(n3609), .CLK(wclk), .R(n10552), .S(1'b1), .Q(
        fifo[139]) );
  DFFSR fifo_reg_27__2_ ( .D(n3610), .CLK(wclk), .R(n10552), .S(1'b1), .Q(
        fifo[138]) );
  DFFSR fifo_reg_27__1_ ( .D(n3611), .CLK(wclk), .R(n10552), .S(1'b1), .Q(
        fifo[137]) );
  DFFSR fifo_reg_27__0_ ( .D(n3612), .CLK(wclk), .R(n10552), .S(1'b1), .Q(
        fifo[136]) );
  DFFSR fifo_reg_28__33_ ( .D(n3613), .CLK(wclk), .R(n10552), .S(1'b1), .Q(
        fifo[135]) );
  DFFSR fifo_reg_28__32_ ( .D(n3614), .CLK(wclk), .R(n10552), .S(1'b1), .Q(
        fifo[134]) );
  DFFSR fifo_reg_28__31_ ( .D(n3615), .CLK(wclk), .R(n10552), .S(1'b1), .Q(
        fifo[133]) );
  DFFSR fifo_reg_28__30_ ( .D(n3616), .CLK(wclk), .R(n10552), .S(1'b1), .Q(
        fifo[132]) );
  DFFSR fifo_reg_28__29_ ( .D(n3617), .CLK(wclk), .R(n10553), .S(1'b1), .Q(
        fifo[131]) );
  DFFSR fifo_reg_28__28_ ( .D(n3618), .CLK(wclk), .R(n10553), .S(1'b1), .Q(
        fifo[130]) );
  DFFSR fifo_reg_28__27_ ( .D(n3619), .CLK(wclk), .R(n10553), .S(1'b1), .Q(
        fifo[129]) );
  DFFSR fifo_reg_28__26_ ( .D(n3620), .CLK(wclk), .R(n10553), .S(1'b1), .Q(
        fifo[128]) );
  DFFSR fifo_reg_28__25_ ( .D(n3621), .CLK(wclk), .R(n10553), .S(1'b1), .Q(
        fifo[127]) );
  DFFSR fifo_reg_28__24_ ( .D(n3622), .CLK(wclk), .R(n10553), .S(1'b1), .Q(
        fifo[126]) );
  DFFSR fifo_reg_28__23_ ( .D(n3623), .CLK(wclk), .R(n10553), .S(1'b1), .Q(
        fifo[125]) );
  DFFSR fifo_reg_28__22_ ( .D(n3624), .CLK(wclk), .R(n10553), .S(1'b1), .Q(
        fifo[124]) );
  DFFSR fifo_reg_28__21_ ( .D(n3625), .CLK(wclk), .R(n10553), .S(1'b1), .Q(
        fifo[123]) );
  DFFSR fifo_reg_28__20_ ( .D(n3626), .CLK(wclk), .R(n10553), .S(1'b1), .Q(
        fifo[122]) );
  DFFSR fifo_reg_28__19_ ( .D(n3627), .CLK(wclk), .R(n10553), .S(1'b1), .Q(
        fifo[121]) );
  DFFSR fifo_reg_28__18_ ( .D(n3628), .CLK(wclk), .R(n10553), .S(1'b1), .Q(
        fifo[120]) );
  DFFSR fifo_reg_28__17_ ( .D(n3629), .CLK(wclk), .R(n10554), .S(1'b1), .Q(
        fifo[119]) );
  DFFSR fifo_reg_28__16_ ( .D(n3630), .CLK(wclk), .R(n10554), .S(1'b1), .Q(
        fifo[118]) );
  DFFSR fifo_reg_28__15_ ( .D(n3631), .CLK(wclk), .R(n10554), .S(1'b1), .Q(
        fifo[117]) );
  DFFSR fifo_reg_28__14_ ( .D(n3632), .CLK(wclk), .R(n10554), .S(1'b1), .Q(
        fifo[116]) );
  DFFSR fifo_reg_28__13_ ( .D(n3633), .CLK(wclk), .R(n10554), .S(1'b1), .Q(
        fifo[115]) );
  DFFSR fifo_reg_28__12_ ( .D(n3634), .CLK(wclk), .R(n10554), .S(1'b1), .Q(
        fifo[114]) );
  DFFSR fifo_reg_28__11_ ( .D(n3635), .CLK(wclk), .R(n10554), .S(1'b1), .Q(
        fifo[113]) );
  DFFSR fifo_reg_28__10_ ( .D(n3636), .CLK(wclk), .R(n10554), .S(1'b1), .Q(
        fifo[112]) );
  DFFSR fifo_reg_28__9_ ( .D(n3637), .CLK(wclk), .R(n10554), .S(1'b1), .Q(
        fifo[111]) );
  DFFSR fifo_reg_28__8_ ( .D(n3638), .CLK(wclk), .R(n10554), .S(1'b1), .Q(
        fifo[110]) );
  DFFSR fifo_reg_28__7_ ( .D(n3639), .CLK(wclk), .R(n10554), .S(1'b1), .Q(
        fifo[109]) );
  DFFSR fifo_reg_28__6_ ( .D(n3640), .CLK(wclk), .R(n10554), .S(1'b1), .Q(
        fifo[108]) );
  DFFSR fifo_reg_28__5_ ( .D(n3641), .CLK(wclk), .R(n10555), .S(1'b1), .Q(
        fifo[107]) );
  DFFSR fifo_reg_28__4_ ( .D(n3642), .CLK(wclk), .R(n10555), .S(1'b1), .Q(
        fifo[106]) );
  DFFSR fifo_reg_28__3_ ( .D(n3643), .CLK(wclk), .R(n10555), .S(1'b1), .Q(
        fifo[105]) );
  DFFSR fifo_reg_28__2_ ( .D(n3644), .CLK(wclk), .R(n10555), .S(1'b1), .Q(
        fifo[104]) );
  DFFSR fifo_reg_28__1_ ( .D(n3645), .CLK(wclk), .R(n10555), .S(1'b1), .Q(
        fifo[103]) );
  DFFSR fifo_reg_28__0_ ( .D(n3646), .CLK(wclk), .R(n10555), .S(1'b1), .Q(
        fifo[102]) );
  DFFSR fifo_reg_29__33_ ( .D(n3647), .CLK(wclk), .R(n10555), .S(1'b1), .Q(
        fifo[101]) );
  DFFSR fifo_reg_29__32_ ( .D(n3648), .CLK(wclk), .R(n10555), .S(1'b1), .Q(
        fifo[100]) );
  DFFSR fifo_reg_29__31_ ( .D(n3649), .CLK(wclk), .R(n10555), .S(1'b1), .Q(
        fifo[99]) );
  DFFSR fifo_reg_29__30_ ( .D(n3650), .CLK(wclk), .R(n10555), .S(1'b1), .Q(
        fifo[98]) );
  DFFSR fifo_reg_29__29_ ( .D(n3651), .CLK(wclk), .R(n10555), .S(1'b1), .Q(
        fifo[97]) );
  DFFSR fifo_reg_29__28_ ( .D(n3652), .CLK(wclk), .R(n10555), .S(1'b1), .Q(
        fifo[96]) );
  DFFSR fifo_reg_29__27_ ( .D(n3653), .CLK(wclk), .R(n10556), .S(1'b1), .Q(
        fifo[95]) );
  DFFSR fifo_reg_29__26_ ( .D(n3654), .CLK(wclk), .R(n10556), .S(1'b1), .Q(
        fifo[94]) );
  DFFSR fifo_reg_29__25_ ( .D(n3655), .CLK(wclk), .R(n10556), .S(1'b1), .Q(
        fifo[93]) );
  DFFSR fifo_reg_29__24_ ( .D(n3656), .CLK(wclk), .R(n10556), .S(1'b1), .Q(
        fifo[92]) );
  DFFSR fifo_reg_29__23_ ( .D(n3657), .CLK(wclk), .R(n10556), .S(1'b1), .Q(
        fifo[91]) );
  DFFSR fifo_reg_29__22_ ( .D(n3658), .CLK(wclk), .R(n10556), .S(1'b1), .Q(
        fifo[90]) );
  DFFSR fifo_reg_29__21_ ( .D(n3659), .CLK(wclk), .R(n10556), .S(1'b1), .Q(
        fifo[89]) );
  DFFSR fifo_reg_29__20_ ( .D(n3660), .CLK(wclk), .R(n10556), .S(1'b1), .Q(
        fifo[88]) );
  DFFSR fifo_reg_29__19_ ( .D(n3661), .CLK(wclk), .R(n10556), .S(1'b1), .Q(
        fifo[87]) );
  DFFSR fifo_reg_29__18_ ( .D(n3662), .CLK(wclk), .R(n10556), .S(1'b1), .Q(
        fifo[86]) );
  DFFSR fifo_reg_29__17_ ( .D(n3663), .CLK(wclk), .R(n10556), .S(1'b1), .Q(
        fifo[85]) );
  DFFSR fifo_reg_29__16_ ( .D(n3664), .CLK(wclk), .R(n10556), .S(1'b1), .Q(
        fifo[84]) );
  DFFSR fifo_reg_29__15_ ( .D(n3665), .CLK(wclk), .R(n10557), .S(1'b1), .Q(
        fifo[83]) );
  DFFSR fifo_reg_29__14_ ( .D(n3666), .CLK(wclk), .R(n10557), .S(1'b1), .Q(
        fifo[82]) );
  DFFSR fifo_reg_29__13_ ( .D(n3667), .CLK(wclk), .R(n10557), .S(1'b1), .Q(
        fifo[81]) );
  DFFSR fifo_reg_29__12_ ( .D(n3668), .CLK(wclk), .R(n10557), .S(1'b1), .Q(
        fifo[80]) );
  DFFSR fifo_reg_29__11_ ( .D(n3669), .CLK(wclk), .R(n10557), .S(1'b1), .Q(
        fifo[79]) );
  DFFSR fifo_reg_29__10_ ( .D(n3670), .CLK(wclk), .R(n10557), .S(1'b1), .Q(
        fifo[78]) );
  DFFSR fifo_reg_29__9_ ( .D(n3671), .CLK(wclk), .R(n10557), .S(1'b1), .Q(
        fifo[77]) );
  DFFSR fifo_reg_29__8_ ( .D(n3672), .CLK(wclk), .R(n10557), .S(1'b1), .Q(
        fifo[76]) );
  DFFSR fifo_reg_29__7_ ( .D(n3673), .CLK(wclk), .R(n10557), .S(1'b1), .Q(
        fifo[75]) );
  DFFSR fifo_reg_29__6_ ( .D(n3674), .CLK(wclk), .R(n10557), .S(1'b1), .Q(
        fifo[74]) );
  DFFSR fifo_reg_29__5_ ( .D(n3675), .CLK(wclk), .R(n10557), .S(1'b1), .Q(
        fifo[73]) );
  DFFSR fifo_reg_29__4_ ( .D(n3676), .CLK(wclk), .R(n10557), .S(1'b1), .Q(
        fifo[72]) );
  DFFSR fifo_reg_29__3_ ( .D(n3677), .CLK(wclk), .R(n10558), .S(1'b1), .Q(
        fifo[71]) );
  DFFSR fifo_reg_29__2_ ( .D(n3678), .CLK(wclk), .R(n10558), .S(1'b1), .Q(
        fifo[70]) );
  DFFSR fifo_reg_29__1_ ( .D(n3679), .CLK(wclk), .R(n10558), .S(1'b1), .Q(
        fifo[69]) );
  DFFSR fifo_reg_29__0_ ( .D(n3680), .CLK(wclk), .R(n10558), .S(1'b1), .Q(
        fifo[68]) );
  DFFSR fifo_reg_30__33_ ( .D(n3681), .CLK(wclk), .R(n10558), .S(1'b1), .Q(
        fifo[67]) );
  DFFSR fifo_reg_30__32_ ( .D(n3682), .CLK(wclk), .R(n10558), .S(1'b1), .Q(
        fifo[66]) );
  DFFSR fifo_reg_30__31_ ( .D(n3683), .CLK(wclk), .R(n10558), .S(1'b1), .Q(
        fifo[65]) );
  DFFSR fifo_reg_30__30_ ( .D(n3684), .CLK(wclk), .R(n10558), .S(1'b1), .Q(
        fifo[64]) );
  DFFSR fifo_reg_30__29_ ( .D(n3685), .CLK(wclk), .R(n10558), .S(1'b1), .Q(
        fifo[63]) );
  DFFSR fifo_reg_30__28_ ( .D(n3686), .CLK(wclk), .R(n10558), .S(1'b1), .Q(
        fifo[62]) );
  DFFSR fifo_reg_30__27_ ( .D(n3687), .CLK(wclk), .R(n10558), .S(1'b1), .Q(
        fifo[61]) );
  DFFSR fifo_reg_30__26_ ( .D(n3688), .CLK(wclk), .R(n10558), .S(1'b1), .Q(
        fifo[60]) );
  DFFSR fifo_reg_30__25_ ( .D(n3689), .CLK(wclk), .R(n10559), .S(1'b1), .Q(
        fifo[59]) );
  DFFSR fifo_reg_30__24_ ( .D(n3690), .CLK(wclk), .R(n10559), .S(1'b1), .Q(
        fifo[58]) );
  DFFSR fifo_reg_30__23_ ( .D(n3691), .CLK(wclk), .R(n10559), .S(1'b1), .Q(
        fifo[57]) );
  DFFSR fifo_reg_30__22_ ( .D(n3692), .CLK(wclk), .R(n10559), .S(1'b1), .Q(
        fifo[56]) );
  DFFSR fifo_reg_30__21_ ( .D(n3693), .CLK(wclk), .R(n10559), .S(1'b1), .Q(
        fifo[55]) );
  DFFSR fifo_reg_30__20_ ( .D(n3694), .CLK(wclk), .R(n10559), .S(1'b1), .Q(
        fifo[54]) );
  DFFSR fifo_reg_30__19_ ( .D(n3695), .CLK(wclk), .R(n10559), .S(1'b1), .Q(
        fifo[53]) );
  DFFSR fifo_reg_30__18_ ( .D(n3696), .CLK(wclk), .R(n10559), .S(1'b1), .Q(
        fifo[52]) );
  DFFSR fifo_reg_30__17_ ( .D(n3697), .CLK(wclk), .R(n10559), .S(1'b1), .Q(
        fifo[51]) );
  DFFSR fifo_reg_30__16_ ( .D(n3698), .CLK(wclk), .R(n10559), .S(1'b1), .Q(
        fifo[50]) );
  DFFSR fifo_reg_30__15_ ( .D(n3699), .CLK(wclk), .R(n10559), .S(1'b1), .Q(
        fifo[49]) );
  DFFSR fifo_reg_30__14_ ( .D(n3700), .CLK(wclk), .R(n10559), .S(1'b1), .Q(
        fifo[48]) );
  DFFSR fifo_reg_30__13_ ( .D(n3701), .CLK(wclk), .R(n10560), .S(1'b1), .Q(
        fifo[47]) );
  DFFSR fifo_reg_30__12_ ( .D(n3702), .CLK(wclk), .R(n10560), .S(1'b1), .Q(
        fifo[46]) );
  DFFSR fifo_reg_30__11_ ( .D(n3703), .CLK(wclk), .R(n10560), .S(1'b1), .Q(
        fifo[45]) );
  DFFSR fifo_reg_30__10_ ( .D(n3704), .CLK(wclk), .R(n10560), .S(1'b1), .Q(
        fifo[44]) );
  DFFSR fifo_reg_30__9_ ( .D(n3705), .CLK(wclk), .R(n10560), .S(1'b1), .Q(
        fifo[43]) );
  DFFSR fifo_reg_30__8_ ( .D(n3706), .CLK(wclk), .R(n10560), .S(1'b1), .Q(
        fifo[42]) );
  DFFSR fifo_reg_30__7_ ( .D(n3707), .CLK(wclk), .R(n10560), .S(1'b1), .Q(
        fifo[41]) );
  DFFSR fifo_reg_30__6_ ( .D(n3708), .CLK(wclk), .R(n10560), .S(1'b1), .Q(
        fifo[40]) );
  DFFSR fifo_reg_30__5_ ( .D(n3709), .CLK(wclk), .R(n10560), .S(1'b1), .Q(
        fifo[39]) );
  DFFSR fifo_reg_30__4_ ( .D(n3710), .CLK(wclk), .R(n10560), .S(1'b1), .Q(
        fifo[38]) );
  DFFSR fifo_reg_30__3_ ( .D(n3711), .CLK(wclk), .R(n10560), .S(1'b1), .Q(
        fifo[37]) );
  DFFSR fifo_reg_30__2_ ( .D(n3712), .CLK(wclk), .R(n10560), .S(1'b1), .Q(
        fifo[36]) );
  DFFSR fifo_reg_30__1_ ( .D(n3713), .CLK(wclk), .R(n10561), .S(1'b1), .Q(
        fifo[35]) );
  DFFSR fifo_reg_30__0_ ( .D(n3714), .CLK(wclk), .R(n10561), .S(1'b1), .Q(
        fifo[34]) );
  DFFSR fifo_reg_31__33_ ( .D(n3715), .CLK(wclk), .R(n10561), .S(1'b1), .Q(
        fifo[33]) );
  DFFSR fifo_reg_31__32_ ( .D(n3716), .CLK(wclk), .R(n10561), .S(1'b1), .Q(
        fifo[32]) );
  DFFSR fifo_reg_31__31_ ( .D(n3717), .CLK(wclk), .R(n10561), .S(1'b1), .Q(
        fifo[31]) );
  DFFSR fifo_reg_31__30_ ( .D(n3718), .CLK(wclk), .R(n10561), .S(1'b1), .Q(
        fifo[30]) );
  DFFSR fifo_reg_31__29_ ( .D(n3719), .CLK(wclk), .R(n10561), .S(1'b1), .Q(
        fifo[29]) );
  DFFSR fifo_reg_31__28_ ( .D(n3720), .CLK(wclk), .R(n10561), .S(1'b1), .Q(
        fifo[28]) );
  DFFSR fifo_reg_31__27_ ( .D(n3721), .CLK(wclk), .R(n10561), .S(1'b1), .Q(
        fifo[27]) );
  DFFSR fifo_reg_31__26_ ( .D(n3722), .CLK(wclk), .R(n10561), .S(1'b1), .Q(
        fifo[26]) );
  DFFSR fifo_reg_31__25_ ( .D(n3723), .CLK(wclk), .R(n10561), .S(1'b1), .Q(
        fifo[25]) );
  DFFSR fifo_reg_31__24_ ( .D(n3724), .CLK(wclk), .R(n10561), .S(1'b1), .Q(
        fifo[24]) );
  DFFSR fifo_reg_31__23_ ( .D(n3725), .CLK(wclk), .R(n10562), .S(1'b1), .Q(
        fifo[23]) );
  DFFSR fifo_reg_31__22_ ( .D(n3726), .CLK(wclk), .R(n10562), .S(1'b1), .Q(
        fifo[22]) );
  DFFSR fifo_reg_31__21_ ( .D(n3727), .CLK(wclk), .R(n10562), .S(1'b1), .Q(
        fifo[21]) );
  DFFSR fifo_reg_31__20_ ( .D(n3728), .CLK(wclk), .R(n10562), .S(1'b1), .Q(
        fifo[20]) );
  DFFSR fifo_reg_31__19_ ( .D(n3729), .CLK(wclk), .R(n10562), .S(1'b1), .Q(
        fifo[19]) );
  DFFSR fifo_reg_31__18_ ( .D(n3730), .CLK(wclk), .R(n10562), .S(1'b1), .Q(
        fifo[18]) );
  DFFSR fifo_reg_31__17_ ( .D(n3731), .CLK(wclk), .R(n10562), .S(1'b1), .Q(
        fifo[17]) );
  DFFSR fifo_reg_31__16_ ( .D(n3732), .CLK(wclk), .R(n10562), .S(1'b1), .Q(
        fifo[16]) );
  DFFSR fifo_reg_31__15_ ( .D(n3733), .CLK(wclk), .R(n10562), .S(1'b1), .Q(
        fifo[15]) );
  DFFSR fifo_reg_31__14_ ( .D(n3734), .CLK(wclk), .R(n10562), .S(1'b1), .Q(
        fifo[14]) );
  DFFSR fifo_reg_31__13_ ( .D(n3735), .CLK(wclk), .R(n10562), .S(1'b1), .Q(
        fifo[13]) );
  DFFSR fifo_reg_31__12_ ( .D(n3736), .CLK(wclk), .R(n10562), .S(1'b1), .Q(
        fifo[12]) );
  DFFSR fifo_reg_31__11_ ( .D(n3737), .CLK(wclk), .R(n10563), .S(1'b1), .Q(
        fifo[11]) );
  DFFSR fifo_reg_31__10_ ( .D(n3738), .CLK(wclk), .R(n10563), .S(1'b1), .Q(
        fifo[10]) );
  DFFSR fifo_reg_31__9_ ( .D(n3739), .CLK(wclk), .R(n10563), .S(1'b1), .Q(
        fifo[9]) );
  DFFSR fifo_reg_31__8_ ( .D(n3740), .CLK(wclk), .R(n10563), .S(1'b1), .Q(
        fifo[8]) );
  DFFSR fifo_reg_31__7_ ( .D(n3741), .CLK(wclk), .R(n10563), .S(1'b1), .Q(
        fifo[7]) );
  DFFSR fifo_reg_31__6_ ( .D(n3742), .CLK(wclk), .R(n10563), .S(1'b1), .Q(
        fifo[6]) );
  DFFSR fifo_reg_31__5_ ( .D(n3743), .CLK(wclk), .R(n10563), .S(1'b1), .Q(
        fifo[5]) );
  DFFSR fifo_reg_31__4_ ( .D(n3744), .CLK(wclk), .R(n10563), .S(1'b1), .Q(
        fifo[4]) );
  DFFSR fifo_reg_31__3_ ( .D(n3745), .CLK(wclk), .R(n10563), .S(1'b1), .Q(
        fifo[3]) );
  DFFSR fifo_reg_31__2_ ( .D(n3746), .CLK(wclk), .R(n10563), .S(1'b1), .Q(
        fifo[2]) );
  DFFSR fifo_reg_31__1_ ( .D(n3747), .CLK(wclk), .R(n10563), .S(1'b1), .Q(
        fifo[1]) );
  DFFSR fifo_reg_31__0_ ( .D(n3748), .CLK(wclk), .R(n10563), .S(1'b1), .Q(
        fifo[0]) );
  XOR2X1 U3 ( .A(rd_ptr_bin_ss[1]), .B(n6693), .Y(rd_ptr_bin_ss[0]) );
  OAI21X1 U9 ( .A(n193), .B(n194), .C(n6678), .Y(n2536) );
  OAI21X1 U12 ( .A(n193), .B(n10536), .C(n6675), .Y(n2541) );
  OAI21X1 U15 ( .A(n193), .B(n10658), .C(n6672), .Y(n2546) );
  OAI21X1 U17 ( .A(n193), .B(n10680), .C(n6669), .Y(n2551) );
  INVX1 U19 ( .A(n202), .Y(n2553) );
  AOI22X1 U20 ( .A(data_out[33]), .B(n10108), .C(n71), .D(n193), .Y(n202) );
  INVX1 U21 ( .A(n204), .Y(n2555) );
  AOI22X1 U22 ( .A(data_out[32]), .B(n10108), .C(n72), .D(n193), .Y(n204) );
  INVX1 U23 ( .A(n205), .Y(n2557) );
  AOI22X1 U24 ( .A(data_out[31]), .B(n10108), .C(n73), .D(n193), .Y(n205) );
  INVX1 U25 ( .A(n206), .Y(n2559) );
  AOI22X1 U26 ( .A(data_out[30]), .B(n10108), .C(n74), .D(n193), .Y(n206) );
  INVX1 U27 ( .A(n207), .Y(n2561) );
  AOI22X1 U28 ( .A(data_out[29]), .B(n10108), .C(n75), .D(n193), .Y(n207) );
  INVX1 U29 ( .A(n208), .Y(n2563) );
  AOI22X1 U30 ( .A(data_out[28]), .B(n10108), .C(n76), .D(n193), .Y(n208) );
  INVX1 U31 ( .A(n209), .Y(n2565) );
  AOI22X1 U32 ( .A(data_out[27]), .B(n10108), .C(n77), .D(n193), .Y(n209) );
  INVX1 U33 ( .A(n210), .Y(n2567) );
  AOI22X1 U34 ( .A(data_out[26]), .B(n10108), .C(n78), .D(n193), .Y(n210) );
  INVX1 U35 ( .A(n211), .Y(n2569) );
  AOI22X1 U36 ( .A(data_out[25]), .B(n10108), .C(n79), .D(n193), .Y(n211) );
  INVX1 U37 ( .A(n212), .Y(n2571) );
  AOI22X1 U38 ( .A(data_out[24]), .B(n10108), .C(n80), .D(n193), .Y(n212) );
  INVX1 U39 ( .A(n213), .Y(n2573) );
  AOI22X1 U40 ( .A(data_out[23]), .B(n10108), .C(n81), .D(n193), .Y(n213) );
  INVX1 U41 ( .A(n214), .Y(n2575) );
  AOI22X1 U42 ( .A(data_out[22]), .B(n10108), .C(n82), .D(n193), .Y(n214) );
  INVX1 U43 ( .A(n215), .Y(n2577) );
  AOI22X1 U44 ( .A(data_out[21]), .B(n10108), .C(n83), .D(n193), .Y(n215) );
  INVX1 U45 ( .A(n216), .Y(n2579) );
  AOI22X1 U46 ( .A(data_out[20]), .B(n10108), .C(n84), .D(n193), .Y(n216) );
  INVX1 U47 ( .A(n217), .Y(n2581) );
  AOI22X1 U48 ( .A(data_out[19]), .B(n10108), .C(n85), .D(n193), .Y(n217) );
  INVX1 U49 ( .A(n218), .Y(n2583) );
  AOI22X1 U50 ( .A(data_out[18]), .B(n10108), .C(n86), .D(n193), .Y(n218) );
  INVX1 U51 ( .A(n219), .Y(n2585) );
  AOI22X1 U52 ( .A(data_out[17]), .B(n10108), .C(n87), .D(n193), .Y(n219) );
  INVX1 U53 ( .A(n220), .Y(n2587) );
  AOI22X1 U54 ( .A(data_out[16]), .B(n10108), .C(n88), .D(n193), .Y(n220) );
  INVX1 U55 ( .A(n221), .Y(n2589) );
  AOI22X1 U56 ( .A(data_out[15]), .B(n10108), .C(n89), .D(n193), .Y(n221) );
  INVX1 U57 ( .A(n222), .Y(n2591) );
  AOI22X1 U58 ( .A(data_out[14]), .B(n10108), .C(n90), .D(n193), .Y(n222) );
  INVX1 U59 ( .A(n223), .Y(n2593) );
  AOI22X1 U60 ( .A(data_out[13]), .B(n10108), .C(n91), .D(n193), .Y(n223) );
  INVX1 U61 ( .A(n224), .Y(n2595) );
  AOI22X1 U62 ( .A(data_out[12]), .B(n10108), .C(n92), .D(n193), .Y(n224) );
  INVX1 U63 ( .A(n225), .Y(n2597) );
  AOI22X1 U64 ( .A(data_out[11]), .B(n10108), .C(n93), .D(n193), .Y(n225) );
  INVX1 U65 ( .A(n226), .Y(n2599) );
  AOI22X1 U66 ( .A(data_out[10]), .B(n10108), .C(n94), .D(n193), .Y(n226) );
  INVX1 U67 ( .A(n227), .Y(n2601) );
  AOI22X1 U68 ( .A(data_out[9]), .B(n10108), .C(n95), .D(n193), .Y(n227) );
  INVX1 U69 ( .A(n228), .Y(n2603) );
  AOI22X1 U70 ( .A(data_out[8]), .B(n10108), .C(n96), .D(n193), .Y(n228) );
  INVX1 U71 ( .A(n229), .Y(n2605) );
  AOI22X1 U72 ( .A(data_out[7]), .B(n10108), .C(n97), .D(n193), .Y(n229) );
  INVX1 U73 ( .A(n230), .Y(n2607) );
  AOI22X1 U74 ( .A(data_out[6]), .B(n10108), .C(n98), .D(n193), .Y(n230) );
  INVX1 U75 ( .A(n231), .Y(n2609) );
  AOI22X1 U76 ( .A(data_out[5]), .B(n10108), .C(n99), .D(n193), .Y(n231) );
  INVX1 U77 ( .A(n232), .Y(n2611) );
  AOI22X1 U78 ( .A(data_out[4]), .B(n10108), .C(n100), .D(n193), .Y(n232) );
  INVX1 U79 ( .A(n233), .Y(n2613) );
  AOI22X1 U80 ( .A(data_out[3]), .B(n10108), .C(n101), .D(n193), .Y(n233) );
  INVX1 U81 ( .A(n234), .Y(n2615) );
  AOI22X1 U82 ( .A(data_out[2]), .B(n10108), .C(n102), .D(n193), .Y(n234) );
  INVX1 U83 ( .A(n235), .Y(n2617) );
  AOI22X1 U84 ( .A(data_out[1]), .B(n10108), .C(n103), .D(n193), .Y(n235) );
  INVX1 U85 ( .A(n236), .Y(n2619) );
  AOI22X1 U86 ( .A(data_out[0]), .B(n10108), .C(n104), .D(n193), .Y(n236) );
  OAI21X1 U87 ( .A(n237), .B(n238), .C(n6666), .Y(n2627) );
  OAI21X1 U89 ( .A(n237), .B(n240), .C(n6663), .Y(n2632) );
  OAI21X1 U91 ( .A(n237), .B(n242), .C(n6660), .Y(n2637) );
  OAI21X1 U93 ( .A(n237), .B(n244), .C(n6657), .Y(n2642) );
  OAI21X1 U95 ( .A(n237), .B(n246), .C(n6654), .Y(n2644) );
  OAI21X1 U97 ( .A(n237), .B(n248), .C(n6651), .Y(n2649) );
  INVX1 U99 ( .A(n10081), .Y(n248) );
  OAI21X1 U100 ( .A(n193), .B(n250), .C(n6648), .Y(n2657) );
  OAI21X1 U103 ( .A(n193), .B(n10722), .C(n6645), .Y(n2660) );
  INVX1 U105 ( .A(n10107), .Y(n193) );
  OAI21X1 U107 ( .A(n10113), .B(n255), .C(n6642), .Y(n2661) );
  OAI21X1 U109 ( .A(n10113), .B(n257), .C(n6639), .Y(n2662) );
  OAI21X1 U111 ( .A(n10113), .B(n259), .C(n6636), .Y(n2663) );
  OAI21X1 U113 ( .A(n10113), .B(n261), .C(n6633), .Y(n2664) );
  OAI21X1 U115 ( .A(n10113), .B(n263), .C(n6630), .Y(n2665) );
  OAI21X1 U117 ( .A(n10113), .B(n265), .C(n6627), .Y(n2666) );
  OAI21X1 U119 ( .A(n10113), .B(n267), .C(n6624), .Y(n2667) );
  OAI21X1 U121 ( .A(n10113), .B(n269), .C(n6621), .Y(n2668) );
  OAI21X1 U123 ( .A(n10113), .B(n271), .C(n6618), .Y(n2669) );
  OAI21X1 U125 ( .A(n10113), .B(n273), .C(n6615), .Y(n2670) );
  OAI21X1 U127 ( .A(n10113), .B(n275), .C(n6612), .Y(n2671) );
  OAI21X1 U129 ( .A(n10113), .B(n277), .C(n6609), .Y(n2672) );
  OAI21X1 U131 ( .A(n10113), .B(n279), .C(n6606), .Y(n2673) );
  OAI21X1 U133 ( .A(n10113), .B(n281), .C(n6603), .Y(n2674) );
  OAI21X1 U135 ( .A(n10113), .B(n283), .C(n6600), .Y(n2675) );
  OAI21X1 U137 ( .A(n10113), .B(n285), .C(n6597), .Y(n2676) );
  OAI21X1 U139 ( .A(n10113), .B(n287), .C(n6594), .Y(n2677) );
  OAI21X1 U141 ( .A(n10113), .B(n289), .C(n6591), .Y(n2678) );
  OAI21X1 U143 ( .A(n10113), .B(n291), .C(n6588), .Y(n2679) );
  OAI21X1 U145 ( .A(n10113), .B(n293), .C(n6585), .Y(n2680) );
  OAI21X1 U147 ( .A(n10113), .B(n295), .C(n6582), .Y(n2681) );
  OAI21X1 U149 ( .A(n10113), .B(n297), .C(n6579), .Y(n2682) );
  OAI21X1 U151 ( .A(n10113), .B(n299), .C(n6576), .Y(n2683) );
  OAI21X1 U153 ( .A(n10113), .B(n301), .C(n6573), .Y(n2684) );
  OAI21X1 U155 ( .A(n10113), .B(n303), .C(n6570), .Y(n2685) );
  OAI21X1 U157 ( .A(n10113), .B(n305), .C(n6567), .Y(n2686) );
  OAI21X1 U159 ( .A(n10113), .B(n307), .C(n6564), .Y(n2687) );
  OAI21X1 U161 ( .A(n10113), .B(n309), .C(n6561), .Y(n2688) );
  OAI21X1 U163 ( .A(n10113), .B(n311), .C(n6558), .Y(n2689) );
  OAI21X1 U165 ( .A(n10113), .B(n313), .C(n6555), .Y(n2690) );
  OAI21X1 U167 ( .A(n10113), .B(n315), .C(n6552), .Y(n2691) );
  OAI21X1 U169 ( .A(n10113), .B(n317), .C(n6549), .Y(n2692) );
  OAI21X1 U171 ( .A(n10113), .B(n319), .C(n6546), .Y(n2693) );
  OAI21X1 U173 ( .A(n10113), .B(n321), .C(n6543), .Y(n2694) );
  OAI21X1 U176 ( .A(n255), .B(n325), .C(n6540), .Y(n2695) );
  OAI21X1 U178 ( .A(n257), .B(n325), .C(n6537), .Y(n2696) );
  OAI21X1 U180 ( .A(n259), .B(n325), .C(n6534), .Y(n2697) );
  OAI21X1 U182 ( .A(n261), .B(n325), .C(n6531), .Y(n2698) );
  OAI21X1 U184 ( .A(n263), .B(n325), .C(n6528), .Y(n2699) );
  OAI21X1 U186 ( .A(n265), .B(n325), .C(n6525), .Y(n2700) );
  OAI21X1 U188 ( .A(n267), .B(n325), .C(n6522), .Y(n2701) );
  OAI21X1 U190 ( .A(n269), .B(n325), .C(n6519), .Y(n2702) );
  OAI21X1 U192 ( .A(n271), .B(n325), .C(n6516), .Y(n2703) );
  OAI21X1 U194 ( .A(n273), .B(n325), .C(n6513), .Y(n2704) );
  OAI21X1 U196 ( .A(n275), .B(n325), .C(n6510), .Y(n2705) );
  OAI21X1 U198 ( .A(n277), .B(n325), .C(n6507), .Y(n2706) );
  OAI21X1 U200 ( .A(n279), .B(n325), .C(n6504), .Y(n2707) );
  OAI21X1 U202 ( .A(n281), .B(n325), .C(n6501), .Y(n2708) );
  OAI21X1 U204 ( .A(n283), .B(n325), .C(n6498), .Y(n2709) );
  OAI21X1 U206 ( .A(n285), .B(n325), .C(n6495), .Y(n2710) );
  OAI21X1 U208 ( .A(n287), .B(n325), .C(n6492), .Y(n2711) );
  OAI21X1 U210 ( .A(n289), .B(n325), .C(n6489), .Y(n2712) );
  OAI21X1 U212 ( .A(n291), .B(n325), .C(n6486), .Y(n2713) );
  OAI21X1 U214 ( .A(n293), .B(n325), .C(n6483), .Y(n2714) );
  OAI21X1 U216 ( .A(n295), .B(n325), .C(n6480), .Y(n2715) );
  OAI21X1 U218 ( .A(n297), .B(n325), .C(n6477), .Y(n2716) );
  OAI21X1 U220 ( .A(n299), .B(n325), .C(n6474), .Y(n2717) );
  OAI21X1 U222 ( .A(n301), .B(n325), .C(n6471), .Y(n2718) );
  OAI21X1 U224 ( .A(n303), .B(n325), .C(n6468), .Y(n2719) );
  OAI21X1 U226 ( .A(n305), .B(n325), .C(n6465), .Y(n2720) );
  OAI21X1 U228 ( .A(n307), .B(n325), .C(n6462), .Y(n2721) );
  OAI21X1 U230 ( .A(n309), .B(n325), .C(n6459), .Y(n2722) );
  OAI21X1 U232 ( .A(n311), .B(n325), .C(n6456), .Y(n2723) );
  OAI21X1 U234 ( .A(n313), .B(n325), .C(n6453), .Y(n2724) );
  OAI21X1 U236 ( .A(n315), .B(n325), .C(n6450), .Y(n2725) );
  OAI21X1 U238 ( .A(n317), .B(n325), .C(n6447), .Y(n2726) );
  OAI21X1 U240 ( .A(n319), .B(n325), .C(n6444), .Y(n2727) );
  OAI21X1 U242 ( .A(n321), .B(n325), .C(n6441), .Y(n2728) );
  OAI21X1 U245 ( .A(n255), .B(n361), .C(n6438), .Y(n2729) );
  OAI21X1 U247 ( .A(n257), .B(n361), .C(n6435), .Y(n2730) );
  OAI21X1 U249 ( .A(n259), .B(n361), .C(n6432), .Y(n2731) );
  OAI21X1 U251 ( .A(n261), .B(n361), .C(n6429), .Y(n2732) );
  OAI21X1 U253 ( .A(n263), .B(n361), .C(n6426), .Y(n2733) );
  OAI21X1 U255 ( .A(n265), .B(n361), .C(n6423), .Y(n2734) );
  OAI21X1 U257 ( .A(n267), .B(n361), .C(n6420), .Y(n2735) );
  OAI21X1 U259 ( .A(n269), .B(n361), .C(n6417), .Y(n2736) );
  OAI21X1 U261 ( .A(n271), .B(n361), .C(n6414), .Y(n2737) );
  OAI21X1 U263 ( .A(n273), .B(n361), .C(n6411), .Y(n2738) );
  OAI21X1 U265 ( .A(n275), .B(n361), .C(n6408), .Y(n2739) );
  OAI21X1 U267 ( .A(n277), .B(n361), .C(n6405), .Y(n2740) );
  OAI21X1 U269 ( .A(n279), .B(n361), .C(n6402), .Y(n2741) );
  OAI21X1 U271 ( .A(n281), .B(n361), .C(n6399), .Y(n2742) );
  OAI21X1 U273 ( .A(n283), .B(n361), .C(n6396), .Y(n2743) );
  OAI21X1 U275 ( .A(n285), .B(n361), .C(n6393), .Y(n2744) );
  OAI21X1 U277 ( .A(n287), .B(n361), .C(n6390), .Y(n2745) );
  OAI21X1 U279 ( .A(n289), .B(n361), .C(n6387), .Y(n2746) );
  OAI21X1 U281 ( .A(n291), .B(n361), .C(n6384), .Y(n2747) );
  OAI21X1 U283 ( .A(n293), .B(n361), .C(n6381), .Y(n2748) );
  OAI21X1 U285 ( .A(n295), .B(n361), .C(n6378), .Y(n2749) );
  OAI21X1 U287 ( .A(n297), .B(n361), .C(n6375), .Y(n2750) );
  OAI21X1 U289 ( .A(n299), .B(n361), .C(n6372), .Y(n2751) );
  OAI21X1 U291 ( .A(n301), .B(n361), .C(n6369), .Y(n2752) );
  OAI21X1 U293 ( .A(n303), .B(n361), .C(n6366), .Y(n2753) );
  OAI21X1 U295 ( .A(n305), .B(n361), .C(n6363), .Y(n2754) );
  OAI21X1 U297 ( .A(n307), .B(n361), .C(n6360), .Y(n2755) );
  OAI21X1 U299 ( .A(n309), .B(n361), .C(n6357), .Y(n2756) );
  OAI21X1 U301 ( .A(n311), .B(n361), .C(n6354), .Y(n2757) );
  OAI21X1 U303 ( .A(n313), .B(n361), .C(n6351), .Y(n2758) );
  OAI21X1 U305 ( .A(n315), .B(n361), .C(n6348), .Y(n2759) );
  OAI21X1 U307 ( .A(n317), .B(n361), .C(n6345), .Y(n2760) );
  OAI21X1 U309 ( .A(n319), .B(n361), .C(n6342), .Y(n2761) );
  OAI21X1 U311 ( .A(n321), .B(n361), .C(n6339), .Y(n2762) );
  OAI21X1 U314 ( .A(n255), .B(n397), .C(n6336), .Y(n2763) );
  OAI21X1 U316 ( .A(n257), .B(n397), .C(n6333), .Y(n2764) );
  OAI21X1 U318 ( .A(n259), .B(n397), .C(n6330), .Y(n2765) );
  OAI21X1 U320 ( .A(n261), .B(n397), .C(n6327), .Y(n2766) );
  OAI21X1 U322 ( .A(n263), .B(n397), .C(n6324), .Y(n2767) );
  OAI21X1 U324 ( .A(n265), .B(n397), .C(n6321), .Y(n2768) );
  OAI21X1 U326 ( .A(n267), .B(n397), .C(n6318), .Y(n2769) );
  OAI21X1 U328 ( .A(n269), .B(n397), .C(n6315), .Y(n2770) );
  OAI21X1 U330 ( .A(n271), .B(n397), .C(n6312), .Y(n2771) );
  OAI21X1 U332 ( .A(n273), .B(n397), .C(n6309), .Y(n2772) );
  OAI21X1 U334 ( .A(n275), .B(n397), .C(n6306), .Y(n2773) );
  OAI21X1 U336 ( .A(n277), .B(n397), .C(n6303), .Y(n2774) );
  OAI21X1 U338 ( .A(n279), .B(n397), .C(n6300), .Y(n2775) );
  OAI21X1 U340 ( .A(n281), .B(n397), .C(n6297), .Y(n2776) );
  OAI21X1 U342 ( .A(n283), .B(n397), .C(n6294), .Y(n2777) );
  OAI21X1 U344 ( .A(n285), .B(n397), .C(n6291), .Y(n2778) );
  OAI21X1 U346 ( .A(n287), .B(n397), .C(n6288), .Y(n2779) );
  OAI21X1 U348 ( .A(n289), .B(n397), .C(n6285), .Y(n2780) );
  OAI21X1 U350 ( .A(n291), .B(n397), .C(n6282), .Y(n2781) );
  OAI21X1 U352 ( .A(n293), .B(n397), .C(n6279), .Y(n2782) );
  OAI21X1 U354 ( .A(n295), .B(n397), .C(n6276), .Y(n2783) );
  OAI21X1 U356 ( .A(n297), .B(n397), .C(n6273), .Y(n2784) );
  OAI21X1 U358 ( .A(n299), .B(n397), .C(n6270), .Y(n2785) );
  OAI21X1 U360 ( .A(n301), .B(n397), .C(n6267), .Y(n2786) );
  OAI21X1 U362 ( .A(n303), .B(n397), .C(n6264), .Y(n2787) );
  OAI21X1 U364 ( .A(n305), .B(n397), .C(n6261), .Y(n2788) );
  OAI21X1 U366 ( .A(n307), .B(n397), .C(n6258), .Y(n2789) );
  OAI21X1 U368 ( .A(n309), .B(n397), .C(n6255), .Y(n2790) );
  OAI21X1 U370 ( .A(n311), .B(n397), .C(n6252), .Y(n2791) );
  OAI21X1 U372 ( .A(n313), .B(n397), .C(n6249), .Y(n2792) );
  OAI21X1 U374 ( .A(n315), .B(n397), .C(n6246), .Y(n2793) );
  OAI21X1 U376 ( .A(n317), .B(n397), .C(n6243), .Y(n2794) );
  OAI21X1 U378 ( .A(n319), .B(n397), .C(n6240), .Y(n2795) );
  OAI21X1 U380 ( .A(n321), .B(n397), .C(n6237), .Y(n2796) );
  OAI21X1 U383 ( .A(n255), .B(n433), .C(n6234), .Y(n2797) );
  OAI21X1 U385 ( .A(n257), .B(n433), .C(n6231), .Y(n2798) );
  OAI21X1 U387 ( .A(n259), .B(n433), .C(n6228), .Y(n2799) );
  OAI21X1 U389 ( .A(n261), .B(n433), .C(n6225), .Y(n2800) );
  OAI21X1 U391 ( .A(n263), .B(n433), .C(n6222), .Y(n2801) );
  OAI21X1 U393 ( .A(n265), .B(n433), .C(n6219), .Y(n2802) );
  OAI21X1 U395 ( .A(n267), .B(n433), .C(n6216), .Y(n2803) );
  OAI21X1 U397 ( .A(n269), .B(n433), .C(n6213), .Y(n2804) );
  OAI21X1 U399 ( .A(n271), .B(n433), .C(n6210), .Y(n2805) );
  OAI21X1 U401 ( .A(n273), .B(n433), .C(n6207), .Y(n2806) );
  OAI21X1 U403 ( .A(n275), .B(n433), .C(n6204), .Y(n2807) );
  OAI21X1 U405 ( .A(n277), .B(n433), .C(n6201), .Y(n2808) );
  OAI21X1 U407 ( .A(n279), .B(n433), .C(n6198), .Y(n2809) );
  OAI21X1 U409 ( .A(n281), .B(n433), .C(n6195), .Y(n2810) );
  OAI21X1 U411 ( .A(n283), .B(n433), .C(n6192), .Y(n2811) );
  OAI21X1 U413 ( .A(n285), .B(n433), .C(n6189), .Y(n2812) );
  OAI21X1 U415 ( .A(n287), .B(n433), .C(n6186), .Y(n2813) );
  OAI21X1 U417 ( .A(n289), .B(n433), .C(n6183), .Y(n2814) );
  OAI21X1 U419 ( .A(n291), .B(n433), .C(n6180), .Y(n2815) );
  OAI21X1 U421 ( .A(n293), .B(n433), .C(n6177), .Y(n2816) );
  OAI21X1 U423 ( .A(n295), .B(n433), .C(n6174), .Y(n2817) );
  OAI21X1 U425 ( .A(n297), .B(n433), .C(n6171), .Y(n2818) );
  OAI21X1 U427 ( .A(n299), .B(n433), .C(n6168), .Y(n2819) );
  OAI21X1 U429 ( .A(n301), .B(n433), .C(n6165), .Y(n2820) );
  OAI21X1 U431 ( .A(n303), .B(n433), .C(n6162), .Y(n2821) );
  OAI21X1 U433 ( .A(n305), .B(n433), .C(n6159), .Y(n2822) );
  OAI21X1 U435 ( .A(n307), .B(n433), .C(n6156), .Y(n2823) );
  OAI21X1 U437 ( .A(n309), .B(n433), .C(n6153), .Y(n2824) );
  OAI21X1 U439 ( .A(n311), .B(n433), .C(n6150), .Y(n2825) );
  OAI21X1 U441 ( .A(n313), .B(n433), .C(n6147), .Y(n2826) );
  OAI21X1 U443 ( .A(n315), .B(n433), .C(n6144), .Y(n2827) );
  OAI21X1 U445 ( .A(n317), .B(n433), .C(n6141), .Y(n2828) );
  OAI21X1 U447 ( .A(n319), .B(n433), .C(n6138), .Y(n2829) );
  OAI21X1 U449 ( .A(n321), .B(n433), .C(n6135), .Y(n2830) );
  OAI21X1 U452 ( .A(n255), .B(n469), .C(n6132), .Y(n2831) );
  OAI21X1 U454 ( .A(n257), .B(n469), .C(n6129), .Y(n2832) );
  OAI21X1 U456 ( .A(n259), .B(n469), .C(n6126), .Y(n2833) );
  OAI21X1 U458 ( .A(n261), .B(n469), .C(n6123), .Y(n2834) );
  OAI21X1 U460 ( .A(n263), .B(n469), .C(n6120), .Y(n2835) );
  OAI21X1 U462 ( .A(n265), .B(n469), .C(n6117), .Y(n2836) );
  OAI21X1 U464 ( .A(n267), .B(n469), .C(n6114), .Y(n2837) );
  OAI21X1 U466 ( .A(n269), .B(n469), .C(n6111), .Y(n2838) );
  OAI21X1 U468 ( .A(n271), .B(n469), .C(n6108), .Y(n2839) );
  OAI21X1 U470 ( .A(n273), .B(n469), .C(n6105), .Y(n2840) );
  OAI21X1 U472 ( .A(n275), .B(n469), .C(n6102), .Y(n2841) );
  OAI21X1 U474 ( .A(n277), .B(n469), .C(n6099), .Y(n2842) );
  OAI21X1 U476 ( .A(n279), .B(n469), .C(n6096), .Y(n2843) );
  OAI21X1 U478 ( .A(n281), .B(n469), .C(n6093), .Y(n2844) );
  OAI21X1 U480 ( .A(n283), .B(n469), .C(n6090), .Y(n2845) );
  OAI21X1 U482 ( .A(n285), .B(n469), .C(n6087), .Y(n2846) );
  OAI21X1 U484 ( .A(n287), .B(n469), .C(n6084), .Y(n2847) );
  OAI21X1 U486 ( .A(n289), .B(n469), .C(n6081), .Y(n2848) );
  OAI21X1 U488 ( .A(n291), .B(n469), .C(n6078), .Y(n2849) );
  OAI21X1 U490 ( .A(n293), .B(n469), .C(n6075), .Y(n2850) );
  OAI21X1 U492 ( .A(n295), .B(n469), .C(n6072), .Y(n2851) );
  OAI21X1 U494 ( .A(n297), .B(n469), .C(n6069), .Y(n2852) );
  OAI21X1 U496 ( .A(n299), .B(n469), .C(n6066), .Y(n2853) );
  OAI21X1 U498 ( .A(n301), .B(n469), .C(n6063), .Y(n2854) );
  OAI21X1 U500 ( .A(n303), .B(n469), .C(n6060), .Y(n2855) );
  OAI21X1 U502 ( .A(n305), .B(n469), .C(n6057), .Y(n2856) );
  OAI21X1 U504 ( .A(n307), .B(n469), .C(n6054), .Y(n2857) );
  OAI21X1 U506 ( .A(n309), .B(n469), .C(n6051), .Y(n2858) );
  OAI21X1 U508 ( .A(n311), .B(n469), .C(n6048), .Y(n2859) );
  OAI21X1 U510 ( .A(n313), .B(n469), .C(n6045), .Y(n2860) );
  OAI21X1 U512 ( .A(n315), .B(n469), .C(n6042), .Y(n2861) );
  OAI21X1 U514 ( .A(n317), .B(n469), .C(n6039), .Y(n2862) );
  OAI21X1 U516 ( .A(n319), .B(n469), .C(n6036), .Y(n2863) );
  OAI21X1 U518 ( .A(n321), .B(n469), .C(n6033), .Y(n2864) );
  OAI21X1 U521 ( .A(n255), .B(n505), .C(n6030), .Y(n2865) );
  OAI21X1 U523 ( .A(n257), .B(n505), .C(n6027), .Y(n2866) );
  OAI21X1 U525 ( .A(n259), .B(n505), .C(n6024), .Y(n2867) );
  OAI21X1 U527 ( .A(n261), .B(n505), .C(n6021), .Y(n2868) );
  OAI21X1 U529 ( .A(n263), .B(n505), .C(n6018), .Y(n2869) );
  OAI21X1 U531 ( .A(n265), .B(n505), .C(n6015), .Y(n2870) );
  OAI21X1 U533 ( .A(n267), .B(n505), .C(n6012), .Y(n2871) );
  OAI21X1 U535 ( .A(n269), .B(n505), .C(n6009), .Y(n2872) );
  OAI21X1 U537 ( .A(n271), .B(n505), .C(n6006), .Y(n2873) );
  OAI21X1 U539 ( .A(n273), .B(n505), .C(n6003), .Y(n2874) );
  OAI21X1 U541 ( .A(n275), .B(n505), .C(n6000), .Y(n2875) );
  OAI21X1 U543 ( .A(n277), .B(n505), .C(n5997), .Y(n2876) );
  OAI21X1 U545 ( .A(n279), .B(n505), .C(n5994), .Y(n2877) );
  OAI21X1 U547 ( .A(n281), .B(n505), .C(n5991), .Y(n2878) );
  OAI21X1 U549 ( .A(n283), .B(n505), .C(n5988), .Y(n2879) );
  OAI21X1 U551 ( .A(n285), .B(n505), .C(n5985), .Y(n2880) );
  OAI21X1 U553 ( .A(n287), .B(n505), .C(n5982), .Y(n2881) );
  OAI21X1 U555 ( .A(n289), .B(n505), .C(n5979), .Y(n2882) );
  OAI21X1 U557 ( .A(n291), .B(n505), .C(n5976), .Y(n2883) );
  OAI21X1 U559 ( .A(n293), .B(n505), .C(n5973), .Y(n2884) );
  OAI21X1 U561 ( .A(n295), .B(n505), .C(n5970), .Y(n2885) );
  OAI21X1 U563 ( .A(n297), .B(n505), .C(n5967), .Y(n2886) );
  OAI21X1 U565 ( .A(n299), .B(n505), .C(n5964), .Y(n2887) );
  OAI21X1 U567 ( .A(n301), .B(n505), .C(n5961), .Y(n2888) );
  OAI21X1 U569 ( .A(n303), .B(n505), .C(n5958), .Y(n2889) );
  OAI21X1 U571 ( .A(n305), .B(n505), .C(n5955), .Y(n2890) );
  OAI21X1 U573 ( .A(n307), .B(n505), .C(n5952), .Y(n2891) );
  OAI21X1 U575 ( .A(n309), .B(n505), .C(n5949), .Y(n2892) );
  OAI21X1 U577 ( .A(n311), .B(n505), .C(n5946), .Y(n2893) );
  OAI21X1 U579 ( .A(n313), .B(n505), .C(n5943), .Y(n2894) );
  OAI21X1 U581 ( .A(n315), .B(n505), .C(n5940), .Y(n2895) );
  OAI21X1 U583 ( .A(n317), .B(n505), .C(n5937), .Y(n2896) );
  OAI21X1 U585 ( .A(n319), .B(n505), .C(n5934), .Y(n2897) );
  OAI21X1 U587 ( .A(n321), .B(n505), .C(n5931), .Y(n2898) );
  OAI21X1 U590 ( .A(n255), .B(n541), .C(n5928), .Y(n2899) );
  OAI21X1 U592 ( .A(n257), .B(n541), .C(n5925), .Y(n2900) );
  OAI21X1 U594 ( .A(n259), .B(n541), .C(n5922), .Y(n2901) );
  OAI21X1 U596 ( .A(n261), .B(n541), .C(n5919), .Y(n2902) );
  OAI21X1 U598 ( .A(n263), .B(n541), .C(n5916), .Y(n2903) );
  OAI21X1 U600 ( .A(n265), .B(n541), .C(n5913), .Y(n2904) );
  OAI21X1 U602 ( .A(n267), .B(n541), .C(n5910), .Y(n2905) );
  OAI21X1 U604 ( .A(n269), .B(n541), .C(n5907), .Y(n2906) );
  OAI21X1 U606 ( .A(n271), .B(n541), .C(n5904), .Y(n2907) );
  OAI21X1 U608 ( .A(n273), .B(n541), .C(n5901), .Y(n2908) );
  OAI21X1 U610 ( .A(n275), .B(n541), .C(n5898), .Y(n2909) );
  OAI21X1 U612 ( .A(n277), .B(n541), .C(n5895), .Y(n2910) );
  OAI21X1 U614 ( .A(n279), .B(n541), .C(n5892), .Y(n2911) );
  OAI21X1 U616 ( .A(n281), .B(n541), .C(n5889), .Y(n2912) );
  OAI21X1 U618 ( .A(n283), .B(n541), .C(n5886), .Y(n2913) );
  OAI21X1 U620 ( .A(n285), .B(n541), .C(n5883), .Y(n2914) );
  OAI21X1 U622 ( .A(n287), .B(n541), .C(n5880), .Y(n2915) );
  OAI21X1 U624 ( .A(n289), .B(n541), .C(n5877), .Y(n2916) );
  OAI21X1 U626 ( .A(n291), .B(n541), .C(n5874), .Y(n2917) );
  OAI21X1 U628 ( .A(n293), .B(n541), .C(n5871), .Y(n2918) );
  OAI21X1 U630 ( .A(n295), .B(n541), .C(n5868), .Y(n2919) );
  OAI21X1 U632 ( .A(n297), .B(n541), .C(n5865), .Y(n2920) );
  OAI21X1 U634 ( .A(n299), .B(n541), .C(n5862), .Y(n2921) );
  OAI21X1 U636 ( .A(n301), .B(n541), .C(n5859), .Y(n2922) );
  OAI21X1 U638 ( .A(n303), .B(n541), .C(n5856), .Y(n2923) );
  OAI21X1 U640 ( .A(n305), .B(n541), .C(n5853), .Y(n2924) );
  OAI21X1 U642 ( .A(n307), .B(n541), .C(n5850), .Y(n2925) );
  OAI21X1 U644 ( .A(n309), .B(n541), .C(n5847), .Y(n2926) );
  OAI21X1 U646 ( .A(n311), .B(n541), .C(n5844), .Y(n2927) );
  OAI21X1 U648 ( .A(n313), .B(n541), .C(n5841), .Y(n2928) );
  OAI21X1 U650 ( .A(n315), .B(n541), .C(n5838), .Y(n2929) );
  OAI21X1 U652 ( .A(n317), .B(n541), .C(n5835), .Y(n2930) );
  OAI21X1 U654 ( .A(n319), .B(n541), .C(n5832), .Y(n2931) );
  OAI21X1 U656 ( .A(n321), .B(n541), .C(n5829), .Y(n2932) );
  NAND3X1 U660 ( .A(n240), .B(n238), .C(n237), .Y(n577) );
  OAI21X1 U661 ( .A(n255), .B(n10506), .C(n5826), .Y(n2933) );
  OAI21X1 U663 ( .A(n257), .B(n10506), .C(n5823), .Y(n2934) );
  OAI21X1 U665 ( .A(n259), .B(n10506), .C(n5820), .Y(n2935) );
  OAI21X1 U667 ( .A(n261), .B(n10506), .C(n5817), .Y(n2936) );
  OAI21X1 U669 ( .A(n263), .B(n10506), .C(n5814), .Y(n2937) );
  OAI21X1 U671 ( .A(n265), .B(n10506), .C(n5811), .Y(n2938) );
  OAI21X1 U673 ( .A(n267), .B(n10506), .C(n5808), .Y(n2939) );
  OAI21X1 U675 ( .A(n269), .B(n10506), .C(n5805), .Y(n2940) );
  OAI21X1 U677 ( .A(n271), .B(n10506), .C(n5802), .Y(n2941) );
  OAI21X1 U679 ( .A(n273), .B(n10506), .C(n5799), .Y(n2942) );
  OAI21X1 U681 ( .A(n275), .B(n10506), .C(n5796), .Y(n2943) );
  OAI21X1 U683 ( .A(n277), .B(n10506), .C(n5793), .Y(n2944) );
  OAI21X1 U685 ( .A(n279), .B(n10506), .C(n5790), .Y(n2945) );
  OAI21X1 U687 ( .A(n281), .B(n10506), .C(n5787), .Y(n2946) );
  OAI21X1 U689 ( .A(n283), .B(n10506), .C(n5784), .Y(n2947) );
  OAI21X1 U691 ( .A(n285), .B(n10506), .C(n5781), .Y(n2948) );
  OAI21X1 U693 ( .A(n287), .B(n10506), .C(n5778), .Y(n2949) );
  OAI21X1 U695 ( .A(n289), .B(n10506), .C(n5775), .Y(n2950) );
  OAI21X1 U697 ( .A(n291), .B(n10506), .C(n5772), .Y(n2951) );
  OAI21X1 U699 ( .A(n293), .B(n10506), .C(n5769), .Y(n2952) );
  OAI21X1 U701 ( .A(n295), .B(n10506), .C(n5766), .Y(n2953) );
  OAI21X1 U703 ( .A(n297), .B(n10506), .C(n5763), .Y(n2954) );
  OAI21X1 U705 ( .A(n299), .B(n10506), .C(n5760), .Y(n2955) );
  OAI21X1 U707 ( .A(n301), .B(n10506), .C(n5757), .Y(n2956) );
  OAI21X1 U709 ( .A(n303), .B(n10506), .C(n5754), .Y(n2957) );
  OAI21X1 U711 ( .A(n305), .B(n10506), .C(n5751), .Y(n2958) );
  OAI21X1 U713 ( .A(n307), .B(n10506), .C(n5748), .Y(n2959) );
  OAI21X1 U715 ( .A(n309), .B(n10506), .C(n5745), .Y(n2960) );
  OAI21X1 U717 ( .A(n311), .B(n10506), .C(n5742), .Y(n2961) );
  OAI21X1 U719 ( .A(n313), .B(n10506), .C(n5739), .Y(n2962) );
  OAI21X1 U721 ( .A(n315), .B(n10506), .C(n5736), .Y(n2963) );
  OAI21X1 U723 ( .A(n317), .B(n10506), .C(n5733), .Y(n2964) );
  OAI21X1 U725 ( .A(n319), .B(n10506), .C(n5730), .Y(n2965) );
  OAI21X1 U727 ( .A(n321), .B(n10506), .C(n5727), .Y(n2966) );
  OAI21X1 U730 ( .A(n255), .B(n10508), .C(n5724), .Y(n2967) );
  OAI21X1 U732 ( .A(n257), .B(n10508), .C(n5721), .Y(n2968) );
  OAI21X1 U734 ( .A(n259), .B(n10508), .C(n5718), .Y(n2969) );
  OAI21X1 U736 ( .A(n261), .B(n10508), .C(n5715), .Y(n2970) );
  OAI21X1 U738 ( .A(n263), .B(n10508), .C(n5712), .Y(n2971) );
  OAI21X1 U740 ( .A(n265), .B(n10508), .C(n5709), .Y(n2972) );
  OAI21X1 U742 ( .A(n267), .B(n10508), .C(n5706), .Y(n2973) );
  OAI21X1 U744 ( .A(n269), .B(n10508), .C(n5703), .Y(n2974) );
  OAI21X1 U746 ( .A(n271), .B(n10508), .C(n5700), .Y(n2975) );
  OAI21X1 U748 ( .A(n273), .B(n10508), .C(n5697), .Y(n2976) );
  OAI21X1 U750 ( .A(n275), .B(n10508), .C(n5694), .Y(n2977) );
  OAI21X1 U752 ( .A(n277), .B(n10508), .C(n5691), .Y(n2978) );
  OAI21X1 U754 ( .A(n279), .B(n10508), .C(n5688), .Y(n2979) );
  OAI21X1 U756 ( .A(n281), .B(n10508), .C(n5685), .Y(n2980) );
  OAI21X1 U758 ( .A(n283), .B(n10508), .C(n5682), .Y(n2981) );
  OAI21X1 U760 ( .A(n285), .B(n10508), .C(n5679), .Y(n2982) );
  OAI21X1 U762 ( .A(n287), .B(n10508), .C(n5676), .Y(n2983) );
  OAI21X1 U764 ( .A(n289), .B(n10508), .C(n5673), .Y(n2984) );
  OAI21X1 U766 ( .A(n291), .B(n10508), .C(n5670), .Y(n2985) );
  OAI21X1 U768 ( .A(n293), .B(n10508), .C(n5667), .Y(n2986) );
  OAI21X1 U770 ( .A(n295), .B(n10508), .C(n5664), .Y(n2987) );
  OAI21X1 U772 ( .A(n297), .B(n10508), .C(n5661), .Y(n2988) );
  OAI21X1 U774 ( .A(n299), .B(n10508), .C(n5658), .Y(n2989) );
  OAI21X1 U776 ( .A(n301), .B(n10508), .C(n5655), .Y(n2990) );
  OAI21X1 U778 ( .A(n303), .B(n10508), .C(n5652), .Y(n2991) );
  OAI21X1 U780 ( .A(n305), .B(n10508), .C(n5649), .Y(n2992) );
  OAI21X1 U782 ( .A(n307), .B(n10508), .C(n5646), .Y(n2993) );
  OAI21X1 U784 ( .A(n309), .B(n10508), .C(n5643), .Y(n2994) );
  OAI21X1 U786 ( .A(n311), .B(n10508), .C(n5640), .Y(n2995) );
  OAI21X1 U788 ( .A(n313), .B(n10508), .C(n5637), .Y(n2996) );
  OAI21X1 U790 ( .A(n315), .B(n10508), .C(n5634), .Y(n2997) );
  OAI21X1 U792 ( .A(n317), .B(n10508), .C(n5631), .Y(n2998) );
  OAI21X1 U794 ( .A(n319), .B(n10508), .C(n5628), .Y(n2999) );
  OAI21X1 U796 ( .A(n321), .B(n10508), .C(n5625), .Y(n3000) );
  OAI21X1 U799 ( .A(n255), .B(n649), .C(n5622), .Y(n3001) );
  OAI21X1 U801 ( .A(n257), .B(n649), .C(n5619), .Y(n3002) );
  OAI21X1 U803 ( .A(n259), .B(n649), .C(n5616), .Y(n3003) );
  OAI21X1 U805 ( .A(n261), .B(n649), .C(n5613), .Y(n3004) );
  OAI21X1 U807 ( .A(n263), .B(n649), .C(n5610), .Y(n3005) );
  OAI21X1 U809 ( .A(n265), .B(n649), .C(n5607), .Y(n3006) );
  OAI21X1 U811 ( .A(n267), .B(n649), .C(n5604), .Y(n3007) );
  OAI21X1 U813 ( .A(n269), .B(n649), .C(n5601), .Y(n3008) );
  OAI21X1 U815 ( .A(n271), .B(n649), .C(n5598), .Y(n3009) );
  OAI21X1 U817 ( .A(n273), .B(n649), .C(n5595), .Y(n3010) );
  OAI21X1 U819 ( .A(n275), .B(n649), .C(n5592), .Y(n3011) );
  OAI21X1 U821 ( .A(n277), .B(n649), .C(n5589), .Y(n3012) );
  OAI21X1 U823 ( .A(n279), .B(n649), .C(n5586), .Y(n3013) );
  OAI21X1 U825 ( .A(n281), .B(n649), .C(n5583), .Y(n3014) );
  OAI21X1 U827 ( .A(n283), .B(n649), .C(n5580), .Y(n3015) );
  OAI21X1 U829 ( .A(n285), .B(n649), .C(n5577), .Y(n3016) );
  OAI21X1 U831 ( .A(n287), .B(n649), .C(n5574), .Y(n3017) );
  OAI21X1 U833 ( .A(n289), .B(n649), .C(n5571), .Y(n3018) );
  OAI21X1 U835 ( .A(n291), .B(n649), .C(n5568), .Y(n3019) );
  OAI21X1 U837 ( .A(n293), .B(n649), .C(n5565), .Y(n3020) );
  OAI21X1 U839 ( .A(n295), .B(n649), .C(n5562), .Y(n3021) );
  OAI21X1 U841 ( .A(n297), .B(n649), .C(n5559), .Y(n3022) );
  OAI21X1 U843 ( .A(n299), .B(n649), .C(n5556), .Y(n3023) );
  OAI21X1 U845 ( .A(n301), .B(n649), .C(n5553), .Y(n3024) );
  OAI21X1 U847 ( .A(n303), .B(n649), .C(n5550), .Y(n3025) );
  OAI21X1 U849 ( .A(n305), .B(n649), .C(n5547), .Y(n3026) );
  OAI21X1 U851 ( .A(n307), .B(n649), .C(n5544), .Y(n3027) );
  OAI21X1 U853 ( .A(n309), .B(n649), .C(n5541), .Y(n3028) );
  OAI21X1 U855 ( .A(n311), .B(n649), .C(n5538), .Y(n3029) );
  OAI21X1 U857 ( .A(n313), .B(n649), .C(n5535), .Y(n3030) );
  OAI21X1 U859 ( .A(n315), .B(n649), .C(n5532), .Y(n3031) );
  OAI21X1 U861 ( .A(n317), .B(n649), .C(n5529), .Y(n3032) );
  OAI21X1 U863 ( .A(n319), .B(n649), .C(n5526), .Y(n3033) );
  OAI21X1 U865 ( .A(n321), .B(n649), .C(n5523), .Y(n3034) );
  OAI21X1 U868 ( .A(n255), .B(n10515), .C(n5520), .Y(n3035) );
  OAI21X1 U870 ( .A(n257), .B(n10515), .C(n5517), .Y(n3036) );
  OAI21X1 U872 ( .A(n259), .B(n10515), .C(n5514), .Y(n3037) );
  OAI21X1 U874 ( .A(n261), .B(n10515), .C(n5511), .Y(n3038) );
  OAI21X1 U876 ( .A(n263), .B(n10515), .C(n5508), .Y(n3039) );
  OAI21X1 U878 ( .A(n265), .B(n10515), .C(n5505), .Y(n3040) );
  OAI21X1 U880 ( .A(n267), .B(n10515), .C(n5502), .Y(n3041) );
  OAI21X1 U882 ( .A(n269), .B(n10515), .C(n5499), .Y(n3042) );
  OAI21X1 U884 ( .A(n271), .B(n10515), .C(n5496), .Y(n3043) );
  OAI21X1 U886 ( .A(n273), .B(n10515), .C(n5493), .Y(n3044) );
  OAI21X1 U888 ( .A(n275), .B(n10515), .C(n5490), .Y(n3045) );
  OAI21X1 U890 ( .A(n277), .B(n10515), .C(n5487), .Y(n3046) );
  OAI21X1 U892 ( .A(n279), .B(n10515), .C(n5484), .Y(n3047) );
  OAI21X1 U894 ( .A(n281), .B(n10515), .C(n5481), .Y(n3048) );
  OAI21X1 U896 ( .A(n283), .B(n10515), .C(n5478), .Y(n3049) );
  OAI21X1 U898 ( .A(n285), .B(n10515), .C(n5475), .Y(n3050) );
  OAI21X1 U900 ( .A(n287), .B(n10515), .C(n5472), .Y(n3051) );
  OAI21X1 U902 ( .A(n289), .B(n10515), .C(n5469), .Y(n3052) );
  OAI21X1 U904 ( .A(n291), .B(n10515), .C(n5466), .Y(n3053) );
  OAI21X1 U906 ( .A(n293), .B(n10515), .C(n5463), .Y(n3054) );
  OAI21X1 U908 ( .A(n295), .B(n10515), .C(n5460), .Y(n3055) );
  OAI21X1 U910 ( .A(n297), .B(n10515), .C(n5457), .Y(n3056) );
  OAI21X1 U912 ( .A(n299), .B(n10515), .C(n5454), .Y(n3057) );
  OAI21X1 U914 ( .A(n301), .B(n10515), .C(n5451), .Y(n3058) );
  OAI21X1 U916 ( .A(n303), .B(n10515), .C(n5448), .Y(n3059) );
  OAI21X1 U918 ( .A(n305), .B(n10515), .C(n5445), .Y(n3060) );
  OAI21X1 U920 ( .A(n307), .B(n10515), .C(n5442), .Y(n3061) );
  OAI21X1 U922 ( .A(n309), .B(n10515), .C(n5439), .Y(n3062) );
  OAI21X1 U924 ( .A(n311), .B(n10515), .C(n5436), .Y(n3063) );
  OAI21X1 U926 ( .A(n313), .B(n10515), .C(n5433), .Y(n3064) );
  OAI21X1 U928 ( .A(n315), .B(n10515), .C(n5430), .Y(n3065) );
  OAI21X1 U930 ( .A(n317), .B(n10515), .C(n5427), .Y(n3066) );
  OAI21X1 U932 ( .A(n319), .B(n10515), .C(n5424), .Y(n3067) );
  OAI21X1 U934 ( .A(n321), .B(n10515), .C(n5421), .Y(n3068) );
  OAI21X1 U937 ( .A(n255), .B(n719), .C(n5418), .Y(n3069) );
  OAI21X1 U939 ( .A(n257), .B(n719), .C(n5415), .Y(n3070) );
  OAI21X1 U941 ( .A(n259), .B(n719), .C(n5412), .Y(n3071) );
  OAI21X1 U943 ( .A(n261), .B(n719), .C(n5409), .Y(n3072) );
  OAI21X1 U945 ( .A(n263), .B(n719), .C(n5406), .Y(n3073) );
  OAI21X1 U947 ( .A(n265), .B(n719), .C(n5403), .Y(n3074) );
  OAI21X1 U949 ( .A(n267), .B(n719), .C(n5400), .Y(n3075) );
  OAI21X1 U951 ( .A(n269), .B(n719), .C(n5397), .Y(n3076) );
  OAI21X1 U953 ( .A(n271), .B(n719), .C(n5394), .Y(n3077) );
  OAI21X1 U955 ( .A(n273), .B(n719), .C(n5391), .Y(n3078) );
  OAI21X1 U957 ( .A(n275), .B(n719), .C(n5388), .Y(n3079) );
  OAI21X1 U959 ( .A(n277), .B(n719), .C(n5385), .Y(n3080) );
  OAI21X1 U961 ( .A(n279), .B(n719), .C(n5382), .Y(n3081) );
  OAI21X1 U963 ( .A(n281), .B(n719), .C(n5379), .Y(n3082) );
  OAI21X1 U965 ( .A(n283), .B(n719), .C(n5376), .Y(n3083) );
  OAI21X1 U967 ( .A(n285), .B(n719), .C(n5373), .Y(n3084) );
  OAI21X1 U969 ( .A(n287), .B(n719), .C(n5370), .Y(n3085) );
  OAI21X1 U971 ( .A(n289), .B(n719), .C(n5367), .Y(n3086) );
  OAI21X1 U973 ( .A(n291), .B(n719), .C(n5364), .Y(n3087) );
  OAI21X1 U975 ( .A(n293), .B(n719), .C(n5361), .Y(n3088) );
  OAI21X1 U977 ( .A(n295), .B(n719), .C(n5358), .Y(n3089) );
  OAI21X1 U979 ( .A(n297), .B(n719), .C(n5355), .Y(n3090) );
  OAI21X1 U981 ( .A(n299), .B(n719), .C(n5352), .Y(n3091) );
  OAI21X1 U983 ( .A(n301), .B(n719), .C(n5349), .Y(n3092) );
  OAI21X1 U985 ( .A(n303), .B(n719), .C(n5346), .Y(n3093) );
  OAI21X1 U987 ( .A(n305), .B(n719), .C(n5343), .Y(n3094) );
  OAI21X1 U989 ( .A(n307), .B(n719), .C(n5340), .Y(n3095) );
  OAI21X1 U991 ( .A(n309), .B(n719), .C(n5337), .Y(n3096) );
  OAI21X1 U993 ( .A(n311), .B(n719), .C(n5334), .Y(n3097) );
  OAI21X1 U995 ( .A(n313), .B(n719), .C(n5331), .Y(n3098) );
  OAI21X1 U997 ( .A(n315), .B(n719), .C(n5328), .Y(n3099) );
  OAI21X1 U999 ( .A(n317), .B(n719), .C(n5325), .Y(n3100) );
  OAI21X1 U1001 ( .A(n319), .B(n719), .C(n5322), .Y(n3101) );
  OAI21X1 U1003 ( .A(n321), .B(n719), .C(n5319), .Y(n3102) );
  OAI21X1 U1006 ( .A(n255), .B(n10517), .C(n5316), .Y(n3103) );
  OAI21X1 U1008 ( .A(n257), .B(n10517), .C(n5313), .Y(n3104) );
  OAI21X1 U1010 ( .A(n259), .B(n10517), .C(n5310), .Y(n3105) );
  OAI21X1 U1012 ( .A(n261), .B(n10517), .C(n5307), .Y(n3106) );
  OAI21X1 U1014 ( .A(n263), .B(n10517), .C(n5304), .Y(n3107) );
  OAI21X1 U1016 ( .A(n265), .B(n10517), .C(n5301), .Y(n3108) );
  OAI21X1 U1018 ( .A(n267), .B(n10517), .C(n5298), .Y(n3109) );
  OAI21X1 U1020 ( .A(n269), .B(n10517), .C(n5295), .Y(n3110) );
  OAI21X1 U1022 ( .A(n271), .B(n10517), .C(n5292), .Y(n3111) );
  OAI21X1 U1024 ( .A(n273), .B(n10517), .C(n5289), .Y(n3112) );
  OAI21X1 U1026 ( .A(n275), .B(n10517), .C(n5286), .Y(n3113) );
  OAI21X1 U1028 ( .A(n277), .B(n10517), .C(n5283), .Y(n3114) );
  OAI21X1 U1030 ( .A(n279), .B(n10517), .C(n5280), .Y(n3115) );
  OAI21X1 U1032 ( .A(n281), .B(n10517), .C(n5277), .Y(n3116) );
  OAI21X1 U1034 ( .A(n283), .B(n10517), .C(n5274), .Y(n3117) );
  OAI21X1 U1036 ( .A(n285), .B(n10517), .C(n5271), .Y(n3118) );
  OAI21X1 U1038 ( .A(n287), .B(n10517), .C(n5268), .Y(n3119) );
  OAI21X1 U1040 ( .A(n289), .B(n10517), .C(n5265), .Y(n3120) );
  OAI21X1 U1042 ( .A(n291), .B(n10517), .C(n5262), .Y(n3121) );
  OAI21X1 U1044 ( .A(n293), .B(n10517), .C(n5259), .Y(n3122) );
  OAI21X1 U1046 ( .A(n295), .B(n10517), .C(n5256), .Y(n3123) );
  OAI21X1 U1048 ( .A(n297), .B(n10517), .C(n5253), .Y(n3124) );
  OAI21X1 U1050 ( .A(n299), .B(n10517), .C(n5250), .Y(n3125) );
  OAI21X1 U1052 ( .A(n301), .B(n10517), .C(n5247), .Y(n3126) );
  OAI21X1 U1054 ( .A(n303), .B(n10517), .C(n5244), .Y(n3127) );
  OAI21X1 U1056 ( .A(n305), .B(n10517), .C(n5241), .Y(n3128) );
  OAI21X1 U1058 ( .A(n307), .B(n10517), .C(n5238), .Y(n3129) );
  OAI21X1 U1060 ( .A(n309), .B(n10517), .C(n5235), .Y(n3130) );
  OAI21X1 U1062 ( .A(n311), .B(n10517), .C(n5232), .Y(n3131) );
  OAI21X1 U1064 ( .A(n313), .B(n10517), .C(n5229), .Y(n3132) );
  OAI21X1 U1066 ( .A(n315), .B(n10517), .C(n5226), .Y(n3133) );
  OAI21X1 U1068 ( .A(n317), .B(n10517), .C(n5223), .Y(n3134) );
  OAI21X1 U1070 ( .A(n319), .B(n10517), .C(n5220), .Y(n3135) );
  OAI21X1 U1072 ( .A(n321), .B(n10517), .C(n5217), .Y(n3136) );
  OAI21X1 U1075 ( .A(n255), .B(n10511), .C(n5214), .Y(n3137) );
  OAI21X1 U1077 ( .A(n257), .B(n10511), .C(n5211), .Y(n3138) );
  OAI21X1 U1079 ( .A(n259), .B(n10511), .C(n5208), .Y(n3139) );
  OAI21X1 U1081 ( .A(n261), .B(n10511), .C(n5205), .Y(n3140) );
  OAI21X1 U1083 ( .A(n263), .B(n10511), .C(n5202), .Y(n3141) );
  OAI21X1 U1085 ( .A(n265), .B(n10511), .C(n5199), .Y(n3142) );
  OAI21X1 U1087 ( .A(n267), .B(n10511), .C(n5196), .Y(n3143) );
  OAI21X1 U1089 ( .A(n269), .B(n10511), .C(n5193), .Y(n3144) );
  OAI21X1 U1091 ( .A(n271), .B(n10511), .C(n5190), .Y(n3145) );
  OAI21X1 U1093 ( .A(n273), .B(n10511), .C(n5187), .Y(n3146) );
  OAI21X1 U1095 ( .A(n275), .B(n10511), .C(n5184), .Y(n3147) );
  OAI21X1 U1097 ( .A(n277), .B(n10511), .C(n5181), .Y(n3148) );
  OAI21X1 U1099 ( .A(n279), .B(n10511), .C(n5178), .Y(n3149) );
  OAI21X1 U1101 ( .A(n281), .B(n10511), .C(n5175), .Y(n3150) );
  OAI21X1 U1103 ( .A(n283), .B(n10511), .C(n5172), .Y(n3151) );
  OAI21X1 U1105 ( .A(n285), .B(n10511), .C(n5169), .Y(n3152) );
  OAI21X1 U1107 ( .A(n287), .B(n10511), .C(n5166), .Y(n3153) );
  OAI21X1 U1109 ( .A(n289), .B(n10511), .C(n5163), .Y(n3154) );
  OAI21X1 U1111 ( .A(n291), .B(n10511), .C(n5160), .Y(n3155) );
  OAI21X1 U1113 ( .A(n293), .B(n10511), .C(n5157), .Y(n3156) );
  OAI21X1 U1115 ( .A(n295), .B(n10511), .C(n5154), .Y(n3157) );
  OAI21X1 U1117 ( .A(n297), .B(n10511), .C(n5151), .Y(n3158) );
  OAI21X1 U1119 ( .A(n299), .B(n10511), .C(n5148), .Y(n3159) );
  OAI21X1 U1121 ( .A(n301), .B(n10511), .C(n5145), .Y(n3160) );
  OAI21X1 U1123 ( .A(n303), .B(n10511), .C(n5142), .Y(n3161) );
  OAI21X1 U1125 ( .A(n305), .B(n10511), .C(n5139), .Y(n3162) );
  OAI21X1 U1127 ( .A(n307), .B(n10511), .C(n5136), .Y(n3163) );
  OAI21X1 U1129 ( .A(n309), .B(n10511), .C(n5133), .Y(n3164) );
  OAI21X1 U1131 ( .A(n311), .B(n10511), .C(n5130), .Y(n3165) );
  OAI21X1 U1133 ( .A(n313), .B(n10511), .C(n5127), .Y(n3166) );
  OAI21X1 U1135 ( .A(n315), .B(n10511), .C(n5124), .Y(n3167) );
  OAI21X1 U1137 ( .A(n317), .B(n10511), .C(n5121), .Y(n3168) );
  OAI21X1 U1139 ( .A(n319), .B(n10511), .C(n5118), .Y(n3169) );
  OAI21X1 U1141 ( .A(n321), .B(n10511), .C(n5115), .Y(n3170) );
  OAI21X1 U1144 ( .A(n255), .B(n824), .C(n5112), .Y(n3171) );
  OAI21X1 U1146 ( .A(n257), .B(n824), .C(n5109), .Y(n3172) );
  OAI21X1 U1148 ( .A(n259), .B(n824), .C(n5106), .Y(n3173) );
  OAI21X1 U1150 ( .A(n261), .B(n824), .C(n5103), .Y(n3174) );
  OAI21X1 U1152 ( .A(n263), .B(n824), .C(n5100), .Y(n3175) );
  OAI21X1 U1154 ( .A(n265), .B(n824), .C(n5097), .Y(n3176) );
  OAI21X1 U1156 ( .A(n267), .B(n824), .C(n5094), .Y(n3177) );
  OAI21X1 U1158 ( .A(n269), .B(n824), .C(n5091), .Y(n3178) );
  OAI21X1 U1160 ( .A(n271), .B(n824), .C(n5088), .Y(n3179) );
  OAI21X1 U1162 ( .A(n273), .B(n824), .C(n5085), .Y(n3180) );
  OAI21X1 U1164 ( .A(n275), .B(n824), .C(n5082), .Y(n3181) );
  OAI21X1 U1166 ( .A(n277), .B(n824), .C(n5079), .Y(n3182) );
  OAI21X1 U1168 ( .A(n279), .B(n824), .C(n5076), .Y(n3183) );
  OAI21X1 U1170 ( .A(n281), .B(n824), .C(n5073), .Y(n3184) );
  OAI21X1 U1172 ( .A(n283), .B(n824), .C(n5070), .Y(n3185) );
  OAI21X1 U1174 ( .A(n285), .B(n824), .C(n5067), .Y(n3186) );
  OAI21X1 U1176 ( .A(n287), .B(n824), .C(n5064), .Y(n3187) );
  OAI21X1 U1178 ( .A(n289), .B(n824), .C(n5061), .Y(n3188) );
  OAI21X1 U1180 ( .A(n291), .B(n824), .C(n5058), .Y(n3189) );
  OAI21X1 U1182 ( .A(n293), .B(n824), .C(n5055), .Y(n3190) );
  OAI21X1 U1184 ( .A(n295), .B(n824), .C(n5052), .Y(n3191) );
  OAI21X1 U1186 ( .A(n297), .B(n824), .C(n5049), .Y(n3192) );
  OAI21X1 U1188 ( .A(n299), .B(n824), .C(n5046), .Y(n3193) );
  OAI21X1 U1190 ( .A(n301), .B(n824), .C(n5043), .Y(n3194) );
  OAI21X1 U1192 ( .A(n303), .B(n824), .C(n5040), .Y(n3195) );
  OAI21X1 U1194 ( .A(n305), .B(n824), .C(n5037), .Y(n3196) );
  OAI21X1 U1196 ( .A(n307), .B(n824), .C(n5034), .Y(n3197) );
  OAI21X1 U1198 ( .A(n309), .B(n824), .C(n5031), .Y(n3198) );
  OAI21X1 U1200 ( .A(n311), .B(n824), .C(n5028), .Y(n3199) );
  OAI21X1 U1202 ( .A(n313), .B(n824), .C(n5025), .Y(n3200) );
  OAI21X1 U1204 ( .A(n315), .B(n824), .C(n5022), .Y(n3201) );
  OAI21X1 U1206 ( .A(n317), .B(n824), .C(n5019), .Y(n3202) );
  OAI21X1 U1208 ( .A(n319), .B(n824), .C(n5016), .Y(n3203) );
  OAI21X1 U1210 ( .A(n321), .B(n824), .C(n5013), .Y(n3204) );
  NAND3X1 U1214 ( .A(n237), .B(n238), .C(n10097), .Y(n859) );
  INVX1 U1215 ( .A(n10104), .Y(n238) );
  OAI21X1 U1216 ( .A(n255), .B(n10137), .C(n5010), .Y(n3205) );
  OAI21X1 U1218 ( .A(n257), .B(n10137), .C(n5007), .Y(n3206) );
  OAI21X1 U1220 ( .A(n259), .B(n10137), .C(n5004), .Y(n3207) );
  OAI21X1 U1222 ( .A(n261), .B(n10137), .C(n5001), .Y(n3208) );
  OAI21X1 U1224 ( .A(n263), .B(n10137), .C(n4998), .Y(n3209) );
  OAI21X1 U1226 ( .A(n265), .B(n10137), .C(n4995), .Y(n3210) );
  OAI21X1 U1228 ( .A(n267), .B(n10137), .C(n4992), .Y(n3211) );
  OAI21X1 U1230 ( .A(n269), .B(n10137), .C(n4989), .Y(n3212) );
  OAI21X1 U1232 ( .A(n271), .B(n10137), .C(n4986), .Y(n3213) );
  OAI21X1 U1234 ( .A(n273), .B(n10137), .C(n4983), .Y(n3214) );
  OAI21X1 U1236 ( .A(n275), .B(n10137), .C(n4980), .Y(n3215) );
  OAI21X1 U1238 ( .A(n277), .B(n10137), .C(n4977), .Y(n3216) );
  OAI21X1 U1240 ( .A(n279), .B(n10137), .C(n4974), .Y(n3217) );
  OAI21X1 U1242 ( .A(n281), .B(n10137), .C(n4971), .Y(n3218) );
  OAI21X1 U1244 ( .A(n283), .B(n10137), .C(n4968), .Y(n3219) );
  OAI21X1 U1246 ( .A(n285), .B(n10137), .C(n4965), .Y(n3220) );
  OAI21X1 U1248 ( .A(n287), .B(n10137), .C(n4962), .Y(n3221) );
  OAI21X1 U1250 ( .A(n289), .B(n10137), .C(n4959), .Y(n3222) );
  OAI21X1 U1252 ( .A(n291), .B(n10137), .C(n4956), .Y(n3223) );
  OAI21X1 U1254 ( .A(n293), .B(n10137), .C(n4953), .Y(n3224) );
  OAI21X1 U1256 ( .A(n295), .B(n10137), .C(n4950), .Y(n3225) );
  OAI21X1 U1258 ( .A(n297), .B(n10137), .C(n4947), .Y(n3226) );
  OAI21X1 U1260 ( .A(n299), .B(n10137), .C(n4944), .Y(n3227) );
  OAI21X1 U1262 ( .A(n301), .B(n10137), .C(n4941), .Y(n3228) );
  OAI21X1 U1264 ( .A(n303), .B(n10137), .C(n4938), .Y(n3229) );
  OAI21X1 U1266 ( .A(n305), .B(n10137), .C(n4935), .Y(n3230) );
  OAI21X1 U1268 ( .A(n307), .B(n10137), .C(n4932), .Y(n3231) );
  OAI21X1 U1270 ( .A(n309), .B(n10137), .C(n4929), .Y(n3232) );
  OAI21X1 U1272 ( .A(n311), .B(n10137), .C(n4926), .Y(n3233) );
  OAI21X1 U1274 ( .A(n313), .B(n10137), .C(n4923), .Y(n3234) );
  OAI21X1 U1276 ( .A(n315), .B(n10137), .C(n4920), .Y(n3235) );
  OAI21X1 U1278 ( .A(n317), .B(n10137), .C(n4917), .Y(n3236) );
  OAI21X1 U1280 ( .A(n319), .B(n10137), .C(n4914), .Y(n3237) );
  OAI21X1 U1282 ( .A(n321), .B(n10137), .C(n4911), .Y(n3238) );
  OAI21X1 U1285 ( .A(n255), .B(n10134), .C(n4908), .Y(n3239) );
  OAI21X1 U1287 ( .A(n257), .B(n10134), .C(n4905), .Y(n3240) );
  OAI21X1 U1289 ( .A(n259), .B(n10134), .C(n4902), .Y(n3241) );
  OAI21X1 U1291 ( .A(n261), .B(n10134), .C(n4899), .Y(n3242) );
  OAI21X1 U1293 ( .A(n263), .B(n10134), .C(n4896), .Y(n3243) );
  OAI21X1 U1295 ( .A(n265), .B(n10134), .C(n4893), .Y(n3244) );
  OAI21X1 U1297 ( .A(n267), .B(n10134), .C(n4890), .Y(n3245) );
  OAI21X1 U1299 ( .A(n269), .B(n10134), .C(n4887), .Y(n3246) );
  OAI21X1 U1301 ( .A(n271), .B(n10134), .C(n4884), .Y(n3247) );
  OAI21X1 U1303 ( .A(n273), .B(n10134), .C(n4881), .Y(n3248) );
  OAI21X1 U1305 ( .A(n275), .B(n10134), .C(n4878), .Y(n3249) );
  OAI21X1 U1307 ( .A(n277), .B(n10134), .C(n4875), .Y(n3250) );
  OAI21X1 U1309 ( .A(n279), .B(n10134), .C(n4872), .Y(n3251) );
  OAI21X1 U1311 ( .A(n281), .B(n10134), .C(n4869), .Y(n3252) );
  OAI21X1 U1313 ( .A(n283), .B(n10134), .C(n4866), .Y(n3253) );
  OAI21X1 U1315 ( .A(n285), .B(n10134), .C(n4863), .Y(n3254) );
  OAI21X1 U1317 ( .A(n287), .B(n10134), .C(n4860), .Y(n3255) );
  OAI21X1 U1319 ( .A(n289), .B(n10134), .C(n4857), .Y(n3256) );
  OAI21X1 U1321 ( .A(n291), .B(n10134), .C(n4854), .Y(n3257) );
  OAI21X1 U1323 ( .A(n293), .B(n10134), .C(n4851), .Y(n3258) );
  OAI21X1 U1325 ( .A(n295), .B(n10134), .C(n4848), .Y(n3259) );
  OAI21X1 U1327 ( .A(n297), .B(n10134), .C(n4845), .Y(n3260) );
  OAI21X1 U1329 ( .A(n299), .B(n10134), .C(n4842), .Y(n3261) );
  OAI21X1 U1331 ( .A(n301), .B(n10134), .C(n4839), .Y(n3262) );
  OAI21X1 U1333 ( .A(n303), .B(n10134), .C(n4836), .Y(n3263) );
  OAI21X1 U1335 ( .A(n305), .B(n10134), .C(n4833), .Y(n3264) );
  OAI21X1 U1337 ( .A(n307), .B(n10134), .C(n4830), .Y(n3265) );
  OAI21X1 U1339 ( .A(n309), .B(n10134), .C(n4827), .Y(n3266) );
  OAI21X1 U1341 ( .A(n311), .B(n10134), .C(n4824), .Y(n3267) );
  OAI21X1 U1343 ( .A(n313), .B(n10134), .C(n4821), .Y(n3268) );
  OAI21X1 U1345 ( .A(n315), .B(n10134), .C(n4818), .Y(n3269) );
  OAI21X1 U1347 ( .A(n317), .B(n10134), .C(n4815), .Y(n3270) );
  OAI21X1 U1349 ( .A(n319), .B(n10134), .C(n4812), .Y(n3271) );
  OAI21X1 U1351 ( .A(n321), .B(n10134), .C(n4809), .Y(n3272) );
  OAI21X1 U1354 ( .A(n255), .B(n10131), .C(n4806), .Y(n3273) );
  OAI21X1 U1356 ( .A(n257), .B(n10131), .C(n4803), .Y(n3274) );
  OAI21X1 U1358 ( .A(n259), .B(n10131), .C(n4800), .Y(n3275) );
  OAI21X1 U1360 ( .A(n261), .B(n10131), .C(n4797), .Y(n3276) );
  OAI21X1 U1362 ( .A(n263), .B(n10131), .C(n4794), .Y(n3277) );
  OAI21X1 U1364 ( .A(n265), .B(n10131), .C(n4791), .Y(n3278) );
  OAI21X1 U1366 ( .A(n267), .B(n10131), .C(n4788), .Y(n3279) );
  OAI21X1 U1368 ( .A(n269), .B(n10131), .C(n4785), .Y(n3280) );
  OAI21X1 U1370 ( .A(n271), .B(n10131), .C(n4782), .Y(n3281) );
  OAI21X1 U1372 ( .A(n273), .B(n10131), .C(n4779), .Y(n3282) );
  OAI21X1 U1374 ( .A(n275), .B(n10131), .C(n4776), .Y(n3283) );
  OAI21X1 U1376 ( .A(n277), .B(n10131), .C(n4773), .Y(n3284) );
  OAI21X1 U1378 ( .A(n279), .B(n10131), .C(n4770), .Y(n3285) );
  OAI21X1 U1380 ( .A(n281), .B(n10131), .C(n4767), .Y(n3286) );
  OAI21X1 U1382 ( .A(n283), .B(n10131), .C(n4764), .Y(n3287) );
  OAI21X1 U1384 ( .A(n285), .B(n10131), .C(n4761), .Y(n3288) );
  OAI21X1 U1386 ( .A(n287), .B(n10131), .C(n4758), .Y(n3289) );
  OAI21X1 U1388 ( .A(n289), .B(n10131), .C(n4755), .Y(n3290) );
  OAI21X1 U1390 ( .A(n291), .B(n10131), .C(n4752), .Y(n3291) );
  OAI21X1 U1392 ( .A(n293), .B(n10131), .C(n4749), .Y(n3292) );
  OAI21X1 U1394 ( .A(n295), .B(n10131), .C(n4746), .Y(n3293) );
  OAI21X1 U1396 ( .A(n297), .B(n10131), .C(n4743), .Y(n3294) );
  OAI21X1 U1398 ( .A(n299), .B(n10131), .C(n4740), .Y(n3295) );
  OAI21X1 U1400 ( .A(n301), .B(n10131), .C(n4737), .Y(n3296) );
  OAI21X1 U1402 ( .A(n303), .B(n10131), .C(n4734), .Y(n3297) );
  OAI21X1 U1404 ( .A(n305), .B(n10131), .C(n4731), .Y(n3298) );
  OAI21X1 U1406 ( .A(n307), .B(n10131), .C(n4728), .Y(n3299) );
  OAI21X1 U1408 ( .A(n309), .B(n10131), .C(n4725), .Y(n3300) );
  OAI21X1 U1410 ( .A(n311), .B(n10131), .C(n4722), .Y(n3301) );
  OAI21X1 U1412 ( .A(n313), .B(n10131), .C(n4719), .Y(n3302) );
  OAI21X1 U1414 ( .A(n315), .B(n10131), .C(n4716), .Y(n3303) );
  OAI21X1 U1416 ( .A(n317), .B(n10131), .C(n4713), .Y(n3304) );
  OAI21X1 U1418 ( .A(n319), .B(n10131), .C(n4710), .Y(n3305) );
  OAI21X1 U1420 ( .A(n321), .B(n10131), .C(n4707), .Y(n3306) );
  OAI21X1 U1423 ( .A(n255), .B(n10128), .C(n4704), .Y(n3307) );
  OAI21X1 U1425 ( .A(n257), .B(n10128), .C(n4701), .Y(n3308) );
  OAI21X1 U1427 ( .A(n259), .B(n10128), .C(n4698), .Y(n3309) );
  OAI21X1 U1429 ( .A(n261), .B(n10128), .C(n4695), .Y(n3310) );
  OAI21X1 U1431 ( .A(n263), .B(n10128), .C(n4692), .Y(n3311) );
  OAI21X1 U1433 ( .A(n265), .B(n10128), .C(n4689), .Y(n3312) );
  OAI21X1 U1435 ( .A(n267), .B(n10128), .C(n4686), .Y(n3313) );
  OAI21X1 U1437 ( .A(n269), .B(n10128), .C(n4683), .Y(n3314) );
  OAI21X1 U1439 ( .A(n271), .B(n10128), .C(n4680), .Y(n3315) );
  OAI21X1 U1441 ( .A(n273), .B(n10128), .C(n4677), .Y(n3316) );
  OAI21X1 U1443 ( .A(n275), .B(n10128), .C(n4674), .Y(n3317) );
  OAI21X1 U1445 ( .A(n277), .B(n10128), .C(n4671), .Y(n3318) );
  OAI21X1 U1447 ( .A(n279), .B(n10128), .C(n4668), .Y(n3319) );
  OAI21X1 U1449 ( .A(n281), .B(n10128), .C(n4665), .Y(n3320) );
  OAI21X1 U1451 ( .A(n283), .B(n10128), .C(n4662), .Y(n3321) );
  OAI21X1 U1453 ( .A(n285), .B(n10128), .C(n4659), .Y(n3322) );
  OAI21X1 U1455 ( .A(n287), .B(n10128), .C(n4656), .Y(n3323) );
  OAI21X1 U1457 ( .A(n289), .B(n10128), .C(n4653), .Y(n3324) );
  OAI21X1 U1459 ( .A(n291), .B(n10128), .C(n4650), .Y(n3325) );
  OAI21X1 U1461 ( .A(n293), .B(n10128), .C(n4647), .Y(n3326) );
  OAI21X1 U1463 ( .A(n295), .B(n10128), .C(n4644), .Y(n3327) );
  OAI21X1 U1465 ( .A(n297), .B(n10128), .C(n4641), .Y(n3328) );
  OAI21X1 U1467 ( .A(n299), .B(n10128), .C(n4638), .Y(n3329) );
  OAI21X1 U1469 ( .A(n301), .B(n10128), .C(n4635), .Y(n3330) );
  OAI21X1 U1471 ( .A(n303), .B(n10128), .C(n4632), .Y(n3331) );
  OAI21X1 U1473 ( .A(n305), .B(n10128), .C(n4629), .Y(n3332) );
  OAI21X1 U1475 ( .A(n307), .B(n10128), .C(n4626), .Y(n3333) );
  OAI21X1 U1477 ( .A(n309), .B(n10128), .C(n4623), .Y(n3334) );
  OAI21X1 U1479 ( .A(n311), .B(n10128), .C(n4620), .Y(n3335) );
  OAI21X1 U1481 ( .A(n313), .B(n10128), .C(n4617), .Y(n3336) );
  OAI21X1 U1483 ( .A(n315), .B(n10128), .C(n4614), .Y(n3337) );
  OAI21X1 U1485 ( .A(n317), .B(n10128), .C(n4611), .Y(n3338) );
  OAI21X1 U1487 ( .A(n319), .B(n10128), .C(n4608), .Y(n3339) );
  OAI21X1 U1489 ( .A(n321), .B(n10128), .C(n4605), .Y(n3340) );
  OAI21X1 U1492 ( .A(n255), .B(n10125), .C(n4602), .Y(n3341) );
  OAI21X1 U1494 ( .A(n257), .B(n10125), .C(n4599), .Y(n3342) );
  OAI21X1 U1496 ( .A(n259), .B(n10125), .C(n4596), .Y(n3343) );
  OAI21X1 U1498 ( .A(n261), .B(n10125), .C(n4593), .Y(n3344) );
  OAI21X1 U1500 ( .A(n263), .B(n10125), .C(n4590), .Y(n3345) );
  OAI21X1 U1502 ( .A(n265), .B(n10125), .C(n4587), .Y(n3346) );
  OAI21X1 U1504 ( .A(n267), .B(n10125), .C(n4584), .Y(n3347) );
  OAI21X1 U1506 ( .A(n269), .B(n10125), .C(n4581), .Y(n3348) );
  OAI21X1 U1508 ( .A(n271), .B(n10125), .C(n4578), .Y(n3349) );
  OAI21X1 U1510 ( .A(n273), .B(n10125), .C(n4575), .Y(n3350) );
  OAI21X1 U1512 ( .A(n275), .B(n10125), .C(n4572), .Y(n3351) );
  OAI21X1 U1514 ( .A(n277), .B(n10125), .C(n4569), .Y(n3352) );
  OAI21X1 U1516 ( .A(n279), .B(n10125), .C(n4566), .Y(n3353) );
  OAI21X1 U1518 ( .A(n281), .B(n10125), .C(n4563), .Y(n3354) );
  OAI21X1 U1520 ( .A(n283), .B(n10125), .C(n4560), .Y(n3355) );
  OAI21X1 U1522 ( .A(n285), .B(n10125), .C(n4557), .Y(n3356) );
  OAI21X1 U1524 ( .A(n287), .B(n10125), .C(n4554), .Y(n3357) );
  OAI21X1 U1526 ( .A(n289), .B(n10125), .C(n4551), .Y(n3358) );
  OAI21X1 U1528 ( .A(n291), .B(n10125), .C(n4548), .Y(n3359) );
  OAI21X1 U1530 ( .A(n293), .B(n10125), .C(n4545), .Y(n3360) );
  OAI21X1 U1532 ( .A(n295), .B(n10125), .C(n4542), .Y(n3361) );
  OAI21X1 U1534 ( .A(n297), .B(n10125), .C(n4539), .Y(n3362) );
  OAI21X1 U1536 ( .A(n299), .B(n10125), .C(n4536), .Y(n3363) );
  OAI21X1 U1538 ( .A(n301), .B(n10125), .C(n4533), .Y(n3364) );
  OAI21X1 U1540 ( .A(n303), .B(n10125), .C(n4530), .Y(n3365) );
  OAI21X1 U1542 ( .A(n305), .B(n10125), .C(n4527), .Y(n3366) );
  OAI21X1 U1544 ( .A(n307), .B(n10125), .C(n4524), .Y(n3367) );
  OAI21X1 U1546 ( .A(n309), .B(n10125), .C(n4521), .Y(n3368) );
  OAI21X1 U1548 ( .A(n311), .B(n10125), .C(n4518), .Y(n3369) );
  OAI21X1 U1550 ( .A(n313), .B(n10125), .C(n4515), .Y(n3370) );
  OAI21X1 U1552 ( .A(n315), .B(n10125), .C(n4512), .Y(n3371) );
  OAI21X1 U1554 ( .A(n317), .B(n10125), .C(n4509), .Y(n3372) );
  OAI21X1 U1556 ( .A(n319), .B(n10125), .C(n4506), .Y(n3373) );
  OAI21X1 U1558 ( .A(n321), .B(n10125), .C(n4503), .Y(n3374) );
  OAI21X1 U1561 ( .A(n255), .B(n10122), .C(n4500), .Y(n3375) );
  OAI21X1 U1563 ( .A(n257), .B(n10122), .C(n4497), .Y(n3376) );
  OAI21X1 U1565 ( .A(n259), .B(n10122), .C(n4494), .Y(n3377) );
  OAI21X1 U1567 ( .A(n261), .B(n10122), .C(n4491), .Y(n3378) );
  OAI21X1 U1569 ( .A(n263), .B(n10122), .C(n4488), .Y(n3379) );
  OAI21X1 U1571 ( .A(n265), .B(n10122), .C(n4485), .Y(n3380) );
  OAI21X1 U1573 ( .A(n267), .B(n10122), .C(n4482), .Y(n3381) );
  OAI21X1 U1575 ( .A(n269), .B(n10122), .C(n4479), .Y(n3382) );
  OAI21X1 U1577 ( .A(n271), .B(n10122), .C(n4476), .Y(n3383) );
  OAI21X1 U1579 ( .A(n273), .B(n10122), .C(n4473), .Y(n3384) );
  OAI21X1 U1581 ( .A(n275), .B(n10122), .C(n4470), .Y(n3385) );
  OAI21X1 U1583 ( .A(n277), .B(n10122), .C(n4467), .Y(n3386) );
  OAI21X1 U1585 ( .A(n279), .B(n10122), .C(n4464), .Y(n3387) );
  OAI21X1 U1587 ( .A(n281), .B(n10122), .C(n4461), .Y(n3388) );
  OAI21X1 U1589 ( .A(n283), .B(n10122), .C(n4458), .Y(n3389) );
  OAI21X1 U1591 ( .A(n285), .B(n10122), .C(n4455), .Y(n3390) );
  OAI21X1 U1593 ( .A(n287), .B(n10122), .C(n4452), .Y(n3391) );
  OAI21X1 U1595 ( .A(n289), .B(n10122), .C(n4449), .Y(n3392) );
  OAI21X1 U1597 ( .A(n291), .B(n10122), .C(n4446), .Y(n3393) );
  OAI21X1 U1599 ( .A(n293), .B(n10122), .C(n4443), .Y(n3394) );
  OAI21X1 U1601 ( .A(n295), .B(n10122), .C(n4440), .Y(n3395) );
  OAI21X1 U1603 ( .A(n297), .B(n10122), .C(n4437), .Y(n3396) );
  OAI21X1 U1605 ( .A(n299), .B(n10122), .C(n4434), .Y(n3397) );
  OAI21X1 U1607 ( .A(n301), .B(n10122), .C(n4431), .Y(n3398) );
  OAI21X1 U1609 ( .A(n303), .B(n10122), .C(n4428), .Y(n3399) );
  OAI21X1 U1611 ( .A(n305), .B(n10122), .C(n4425), .Y(n3400) );
  OAI21X1 U1613 ( .A(n307), .B(n10122), .C(n4422), .Y(n3401) );
  OAI21X1 U1615 ( .A(n309), .B(n10122), .C(n4419), .Y(n3402) );
  OAI21X1 U1617 ( .A(n311), .B(n10122), .C(n4416), .Y(n3403) );
  OAI21X1 U1619 ( .A(n313), .B(n10122), .C(n4413), .Y(n3404) );
  OAI21X1 U1621 ( .A(n315), .B(n10122), .C(n4410), .Y(n3405) );
  OAI21X1 U1623 ( .A(n317), .B(n10122), .C(n4407), .Y(n3406) );
  OAI21X1 U1625 ( .A(n319), .B(n10122), .C(n4404), .Y(n3407) );
  OAI21X1 U1627 ( .A(n321), .B(n10122), .C(n4401), .Y(n3408) );
  OAI21X1 U1630 ( .A(n255), .B(n10119), .C(n4398), .Y(n3409) );
  OAI21X1 U1632 ( .A(n257), .B(n10119), .C(n4395), .Y(n3410) );
  OAI21X1 U1634 ( .A(n259), .B(n10119), .C(n4392), .Y(n3411) );
  OAI21X1 U1636 ( .A(n261), .B(n10119), .C(n4389), .Y(n3412) );
  OAI21X1 U1638 ( .A(n263), .B(n10119), .C(n4386), .Y(n3413) );
  OAI21X1 U1640 ( .A(n265), .B(n10119), .C(n4383), .Y(n3414) );
  OAI21X1 U1642 ( .A(n267), .B(n10119), .C(n4380), .Y(n3415) );
  OAI21X1 U1644 ( .A(n269), .B(n10119), .C(n4377), .Y(n3416) );
  OAI21X1 U1646 ( .A(n271), .B(n10119), .C(n4374), .Y(n3417) );
  OAI21X1 U1648 ( .A(n273), .B(n10119), .C(n4371), .Y(n3418) );
  OAI21X1 U1650 ( .A(n275), .B(n10119), .C(n4368), .Y(n3419) );
  OAI21X1 U1652 ( .A(n277), .B(n10119), .C(n4365), .Y(n3420) );
  OAI21X1 U1654 ( .A(n279), .B(n10119), .C(n4362), .Y(n3421) );
  OAI21X1 U1656 ( .A(n281), .B(n10119), .C(n4359), .Y(n3422) );
  OAI21X1 U1658 ( .A(n283), .B(n10119), .C(n4356), .Y(n3423) );
  OAI21X1 U1660 ( .A(n285), .B(n10119), .C(n4353), .Y(n3424) );
  OAI21X1 U1662 ( .A(n287), .B(n10119), .C(n4350), .Y(n3425) );
  OAI21X1 U1664 ( .A(n289), .B(n10119), .C(n4347), .Y(n3426) );
  OAI21X1 U1666 ( .A(n291), .B(n10119), .C(n4344), .Y(n3427) );
  OAI21X1 U1668 ( .A(n293), .B(n10119), .C(n4341), .Y(n3428) );
  OAI21X1 U1670 ( .A(n295), .B(n10119), .C(n4338), .Y(n3429) );
  OAI21X1 U1672 ( .A(n297), .B(n10119), .C(n4335), .Y(n3430) );
  OAI21X1 U1674 ( .A(n299), .B(n10119), .C(n4332), .Y(n3431) );
  OAI21X1 U1676 ( .A(n301), .B(n10119), .C(n4329), .Y(n3432) );
  OAI21X1 U1678 ( .A(n303), .B(n10119), .C(n4326), .Y(n3433) );
  OAI21X1 U1680 ( .A(n305), .B(n10119), .C(n4323), .Y(n3434) );
  OAI21X1 U1682 ( .A(n307), .B(n10119), .C(n4320), .Y(n3435) );
  OAI21X1 U1684 ( .A(n309), .B(n10119), .C(n4317), .Y(n3436) );
  OAI21X1 U1686 ( .A(n311), .B(n10119), .C(n4314), .Y(n3437) );
  OAI21X1 U1688 ( .A(n313), .B(n10119), .C(n4311), .Y(n3438) );
  OAI21X1 U1690 ( .A(n315), .B(n10119), .C(n4308), .Y(n3439) );
  OAI21X1 U1692 ( .A(n317), .B(n10119), .C(n4305), .Y(n3440) );
  OAI21X1 U1694 ( .A(n319), .B(n10119), .C(n4302), .Y(n3441) );
  OAI21X1 U1696 ( .A(n321), .B(n10119), .C(n4299), .Y(n3442) );
  OAI21X1 U1699 ( .A(n255), .B(n10116), .C(n4296), .Y(n3443) );
  OAI21X1 U1701 ( .A(n257), .B(n10116), .C(n4293), .Y(n3444) );
  OAI21X1 U1703 ( .A(n259), .B(n10116), .C(n4290), .Y(n3445) );
  OAI21X1 U1705 ( .A(n261), .B(n10116), .C(n4287), .Y(n3446) );
  OAI21X1 U1707 ( .A(n263), .B(n10116), .C(n4284), .Y(n3447) );
  OAI21X1 U1709 ( .A(n265), .B(n10116), .C(n4281), .Y(n3448) );
  OAI21X1 U1711 ( .A(n267), .B(n10116), .C(n4278), .Y(n3449) );
  OAI21X1 U1713 ( .A(n269), .B(n10116), .C(n4275), .Y(n3450) );
  OAI21X1 U1715 ( .A(n271), .B(n10116), .C(n4272), .Y(n3451) );
  OAI21X1 U1717 ( .A(n273), .B(n10116), .C(n4269), .Y(n3452) );
  OAI21X1 U1719 ( .A(n275), .B(n10116), .C(n4266), .Y(n3453) );
  OAI21X1 U1721 ( .A(n277), .B(n10116), .C(n4263), .Y(n3454) );
  OAI21X1 U1723 ( .A(n279), .B(n10116), .C(n4260), .Y(n3455) );
  OAI21X1 U1725 ( .A(n281), .B(n10116), .C(n4257), .Y(n3456) );
  OAI21X1 U1727 ( .A(n283), .B(n10116), .C(n4254), .Y(n3457) );
  OAI21X1 U1729 ( .A(n285), .B(n10116), .C(n4251), .Y(n3458) );
  OAI21X1 U1731 ( .A(n287), .B(n10116), .C(n4248), .Y(n3459) );
  OAI21X1 U1733 ( .A(n289), .B(n10116), .C(n4245), .Y(n3460) );
  OAI21X1 U1735 ( .A(n291), .B(n10116), .C(n4242), .Y(n3461) );
  OAI21X1 U1737 ( .A(n293), .B(n10116), .C(n4239), .Y(n3462) );
  OAI21X1 U1739 ( .A(n295), .B(n10116), .C(n4236), .Y(n3463) );
  OAI21X1 U1741 ( .A(n297), .B(n10116), .C(n4233), .Y(n3464) );
  OAI21X1 U1743 ( .A(n299), .B(n10116), .C(n4230), .Y(n3465) );
  OAI21X1 U1745 ( .A(n301), .B(n10116), .C(n4227), .Y(n3466) );
  OAI21X1 U1747 ( .A(n303), .B(n10116), .C(n4224), .Y(n3467) );
  OAI21X1 U1749 ( .A(n305), .B(n10116), .C(n4221), .Y(n3468) );
  OAI21X1 U1751 ( .A(n307), .B(n10116), .C(n4218), .Y(n3469) );
  OAI21X1 U1753 ( .A(n309), .B(n10116), .C(n4215), .Y(n3470) );
  OAI21X1 U1755 ( .A(n311), .B(n10116), .C(n4212), .Y(n3471) );
  OAI21X1 U1757 ( .A(n313), .B(n10116), .C(n4209), .Y(n3472) );
  OAI21X1 U1759 ( .A(n315), .B(n10116), .C(n4206), .Y(n3473) );
  OAI21X1 U1761 ( .A(n317), .B(n10116), .C(n4203), .Y(n3474) );
  OAI21X1 U1763 ( .A(n319), .B(n10116), .C(n4200), .Y(n3475) );
  OAI21X1 U1765 ( .A(n321), .B(n10116), .C(n4197), .Y(n3476) );
  INVX1 U1770 ( .A(n10097), .Y(n240) );
  OAI21X1 U1771 ( .A(n255), .B(n1142), .C(n4194), .Y(n3477) );
  OAI21X1 U1773 ( .A(n257), .B(n1142), .C(n4191), .Y(n3478) );
  OAI21X1 U1775 ( .A(n259), .B(n1142), .C(n4188), .Y(n3479) );
  OAI21X1 U1777 ( .A(n261), .B(n1142), .C(n4185), .Y(n3480) );
  OAI21X1 U1779 ( .A(n263), .B(n1142), .C(n4182), .Y(n3481) );
  OAI21X1 U1781 ( .A(n265), .B(n1142), .C(n4179), .Y(n3482) );
  OAI21X1 U1783 ( .A(n267), .B(n1142), .C(n4176), .Y(n3483) );
  OAI21X1 U1785 ( .A(n269), .B(n1142), .C(n4173), .Y(n3484) );
  OAI21X1 U1787 ( .A(n271), .B(n1142), .C(n4170), .Y(n3485) );
  OAI21X1 U1789 ( .A(n273), .B(n1142), .C(n4167), .Y(n3486) );
  OAI21X1 U1791 ( .A(n275), .B(n1142), .C(n4164), .Y(n3487) );
  OAI21X1 U1793 ( .A(n277), .B(n1142), .C(n4161), .Y(n3488) );
  OAI21X1 U1795 ( .A(n279), .B(n1142), .C(n4158), .Y(n3489) );
  OAI21X1 U1797 ( .A(n281), .B(n1142), .C(n4155), .Y(n3490) );
  OAI21X1 U1799 ( .A(n283), .B(n1142), .C(n4152), .Y(n3491) );
  OAI21X1 U1801 ( .A(n285), .B(n1142), .C(n4149), .Y(n3492) );
  OAI21X1 U1803 ( .A(n287), .B(n1142), .C(n4146), .Y(n3493) );
  OAI21X1 U1805 ( .A(n289), .B(n1142), .C(n4143), .Y(n3494) );
  OAI21X1 U1807 ( .A(n291), .B(n1142), .C(n4140), .Y(n3495) );
  OAI21X1 U1809 ( .A(n293), .B(n1142), .C(n4137), .Y(n3496) );
  OAI21X1 U1811 ( .A(n295), .B(n1142), .C(n4134), .Y(n3497) );
  OAI21X1 U1813 ( .A(n297), .B(n1142), .C(n4131), .Y(n3498) );
  OAI21X1 U1815 ( .A(n299), .B(n1142), .C(n4128), .Y(n3499) );
  OAI21X1 U1817 ( .A(n301), .B(n1142), .C(n4125), .Y(n3500) );
  OAI21X1 U1819 ( .A(n303), .B(n1142), .C(n4122), .Y(n3501) );
  OAI21X1 U1821 ( .A(n305), .B(n1142), .C(n4119), .Y(n3502) );
  OAI21X1 U1823 ( .A(n307), .B(n1142), .C(n4116), .Y(n3503) );
  OAI21X1 U1825 ( .A(n309), .B(n1142), .C(n4113), .Y(n3504) );
  OAI21X1 U1827 ( .A(n311), .B(n1142), .C(n4110), .Y(n3505) );
  OAI21X1 U1829 ( .A(n313), .B(n1142), .C(n4107), .Y(n3506) );
  OAI21X1 U1831 ( .A(n315), .B(n1142), .C(n4104), .Y(n3507) );
  OAI21X1 U1833 ( .A(n317), .B(n1142), .C(n4101), .Y(n3508) );
  OAI21X1 U1835 ( .A(n319), .B(n1142), .C(n4098), .Y(n3509) );
  OAI21X1 U1837 ( .A(n321), .B(n1142), .C(n4095), .Y(n3510) );
  NOR3X1 U1840 ( .A(n10087), .B(n10091), .C(n10101), .Y(n323) );
  OAI21X1 U1841 ( .A(n255), .B(n1178), .C(n4092), .Y(n3511) );
  OAI21X1 U1843 ( .A(n257), .B(n1178), .C(n4089), .Y(n3512) );
  OAI21X1 U1845 ( .A(n259), .B(n1178), .C(n4086), .Y(n3513) );
  OAI21X1 U1847 ( .A(n261), .B(n1178), .C(n4083), .Y(n3514) );
  OAI21X1 U1849 ( .A(n263), .B(n1178), .C(n4080), .Y(n3515) );
  OAI21X1 U1851 ( .A(n265), .B(n1178), .C(n4077), .Y(n3516) );
  OAI21X1 U1853 ( .A(n267), .B(n1178), .C(n4074), .Y(n3517) );
  OAI21X1 U1855 ( .A(n269), .B(n1178), .C(n4071), .Y(n3518) );
  OAI21X1 U1857 ( .A(n271), .B(n1178), .C(n4068), .Y(n3519) );
  OAI21X1 U1859 ( .A(n273), .B(n1178), .C(n4065), .Y(n3520) );
  OAI21X1 U1861 ( .A(n275), .B(n1178), .C(n4062), .Y(n3521) );
  OAI21X1 U1863 ( .A(n277), .B(n1178), .C(n4059), .Y(n3522) );
  OAI21X1 U1865 ( .A(n279), .B(n1178), .C(n4056), .Y(n3523) );
  OAI21X1 U1867 ( .A(n281), .B(n1178), .C(n4053), .Y(n3524) );
  OAI21X1 U1869 ( .A(n283), .B(n1178), .C(n4050), .Y(n3525) );
  OAI21X1 U1871 ( .A(n285), .B(n1178), .C(n4047), .Y(n3526) );
  OAI21X1 U1873 ( .A(n287), .B(n1178), .C(n4044), .Y(n3527) );
  OAI21X1 U1875 ( .A(n289), .B(n1178), .C(n4041), .Y(n3528) );
  OAI21X1 U1877 ( .A(n291), .B(n1178), .C(n4038), .Y(n3529) );
  OAI21X1 U1879 ( .A(n293), .B(n1178), .C(n4035), .Y(n3530) );
  OAI21X1 U1881 ( .A(n295), .B(n1178), .C(n4032), .Y(n3531) );
  OAI21X1 U1883 ( .A(n297), .B(n1178), .C(n4029), .Y(n3532) );
  OAI21X1 U1885 ( .A(n299), .B(n1178), .C(n4026), .Y(n3533) );
  OAI21X1 U1887 ( .A(n301), .B(n1178), .C(n4023), .Y(n3534) );
  OAI21X1 U1889 ( .A(n303), .B(n1178), .C(n4020), .Y(n3535) );
  OAI21X1 U1891 ( .A(n305), .B(n1178), .C(n4017), .Y(n3536) );
  OAI21X1 U1893 ( .A(n307), .B(n1178), .C(n4014), .Y(n3537) );
  OAI21X1 U1895 ( .A(n309), .B(n1178), .C(n4011), .Y(n3538) );
  OAI21X1 U1897 ( .A(n311), .B(n1178), .C(n4008), .Y(n3539) );
  OAI21X1 U1899 ( .A(n313), .B(n1178), .C(n4005), .Y(n3540) );
  OAI21X1 U1901 ( .A(n315), .B(n1178), .C(n4002), .Y(n3541) );
  OAI21X1 U1903 ( .A(n317), .B(n1178), .C(n3999), .Y(n3542) );
  OAI21X1 U1905 ( .A(n319), .B(n1178), .C(n3996), .Y(n3543) );
  OAI21X1 U1907 ( .A(n321), .B(n1178), .C(n3993), .Y(n3544) );
  NOR3X1 U1910 ( .A(n10088), .B(n10091), .C(n246), .Y(n360) );
  OAI21X1 U1911 ( .A(n255), .B(n10500), .C(n3990), .Y(n3545) );
  OAI21X1 U1913 ( .A(n257), .B(n10500), .C(n3987), .Y(n3546) );
  OAI21X1 U1915 ( .A(n259), .B(n10500), .C(n3984), .Y(n3547) );
  OAI21X1 U1917 ( .A(n261), .B(n10500), .C(n3981), .Y(n3548) );
  OAI21X1 U1919 ( .A(n263), .B(n10500), .C(n3978), .Y(n3549) );
  OAI21X1 U1921 ( .A(n265), .B(n10500), .C(n3975), .Y(n3550) );
  OAI21X1 U1923 ( .A(n267), .B(n10500), .C(n3972), .Y(n3551) );
  OAI21X1 U1925 ( .A(n269), .B(n10500), .C(n3969), .Y(n3552) );
  OAI21X1 U1927 ( .A(n271), .B(n10500), .C(n3966), .Y(n3553) );
  OAI21X1 U1929 ( .A(n273), .B(n10500), .C(n3963), .Y(n3554) );
  OAI21X1 U1931 ( .A(n275), .B(n10500), .C(n3960), .Y(n3555) );
  OAI21X1 U1933 ( .A(n277), .B(n10500), .C(n3957), .Y(n3556) );
  OAI21X1 U1935 ( .A(n279), .B(n10500), .C(n3954), .Y(n3557) );
  OAI21X1 U1937 ( .A(n281), .B(n10500), .C(n3951), .Y(n3558) );
  OAI21X1 U1939 ( .A(n283), .B(n10500), .C(n3948), .Y(n3559) );
  OAI21X1 U1941 ( .A(n285), .B(n10500), .C(n3945), .Y(n3560) );
  OAI21X1 U1943 ( .A(n287), .B(n10500), .C(n3942), .Y(n3561) );
  OAI21X1 U1945 ( .A(n289), .B(n10500), .C(n3939), .Y(n3562) );
  OAI21X1 U1947 ( .A(n291), .B(n10500), .C(n3936), .Y(n3563) );
  OAI21X1 U1949 ( .A(n293), .B(n10500), .C(n3933), .Y(n3564) );
  OAI21X1 U1951 ( .A(n295), .B(n10500), .C(n3930), .Y(n3565) );
  OAI21X1 U1953 ( .A(n297), .B(n10500), .C(n3927), .Y(n3566) );
  OAI21X1 U1955 ( .A(n299), .B(n10500), .C(n3924), .Y(n3567) );
  OAI21X1 U1957 ( .A(n301), .B(n10500), .C(n3921), .Y(n3568) );
  OAI21X1 U1959 ( .A(n303), .B(n10500), .C(n3918), .Y(n3569) );
  OAI21X1 U1961 ( .A(n305), .B(n10500), .C(n3915), .Y(n3570) );
  OAI21X1 U1963 ( .A(n307), .B(n10500), .C(n3912), .Y(n3571) );
  OAI21X1 U1965 ( .A(n309), .B(n10500), .C(n3909), .Y(n3572) );
  OAI21X1 U1967 ( .A(n311), .B(n10500), .C(n3906), .Y(n3573) );
  OAI21X1 U1969 ( .A(n313), .B(n10500), .C(n3903), .Y(n3574) );
  OAI21X1 U1971 ( .A(n315), .B(n10500), .C(n3900), .Y(n3575) );
  OAI21X1 U1973 ( .A(n317), .B(n10500), .C(n3897), .Y(n3576) );
  OAI21X1 U1975 ( .A(n319), .B(n10500), .C(n3894), .Y(n3577) );
  OAI21X1 U1977 ( .A(n321), .B(n10500), .C(n3891), .Y(n3578) );
  OAI21X1 U1981 ( .A(n255), .B(n1249), .C(n3888), .Y(n3579) );
  OAI21X1 U1983 ( .A(n257), .B(n1249), .C(n3885), .Y(n3580) );
  OAI21X1 U1985 ( .A(n259), .B(n1249), .C(n3882), .Y(n3581) );
  OAI21X1 U1987 ( .A(n261), .B(n1249), .C(n3879), .Y(n3582) );
  OAI21X1 U1989 ( .A(n263), .B(n1249), .C(n3876), .Y(n3583) );
  OAI21X1 U1991 ( .A(n265), .B(n1249), .C(n3873), .Y(n3584) );
  OAI21X1 U1993 ( .A(n267), .B(n1249), .C(n3870), .Y(n3585) );
  OAI21X1 U1995 ( .A(n269), .B(n1249), .C(n3867), .Y(n3586) );
  OAI21X1 U1997 ( .A(n271), .B(n1249), .C(n3864), .Y(n3587) );
  OAI21X1 U1999 ( .A(n273), .B(n1249), .C(n3861), .Y(n3588) );
  OAI21X1 U2001 ( .A(n275), .B(n1249), .C(n3858), .Y(n3589) );
  OAI21X1 U2003 ( .A(n277), .B(n1249), .C(n3855), .Y(n3590) );
  OAI21X1 U2005 ( .A(n279), .B(n1249), .C(n3852), .Y(n3591) );
  OAI21X1 U2007 ( .A(n281), .B(n1249), .C(n3849), .Y(n3592) );
  OAI21X1 U2009 ( .A(n283), .B(n1249), .C(n3846), .Y(n3593) );
  OAI21X1 U2011 ( .A(n285), .B(n1249), .C(n3843), .Y(n3594) );
  OAI21X1 U2013 ( .A(n287), .B(n1249), .C(n3840), .Y(n3595) );
  OAI21X1 U2015 ( .A(n289), .B(n1249), .C(n3837), .Y(n3596) );
  OAI21X1 U2017 ( .A(n291), .B(n1249), .C(n3834), .Y(n3597) );
  OAI21X1 U2019 ( .A(n293), .B(n1249), .C(n3831), .Y(n3598) );
  OAI21X1 U2021 ( .A(n295), .B(n1249), .C(n3828), .Y(n3599) );
  OAI21X1 U2023 ( .A(n297), .B(n1249), .C(n3825), .Y(n3600) );
  OAI21X1 U2025 ( .A(n299), .B(n1249), .C(n3822), .Y(n3601) );
  OAI21X1 U2027 ( .A(n301), .B(n1249), .C(n3819), .Y(n3602) );
  OAI21X1 U2029 ( .A(n303), .B(n1249), .C(n3816), .Y(n3603) );
  OAI21X1 U2031 ( .A(n305), .B(n1249), .C(n3813), .Y(n3604) );
  OAI21X1 U2033 ( .A(n307), .B(n1249), .C(n3810), .Y(n3605) );
  OAI21X1 U2035 ( .A(n309), .B(n1249), .C(n3807), .Y(n3606) );
  OAI21X1 U2037 ( .A(n311), .B(n1249), .C(n3804), .Y(n3607) );
  OAI21X1 U2039 ( .A(n313), .B(n1249), .C(n3801), .Y(n3608) );
  OAI21X1 U2041 ( .A(n315), .B(n1249), .C(n3798), .Y(n3609) );
  OAI21X1 U2043 ( .A(n317), .B(n1249), .C(n3795), .Y(n3610) );
  OAI21X1 U2045 ( .A(n319), .B(n1249), .C(n3792), .Y(n3611) );
  OAI21X1 U2047 ( .A(n321), .B(n1249), .C(n3789), .Y(n3612) );
  OAI21X1 U2051 ( .A(n255), .B(n1284), .C(n3786), .Y(n3613) );
  OAI21X1 U2053 ( .A(n257), .B(n1284), .C(n3783), .Y(n3614) );
  OAI21X1 U2055 ( .A(n259), .B(n1284), .C(n3780), .Y(n3615) );
  OAI21X1 U2057 ( .A(n261), .B(n1284), .C(n3777), .Y(n3616) );
  OAI21X1 U2059 ( .A(n263), .B(n1284), .C(n3774), .Y(n3617) );
  OAI21X1 U2061 ( .A(n265), .B(n1284), .C(n3771), .Y(n3618) );
  OAI21X1 U2063 ( .A(n267), .B(n1284), .C(n3768), .Y(n3619) );
  OAI21X1 U2065 ( .A(n269), .B(n1284), .C(n3765), .Y(n3620) );
  OAI21X1 U2067 ( .A(n271), .B(n1284), .C(n3762), .Y(n3621) );
  OAI21X1 U2069 ( .A(n273), .B(n1284), .C(n3759), .Y(n3622) );
  OAI21X1 U2071 ( .A(n275), .B(n1284), .C(n3756), .Y(n3623) );
  OAI21X1 U2073 ( .A(n277), .B(n1284), .C(n3753), .Y(n3624) );
  OAI21X1 U2075 ( .A(n279), .B(n1284), .C(n3750), .Y(n3625) );
  OAI21X1 U2077 ( .A(n281), .B(n1284), .C(n2656), .Y(n3626) );
  OAI21X1 U2079 ( .A(n283), .B(n1284), .C(n2618), .Y(n3627) );
  OAI21X1 U2081 ( .A(n285), .B(n1284), .C(n2612), .Y(n3628) );
  OAI21X1 U2083 ( .A(n287), .B(n1284), .C(n2606), .Y(n3629) );
  OAI21X1 U2085 ( .A(n289), .B(n1284), .C(n2600), .Y(n3630) );
  OAI21X1 U2087 ( .A(n291), .B(n1284), .C(n2594), .Y(n3631) );
  OAI21X1 U2089 ( .A(n293), .B(n1284), .C(n2588), .Y(n3632) );
  OAI21X1 U2091 ( .A(n295), .B(n1284), .C(n2582), .Y(n3633) );
  OAI21X1 U2093 ( .A(n297), .B(n1284), .C(n2576), .Y(n3634) );
  OAI21X1 U2095 ( .A(n299), .B(n1284), .C(n2570), .Y(n3635) );
  OAI21X1 U2097 ( .A(n301), .B(n1284), .C(n2564), .Y(n3636) );
  OAI21X1 U2099 ( .A(n303), .B(n1284), .C(n2558), .Y(n3637) );
  OAI21X1 U2101 ( .A(n305), .B(n1284), .C(n2545), .Y(n3638) );
  OAI21X1 U2103 ( .A(n307), .B(n1284), .C(n2531), .Y(n3639) );
  OAI21X1 U2105 ( .A(n309), .B(n1284), .C(n2528), .Y(n3640) );
  OAI21X1 U2107 ( .A(n311), .B(n1284), .C(n2525), .Y(n3641) );
  OAI21X1 U2109 ( .A(n313), .B(n1284), .C(n2522), .Y(n3642) );
  OAI21X1 U2111 ( .A(n315), .B(n1284), .C(n2519), .Y(n3643) );
  OAI21X1 U2113 ( .A(n317), .B(n1284), .C(n2516), .Y(n3644) );
  OAI21X1 U2115 ( .A(n319), .B(n1284), .C(n2513), .Y(n3645) );
  OAI21X1 U2117 ( .A(n321), .B(n1284), .C(n2510), .Y(n3646) );
  OAI21X1 U2121 ( .A(n255), .B(n10504), .C(n2507), .Y(n3647) );
  OAI21X1 U2123 ( .A(n257), .B(n10504), .C(n2504), .Y(n3648) );
  OAI21X1 U2125 ( .A(n259), .B(n10504), .C(n2501), .Y(n3649) );
  OAI21X1 U2127 ( .A(n261), .B(n10504), .C(n2498), .Y(n3650) );
  OAI21X1 U2129 ( .A(n263), .B(n10504), .C(n1985), .Y(n3651) );
  OAI21X1 U2131 ( .A(n265), .B(n10504), .C(n1982), .Y(n3652) );
  OAI21X1 U2133 ( .A(n267), .B(n10504), .C(n1979), .Y(n3653) );
  OAI21X1 U2135 ( .A(n269), .B(n10504), .C(n1976), .Y(n3654) );
  OAI21X1 U2137 ( .A(n271), .B(n10504), .C(n1973), .Y(n3655) );
  OAI21X1 U2139 ( .A(n273), .B(n10504), .C(n1970), .Y(n3656) );
  OAI21X1 U2141 ( .A(n275), .B(n10504), .C(n1967), .Y(n3657) );
  OAI21X1 U2143 ( .A(n277), .B(n10504), .C(n1964), .Y(n3658) );
  OAI21X1 U2145 ( .A(n279), .B(n10504), .C(n1961), .Y(n3659) );
  OAI21X1 U2147 ( .A(n281), .B(n10504), .C(n1958), .Y(n3660) );
  OAI21X1 U2149 ( .A(n283), .B(n10504), .C(n1955), .Y(n3661) );
  OAI21X1 U2151 ( .A(n285), .B(n10504), .C(n1952), .Y(n3662) );
  OAI21X1 U2153 ( .A(n287), .B(n10504), .C(n1949), .Y(n3663) );
  OAI21X1 U2155 ( .A(n289), .B(n10504), .C(n1946), .Y(n3664) );
  OAI21X1 U2157 ( .A(n291), .B(n10504), .C(n1943), .Y(n3665) );
  OAI21X1 U2159 ( .A(n293), .B(n10504), .C(n1940), .Y(n3666) );
  OAI21X1 U2161 ( .A(n295), .B(n10504), .C(n1937), .Y(n3667) );
  OAI21X1 U2163 ( .A(n297), .B(n10504), .C(n1934), .Y(n3668) );
  OAI21X1 U2165 ( .A(n299), .B(n10504), .C(n1931), .Y(n3669) );
  OAI21X1 U2167 ( .A(n301), .B(n10504), .C(n1928), .Y(n3670) );
  OAI21X1 U2169 ( .A(n303), .B(n10504), .C(n1925), .Y(n3671) );
  OAI21X1 U2171 ( .A(n305), .B(n10504), .C(n1922), .Y(n3672) );
  OAI21X1 U2173 ( .A(n307), .B(n10504), .C(n1919), .Y(n3673) );
  OAI21X1 U2175 ( .A(n309), .B(n10504), .C(n1916), .Y(n3674) );
  OAI21X1 U2177 ( .A(n311), .B(n10504), .C(n1913), .Y(n3675) );
  OAI21X1 U2179 ( .A(n313), .B(n10504), .C(n1910), .Y(n3676) );
  OAI21X1 U2181 ( .A(n315), .B(n10504), .C(n1907), .Y(n3677) );
  OAI21X1 U2183 ( .A(n317), .B(n10504), .C(n1904), .Y(n3678) );
  OAI21X1 U2185 ( .A(n319), .B(n10504), .C(n1901), .Y(n3679) );
  OAI21X1 U2187 ( .A(n321), .B(n10504), .C(n1898), .Y(n3680) );
  OAI21X1 U2191 ( .A(n255), .B(n10496), .C(n1895), .Y(n3681) );
  OAI21X1 U2193 ( .A(n257), .B(n10496), .C(n1892), .Y(n3682) );
  OAI21X1 U2195 ( .A(n259), .B(n10496), .C(n1889), .Y(n3683) );
  OAI21X1 U2197 ( .A(n261), .B(n10496), .C(n1886), .Y(n3684) );
  OAI21X1 U2199 ( .A(n263), .B(n10496), .C(n1883), .Y(n3685) );
  OAI21X1 U2201 ( .A(n265), .B(n10496), .C(n1880), .Y(n3686) );
  OAI21X1 U2203 ( .A(n267), .B(n10496), .C(n1877), .Y(n3687) );
  OAI21X1 U2205 ( .A(n269), .B(n10496), .C(n1874), .Y(n3688) );
  OAI21X1 U2207 ( .A(n271), .B(n10496), .C(n1871), .Y(n3689) );
  OAI21X1 U2209 ( .A(n273), .B(n10496), .C(n1868), .Y(n3690) );
  OAI21X1 U2211 ( .A(n275), .B(n10496), .C(n1865), .Y(n3691) );
  OAI21X1 U2213 ( .A(n277), .B(n10496), .C(n1862), .Y(n3692) );
  OAI21X1 U2215 ( .A(n279), .B(n10496), .C(n1859), .Y(n3693) );
  OAI21X1 U2217 ( .A(n281), .B(n10496), .C(n1856), .Y(n3694) );
  OAI21X1 U2219 ( .A(n283), .B(n10496), .C(n1853), .Y(n3695) );
  OAI21X1 U2221 ( .A(n285), .B(n10496), .C(n1850), .Y(n3696) );
  OAI21X1 U2223 ( .A(n287), .B(n10496), .C(n1847), .Y(n3697) );
  OAI21X1 U2225 ( .A(n289), .B(n10496), .C(n1844), .Y(n3698) );
  OAI21X1 U2227 ( .A(n291), .B(n10496), .C(n1841), .Y(n3699) );
  OAI21X1 U2229 ( .A(n293), .B(n10496), .C(n1838), .Y(n3700) );
  OAI21X1 U2231 ( .A(n295), .B(n10496), .C(n1835), .Y(n3701) );
  OAI21X1 U2233 ( .A(n297), .B(n10496), .C(n1832), .Y(n3702) );
  OAI21X1 U2235 ( .A(n299), .B(n10496), .C(n1829), .Y(n3703) );
  OAI21X1 U2237 ( .A(n301), .B(n10496), .C(n1826), .Y(n3704) );
  OAI21X1 U2239 ( .A(n303), .B(n10496), .C(n1823), .Y(n3705) );
  OAI21X1 U2241 ( .A(n305), .B(n10496), .C(n1820), .Y(n3706) );
  OAI21X1 U2243 ( .A(n307), .B(n10496), .C(n1817), .Y(n3707) );
  OAI21X1 U2245 ( .A(n309), .B(n10496), .C(n1814), .Y(n3708) );
  OAI21X1 U2247 ( .A(n311), .B(n10496), .C(n1811), .Y(n3709) );
  OAI21X1 U2249 ( .A(n313), .B(n10496), .C(n1808), .Y(n3710) );
  OAI21X1 U2251 ( .A(n315), .B(n10496), .C(n1805), .Y(n3711) );
  OAI21X1 U2253 ( .A(n317), .B(n10496), .C(n1802), .Y(n3712) );
  OAI21X1 U2255 ( .A(n319), .B(n10496), .C(n1799), .Y(n3713) );
  OAI21X1 U2257 ( .A(n321), .B(n10496), .C(n1796), .Y(n3714) );
  NOR3X1 U2260 ( .A(n242), .B(n10101), .C(n244), .Y(n540) );
  OAI21X1 U2261 ( .A(n255), .B(n10498), .C(n1793), .Y(n3715) );
  INVX1 U2263 ( .A(data_in[33]), .Y(n255) );
  OAI21X1 U2264 ( .A(n257), .B(n10498), .C(n1790), .Y(n3716) );
  INVX1 U2266 ( .A(data_in[32]), .Y(n257) );
  OAI21X1 U2267 ( .A(n259), .B(n10498), .C(n1787), .Y(n3717) );
  INVX1 U2269 ( .A(data_in[31]), .Y(n259) );
  OAI21X1 U2270 ( .A(n261), .B(n10498), .C(n1784), .Y(n3718) );
  INVX1 U2272 ( .A(data_in[30]), .Y(n261) );
  OAI21X1 U2273 ( .A(n263), .B(n10498), .C(n1781), .Y(n3719) );
  INVX1 U2275 ( .A(data_in[29]), .Y(n263) );
  OAI21X1 U2276 ( .A(n265), .B(n10498), .C(n1778), .Y(n3720) );
  INVX1 U2278 ( .A(data_in[28]), .Y(n265) );
  OAI21X1 U2279 ( .A(n267), .B(n10498), .C(n1775), .Y(n3721) );
  INVX1 U2281 ( .A(data_in[27]), .Y(n267) );
  OAI21X1 U2282 ( .A(n269), .B(n10498), .C(n1772), .Y(n3722) );
  INVX1 U2284 ( .A(data_in[26]), .Y(n269) );
  OAI21X1 U2285 ( .A(n271), .B(n10498), .C(n1769), .Y(n3723) );
  INVX1 U2287 ( .A(data_in[25]), .Y(n271) );
  OAI21X1 U2288 ( .A(n273), .B(n10498), .C(n1766), .Y(n3724) );
  INVX1 U2290 ( .A(data_in[24]), .Y(n273) );
  OAI21X1 U2291 ( .A(n275), .B(n10498), .C(n1763), .Y(n3725) );
  INVX1 U2293 ( .A(data_in[23]), .Y(n275) );
  OAI21X1 U2294 ( .A(n277), .B(n10498), .C(n1760), .Y(n3726) );
  INVX1 U2296 ( .A(data_in[22]), .Y(n277) );
  OAI21X1 U2297 ( .A(n279), .B(n10498), .C(n1757), .Y(n3727) );
  INVX1 U2299 ( .A(data_in[21]), .Y(n279) );
  OAI21X1 U2300 ( .A(n281), .B(n10498), .C(n1754), .Y(n3728) );
  INVX1 U2302 ( .A(data_in[20]), .Y(n281) );
  OAI21X1 U2303 ( .A(n283), .B(n10498), .C(n1751), .Y(n3729) );
  INVX1 U2305 ( .A(data_in[19]), .Y(n283) );
  OAI21X1 U2306 ( .A(n285), .B(n10498), .C(n1748), .Y(n3730) );
  INVX1 U2308 ( .A(data_in[18]), .Y(n285) );
  OAI21X1 U2309 ( .A(n287), .B(n10498), .C(n1745), .Y(n3731) );
  INVX1 U2311 ( .A(data_in[17]), .Y(n287) );
  OAI21X1 U2312 ( .A(n289), .B(n10498), .C(n1742), .Y(n3732) );
  INVX1 U2314 ( .A(data_in[16]), .Y(n289) );
  OAI21X1 U2315 ( .A(n291), .B(n10498), .C(n1739), .Y(n3733) );
  INVX1 U2317 ( .A(data_in[15]), .Y(n291) );
  OAI21X1 U2318 ( .A(n293), .B(n10498), .C(n1736), .Y(n3734) );
  INVX1 U2320 ( .A(data_in[14]), .Y(n293) );
  OAI21X1 U2321 ( .A(n295), .B(n10498), .C(n1733), .Y(n3735) );
  INVX1 U2323 ( .A(data_in[13]), .Y(n295) );
  OAI21X1 U2324 ( .A(n297), .B(n10498), .C(n1730), .Y(n3736) );
  INVX1 U2326 ( .A(data_in[12]), .Y(n297) );
  OAI21X1 U2327 ( .A(n299), .B(n10498), .C(n1727), .Y(n3737) );
  INVX1 U2329 ( .A(data_in[11]), .Y(n299) );
  OAI21X1 U2330 ( .A(n301), .B(n10498), .C(n1724), .Y(n3738) );
  INVX1 U2332 ( .A(data_in[10]), .Y(n301) );
  OAI21X1 U2333 ( .A(n303), .B(n10498), .C(n1721), .Y(n3739) );
  INVX1 U2335 ( .A(data_in[9]), .Y(n303) );
  OAI21X1 U2336 ( .A(n305), .B(n10498), .C(n1718), .Y(n3740) );
  INVX1 U2338 ( .A(data_in[8]), .Y(n305) );
  OAI21X1 U2339 ( .A(n307), .B(n10498), .C(n1432), .Y(n3741) );
  INVX1 U2341 ( .A(data_in[7]), .Y(n307) );
  OAI21X1 U2342 ( .A(n309), .B(n10498), .C(n252), .Y(n3742) );
  INVX1 U2344 ( .A(data_in[6]), .Y(n309) );
  OAI21X1 U2345 ( .A(n311), .B(n10498), .C(n192), .Y(n3743) );
  INVX1 U2347 ( .A(data_in[5]), .Y(n311) );
  OAI21X1 U2348 ( .A(n313), .B(n10498), .C(n189), .Y(n3744) );
  INVX1 U2350 ( .A(data_in[4]), .Y(n313) );
  OAI21X1 U2351 ( .A(n315), .B(n10498), .C(n186), .Y(n3745) );
  INVX1 U2353 ( .A(data_in[3]), .Y(n315) );
  OAI21X1 U2354 ( .A(n317), .B(n10498), .C(n183), .Y(n3746) );
  INVX1 U2356 ( .A(data_in[2]), .Y(n317) );
  OAI21X1 U2357 ( .A(n319), .B(n10498), .C(n180), .Y(n3747) );
  INVX1 U2359 ( .A(data_in[1]), .Y(n319) );
  OAI21X1 U2360 ( .A(n321), .B(n10498), .C(n177), .Y(n3748) );
  NOR3X1 U2363 ( .A(n244), .B(n242), .C(n246), .Y(n576) );
  INVX1 U2364 ( .A(n10101), .Y(n246) );
  NAND3X1 U2366 ( .A(n10104), .B(n237), .C(n10097), .Y(n1425) );
  INVX1 U2368 ( .A(data_in[0]), .Y(n321) );
  XOR2X1 U2369 ( .A(n10087), .B(n10101), .Y(n24) );
  INVX1 U2372 ( .A(n10091), .Y(n242) );
  INVX1 U2374 ( .A(n10088), .Y(n244) );
  XOR2X1 U2375 ( .A(n10097), .B(n10091), .Y(n22) );
  XOR2X1 U2376 ( .A(n10104), .B(n10097), .Y(n21) );
  XOR2X1 U2377 ( .A(n10081), .B(n10104), .Y(n20) );
  XOR2X1 U2378 ( .A(n10663), .B(n10689), .Y(n19) );
  XOR2X1 U2379 ( .A(n10649), .B(n10663), .Y(n18) );
  XOR2X1 U2380 ( .A(n10111), .B(n10649), .Y(n17) );
  XOR2X1 U2381 ( .A(n10529), .B(n10111), .Y(n16) );
  XOR2X1 U2382 ( .A(n10047), .B(n10529), .Y(n15) );
  NAND3X1 U2383 ( .A(n6681), .B(fillcount[5]), .C(n1427), .Y(full_bar) );
  NOR3X1 U2384 ( .A(fillcount[2]), .B(fillcount[4]), .C(fillcount[3]), .Y(
        n1427) );
  NAND3X1 U2386 ( .A(n8), .B(n1429), .C(n6690), .Y(n11796) );
  XOR2X1 U2390 ( .A(n250), .B(n10017), .Y(n1429) );
  INVX1 U2391 ( .A(n10046), .Y(n250) );
  AOI22X1 U2392 ( .A(n1435), .B(n152), .C(n1437), .D(n6684), .Y(n1428) );
  NAND3X1 U2393 ( .A(n1439), .B(n10659), .C(n1440), .Y(n1438) );
  XOR2X1 U2394 ( .A(n10733), .B(n1441), .Y(n1440) );
  XOR2X1 U2397 ( .A(n10044), .B(n10685), .Y(n1439) );
  NAND3X1 U2399 ( .A(n1442), .B(n1443), .C(n10657), .Y(n1436) );
  XOR2X1 U2400 ( .A(n10044), .B(n10663), .Y(n1443) );
  XOR2X1 U2401 ( .A(n10689), .B(n1441), .Y(n1442) );
  XOR2X1 U2402 ( .A(n10043), .B(n26), .Y(n1441) );
  XNOR2X1 U2404 ( .A(n1434), .B(n6696), .Y(n1437) );
  XOR2X1 U2405 ( .A(n1433), .B(n6699), .Y(n1434) );
  XOR2X1 U2406 ( .A(n10016), .B(n25), .Y(n1433) );
  HAX1 add_176_U1_1_1 ( .A(n10663), .B(n10721), .YC(add_176_carry[2]), .YS(
        n106) );
  HAX1 add_176_U1_1_2 ( .A(n10649), .B(add_176_carry[2]), .YC(add_176_carry[3]), .YS(n107) );
  HAX1 add_176_U1_1_3 ( .A(n10111), .B(add_176_carry[3]), .YC(add_176_carry[4]), .YS(n108) );
  HAX1 add_176_U1_1_4 ( .A(n10529), .B(add_176_carry[4]), .YC(add_176_carry[5]), .YS(n109) );
  HAX1 add_158_U1_1_1 ( .A(n10087), .B(n10101), .YC(add_158_carry[2]), .YS(n34) );
  HAX1 add_158_U1_1_2 ( .A(n10091), .B(add_158_carry[2]), .YC(add_158_carry[3]), .YS(n35) );
  HAX1 add_158_U1_1_3 ( .A(n10097), .B(add_158_carry[3]), .YC(add_158_carry[4]), .YS(n36) );
  HAX1 add_158_U1_1_4 ( .A(n10104), .B(add_158_carry[4]), .YC(add_158_carry[5]), .YS(n37) );
  FAX1 r301_U2_1 ( .A(n10087), .B(r301_B_not_1_), .C(n32), .YC(r301_carry[2]), 
        .YS(fillcount[1]) );
  FAX1 r301_U2_2 ( .A(n10091), .B(r301_B_not_2_), .C(r301_carry[2]), .YC(
        r301_carry[3]), .YS(fillcount[2]) );
  FAX1 r301_U2_3 ( .A(n10097), .B(r301_B_not_3_), .C(r301_carry[3]), .YC(
        r301_carry[4]), .YS(fillcount[3]) );
  FAX1 r301_U2_5 ( .A(n10081), .B(r301_B_not_5_), .C(n28), .YC(), .YS(
        fillcount[5]) );
  DFFSR data_out_reg_33_ ( .D(n2553), .CLK(rclk), .R(n10634), .S(1'b1), .Q(
        n11797) );
  DFFSR data_out_reg_30_ ( .D(n2559), .CLK(rclk), .R(n10634), .S(1'b1), .Q(
        n11800) );
  DFFSR data_out_reg_29_ ( .D(n2561), .CLK(rclk), .R(n10634), .S(1'b1), .Q(
        n11801) );
  DFFSR data_out_reg_28_ ( .D(n2563), .CLK(rclk), .R(n10634), .S(1'b1), .Q(
        n11802) );
  DFFSR data_out_reg_27_ ( .D(n2565), .CLK(rclk), .R(n10634), .S(1'b1), .Q(
        n11803) );
  DFFSR data_out_reg_26_ ( .D(n2567), .CLK(rclk), .R(n10634), .S(1'b1), .Q(
        n11804) );
  DFFSR data_out_reg_25_ ( .D(n2569), .CLK(rclk), .R(n10634), .S(1'b1), .Q(
        n11805) );
  DFFSR data_out_reg_24_ ( .D(n2571), .CLK(rclk), .R(n10634), .S(1'b1), .Q(
        n11806) );
  DFFSR data_out_reg_23_ ( .D(n2573), .CLK(rclk), .R(n10634), .S(1'b1), .Q(
        n11807) );
  DFFSR data_out_reg_22_ ( .D(n2575), .CLK(rclk), .R(n10634), .S(1'b1), .Q(
        n11808) );
  DFFSR data_out_reg_21_ ( .D(n2577), .CLK(rclk), .R(n10634), .S(1'b1), .Q(
        n11809) );
  DFFSR data_out_reg_20_ ( .D(n2579), .CLK(rclk), .R(n10634), .S(1'b1), .Q(
        n11810) );
  DFFSR data_out_reg_19_ ( .D(n2581), .CLK(rclk), .R(n10634), .S(1'b1), .Q(
        n11811) );
  DFFSR data_out_reg_18_ ( .D(n2583), .CLK(rclk), .R(n10634), .S(1'b1), .Q(
        n11812) );
  DFFSR data_out_reg_17_ ( .D(n2585), .CLK(rclk), .R(n10634), .S(1'b1), .Q(
        n11813) );
  DFFSR data_out_reg_16_ ( .D(n2587), .CLK(rclk), .R(n10634), .S(1'b1), .Q(
        n11814) );
  DFFSR data_out_reg_15_ ( .D(n2589), .CLK(rclk), .R(n10634), .S(1'b1), .Q(
        n11815) );
  DFFSR data_out_reg_14_ ( .D(n2591), .CLK(rclk), .R(n10634), .S(1'b1), .Q(
        n11816) );
  DFFSR data_out_reg_13_ ( .D(n2593), .CLK(rclk), .R(n10634), .S(1'b1), .Q(
        n11817) );
  DFFSR data_out_reg_12_ ( .D(n2595), .CLK(rclk), .R(n10634), .S(1'b1), .Q(
        n11818) );
  DFFSR data_out_reg_11_ ( .D(n2597), .CLK(rclk), .R(n10634), .S(1'b1), .Q(
        n11819) );
  DFFSR data_out_reg_10_ ( .D(n2599), .CLK(rclk), .R(n10634), .S(1'b1), .Q(
        n11820) );
  DFFSR data_out_reg_9_ ( .D(n2601), .CLK(rclk), .R(n10634), .S(1'b1), .Q(
        n11821) );
  DFFSR data_out_reg_8_ ( .D(n2603), .CLK(rclk), .R(n10634), .S(1'b1), .Q(
        n11822) );
  DFFSR data_out_reg_7_ ( .D(n2605), .CLK(rclk), .R(n10634), .S(1'b1), .Q(
        n11823) );
  DFFSR data_out_reg_6_ ( .D(n2607), .CLK(rclk), .R(n10634), .S(1'b1), .Q(
        n11824) );
  DFFSR data_out_reg_5_ ( .D(n2609), .CLK(rclk), .R(n10634), .S(1'b1), .Q(
        n11825) );
  DFFSR data_out_reg_4_ ( .D(n2611), .CLK(rclk), .R(n10634), .S(1'b1), .Q(
        n11826) );
  DFFSR data_out_reg_3_ ( .D(n2613), .CLK(rclk), .R(n10634), .S(1'b1), .Q(
        n11827) );
  DFFSR data_out_reg_2_ ( .D(n2615), .CLK(rclk), .R(n10634), .S(1'b1), .Q(
        n11828) );
  DFFSR data_out_reg_1_ ( .D(n2617), .CLK(rclk), .R(n10634), .S(1'b1), .Q(
        n11829) );
  DFFSR data_out_reg_0_ ( .D(n2619), .CLK(rclk), .R(n10634), .S(1'b1), .Q(
        n11830) );
  DFFSR rd_ptr_bin_reg_5_ ( .D(n2657), .CLK(rclk), .R(n10634), .S(1'b1), .Q(
        rd_ptr_bin_5_) );
  DFFSR rd_ptr_bin_reg_4_ ( .D(n2536), .CLK(rclk), .R(n10634), .S(1'b1), .Q(
        n14) );
  DFFSR rd_ptr_bin_reg_3_ ( .D(n2541), .CLK(rclk), .R(n10634), .S(1'b1), .Q(
        n13) );
  DFFSR rd_ptr_bin_reg_2_ ( .D(n2546), .CLK(rclk), .R(n10634), .S(1'b1), .Q(
        n12) );
  DFFSR rd_ptr_bin_reg_1_ ( .D(n2551), .CLK(rclk), .R(n10634), .S(1'b1), .Q(
        n11) );
  DFFSR fifo_reg_0__33_ ( .D(n2661), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[1087]) );
  DFFSR fifo_reg_0__32_ ( .D(n2662), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[1086]) );
  DFFSR fifo_reg_0__31_ ( .D(n2663), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[1085]) );
  DFFSR fifo_reg_0__30_ ( .D(n2664), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[1084]) );
  DFFSR fifo_reg_0__29_ ( .D(n2665), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[1083]) );
  DFFSR fifo_reg_0__28_ ( .D(n2666), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[1082]) );
  DFFSR fifo_reg_0__27_ ( .D(n2667), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[1081]) );
  DFFSR fifo_reg_0__26_ ( .D(n2668), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[1080]) );
  DFFSR fifo_reg_0__25_ ( .D(n2669), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[1079]) );
  DFFSR fifo_reg_0__24_ ( .D(n2670), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[1078]) );
  DFFSR fifo_reg_0__23_ ( .D(n2671), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[1077]) );
  DFFSR fifo_reg_0__22_ ( .D(n2672), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[1076]) );
  DFFSR fifo_reg_0__21_ ( .D(n2673), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[1075]) );
  DFFSR fifo_reg_0__20_ ( .D(n2674), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[1074]) );
  DFFSR fifo_reg_0__19_ ( .D(n2675), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[1073]) );
  DFFSR fifo_reg_0__18_ ( .D(n2676), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[1072]) );
  DFFSR fifo_reg_0__17_ ( .D(n2677), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[1071]) );
  DFFSR fifo_reg_0__16_ ( .D(n2678), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[1070]) );
  DFFSR fifo_reg_0__15_ ( .D(n2679), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[1069]) );
  DFFSR fifo_reg_0__14_ ( .D(n2680), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[1068]) );
  DFFSR fifo_reg_0__13_ ( .D(n2681), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[1067]) );
  DFFSR fifo_reg_0__12_ ( .D(n2682), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[1066]) );
  DFFSR fifo_reg_0__11_ ( .D(n2683), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[1065]) );
  DFFSR fifo_reg_0__10_ ( .D(n2684), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[1064]) );
  DFFSR fifo_reg_0__9_ ( .D(n2685), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[1063]) );
  DFFSR fifo_reg_0__8_ ( .D(n2686), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[1062]) );
  DFFSR fifo_reg_0__7_ ( .D(n2687), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[1061]) );
  DFFSR fifo_reg_0__6_ ( .D(n2688), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[1060]) );
  DFFSR fifo_reg_0__5_ ( .D(n2689), .CLK(wclk), .R(n10640), .S(1'b1), .Q(
        fifo[1059]) );
  DFFSR fifo_reg_0__4_ ( .D(n2690), .CLK(wclk), .R(n10640), .S(1'b1), .Q(
        fifo[1058]) );
  DFFSR fifo_reg_0__3_ ( .D(n2691), .CLK(wclk), .R(n10640), .S(1'b1), .Q(
        fifo[1057]) );
  DFFSR fifo_reg_0__2_ ( .D(n2692), .CLK(wclk), .R(n10640), .S(1'b1), .Q(
        fifo[1056]) );
  DFFSR fifo_reg_0__1_ ( .D(n2693), .CLK(wclk), .R(n10640), .S(1'b1), .Q(
        fifo[1055]) );
  DFFSR fifo_reg_0__0_ ( .D(n2694), .CLK(wclk), .R(n10640), .S(1'b1), .Q(
        fifo[1054]) );
  DFFSR fifo_reg_16__33_ ( .D(n3205), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[543]) );
  DFFSR fifo_reg_16__32_ ( .D(n3206), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[542]) );
  DFFSR fifo_reg_16__31_ ( .D(n3207), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[541]) );
  DFFSR fifo_reg_16__30_ ( .D(n3208), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[540]) );
  DFFSR fifo_reg_16__29_ ( .D(n3209), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[539]) );
  DFFSR fifo_reg_16__28_ ( .D(n3210), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[538]) );
  DFFSR fifo_reg_16__27_ ( .D(n3211), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[537]) );
  DFFSR fifo_reg_16__26_ ( .D(n3212), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[536]) );
  DFFSR fifo_reg_16__25_ ( .D(n3213), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[535]) );
  DFFSR fifo_reg_16__24_ ( .D(n3214), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[534]) );
  DFFSR fifo_reg_16__23_ ( .D(n3215), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[533]) );
  DFFSR fifo_reg_16__22_ ( .D(n3216), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[532]) );
  DFFSR fifo_reg_16__21_ ( .D(n3217), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[531]) );
  DFFSR fifo_reg_16__20_ ( .D(n3218), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[530]) );
  DFFSR fifo_reg_16__19_ ( .D(n3219), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[529]) );
  DFFSR fifo_reg_16__18_ ( .D(n3220), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[528]) );
  DFFSR fifo_reg_16__17_ ( .D(n3221), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[527]) );
  DFFSR fifo_reg_16__16_ ( .D(n3222), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[526]) );
  DFFSR fifo_reg_16__15_ ( .D(n3223), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[525]) );
  DFFSR fifo_reg_16__14_ ( .D(n3224), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[524]) );
  DFFSR fifo_reg_16__13_ ( .D(n3225), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[523]) );
  DFFSR fifo_reg_16__12_ ( .D(n3226), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[522]) );
  DFFSR fifo_reg_16__11_ ( .D(n3227), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[521]) );
  DFFSR fifo_reg_16__10_ ( .D(n3228), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[520]) );
  DFFSR fifo_reg_16__9_ ( .D(n3229), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[519]) );
  DFFSR fifo_reg_16__8_ ( .D(n3230), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[518]) );
  DFFSR fifo_reg_16__7_ ( .D(n3231), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[517]) );
  DFFSR fifo_reg_16__6_ ( .D(n3232), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[516]) );
  DFFSR fifo_reg_16__5_ ( .D(n3233), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[515]) );
  DFFSR fifo_reg_16__4_ ( .D(n3234), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[514]) );
  DFFSR fifo_reg_16__3_ ( .D(n3235), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[513]) );
  DFFSR fifo_reg_16__2_ ( .D(n3236), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[512]) );
  DFFSR fifo_reg_16__1_ ( .D(n3237), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[511]) );
  DFFSR fifo_reg_16__0_ ( .D(n3238), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[510]) );
  DFFSR fifo_reg_17__33_ ( .D(n3239), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[509]) );
  DFFSR fifo_reg_17__32_ ( .D(n3240), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[508]) );
  DFFSR fifo_reg_17__31_ ( .D(n3241), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[507]) );
  DFFSR fifo_reg_17__30_ ( .D(n3242), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[506]) );
  DFFSR fifo_reg_17__29_ ( .D(n3243), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[505]) );
  DFFSR fifo_reg_17__28_ ( .D(n3244), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[504]) );
  DFFSR fifo_reg_17__27_ ( .D(n3245), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[503]) );
  DFFSR fifo_reg_17__26_ ( .D(n3246), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[502]) );
  DFFSR fifo_reg_17__25_ ( .D(n3247), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[501]) );
  DFFSR fifo_reg_17__24_ ( .D(n3248), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[500]) );
  DFFSR fifo_reg_17__23_ ( .D(n3249), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[499]) );
  DFFSR fifo_reg_17__22_ ( .D(n3250), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[498]) );
  DFFSR fifo_reg_17__21_ ( .D(n3251), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[497]) );
  DFFSR fifo_reg_17__20_ ( .D(n3252), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[496]) );
  DFFSR fifo_reg_17__19_ ( .D(n3253), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[495]) );
  DFFSR fifo_reg_17__18_ ( .D(n3254), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[494]) );
  DFFSR fifo_reg_17__17_ ( .D(n3255), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[493]) );
  DFFSR fifo_reg_17__16_ ( .D(n3256), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[492]) );
  DFFSR fifo_reg_17__15_ ( .D(n3257), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[491]) );
  DFFSR fifo_reg_17__14_ ( .D(n3258), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[490]) );
  DFFSR fifo_reg_17__13_ ( .D(n3259), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[489]) );
  DFFSR fifo_reg_17__12_ ( .D(n3260), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[488]) );
  DFFSR fifo_reg_17__11_ ( .D(n3261), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[487]) );
  DFFSR fifo_reg_17__10_ ( .D(n3262), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[486]) );
  DFFSR fifo_reg_17__9_ ( .D(n3263), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[485]) );
  DFFSR fifo_reg_17__8_ ( .D(n3264), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[484]) );
  DFFSR fifo_reg_17__7_ ( .D(n3265), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[483]) );
  DFFSR fifo_reg_17__6_ ( .D(n3266), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[482]) );
  DFFSR fifo_reg_17__5_ ( .D(n3267), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[481]) );
  DFFSR fifo_reg_17__4_ ( .D(n3268), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[480]) );
  DFFSR fifo_reg_17__3_ ( .D(n3269), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[479]) );
  DFFSR fifo_reg_17__2_ ( .D(n3270), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[478]) );
  DFFSR fifo_reg_17__1_ ( .D(n3271), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[477]) );
  DFFSR fifo_reg_17__0_ ( .D(n3272), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[476]) );
  DFFSR fifo_reg_22__33_ ( .D(n3409), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[339]) );
  DFFSR fifo_reg_22__32_ ( .D(n3410), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[338]) );
  DFFSR fifo_reg_22__31_ ( .D(n3411), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[337]) );
  DFFSR fifo_reg_22__30_ ( .D(n3412), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[336]) );
  DFFSR fifo_reg_22__29_ ( .D(n3413), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[335]) );
  DFFSR fifo_reg_22__28_ ( .D(n3414), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[334]) );
  DFFSR fifo_reg_22__27_ ( .D(n3415), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[333]) );
  DFFSR fifo_reg_22__26_ ( .D(n3416), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[332]) );
  DFFSR fifo_reg_22__25_ ( .D(n3417), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[331]) );
  DFFSR fifo_reg_22__24_ ( .D(n3418), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[330]) );
  DFFSR fifo_reg_22__23_ ( .D(n3419), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[329]) );
  DFFSR fifo_reg_22__22_ ( .D(n3420), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[328]) );
  DFFSR fifo_reg_22__21_ ( .D(n3421), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[327]) );
  DFFSR fifo_reg_22__20_ ( .D(n3422), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[326]) );
  DFFSR fifo_reg_22__19_ ( .D(n3423), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[325]) );
  DFFSR fifo_reg_22__18_ ( .D(n3424), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[324]) );
  DFFSR fifo_reg_22__17_ ( .D(n3425), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[323]) );
  DFFSR fifo_reg_22__16_ ( .D(n3426), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[322]) );
  DFFSR fifo_reg_22__15_ ( .D(n3427), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[321]) );
  DFFSR fifo_reg_22__14_ ( .D(n3428), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[320]) );
  DFFSR fifo_reg_22__13_ ( .D(n3429), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[319]) );
  DFFSR fifo_reg_22__12_ ( .D(n3430), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[318]) );
  DFFSR fifo_reg_22__11_ ( .D(n3431), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[317]) );
  DFFSR fifo_reg_22__10_ ( .D(n3432), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[316]) );
  DFFSR fifo_reg_22__9_ ( .D(n3433), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[315]) );
  DFFSR fifo_reg_22__8_ ( .D(n3434), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[314]) );
  DFFSR fifo_reg_22__7_ ( .D(n3435), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[313]) );
  DFFSR fifo_reg_22__6_ ( .D(n3436), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[312]) );
  DFFSR fifo_reg_22__5_ ( .D(n3437), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[311]) );
  DFFSR fifo_reg_22__4_ ( .D(n3438), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[310]) );
  DFFSR fifo_reg_22__3_ ( .D(n3439), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[309]) );
  DFFSR fifo_reg_22__2_ ( .D(n3440), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[308]) );
  DFFSR fifo_reg_22__1_ ( .D(n3441), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[307]) );
  DFFSR fifo_reg_22__0_ ( .D(n3442), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[306]) );
  DFFSR fifo_reg_23__33_ ( .D(n3443), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[305]) );
  DFFSR fifo_reg_23__32_ ( .D(n3444), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[304]) );
  DFFSR fifo_reg_23__31_ ( .D(n3445), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[303]) );
  DFFSR fifo_reg_23__30_ ( .D(n3446), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[302]) );
  DFFSR fifo_reg_23__29_ ( .D(n3447), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[301]) );
  DFFSR fifo_reg_23__28_ ( .D(n3448), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[300]) );
  DFFSR fifo_reg_23__27_ ( .D(n3449), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[299]) );
  DFFSR fifo_reg_23__26_ ( .D(n3450), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[298]) );
  DFFSR fifo_reg_23__25_ ( .D(n3451), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[297]) );
  DFFSR fifo_reg_23__24_ ( .D(n3452), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[296]) );
  DFFSR fifo_reg_23__23_ ( .D(n3453), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[295]) );
  DFFSR fifo_reg_23__22_ ( .D(n3454), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[294]) );
  DFFSR fifo_reg_23__21_ ( .D(n3455), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[293]) );
  DFFSR fifo_reg_23__20_ ( .D(n3456), .CLK(wclk), .R(n10639), .S(1'b1), .Q(
        fifo[292]) );
  DFFSR fifo_reg_23__19_ ( .D(n3457), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[291]) );
  DFFSR fifo_reg_23__18_ ( .D(n3458), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[290]) );
  DFFSR fifo_reg_23__17_ ( .D(n3459), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[289]) );
  DFFSR fifo_reg_23__16_ ( .D(n3460), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[288]) );
  DFFSR fifo_reg_23__15_ ( .D(n3461), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[287]) );
  DFFSR fifo_reg_23__14_ ( .D(n3462), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[286]) );
  DFFSR fifo_reg_23__13_ ( .D(n3463), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[285]) );
  DFFSR fifo_reg_23__12_ ( .D(n3464), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[284]) );
  DFFSR fifo_reg_23__11_ ( .D(n3465), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[283]) );
  DFFSR fifo_reg_23__10_ ( .D(n3466), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[282]) );
  DFFSR fifo_reg_23__9_ ( .D(n3467), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[281]) );
  DFFSR fifo_reg_23__8_ ( .D(n3468), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[280]) );
  DFFSR fifo_reg_23__7_ ( .D(n3469), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[279]) );
  DFFSR fifo_reg_23__6_ ( .D(n3470), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[278]) );
  DFFSR fifo_reg_23__5_ ( .D(n3471), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[277]) );
  DFFSR fifo_reg_23__4_ ( .D(n3472), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[276]) );
  DFFSR fifo_reg_23__3_ ( .D(n3473), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[275]) );
  DFFSR fifo_reg_23__2_ ( .D(n3474), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[274]) );
  DFFSR fifo_reg_23__1_ ( .D(n3475), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[273]) );
  DFFSR fifo_reg_23__0_ ( .D(n3476), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[272]) );
  DFFSR fifo_reg_18__33_ ( .D(n3273), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[475]) );
  DFFSR fifo_reg_18__32_ ( .D(n3274), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[474]) );
  DFFSR fifo_reg_18__31_ ( .D(n3275), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[473]) );
  DFFSR fifo_reg_18__30_ ( .D(n3276), .CLK(wclk), .R(n10637), .S(1'b1), .Q(
        fifo[472]) );
  DFFSR fifo_reg_18__29_ ( .D(n3277), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[471]) );
  DFFSR fifo_reg_18__28_ ( .D(n3278), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[470]) );
  DFFSR fifo_reg_18__27_ ( .D(n3279), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[469]) );
  DFFSR fifo_reg_18__26_ ( .D(n3280), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[468]) );
  DFFSR fifo_reg_18__25_ ( .D(n3281), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[467]) );
  DFFSR fifo_reg_18__24_ ( .D(n3282), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[466]) );
  DFFSR fifo_reg_18__23_ ( .D(n3283), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[465]) );
  DFFSR fifo_reg_18__22_ ( .D(n3284), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[464]) );
  DFFSR fifo_reg_18__21_ ( .D(n3285), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[463]) );
  DFFSR fifo_reg_18__20_ ( .D(n3286), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[462]) );
  DFFSR fifo_reg_18__19_ ( .D(n3287), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[461]) );
  DFFSR fifo_reg_18__18_ ( .D(n3288), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[460]) );
  DFFSR fifo_reg_18__17_ ( .D(n3289), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[459]) );
  DFFSR fifo_reg_18__16_ ( .D(n3290), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[458]) );
  DFFSR fifo_reg_18__15_ ( .D(n3291), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[457]) );
  DFFSR fifo_reg_18__14_ ( .D(n3292), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[456]) );
  DFFSR fifo_reg_18__13_ ( .D(n3293), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[455]) );
  DFFSR fifo_reg_18__12_ ( .D(n3294), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[454]) );
  DFFSR fifo_reg_18__11_ ( .D(n3295), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[453]) );
  DFFSR fifo_reg_18__10_ ( .D(n3296), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[452]) );
  DFFSR fifo_reg_18__9_ ( .D(n3297), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[451]) );
  DFFSR fifo_reg_18__8_ ( .D(n3298), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[450]) );
  DFFSR fifo_reg_18__7_ ( .D(n3299), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[449]) );
  DFFSR fifo_reg_18__6_ ( .D(n3300), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[448]) );
  DFFSR fifo_reg_18__5_ ( .D(n3301), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[447]) );
  DFFSR fifo_reg_18__4_ ( .D(n3302), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[446]) );
  DFFSR fifo_reg_18__3_ ( .D(n3303), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[445]) );
  DFFSR fifo_reg_18__2_ ( .D(n3304), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[444]) );
  DFFSR fifo_reg_18__1_ ( .D(n3305), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[443]) );
  DFFSR fifo_reg_18__0_ ( .D(n3306), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[442]) );
  DFFSR fifo_reg_20__33_ ( .D(n3341), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[407]) );
  DFFSR fifo_reg_20__32_ ( .D(n3342), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[406]) );
  DFFSR fifo_reg_20__31_ ( .D(n3343), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[405]) );
  DFFSR fifo_reg_20__30_ ( .D(n3344), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[404]) );
  DFFSR fifo_reg_20__29_ ( .D(n3345), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[403]) );
  DFFSR fifo_reg_20__28_ ( .D(n3346), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[402]) );
  DFFSR fifo_reg_20__27_ ( .D(n3347), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[401]) );
  DFFSR fifo_reg_20__26_ ( .D(n3348), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[400]) );
  DFFSR fifo_reg_20__25_ ( .D(n3349), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[399]) );
  DFFSR fifo_reg_20__24_ ( .D(n3350), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[398]) );
  DFFSR fifo_reg_20__23_ ( .D(n3351), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[397]) );
  DFFSR fifo_reg_20__22_ ( .D(n3352), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[396]) );
  DFFSR fifo_reg_20__21_ ( .D(n3353), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[395]) );
  DFFSR fifo_reg_20__20_ ( .D(n3354), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[394]) );
  DFFSR fifo_reg_20__19_ ( .D(n3355), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[393]) );
  DFFSR fifo_reg_20__18_ ( .D(n3356), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[392]) );
  DFFSR fifo_reg_20__17_ ( .D(n3357), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[391]) );
  DFFSR fifo_reg_20__16_ ( .D(n3358), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[390]) );
  DFFSR fifo_reg_20__15_ ( .D(n3359), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[389]) );
  DFFSR fifo_reg_20__14_ ( .D(n3360), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[388]) );
  DFFSR fifo_reg_20__13_ ( .D(n3361), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[387]) );
  DFFSR fifo_reg_20__12_ ( .D(n3362), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[386]) );
  DFFSR fifo_reg_20__11_ ( .D(n3363), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[385]) );
  DFFSR fifo_reg_20__10_ ( .D(n3364), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[384]) );
  DFFSR fifo_reg_20__9_ ( .D(n3365), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[383]) );
  DFFSR fifo_reg_20__8_ ( .D(n3366), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[382]) );
  DFFSR fifo_reg_20__7_ ( .D(n3367), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[381]) );
  DFFSR fifo_reg_20__6_ ( .D(n3368), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[380]) );
  DFFSR fifo_reg_20__5_ ( .D(n3369), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[379]) );
  DFFSR fifo_reg_20__4_ ( .D(n3370), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[378]) );
  DFFSR fifo_reg_20__3_ ( .D(n3371), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[377]) );
  DFFSR fifo_reg_20__2_ ( .D(n3372), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[376]) );
  DFFSR fifo_reg_20__1_ ( .D(n3373), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[375]) );
  DFFSR fifo_reg_20__0_ ( .D(n3374), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[374]) );
  DFFSR fifo_reg_21__33_ ( .D(n3375), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[373]) );
  DFFSR fifo_reg_21__32_ ( .D(n3376), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[372]) );
  DFFSR fifo_reg_21__31_ ( .D(n3377), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[371]) );
  DFFSR fifo_reg_21__30_ ( .D(n3378), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[370]) );
  DFFSR fifo_reg_21__29_ ( .D(n3379), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[369]) );
  DFFSR fifo_reg_21__28_ ( .D(n3380), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[368]) );
  DFFSR fifo_reg_21__27_ ( .D(n3381), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[367]) );
  DFFSR fifo_reg_21__26_ ( .D(n3382), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[366]) );
  DFFSR fifo_reg_21__25_ ( .D(n3383), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[365]) );
  DFFSR fifo_reg_21__24_ ( .D(n3384), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[364]) );
  DFFSR fifo_reg_21__23_ ( .D(n3385), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[363]) );
  DFFSR fifo_reg_21__22_ ( .D(n3386), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[362]) );
  DFFSR fifo_reg_21__21_ ( .D(n3387), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[361]) );
  DFFSR fifo_reg_21__20_ ( .D(n3388), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[360]) );
  DFFSR fifo_reg_21__19_ ( .D(n3389), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[359]) );
  DFFSR fifo_reg_21__18_ ( .D(n3390), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[358]) );
  DFFSR fifo_reg_21__17_ ( .D(n3391), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[357]) );
  DFFSR fifo_reg_21__16_ ( .D(n3392), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[356]) );
  DFFSR fifo_reg_21__15_ ( .D(n3393), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[355]) );
  DFFSR fifo_reg_21__14_ ( .D(n3394), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[354]) );
  DFFSR fifo_reg_21__13_ ( .D(n3395), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[353]) );
  DFFSR fifo_reg_21__12_ ( .D(n3396), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[352]) );
  DFFSR fifo_reg_21__11_ ( .D(n3397), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[351]) );
  DFFSR fifo_reg_21__10_ ( .D(n3398), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[350]) );
  DFFSR fifo_reg_21__9_ ( .D(n3399), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[349]) );
  DFFSR fifo_reg_21__8_ ( .D(n3400), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[348]) );
  DFFSR fifo_reg_21__7_ ( .D(n3401), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[347]) );
  DFFSR fifo_reg_21__6_ ( .D(n3402), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[346]) );
  DFFSR fifo_reg_21__5_ ( .D(n3403), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[345]) );
  DFFSR fifo_reg_21__4_ ( .D(n3404), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[344]) );
  DFFSR fifo_reg_21__3_ ( .D(n3405), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[343]) );
  DFFSR fifo_reg_21__2_ ( .D(n3406), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[342]) );
  DFFSR fifo_reg_21__1_ ( .D(n3407), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[341]) );
  DFFSR fifo_reg_21__0_ ( .D(n3408), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[340]) );
  DFFSR fifo_reg_19__33_ ( .D(n3307), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[441]) );
  DFFSR fifo_reg_19__32_ ( .D(n3308), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[440]) );
  DFFSR fifo_reg_19__31_ ( .D(n3309), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[439]) );
  DFFSR fifo_reg_19__30_ ( .D(n3310), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[438]) );
  DFFSR fifo_reg_19__29_ ( .D(n3311), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[437]) );
  DFFSR fifo_reg_19__28_ ( .D(n3312), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[436]) );
  DFFSR fifo_reg_19__27_ ( .D(n3313), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[435]) );
  DFFSR fifo_reg_19__26_ ( .D(n3314), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[434]) );
  DFFSR fifo_reg_19__25_ ( .D(n3315), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[433]) );
  DFFSR fifo_reg_19__24_ ( .D(n3316), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[432]) );
  DFFSR fifo_reg_19__23_ ( .D(n3317), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[431]) );
  DFFSR fifo_reg_19__22_ ( .D(n3318), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[430]) );
  DFFSR fifo_reg_19__21_ ( .D(n3319), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[429]) );
  DFFSR fifo_reg_19__20_ ( .D(n3320), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[428]) );
  DFFSR fifo_reg_19__19_ ( .D(n3321), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[427]) );
  DFFSR fifo_reg_19__18_ ( .D(n3322), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[426]) );
  DFFSR fifo_reg_19__17_ ( .D(n3323), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[425]) );
  DFFSR fifo_reg_19__16_ ( .D(n3324), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[424]) );
  DFFSR fifo_reg_19__15_ ( .D(n3325), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[423]) );
  DFFSR fifo_reg_19__14_ ( .D(n3326), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[422]) );
  DFFSR fifo_reg_19__13_ ( .D(n3327), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[421]) );
  DFFSR fifo_reg_19__12_ ( .D(n3328), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[420]) );
  DFFSR fifo_reg_19__11_ ( .D(n3329), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[419]) );
  DFFSR fifo_reg_19__10_ ( .D(n3330), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[418]) );
  DFFSR fifo_reg_19__9_ ( .D(n3331), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[417]) );
  DFFSR fifo_reg_19__8_ ( .D(n3332), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[416]) );
  DFFSR fifo_reg_19__7_ ( .D(n3333), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[415]) );
  DFFSR fifo_reg_19__6_ ( .D(n3334), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[414]) );
  DFFSR fifo_reg_19__5_ ( .D(n3335), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[413]) );
  DFFSR fifo_reg_19__4_ ( .D(n3336), .CLK(wclk), .R(n10638), .S(1'b1), .Q(
        fifo[412]) );
  DFFSR fifo_reg_19__3_ ( .D(n3337), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[411]) );
  DFFSR fifo_reg_19__2_ ( .D(n3338), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[410]) );
  DFFSR fifo_reg_19__1_ ( .D(n3339), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[409]) );
  DFFSR fifo_reg_19__0_ ( .D(n3340), .CLK(wclk), .R(n2658), .S(1'b1), .Q(
        fifo[408]) );
  DFFSR rd_ptr_bin_reg_0_ ( .D(n2660), .CLK(rclk), .R(n10634), .S(1'b1), .Q(
        n10) );
  DFFSR wr_ptr_gray_ss_reg_4_ ( .D(n65), .CLK(rclk), .R(n10634), .S(1'b1), .Q(
        wr_ptr_gray_ss[4]) );
  DFFSR wr_ptr_gray_ss_reg_5_ ( .D(n134), .CLK(rclk), .R(n10644), .S(1'b1), 
        .Q(wr_ptr_gray_ss[5]) );
  INVX1 U4 ( .A(r301_carry[4]), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
  XNOR2X1 U6 ( .A(n27), .B(n9965), .Y(rd_ptr_bin_ss[4]) );
  BUFX2 U7 ( .A(rd_ptr_bin_ss[1]), .Y(n3) );
  BUFX2 U8 ( .A(n9966), .Y(n4) );
  AND2X2 U10 ( .A(n10104), .B(r301_carry[4]), .Y(n10522) );
  BUFX2 U11 ( .A(rd_ptr_bin_ss[3]), .Y(n5) );
  BUFX2 U13 ( .A(rd_ptr_bin_ss[4]), .Y(n6) );
  INVX2 U14 ( .A(n10740), .Y(n10739) );
  INVX4 U16 ( .A(n10741), .Y(n10740) );
  INVX1 U18 ( .A(n1437), .Y(n1435) );
  OR2X2 U88 ( .A(n31), .B(n30), .Y(n28) );
  OR2X2 U90 ( .A(n10522), .B(n29), .Y(n31) );
  AND2X2 U92 ( .A(r301_B_not_4_), .B(r301_carry[4]), .Y(n10521) );
  INVX1 U94 ( .A(n10521), .Y(n7) );
  BUFX2 U96 ( .A(n1428), .Y(n8) );
  BUFX2 U98 ( .A(n11796), .Y(empty_bar) );
  BUFX2 U101 ( .A(wr_ptr_gray_ss[4]), .Y(n25) );
  BUFX2 U102 ( .A(wr_ptr_gray_ss[0]), .Y(n26) );
  BUFX2 U104 ( .A(rd_ptr_gray_ss[4]), .Y(n27) );
  INVX1 U106 ( .A(n6687), .Y(n29) );
  INVX1 U108 ( .A(n7), .Y(n30) );
  AND2X2 U110 ( .A(n33), .B(rd_ptr_bin_ss[0]), .Y(n10485) );
  INVX1 U112 ( .A(n10485), .Y(n32) );
  INVX1 U114 ( .A(n10686), .Y(n10683) );
  INVX1 U116 ( .A(n10532), .Y(n196) );
  INVX2 U118 ( .A(n1434), .Y(n10534) );
  AND2X1 U120 ( .A(n1177), .B(n10022), .Y(n10502) );
  AND2X1 U122 ( .A(n1177), .B(n10019), .Y(n10501) );
  AND2X1 U124 ( .A(n1177), .B(n360), .Y(n10494) );
  AND2X1 U126 ( .A(n613), .B(n10019), .Y(n10513) );
  AND2X1 U128 ( .A(n613), .B(n10025), .Y(n10512) );
  AND2X1 U130 ( .A(n613), .B(n576), .Y(n10509) );
  BUFX2 U132 ( .A(full_bar), .Y(n39) );
  INVX1 U134 ( .A(n42), .Y(n40) );
  INVX1 U136 ( .A(n40), .Y(n41) );
  BUFX2 U138 ( .A(rd_ptr_gray_s[3]), .Y(n42) );
  INVX1 U140 ( .A(n45), .Y(n43) );
  INVX1 U142 ( .A(n43), .Y(n44) );
  BUFX2 U144 ( .A(rd_ptr_gray[3]), .Y(n45) );
  INVX1 U146 ( .A(n48), .Y(n46) );
  INVX1 U148 ( .A(n46), .Y(n47) );
  BUFX2 U150 ( .A(rd_ptr_gray_s[2]), .Y(n48) );
  INVX1 U152 ( .A(n51), .Y(n49) );
  INVX1 U154 ( .A(n49), .Y(n50) );
  BUFX2 U156 ( .A(rd_ptr_gray[2]), .Y(n51) );
  INVX1 U158 ( .A(n54), .Y(n52) );
  INVX1 U160 ( .A(n52), .Y(n53) );
  BUFX2 U162 ( .A(rd_ptr_gray_s[1]), .Y(n54) );
  INVX1 U164 ( .A(n57), .Y(n55) );
  INVX1 U166 ( .A(n55), .Y(n56) );
  BUFX2 U168 ( .A(rd_ptr_gray[1]), .Y(n57) );
  INVX1 U170 ( .A(n60), .Y(n58) );
  INVX1 U172 ( .A(n58), .Y(n59) );
  BUFX2 U174 ( .A(rd_ptr_gray_s[0]), .Y(n60) );
  INVX1 U175 ( .A(n63), .Y(n61) );
  INVX1 U177 ( .A(n61), .Y(n62) );
  BUFX2 U179 ( .A(rd_ptr_gray[0]), .Y(n63) );
  INVX1 U181 ( .A(n66), .Y(n64) );
  INVX1 U183 ( .A(n64), .Y(n65) );
  BUFX2 U185 ( .A(wr_ptr_gray_s[4]), .Y(n66) );
  INVX1 U187 ( .A(n69), .Y(n67) );
  INVX1 U189 ( .A(n67), .Y(n68) );
  BUFX2 U191 ( .A(wr_ptr_gray[4]), .Y(n69) );
  INVX1 U193 ( .A(n111), .Y(n70) );
  INVX1 U195 ( .A(n70), .Y(n105) );
  BUFX2 U197 ( .A(wr_ptr_gray_s[3]), .Y(n111) );
  INVX1 U199 ( .A(n114), .Y(n112) );
  INVX1 U201 ( .A(n112), .Y(n113) );
  BUFX2 U203 ( .A(wr_ptr_gray[3]), .Y(n114) );
  INVX1 U205 ( .A(n117), .Y(n115) );
  INVX1 U207 ( .A(n115), .Y(n116) );
  BUFX2 U209 ( .A(wr_ptr_gray_s[2]), .Y(n117) );
  INVX1 U211 ( .A(n120), .Y(n118) );
  INVX1 U213 ( .A(n118), .Y(n119) );
  BUFX2 U215 ( .A(wr_ptr_gray[2]), .Y(n120) );
  INVX1 U217 ( .A(n123), .Y(n121) );
  INVX1 U219 ( .A(n121), .Y(n122) );
  BUFX2 U221 ( .A(wr_ptr_gray_s[1]), .Y(n123) );
  INVX1 U223 ( .A(n126), .Y(n124) );
  INVX1 U225 ( .A(n124), .Y(n125) );
  BUFX2 U227 ( .A(wr_ptr_gray[1]), .Y(n126) );
  INVX1 U229 ( .A(n129), .Y(n127) );
  INVX1 U231 ( .A(n127), .Y(n128) );
  BUFX2 U233 ( .A(wr_ptr_gray_s[0]), .Y(n129) );
  INVX1 U235 ( .A(n132), .Y(n130) );
  INVX1 U237 ( .A(n130), .Y(n131) );
  BUFX2 U239 ( .A(wr_ptr_gray[0]), .Y(n132) );
  INVX1 U241 ( .A(n135), .Y(n133) );
  INVX1 U243 ( .A(n133), .Y(n134) );
  BUFX2 U244 ( .A(wr_ptr_gray_s[5]), .Y(n135) );
  INVX1 U246 ( .A(n138), .Y(n136) );
  INVX1 U248 ( .A(n136), .Y(n137) );
  BUFX2 U250 ( .A(wr_ptr_gray[5]), .Y(n138) );
  INVX1 U252 ( .A(n141), .Y(n139) );
  INVX1 U254 ( .A(n139), .Y(n140) );
  BUFX2 U256 ( .A(rd_ptr_gray_s[4]), .Y(n141) );
  INVX1 U258 ( .A(n144), .Y(n142) );
  INVX1 U260 ( .A(n142), .Y(n143) );
  BUFX2 U262 ( .A(rd_ptr_gray[4]), .Y(n144) );
  INVX1 U264 ( .A(n147), .Y(n145) );
  INVX1 U266 ( .A(n145), .Y(n146) );
  BUFX2 U268 ( .A(rd_ptr_gray_s[5]), .Y(n147) );
  INVX1 U270 ( .A(n150), .Y(n148) );
  INVX1 U272 ( .A(n148), .Y(n149) );
  BUFX2 U274 ( .A(rd_ptr_gray[5]), .Y(n150) );
  INVX1 U276 ( .A(n1436), .Y(n151) );
  INVX1 U278 ( .A(n151), .Y(n152) );
  INVX1 U280 ( .A(n155), .Y(n153) );
  INVX1 U282 ( .A(n153), .Y(data_out[26]) );
  BUFX2 U284 ( .A(n11804), .Y(n155) );
  INVX1 U286 ( .A(n158), .Y(n156) );
  INVX1 U288 ( .A(n156), .Y(data_out[27]) );
  BUFX2 U290 ( .A(n11803), .Y(n158) );
  INVX1 U292 ( .A(n161), .Y(n159) );
  INVX1 U294 ( .A(n159), .Y(data_out[28]) );
  BUFX2 U296 ( .A(n11802), .Y(n161) );
  BUFX2 U298 ( .A(empty_bar), .Y(n162) );
  AND2X1 U300 ( .A(n10104), .B(n240), .Y(n10518) );
  INVX1 U302 ( .A(n10518), .Y(n163) );
  AND2X1 U304 ( .A(n1177), .B(n576), .Y(n1390) );
  INVX1 U306 ( .A(n1390), .Y(n164) );
  AND2X1 U308 ( .A(n1177), .B(n540), .Y(n1355) );
  INVX1 U310 ( .A(n1355), .Y(n165) );
  AND2X1 U312 ( .A(n1177), .B(n10031), .Y(n1320) );
  INVX1 U313 ( .A(n1320), .Y(n166) );
  AND2X1 U315 ( .A(n1177), .B(n10025), .Y(n1213) );
  INVX1 U317 ( .A(n1213), .Y(n167) );
  INVX1 U319 ( .A(n1425), .Y(n1177) );
  AND2X1 U321 ( .A(n613), .B(n540), .Y(n789) );
  INVX1 U323 ( .A(n789), .Y(n168) );
  AND2X1 U325 ( .A(n613), .B(n10031), .Y(n754) );
  INVX1 U327 ( .A(n754), .Y(n169) );
  AND2X1 U329 ( .A(n613), .B(n10022), .Y(n684) );
  INVX1 U331 ( .A(n684), .Y(n170) );
  AND2X1 U333 ( .A(n613), .B(n360), .Y(n614) );
  INVX1 U335 ( .A(n614), .Y(n171) );
  AND2X1 U337 ( .A(n613), .B(n323), .Y(n578) );
  INVX1 U339 ( .A(n578), .Y(n172) );
  INVX1 U341 ( .A(n859), .Y(n613) );
  INVX1 U343 ( .A(n175), .Y(n173) );
  INVX1 U345 ( .A(n173), .Y(n174) );
  AND2X1 U347 ( .A(n10001), .B(n9998), .Y(n23) );
  INVX1 U349 ( .A(n23), .Y(n175) );
  INVX1 U351 ( .A(n178), .Y(n176) );
  INVX1 U353 ( .A(n176), .Y(n177) );
  AND2X1 U355 ( .A(n8742), .B(n10498), .Y(n1424) );
  INVX1 U357 ( .A(n1424), .Y(n178) );
  INVX1 U359 ( .A(n181), .Y(n179) );
  INVX1 U361 ( .A(n179), .Y(n180) );
  AND2X1 U363 ( .A(n8745), .B(n10498), .Y(n1423) );
  INVX1 U365 ( .A(n1423), .Y(n181) );
  INVX1 U367 ( .A(n184), .Y(n182) );
  INVX1 U369 ( .A(n182), .Y(n183) );
  AND2X1 U371 ( .A(n8748), .B(n10498), .Y(n1422) );
  INVX1 U373 ( .A(n1422), .Y(n184) );
  INVX1 U375 ( .A(n187), .Y(n185) );
  INVX1 U377 ( .A(n185), .Y(n186) );
  AND2X1 U379 ( .A(n8751), .B(n10498), .Y(n1421) );
  INVX1 U381 ( .A(n1421), .Y(n187) );
  INVX1 U382 ( .A(n190), .Y(n188) );
  INVX1 U384 ( .A(n188), .Y(n189) );
  AND2X1 U386 ( .A(n8754), .B(n10498), .Y(n1420) );
  INVX1 U388 ( .A(n1420), .Y(n190) );
  INVX1 U390 ( .A(n198), .Y(n191) );
  INVX1 U392 ( .A(n191), .Y(n192) );
  AND2X1 U394 ( .A(n8757), .B(n10498), .Y(n1419) );
  INVX1 U396 ( .A(n1419), .Y(n198) );
  INVX1 U398 ( .A(n1141), .Y(n200) );
  INVX1 U400 ( .A(n200), .Y(n252) );
  AND2X1 U402 ( .A(n8760), .B(n10498), .Y(n1418) );
  INVX1 U404 ( .A(n1418), .Y(n1141) );
  INVX1 U406 ( .A(n1716), .Y(n1431) );
  INVX1 U408 ( .A(n1431), .Y(n1432) );
  AND2X1 U410 ( .A(n8763), .B(n10498), .Y(n1417) );
  INVX1 U412 ( .A(n1417), .Y(n1716) );
  INVX1 U414 ( .A(n1719), .Y(n1717) );
  INVX1 U416 ( .A(n1717), .Y(n1718) );
  AND2X1 U418 ( .A(n8766), .B(n10498), .Y(n1416) );
  INVX1 U420 ( .A(n1416), .Y(n1719) );
  INVX1 U422 ( .A(n1722), .Y(n1720) );
  INVX1 U424 ( .A(n1720), .Y(n1721) );
  AND2X1 U426 ( .A(n8769), .B(n10498), .Y(n1415) );
  INVX1 U428 ( .A(n1415), .Y(n1722) );
  INVX1 U430 ( .A(n1725), .Y(n1723) );
  INVX1 U432 ( .A(n1723), .Y(n1724) );
  AND2X1 U434 ( .A(n8772), .B(n10498), .Y(n1414) );
  INVX1 U436 ( .A(n1414), .Y(n1725) );
  INVX1 U438 ( .A(n1728), .Y(n1726) );
  INVX1 U440 ( .A(n1726), .Y(n1727) );
  AND2X1 U442 ( .A(n8775), .B(n10498), .Y(n1413) );
  INVX1 U444 ( .A(n1413), .Y(n1728) );
  INVX1 U446 ( .A(n1731), .Y(n1729) );
  INVX1 U448 ( .A(n1729), .Y(n1730) );
  AND2X1 U450 ( .A(n8778), .B(n10498), .Y(n1412) );
  INVX1 U451 ( .A(n1412), .Y(n1731) );
  INVX1 U453 ( .A(n1734), .Y(n1732) );
  INVX1 U455 ( .A(n1732), .Y(n1733) );
  AND2X1 U457 ( .A(n8781), .B(n10498), .Y(n1411) );
  INVX1 U459 ( .A(n1411), .Y(n1734) );
  INVX1 U461 ( .A(n1737), .Y(n1735) );
  INVX1 U463 ( .A(n1735), .Y(n1736) );
  AND2X1 U465 ( .A(n8784), .B(n10498), .Y(n1410) );
  INVX1 U467 ( .A(n1410), .Y(n1737) );
  INVX1 U469 ( .A(n1740), .Y(n1738) );
  INVX1 U471 ( .A(n1738), .Y(n1739) );
  AND2X1 U473 ( .A(n8787), .B(n10498), .Y(n1409) );
  INVX1 U475 ( .A(n1409), .Y(n1740) );
  INVX1 U477 ( .A(n1743), .Y(n1741) );
  INVX1 U479 ( .A(n1741), .Y(n1742) );
  AND2X1 U481 ( .A(n8790), .B(n10498), .Y(n1408) );
  INVX1 U483 ( .A(n1408), .Y(n1743) );
  INVX1 U485 ( .A(n1746), .Y(n1744) );
  INVX1 U487 ( .A(n1744), .Y(n1745) );
  AND2X1 U489 ( .A(n8793), .B(n10498), .Y(n1407) );
  INVX1 U491 ( .A(n1407), .Y(n1746) );
  INVX1 U493 ( .A(n1749), .Y(n1747) );
  INVX1 U495 ( .A(n1747), .Y(n1748) );
  AND2X1 U497 ( .A(n8796), .B(n10498), .Y(n1406) );
  INVX1 U499 ( .A(n1406), .Y(n1749) );
  INVX1 U501 ( .A(n1752), .Y(n1750) );
  INVX1 U503 ( .A(n1750), .Y(n1751) );
  AND2X1 U505 ( .A(n8799), .B(n10498), .Y(n1405) );
  INVX1 U507 ( .A(n1405), .Y(n1752) );
  INVX1 U509 ( .A(n1755), .Y(n1753) );
  INVX1 U511 ( .A(n1753), .Y(n1754) );
  AND2X1 U513 ( .A(n8802), .B(n10498), .Y(n1404) );
  INVX1 U515 ( .A(n1404), .Y(n1755) );
  INVX1 U517 ( .A(n1758), .Y(n1756) );
  INVX1 U519 ( .A(n1756), .Y(n1757) );
  AND2X1 U520 ( .A(n8805), .B(n10498), .Y(n1403) );
  INVX1 U522 ( .A(n1403), .Y(n1758) );
  INVX1 U524 ( .A(n1761), .Y(n1759) );
  INVX1 U526 ( .A(n1759), .Y(n1760) );
  AND2X1 U528 ( .A(n8808), .B(n10498), .Y(n1402) );
  INVX1 U530 ( .A(n1402), .Y(n1761) );
  INVX1 U532 ( .A(n1764), .Y(n1762) );
  INVX1 U534 ( .A(n1762), .Y(n1763) );
  AND2X1 U536 ( .A(n8811), .B(n10498), .Y(n1401) );
  INVX1 U538 ( .A(n1401), .Y(n1764) );
  INVX1 U540 ( .A(n1767), .Y(n1765) );
  INVX1 U542 ( .A(n1765), .Y(n1766) );
  AND2X1 U544 ( .A(n8814), .B(n10498), .Y(n1400) );
  INVX1 U546 ( .A(n1400), .Y(n1767) );
  INVX1 U548 ( .A(n1770), .Y(n1768) );
  INVX1 U550 ( .A(n1768), .Y(n1769) );
  AND2X1 U552 ( .A(n8817), .B(n10498), .Y(n1399) );
  INVX1 U554 ( .A(n1399), .Y(n1770) );
  INVX1 U556 ( .A(n1773), .Y(n1771) );
  INVX1 U558 ( .A(n1771), .Y(n1772) );
  AND2X1 U560 ( .A(n8820), .B(n10498), .Y(n1398) );
  INVX1 U562 ( .A(n1398), .Y(n1773) );
  INVX1 U564 ( .A(n1776), .Y(n1774) );
  INVX1 U566 ( .A(n1774), .Y(n1775) );
  AND2X1 U568 ( .A(n8823), .B(n10498), .Y(n1397) );
  INVX1 U570 ( .A(n1397), .Y(n1776) );
  INVX1 U572 ( .A(n1779), .Y(n1777) );
  INVX1 U574 ( .A(n1777), .Y(n1778) );
  AND2X1 U576 ( .A(n8826), .B(n10498), .Y(n1396) );
  INVX1 U578 ( .A(n1396), .Y(n1779) );
  INVX1 U580 ( .A(n1782), .Y(n1780) );
  INVX1 U582 ( .A(n1780), .Y(n1781) );
  AND2X1 U584 ( .A(n8829), .B(n10498), .Y(n1395) );
  INVX1 U586 ( .A(n1395), .Y(n1782) );
  INVX1 U588 ( .A(n1785), .Y(n1783) );
  INVX1 U589 ( .A(n1783), .Y(n1784) );
  AND2X1 U591 ( .A(n8832), .B(n10498), .Y(n1394) );
  INVX1 U593 ( .A(n1394), .Y(n1785) );
  INVX1 U595 ( .A(n1788), .Y(n1786) );
  INVX1 U597 ( .A(n1786), .Y(n1787) );
  AND2X1 U599 ( .A(n8835), .B(n10498), .Y(n1393) );
  INVX1 U601 ( .A(n1393), .Y(n1788) );
  INVX1 U603 ( .A(n1791), .Y(n1789) );
  INVX1 U605 ( .A(n1789), .Y(n1790) );
  AND2X1 U607 ( .A(n8838), .B(n10498), .Y(n1392) );
  INVX1 U609 ( .A(n1392), .Y(n1791) );
  INVX1 U611 ( .A(n1794), .Y(n1792) );
  INVX1 U613 ( .A(n1792), .Y(n1793) );
  AND2X1 U615 ( .A(n8841), .B(n10498), .Y(n1391) );
  INVX1 U617 ( .A(n1391), .Y(n1794) );
  INVX1 U619 ( .A(n1797), .Y(n1795) );
  INVX1 U621 ( .A(n1795), .Y(n1796) );
  AND2X1 U623 ( .A(n7212), .B(n10496), .Y(n1389) );
  INVX1 U625 ( .A(n1389), .Y(n1797) );
  INVX1 U627 ( .A(n1800), .Y(n1798) );
  INVX1 U629 ( .A(n1798), .Y(n1799) );
  AND2X1 U631 ( .A(n7215), .B(n10496), .Y(n1388) );
  INVX1 U633 ( .A(n1388), .Y(n1800) );
  INVX1 U635 ( .A(n1803), .Y(n1801) );
  INVX1 U637 ( .A(n1801), .Y(n1802) );
  AND2X1 U639 ( .A(n7218), .B(n10496), .Y(n1387) );
  INVX1 U641 ( .A(n1387), .Y(n1803) );
  INVX1 U643 ( .A(n1806), .Y(n1804) );
  INVX1 U645 ( .A(n1804), .Y(n1805) );
  AND2X1 U647 ( .A(n7221), .B(n10496), .Y(n1386) );
  INVX1 U649 ( .A(n1386), .Y(n1806) );
  INVX1 U651 ( .A(n1809), .Y(n1807) );
  INVX1 U653 ( .A(n1807), .Y(n1808) );
  AND2X1 U655 ( .A(n7224), .B(n10496), .Y(n1385) );
  INVX1 U657 ( .A(n1385), .Y(n1809) );
  INVX1 U658 ( .A(n1812), .Y(n1810) );
  INVX1 U659 ( .A(n1810), .Y(n1811) );
  AND2X1 U662 ( .A(n7227), .B(n10496), .Y(n1384) );
  INVX1 U664 ( .A(n1384), .Y(n1812) );
  INVX1 U666 ( .A(n1815), .Y(n1813) );
  INVX1 U668 ( .A(n1813), .Y(n1814) );
  AND2X1 U670 ( .A(n7230), .B(n10496), .Y(n1383) );
  INVX1 U672 ( .A(n1383), .Y(n1815) );
  INVX1 U674 ( .A(n1818), .Y(n1816) );
  INVX1 U676 ( .A(n1816), .Y(n1817) );
  AND2X1 U678 ( .A(n7233), .B(n10496), .Y(n1382) );
  INVX1 U680 ( .A(n1382), .Y(n1818) );
  INVX1 U682 ( .A(n1821), .Y(n1819) );
  INVX1 U684 ( .A(n1819), .Y(n1820) );
  AND2X1 U686 ( .A(n7236), .B(n10496), .Y(n1381) );
  INVX1 U688 ( .A(n1381), .Y(n1821) );
  INVX1 U690 ( .A(n1824), .Y(n1822) );
  INVX1 U692 ( .A(n1822), .Y(n1823) );
  AND2X1 U694 ( .A(n7239), .B(n10496), .Y(n1380) );
  INVX1 U696 ( .A(n1380), .Y(n1824) );
  INVX1 U698 ( .A(n1827), .Y(n1825) );
  INVX1 U700 ( .A(n1825), .Y(n1826) );
  AND2X1 U702 ( .A(n7242), .B(n10496), .Y(n1379) );
  INVX1 U704 ( .A(n1379), .Y(n1827) );
  INVX1 U706 ( .A(n1830), .Y(n1828) );
  INVX1 U708 ( .A(n1828), .Y(n1829) );
  AND2X1 U710 ( .A(n7245), .B(n10496), .Y(n1378) );
  INVX1 U712 ( .A(n1378), .Y(n1830) );
  INVX1 U714 ( .A(n1833), .Y(n1831) );
  INVX1 U716 ( .A(n1831), .Y(n1832) );
  AND2X1 U718 ( .A(n7248), .B(n10496), .Y(n1377) );
  INVX1 U720 ( .A(n1377), .Y(n1833) );
  INVX1 U722 ( .A(n1836), .Y(n1834) );
  INVX1 U724 ( .A(n1834), .Y(n1835) );
  AND2X1 U726 ( .A(n7251), .B(n10496), .Y(n1376) );
  INVX1 U728 ( .A(n1376), .Y(n1836) );
  INVX1 U729 ( .A(n1839), .Y(n1837) );
  INVX1 U731 ( .A(n1837), .Y(n1838) );
  AND2X1 U733 ( .A(n7254), .B(n10496), .Y(n1375) );
  INVX1 U735 ( .A(n1375), .Y(n1839) );
  INVX1 U737 ( .A(n1842), .Y(n1840) );
  INVX1 U739 ( .A(n1840), .Y(n1841) );
  AND2X1 U741 ( .A(n7257), .B(n10496), .Y(n1374) );
  INVX1 U743 ( .A(n1374), .Y(n1842) );
  INVX1 U745 ( .A(n1845), .Y(n1843) );
  INVX1 U747 ( .A(n1843), .Y(n1844) );
  AND2X1 U749 ( .A(n7260), .B(n10496), .Y(n1373) );
  INVX1 U751 ( .A(n1373), .Y(n1845) );
  INVX1 U753 ( .A(n1848), .Y(n1846) );
  INVX1 U755 ( .A(n1846), .Y(n1847) );
  AND2X1 U757 ( .A(n7263), .B(n10496), .Y(n1372) );
  INVX1 U759 ( .A(n1372), .Y(n1848) );
  INVX1 U761 ( .A(n1851), .Y(n1849) );
  INVX1 U763 ( .A(n1849), .Y(n1850) );
  AND2X1 U765 ( .A(n7266), .B(n10496), .Y(n1371) );
  INVX1 U767 ( .A(n1371), .Y(n1851) );
  INVX1 U769 ( .A(n1854), .Y(n1852) );
  INVX1 U771 ( .A(n1852), .Y(n1853) );
  AND2X1 U773 ( .A(n7269), .B(n10496), .Y(n1370) );
  INVX1 U775 ( .A(n1370), .Y(n1854) );
  INVX1 U777 ( .A(n1857), .Y(n1855) );
  INVX1 U779 ( .A(n1855), .Y(n1856) );
  AND2X1 U781 ( .A(n7272), .B(n10496), .Y(n1369) );
  INVX1 U783 ( .A(n1369), .Y(n1857) );
  INVX1 U785 ( .A(n1860), .Y(n1858) );
  INVX1 U787 ( .A(n1858), .Y(n1859) );
  AND2X1 U789 ( .A(n7275), .B(n10496), .Y(n1368) );
  INVX1 U791 ( .A(n1368), .Y(n1860) );
  INVX1 U793 ( .A(n1863), .Y(n1861) );
  INVX1 U795 ( .A(n1861), .Y(n1862) );
  AND2X1 U797 ( .A(n7278), .B(n10496), .Y(n1367) );
  INVX1 U798 ( .A(n1367), .Y(n1863) );
  INVX1 U800 ( .A(n1866), .Y(n1864) );
  INVX1 U802 ( .A(n1864), .Y(n1865) );
  AND2X1 U804 ( .A(n7281), .B(n10496), .Y(n1366) );
  INVX1 U806 ( .A(n1366), .Y(n1866) );
  INVX1 U808 ( .A(n1869), .Y(n1867) );
  INVX1 U810 ( .A(n1867), .Y(n1868) );
  AND2X1 U812 ( .A(n7284), .B(n10496), .Y(n1365) );
  INVX1 U814 ( .A(n1365), .Y(n1869) );
  INVX1 U816 ( .A(n1872), .Y(n1870) );
  INVX1 U818 ( .A(n1870), .Y(n1871) );
  AND2X1 U820 ( .A(n7287), .B(n10496), .Y(n1364) );
  INVX1 U822 ( .A(n1364), .Y(n1872) );
  INVX1 U824 ( .A(n1875), .Y(n1873) );
  INVX1 U826 ( .A(n1873), .Y(n1874) );
  AND2X1 U828 ( .A(n7290), .B(n10496), .Y(n1363) );
  INVX1 U830 ( .A(n1363), .Y(n1875) );
  INVX1 U832 ( .A(n1878), .Y(n1876) );
  INVX1 U834 ( .A(n1876), .Y(n1877) );
  AND2X1 U836 ( .A(n7293), .B(n10496), .Y(n1362) );
  INVX1 U838 ( .A(n1362), .Y(n1878) );
  INVX1 U840 ( .A(n1881), .Y(n1879) );
  INVX1 U842 ( .A(n1879), .Y(n1880) );
  AND2X1 U844 ( .A(n7296), .B(n10496), .Y(n1361) );
  INVX1 U846 ( .A(n1361), .Y(n1881) );
  INVX1 U848 ( .A(n1884), .Y(n1882) );
  INVX1 U850 ( .A(n1882), .Y(n1883) );
  AND2X1 U852 ( .A(n7299), .B(n10496), .Y(n1360) );
  INVX1 U854 ( .A(n1360), .Y(n1884) );
  INVX1 U856 ( .A(n1887), .Y(n1885) );
  INVX1 U858 ( .A(n1885), .Y(n1886) );
  AND2X1 U860 ( .A(n7302), .B(n10496), .Y(n1359) );
  INVX1 U862 ( .A(n1359), .Y(n1887) );
  INVX1 U864 ( .A(n1890), .Y(n1888) );
  INVX1 U866 ( .A(n1888), .Y(n1889) );
  AND2X1 U867 ( .A(n7305), .B(n10496), .Y(n1358) );
  INVX1 U869 ( .A(n1358), .Y(n1890) );
  INVX1 U871 ( .A(n1893), .Y(n1891) );
  INVX1 U873 ( .A(n1891), .Y(n1892) );
  AND2X1 U875 ( .A(n7308), .B(n10496), .Y(n1357) );
  INVX1 U877 ( .A(n1357), .Y(n1893) );
  INVX1 U879 ( .A(n1896), .Y(n1894) );
  INVX1 U881 ( .A(n1894), .Y(n1895) );
  AND2X1 U883 ( .A(n7311), .B(n10496), .Y(n1356) );
  INVX1 U885 ( .A(n1356), .Y(n1896) );
  INVX1 U887 ( .A(n1899), .Y(n1897) );
  INVX1 U889 ( .A(n1897), .Y(n1898) );
  AND2X1 U891 ( .A(n8844), .B(n10504), .Y(n1354) );
  INVX1 U893 ( .A(n1354), .Y(n1899) );
  INVX1 U895 ( .A(n1902), .Y(n1900) );
  INVX1 U897 ( .A(n1900), .Y(n1901) );
  AND2X1 U899 ( .A(n8847), .B(n10504), .Y(n1353) );
  INVX1 U901 ( .A(n1353), .Y(n1902) );
  INVX1 U903 ( .A(n1905), .Y(n1903) );
  INVX1 U905 ( .A(n1903), .Y(n1904) );
  AND2X1 U907 ( .A(n8850), .B(n10504), .Y(n1352) );
  INVX1 U909 ( .A(n1352), .Y(n1905) );
  INVX1 U911 ( .A(n1908), .Y(n1906) );
  INVX1 U913 ( .A(n1906), .Y(n1907) );
  AND2X1 U915 ( .A(n8853), .B(n10504), .Y(n1351) );
  INVX1 U917 ( .A(n1351), .Y(n1908) );
  INVX1 U919 ( .A(n1911), .Y(n1909) );
  INVX1 U921 ( .A(n1909), .Y(n1910) );
  AND2X1 U923 ( .A(n8856), .B(n10504), .Y(n1350) );
  INVX1 U925 ( .A(n1350), .Y(n1911) );
  INVX1 U927 ( .A(n1914), .Y(n1912) );
  INVX1 U929 ( .A(n1912), .Y(n1913) );
  AND2X1 U931 ( .A(n8859), .B(n10504), .Y(n1349) );
  INVX1 U933 ( .A(n1349), .Y(n1914) );
  INVX1 U935 ( .A(n1917), .Y(n1915) );
  INVX1 U936 ( .A(n1915), .Y(n1916) );
  AND2X1 U938 ( .A(n8862), .B(n10504), .Y(n1348) );
  INVX1 U940 ( .A(n1348), .Y(n1917) );
  INVX1 U942 ( .A(n1920), .Y(n1918) );
  INVX1 U944 ( .A(n1918), .Y(n1919) );
  AND2X1 U946 ( .A(n8865), .B(n10504), .Y(n1347) );
  INVX1 U948 ( .A(n1347), .Y(n1920) );
  INVX1 U950 ( .A(n1923), .Y(n1921) );
  INVX1 U952 ( .A(n1921), .Y(n1922) );
  AND2X1 U954 ( .A(n8868), .B(n10504), .Y(n1346) );
  INVX1 U956 ( .A(n1346), .Y(n1923) );
  INVX1 U958 ( .A(n1926), .Y(n1924) );
  INVX1 U960 ( .A(n1924), .Y(n1925) );
  AND2X1 U962 ( .A(n8871), .B(n10504), .Y(n1345) );
  INVX1 U964 ( .A(n1345), .Y(n1926) );
  INVX1 U966 ( .A(n1929), .Y(n1927) );
  INVX1 U968 ( .A(n1927), .Y(n1928) );
  AND2X1 U970 ( .A(n8874), .B(n10504), .Y(n1344) );
  INVX1 U972 ( .A(n1344), .Y(n1929) );
  INVX1 U974 ( .A(n1932), .Y(n1930) );
  INVX1 U976 ( .A(n1930), .Y(n1931) );
  AND2X1 U978 ( .A(n8877), .B(n10504), .Y(n1343) );
  INVX1 U980 ( .A(n1343), .Y(n1932) );
  INVX1 U982 ( .A(n1935), .Y(n1933) );
  INVX1 U984 ( .A(n1933), .Y(n1934) );
  AND2X1 U986 ( .A(n8880), .B(n10504), .Y(n1342) );
  INVX1 U988 ( .A(n1342), .Y(n1935) );
  INVX1 U990 ( .A(n1938), .Y(n1936) );
  INVX1 U992 ( .A(n1936), .Y(n1937) );
  AND2X1 U994 ( .A(n8883), .B(n10504), .Y(n1341) );
  INVX1 U996 ( .A(n1341), .Y(n1938) );
  INVX1 U998 ( .A(n1941), .Y(n1939) );
  INVX1 U1000 ( .A(n1939), .Y(n1940) );
  AND2X1 U1002 ( .A(n8886), .B(n10504), .Y(n1340) );
  INVX1 U1004 ( .A(n1340), .Y(n1941) );
  INVX1 U1005 ( .A(n1944), .Y(n1942) );
  INVX1 U1007 ( .A(n1942), .Y(n1943) );
  AND2X1 U1009 ( .A(n8889), .B(n10504), .Y(n1339) );
  INVX1 U1011 ( .A(n1339), .Y(n1944) );
  INVX1 U1013 ( .A(n1947), .Y(n1945) );
  INVX1 U1015 ( .A(n1945), .Y(n1946) );
  AND2X1 U1017 ( .A(n8892), .B(n10504), .Y(n1338) );
  INVX1 U1019 ( .A(n1338), .Y(n1947) );
  INVX1 U1021 ( .A(n1950), .Y(n1948) );
  INVX1 U1023 ( .A(n1948), .Y(n1949) );
  AND2X1 U1025 ( .A(n8895), .B(n10504), .Y(n1337) );
  INVX1 U1027 ( .A(n1337), .Y(n1950) );
  INVX1 U1029 ( .A(n1953), .Y(n1951) );
  INVX1 U1031 ( .A(n1951), .Y(n1952) );
  AND2X1 U1033 ( .A(n8898), .B(n10504), .Y(n1336) );
  INVX1 U1035 ( .A(n1336), .Y(n1953) );
  INVX1 U1037 ( .A(n1956), .Y(n1954) );
  INVX1 U1039 ( .A(n1954), .Y(n1955) );
  AND2X1 U1041 ( .A(n8901), .B(n10504), .Y(n1335) );
  INVX1 U1043 ( .A(n1335), .Y(n1956) );
  INVX1 U1045 ( .A(n1959), .Y(n1957) );
  INVX1 U1047 ( .A(n1957), .Y(n1958) );
  AND2X1 U1049 ( .A(n8904), .B(n10504), .Y(n1334) );
  INVX1 U1051 ( .A(n1334), .Y(n1959) );
  INVX1 U1053 ( .A(n1962), .Y(n1960) );
  INVX1 U1055 ( .A(n1960), .Y(n1961) );
  AND2X1 U1057 ( .A(n8907), .B(n10504), .Y(n1333) );
  INVX1 U1059 ( .A(n1333), .Y(n1962) );
  INVX1 U1061 ( .A(n1965), .Y(n1963) );
  INVX1 U1063 ( .A(n1963), .Y(n1964) );
  AND2X1 U1065 ( .A(n8910), .B(n10504), .Y(n1332) );
  INVX1 U1067 ( .A(n1332), .Y(n1965) );
  INVX1 U1069 ( .A(n1968), .Y(n1966) );
  INVX1 U1071 ( .A(n1966), .Y(n1967) );
  AND2X1 U1073 ( .A(n8913), .B(n10504), .Y(n1331) );
  INVX1 U1074 ( .A(n1331), .Y(n1968) );
  INVX1 U1076 ( .A(n1971), .Y(n1969) );
  INVX1 U1078 ( .A(n1969), .Y(n1970) );
  AND2X1 U1080 ( .A(n8916), .B(n10504), .Y(n1330) );
  INVX1 U1082 ( .A(n1330), .Y(n1971) );
  INVX1 U1084 ( .A(n1974), .Y(n1972) );
  INVX1 U1086 ( .A(n1972), .Y(n1973) );
  AND2X1 U1088 ( .A(n8919), .B(n10504), .Y(n1329) );
  INVX1 U1090 ( .A(n1329), .Y(n1974) );
  INVX1 U1092 ( .A(n1977), .Y(n1975) );
  INVX1 U1094 ( .A(n1975), .Y(n1976) );
  AND2X1 U1096 ( .A(n8922), .B(n10504), .Y(n1328) );
  INVX1 U1098 ( .A(n1328), .Y(n1977) );
  INVX1 U1100 ( .A(n1980), .Y(n1978) );
  INVX1 U1102 ( .A(n1978), .Y(n1979) );
  AND2X1 U1104 ( .A(n8925), .B(n10504), .Y(n1327) );
  INVX1 U1106 ( .A(n1327), .Y(n1980) );
  INVX1 U1108 ( .A(n1983), .Y(n1981) );
  INVX1 U1110 ( .A(n1981), .Y(n1982) );
  AND2X1 U1112 ( .A(n8928), .B(n10504), .Y(n1326) );
  INVX1 U1114 ( .A(n1326), .Y(n1983) );
  INVX1 U1116 ( .A(n1986), .Y(n1984) );
  INVX1 U1118 ( .A(n1984), .Y(n1985) );
  AND2X1 U1120 ( .A(n8931), .B(n10504), .Y(n1325) );
  INVX1 U1122 ( .A(n1325), .Y(n1986) );
  INVX1 U1124 ( .A(n2499), .Y(n1987) );
  INVX1 U1126 ( .A(n1987), .Y(n2498) );
  AND2X1 U1128 ( .A(n8934), .B(n10504), .Y(n1324) );
  INVX1 U1130 ( .A(n1324), .Y(n2499) );
  INVX1 U1132 ( .A(n2502), .Y(n2500) );
  INVX1 U1134 ( .A(n2500), .Y(n2501) );
  AND2X1 U1136 ( .A(n8937), .B(n10504), .Y(n1323) );
  INVX1 U1138 ( .A(n1323), .Y(n2502) );
  INVX1 U1140 ( .A(n2505), .Y(n2503) );
  INVX1 U1142 ( .A(n2503), .Y(n2504) );
  AND2X1 U1143 ( .A(n8940), .B(n10504), .Y(n1322) );
  INVX1 U1145 ( .A(n1322), .Y(n2505) );
  INVX1 U1147 ( .A(n2508), .Y(n2506) );
  INVX1 U1149 ( .A(n2506), .Y(n2507) );
  AND2X1 U1151 ( .A(n8943), .B(n10504), .Y(n1321) );
  INVX1 U1153 ( .A(n1321), .Y(n2508) );
  INVX1 U1155 ( .A(n2511), .Y(n2509) );
  INVX1 U1157 ( .A(n2509), .Y(n2510) );
  AND2X1 U1159 ( .A(n7314), .B(n1284), .Y(n1318) );
  INVX1 U1161 ( .A(n1318), .Y(n2511) );
  INVX1 U1163 ( .A(n2514), .Y(n2512) );
  INVX1 U1165 ( .A(n2512), .Y(n2513) );
  AND2X1 U1167 ( .A(n7317), .B(n1284), .Y(n1317) );
  INVX1 U1169 ( .A(n1317), .Y(n2514) );
  INVX1 U1171 ( .A(n2517), .Y(n2515) );
  INVX1 U1173 ( .A(n2515), .Y(n2516) );
  AND2X1 U1175 ( .A(n7320), .B(n1284), .Y(n1316) );
  INVX1 U1177 ( .A(n1316), .Y(n2517) );
  INVX1 U1179 ( .A(n2520), .Y(n2518) );
  INVX1 U1181 ( .A(n2518), .Y(n2519) );
  AND2X1 U1183 ( .A(n7323), .B(n1284), .Y(n1315) );
  INVX1 U1185 ( .A(n1315), .Y(n2520) );
  INVX1 U1187 ( .A(n2523), .Y(n2521) );
  INVX1 U1189 ( .A(n2521), .Y(n2522) );
  AND2X1 U1191 ( .A(n7326), .B(n1284), .Y(n1314) );
  INVX1 U1193 ( .A(n1314), .Y(n2523) );
  INVX1 U1195 ( .A(n2526), .Y(n2524) );
  INVX1 U1197 ( .A(n2524), .Y(n2525) );
  AND2X1 U1199 ( .A(n7329), .B(n1284), .Y(n1313) );
  INVX1 U1201 ( .A(n1313), .Y(n2526) );
  INVX1 U1203 ( .A(n2529), .Y(n2527) );
  INVX1 U1205 ( .A(n2527), .Y(n2528) );
  AND2X1 U1207 ( .A(n7332), .B(n1284), .Y(n1312) );
  INVX1 U1209 ( .A(n1312), .Y(n2529) );
  INVX1 U1211 ( .A(n2535), .Y(n2530) );
  INVX1 U1212 ( .A(n2530), .Y(n2531) );
  AND2X1 U1213 ( .A(n7335), .B(n1284), .Y(n1311) );
  INVX1 U1217 ( .A(n1311), .Y(n2535) );
  INVX1 U1219 ( .A(n2550), .Y(n2540) );
  INVX1 U1221 ( .A(n2540), .Y(n2545) );
  AND2X1 U1223 ( .A(n7338), .B(n1284), .Y(n1310) );
  INVX1 U1225 ( .A(n1310), .Y(n2550) );
  INVX1 U1227 ( .A(n2560), .Y(n2552) );
  INVX1 U1229 ( .A(n2552), .Y(n2558) );
  AND2X1 U1231 ( .A(n7341), .B(n1284), .Y(n1309) );
  INVX1 U1233 ( .A(n1309), .Y(n2560) );
  INVX1 U1235 ( .A(n2566), .Y(n2562) );
  INVX1 U1237 ( .A(n2562), .Y(n2564) );
  AND2X1 U1239 ( .A(n7344), .B(n1284), .Y(n1308) );
  INVX1 U1241 ( .A(n1308), .Y(n2566) );
  INVX1 U1243 ( .A(n2572), .Y(n2568) );
  INVX1 U1245 ( .A(n2568), .Y(n2570) );
  AND2X1 U1247 ( .A(n7347), .B(n1284), .Y(n1307) );
  INVX1 U1249 ( .A(n1307), .Y(n2572) );
  INVX1 U1251 ( .A(n2578), .Y(n2574) );
  INVX1 U1253 ( .A(n2574), .Y(n2576) );
  AND2X1 U1255 ( .A(n7350), .B(n1284), .Y(n1306) );
  INVX1 U1257 ( .A(n1306), .Y(n2578) );
  INVX1 U1259 ( .A(n2584), .Y(n2580) );
  INVX1 U1261 ( .A(n2580), .Y(n2582) );
  AND2X1 U1263 ( .A(n7353), .B(n1284), .Y(n1305) );
  INVX1 U1265 ( .A(n1305), .Y(n2584) );
  INVX1 U1267 ( .A(n2590), .Y(n2586) );
  INVX1 U1269 ( .A(n2586), .Y(n2588) );
  AND2X1 U1271 ( .A(n7356), .B(n1284), .Y(n1304) );
  INVX1 U1273 ( .A(n1304), .Y(n2590) );
  INVX1 U1275 ( .A(n2596), .Y(n2592) );
  INVX1 U1277 ( .A(n2592), .Y(n2594) );
  AND2X1 U1279 ( .A(n7359), .B(n1284), .Y(n1303) );
  INVX1 U1281 ( .A(n1303), .Y(n2596) );
  INVX1 U1283 ( .A(n2602), .Y(n2598) );
  INVX1 U1284 ( .A(n2598), .Y(n2600) );
  AND2X1 U1286 ( .A(n7362), .B(n1284), .Y(n1302) );
  INVX1 U1288 ( .A(n1302), .Y(n2602) );
  INVX1 U1290 ( .A(n2608), .Y(n2604) );
  INVX1 U1292 ( .A(n2604), .Y(n2606) );
  AND2X1 U1294 ( .A(n7365), .B(n1284), .Y(n1301) );
  INVX1 U1296 ( .A(n1301), .Y(n2608) );
  INVX1 U1298 ( .A(n2614), .Y(n2610) );
  INVX1 U1300 ( .A(n2610), .Y(n2612) );
  AND2X1 U1302 ( .A(n7368), .B(n1284), .Y(n1300) );
  INVX1 U1304 ( .A(n1300), .Y(n2614) );
  INVX1 U1306 ( .A(n2620), .Y(n2616) );
  INVX1 U1308 ( .A(n2616), .Y(n2618) );
  AND2X1 U1310 ( .A(n7371), .B(n1284), .Y(n1299) );
  INVX1 U1312 ( .A(n1299), .Y(n2620) );
  INVX1 U1314 ( .A(n2659), .Y(n2645) );
  INVX1 U1316 ( .A(n2645), .Y(n2656) );
  AND2X1 U1318 ( .A(n7374), .B(n1284), .Y(n1298) );
  INVX1 U1320 ( .A(n1298), .Y(n2659) );
  INVX1 U1322 ( .A(n3751), .Y(n3749) );
  INVX1 U1324 ( .A(n3749), .Y(n3750) );
  AND2X1 U1326 ( .A(n7377), .B(n1284), .Y(n1297) );
  INVX1 U1328 ( .A(n1297), .Y(n3751) );
  INVX1 U1330 ( .A(n3754), .Y(n3752) );
  INVX1 U1332 ( .A(n3752), .Y(n3753) );
  AND2X1 U1334 ( .A(n7380), .B(n1284), .Y(n1296) );
  INVX1 U1336 ( .A(n1296), .Y(n3754) );
  INVX1 U1338 ( .A(n3757), .Y(n3755) );
  INVX1 U1340 ( .A(n3755), .Y(n3756) );
  AND2X1 U1342 ( .A(n7383), .B(n1284), .Y(n1295) );
  INVX1 U1344 ( .A(n1295), .Y(n3757) );
  INVX1 U1346 ( .A(n3760), .Y(n3758) );
  INVX1 U1348 ( .A(n3758), .Y(n3759) );
  AND2X1 U1350 ( .A(n7386), .B(n1284), .Y(n1294) );
  INVX1 U1352 ( .A(n1294), .Y(n3760) );
  INVX1 U1353 ( .A(n3763), .Y(n3761) );
  INVX1 U1355 ( .A(n3761), .Y(n3762) );
  AND2X1 U1357 ( .A(n7389), .B(n1284), .Y(n1293) );
  INVX1 U1359 ( .A(n1293), .Y(n3763) );
  INVX1 U1361 ( .A(n3766), .Y(n3764) );
  INVX1 U1363 ( .A(n3764), .Y(n3765) );
  AND2X1 U1365 ( .A(n7392), .B(n1284), .Y(n1292) );
  INVX1 U1367 ( .A(n1292), .Y(n3766) );
  INVX1 U1369 ( .A(n3769), .Y(n3767) );
  INVX1 U1371 ( .A(n3767), .Y(n3768) );
  AND2X1 U1373 ( .A(n7395), .B(n1284), .Y(n1291) );
  INVX1 U1375 ( .A(n1291), .Y(n3769) );
  INVX1 U1377 ( .A(n3772), .Y(n3770) );
  INVX1 U1379 ( .A(n3770), .Y(n3771) );
  AND2X1 U1381 ( .A(n7398), .B(n1284), .Y(n1290) );
  INVX1 U1383 ( .A(n1290), .Y(n3772) );
  INVX1 U1385 ( .A(n3775), .Y(n3773) );
  INVX1 U1387 ( .A(n3773), .Y(n3774) );
  AND2X1 U1389 ( .A(n7401), .B(n1284), .Y(n1289) );
  INVX1 U1391 ( .A(n1289), .Y(n3775) );
  INVX1 U1393 ( .A(n3778), .Y(n3776) );
  INVX1 U1395 ( .A(n3776), .Y(n3777) );
  AND2X1 U1397 ( .A(n7404), .B(n1284), .Y(n1288) );
  INVX1 U1399 ( .A(n1288), .Y(n3778) );
  INVX1 U1401 ( .A(n3781), .Y(n3779) );
  INVX1 U1403 ( .A(n3779), .Y(n3780) );
  AND2X1 U1405 ( .A(n7407), .B(n1284), .Y(n1287) );
  INVX1 U1407 ( .A(n1287), .Y(n3781) );
  INVX1 U1409 ( .A(n3784), .Y(n3782) );
  INVX1 U1411 ( .A(n3782), .Y(n3783) );
  AND2X1 U1413 ( .A(n7410), .B(n1284), .Y(n1286) );
  INVX1 U1415 ( .A(n1286), .Y(n3784) );
  INVX1 U1417 ( .A(n3787), .Y(n3785) );
  INVX1 U1419 ( .A(n3785), .Y(n3786) );
  AND2X1 U1421 ( .A(n7413), .B(n1284), .Y(n1285) );
  INVX1 U1422 ( .A(n1285), .Y(n3787) );
  INVX1 U1424 ( .A(n3790), .Y(n3788) );
  INVX1 U1426 ( .A(n3788), .Y(n3789) );
  AND2X1 U1428 ( .A(n8946), .B(n1249), .Y(n1283) );
  INVX1 U1430 ( .A(n1283), .Y(n3790) );
  INVX1 U1432 ( .A(n3793), .Y(n3791) );
  INVX1 U1434 ( .A(n3791), .Y(n3792) );
  AND2X1 U1436 ( .A(n8949), .B(n1249), .Y(n1282) );
  INVX1 U1438 ( .A(n1282), .Y(n3793) );
  INVX1 U1440 ( .A(n3796), .Y(n3794) );
  INVX1 U1442 ( .A(n3794), .Y(n3795) );
  AND2X1 U1444 ( .A(n8952), .B(n1249), .Y(n1281) );
  INVX1 U1446 ( .A(n1281), .Y(n3796) );
  INVX1 U1448 ( .A(n3799), .Y(n3797) );
  INVX1 U1450 ( .A(n3797), .Y(n3798) );
  AND2X1 U1452 ( .A(n8955), .B(n1249), .Y(n1280) );
  INVX1 U1454 ( .A(n1280), .Y(n3799) );
  INVX1 U1456 ( .A(n3802), .Y(n3800) );
  INVX1 U1458 ( .A(n3800), .Y(n3801) );
  AND2X1 U1460 ( .A(n8958), .B(n1249), .Y(n1279) );
  INVX1 U1462 ( .A(n1279), .Y(n3802) );
  INVX1 U1464 ( .A(n3805), .Y(n3803) );
  INVX1 U1466 ( .A(n3803), .Y(n3804) );
  AND2X1 U1468 ( .A(n8961), .B(n1249), .Y(n1278) );
  INVX1 U1470 ( .A(n1278), .Y(n3805) );
  INVX1 U1472 ( .A(n3808), .Y(n3806) );
  INVX1 U1474 ( .A(n3806), .Y(n3807) );
  AND2X1 U1476 ( .A(n8964), .B(n1249), .Y(n1277) );
  INVX1 U1478 ( .A(n1277), .Y(n3808) );
  INVX1 U1480 ( .A(n3811), .Y(n3809) );
  INVX1 U1482 ( .A(n3809), .Y(n3810) );
  AND2X1 U1484 ( .A(n8967), .B(n1249), .Y(n1276) );
  INVX1 U1486 ( .A(n1276), .Y(n3811) );
  INVX1 U1488 ( .A(n3814), .Y(n3812) );
  INVX1 U1490 ( .A(n3812), .Y(n3813) );
  AND2X1 U1491 ( .A(n8970), .B(n1249), .Y(n1275) );
  INVX1 U1493 ( .A(n1275), .Y(n3814) );
  INVX1 U1495 ( .A(n3817), .Y(n3815) );
  INVX1 U1497 ( .A(n3815), .Y(n3816) );
  AND2X1 U1499 ( .A(n8973), .B(n1249), .Y(n1274) );
  INVX1 U1501 ( .A(n1274), .Y(n3817) );
  INVX1 U1503 ( .A(n3820), .Y(n3818) );
  INVX1 U1505 ( .A(n3818), .Y(n3819) );
  AND2X1 U1507 ( .A(n8976), .B(n1249), .Y(n1273) );
  INVX1 U1509 ( .A(n1273), .Y(n3820) );
  INVX1 U1511 ( .A(n3823), .Y(n3821) );
  INVX1 U1513 ( .A(n3821), .Y(n3822) );
  AND2X1 U1515 ( .A(n8979), .B(n1249), .Y(n1272) );
  INVX1 U1517 ( .A(n1272), .Y(n3823) );
  INVX1 U1519 ( .A(n3826), .Y(n3824) );
  INVX1 U1521 ( .A(n3824), .Y(n3825) );
  AND2X1 U1523 ( .A(n8982), .B(n1249), .Y(n1271) );
  INVX1 U1525 ( .A(n1271), .Y(n3826) );
  INVX1 U1527 ( .A(n3829), .Y(n3827) );
  INVX1 U1529 ( .A(n3827), .Y(n3828) );
  AND2X1 U1531 ( .A(n8985), .B(n1249), .Y(n1270) );
  INVX1 U1533 ( .A(n1270), .Y(n3829) );
  INVX1 U1535 ( .A(n3832), .Y(n3830) );
  INVX1 U1537 ( .A(n3830), .Y(n3831) );
  AND2X1 U1539 ( .A(n8988), .B(n1249), .Y(n1269) );
  INVX1 U1541 ( .A(n1269), .Y(n3832) );
  INVX1 U1543 ( .A(n3835), .Y(n3833) );
  INVX1 U1545 ( .A(n3833), .Y(n3834) );
  AND2X1 U1547 ( .A(n8991), .B(n1249), .Y(n1268) );
  INVX1 U1549 ( .A(n1268), .Y(n3835) );
  INVX1 U1551 ( .A(n3838), .Y(n3836) );
  INVX1 U1553 ( .A(n3836), .Y(n3837) );
  AND2X1 U1555 ( .A(n8994), .B(n1249), .Y(n1267) );
  INVX1 U1557 ( .A(n1267), .Y(n3838) );
  INVX1 U1559 ( .A(n3841), .Y(n3839) );
  INVX1 U1560 ( .A(n3839), .Y(n3840) );
  AND2X1 U1562 ( .A(n8997), .B(n1249), .Y(n1266) );
  INVX1 U1564 ( .A(n1266), .Y(n3841) );
  INVX1 U1566 ( .A(n3844), .Y(n3842) );
  INVX1 U1568 ( .A(n3842), .Y(n3843) );
  AND2X1 U1570 ( .A(n9000), .B(n1249), .Y(n1265) );
  INVX1 U1572 ( .A(n1265), .Y(n3844) );
  INVX1 U1574 ( .A(n3847), .Y(n3845) );
  INVX1 U1576 ( .A(n3845), .Y(n3846) );
  AND2X1 U1578 ( .A(n9003), .B(n1249), .Y(n1264) );
  INVX1 U1580 ( .A(n1264), .Y(n3847) );
  INVX1 U1582 ( .A(n3850), .Y(n3848) );
  INVX1 U1584 ( .A(n3848), .Y(n3849) );
  AND2X1 U1586 ( .A(n9006), .B(n1249), .Y(n1263) );
  INVX1 U1588 ( .A(n1263), .Y(n3850) );
  INVX1 U1590 ( .A(n3853), .Y(n3851) );
  INVX1 U1592 ( .A(n3851), .Y(n3852) );
  AND2X1 U1594 ( .A(n9009), .B(n1249), .Y(n1262) );
  INVX1 U1596 ( .A(n1262), .Y(n3853) );
  INVX1 U1598 ( .A(n3856), .Y(n3854) );
  INVX1 U1600 ( .A(n3854), .Y(n3855) );
  AND2X1 U1602 ( .A(n9012), .B(n1249), .Y(n1261) );
  INVX1 U1604 ( .A(n1261), .Y(n3856) );
  INVX1 U1606 ( .A(n3859), .Y(n3857) );
  INVX1 U1608 ( .A(n3857), .Y(n3858) );
  AND2X1 U1610 ( .A(n9015), .B(n1249), .Y(n1260) );
  INVX1 U1612 ( .A(n1260), .Y(n3859) );
  INVX1 U1614 ( .A(n3862), .Y(n3860) );
  INVX1 U1616 ( .A(n3860), .Y(n3861) );
  AND2X1 U1618 ( .A(n9018), .B(n1249), .Y(n1259) );
  INVX1 U1620 ( .A(n1259), .Y(n3862) );
  INVX1 U1622 ( .A(n3865), .Y(n3863) );
  INVX1 U1624 ( .A(n3863), .Y(n3864) );
  AND2X1 U1626 ( .A(n9021), .B(n1249), .Y(n1258) );
  INVX1 U1628 ( .A(n1258), .Y(n3865) );
  INVX1 U1629 ( .A(n3868), .Y(n3866) );
  INVX1 U1631 ( .A(n3866), .Y(n3867) );
  AND2X1 U1633 ( .A(n9024), .B(n1249), .Y(n1257) );
  INVX1 U1635 ( .A(n1257), .Y(n3868) );
  INVX1 U1637 ( .A(n3871), .Y(n3869) );
  INVX1 U1639 ( .A(n3869), .Y(n3870) );
  AND2X1 U1641 ( .A(n9027), .B(n1249), .Y(n1256) );
  INVX1 U1643 ( .A(n1256), .Y(n3871) );
  INVX1 U1645 ( .A(n3874), .Y(n3872) );
  INVX1 U1647 ( .A(n3872), .Y(n3873) );
  AND2X1 U1649 ( .A(n9030), .B(n1249), .Y(n1255) );
  INVX1 U1651 ( .A(n1255), .Y(n3874) );
  INVX1 U1653 ( .A(n3877), .Y(n3875) );
  INVX1 U1655 ( .A(n3875), .Y(n3876) );
  AND2X1 U1657 ( .A(n9033), .B(n1249), .Y(n1254) );
  INVX1 U1659 ( .A(n1254), .Y(n3877) );
  INVX1 U1661 ( .A(n3880), .Y(n3878) );
  INVX1 U1663 ( .A(n3878), .Y(n3879) );
  AND2X1 U1665 ( .A(n9036), .B(n1249), .Y(n1253) );
  INVX1 U1667 ( .A(n1253), .Y(n3880) );
  INVX1 U1669 ( .A(n3883), .Y(n3881) );
  INVX1 U1671 ( .A(n3881), .Y(n3882) );
  AND2X1 U1673 ( .A(n9039), .B(n1249), .Y(n1252) );
  INVX1 U1675 ( .A(n1252), .Y(n3883) );
  INVX1 U1677 ( .A(n3886), .Y(n3884) );
  INVX1 U1679 ( .A(n3884), .Y(n3885) );
  AND2X1 U1681 ( .A(n9042), .B(n1249), .Y(n1251) );
  INVX1 U1683 ( .A(n1251), .Y(n3886) );
  INVX1 U1685 ( .A(n3889), .Y(n3887) );
  INVX1 U1687 ( .A(n3887), .Y(n3888) );
  AND2X1 U1689 ( .A(n9045), .B(n1249), .Y(n1250) );
  INVX1 U1691 ( .A(n1250), .Y(n3889) );
  INVX1 U1693 ( .A(n3892), .Y(n3890) );
  INVX1 U1695 ( .A(n3890), .Y(n3891) );
  AND2X1 U1697 ( .A(n7416), .B(n10500), .Y(n1247) );
  INVX1 U1698 ( .A(n1247), .Y(n3892) );
  INVX1 U1700 ( .A(n3895), .Y(n3893) );
  INVX1 U1702 ( .A(n3893), .Y(n3894) );
  AND2X1 U1704 ( .A(n7419), .B(n10500), .Y(n1246) );
  INVX1 U1706 ( .A(n1246), .Y(n3895) );
  INVX1 U1708 ( .A(n3898), .Y(n3896) );
  INVX1 U1710 ( .A(n3896), .Y(n3897) );
  AND2X1 U1712 ( .A(n7422), .B(n10500), .Y(n1245) );
  INVX1 U1714 ( .A(n1245), .Y(n3898) );
  INVX1 U1716 ( .A(n3901), .Y(n3899) );
  INVX1 U1718 ( .A(n3899), .Y(n3900) );
  AND2X1 U1720 ( .A(n7425), .B(n10500), .Y(n1244) );
  INVX1 U1722 ( .A(n1244), .Y(n3901) );
  INVX1 U1724 ( .A(n3904), .Y(n3902) );
  INVX1 U1726 ( .A(n3902), .Y(n3903) );
  AND2X1 U1728 ( .A(n7428), .B(n10500), .Y(n1243) );
  INVX1 U1730 ( .A(n1243), .Y(n3904) );
  INVX1 U1732 ( .A(n3907), .Y(n3905) );
  INVX1 U1734 ( .A(n3905), .Y(n3906) );
  AND2X1 U1736 ( .A(n7431), .B(n10500), .Y(n1242) );
  INVX1 U1738 ( .A(n1242), .Y(n3907) );
  INVX1 U1740 ( .A(n3910), .Y(n3908) );
  INVX1 U1742 ( .A(n3908), .Y(n3909) );
  AND2X1 U1744 ( .A(n7434), .B(n10500), .Y(n1241) );
  INVX1 U1746 ( .A(n1241), .Y(n3910) );
  INVX1 U1748 ( .A(n3913), .Y(n3911) );
  INVX1 U1750 ( .A(n3911), .Y(n3912) );
  AND2X1 U1752 ( .A(n7437), .B(n10500), .Y(n1240) );
  INVX1 U1754 ( .A(n1240), .Y(n3913) );
  INVX1 U1756 ( .A(n3916), .Y(n3914) );
  INVX1 U1758 ( .A(n3914), .Y(n3915) );
  AND2X1 U1760 ( .A(n7440), .B(n10500), .Y(n1239) );
  INVX1 U1762 ( .A(n1239), .Y(n3916) );
  INVX1 U1764 ( .A(n3919), .Y(n3917) );
  INVX1 U1766 ( .A(n3917), .Y(n3918) );
  AND2X1 U1767 ( .A(n7443), .B(n10500), .Y(n1238) );
  INVX1 U1768 ( .A(n1238), .Y(n3919) );
  INVX1 U1769 ( .A(n3922), .Y(n3920) );
  INVX1 U1772 ( .A(n3920), .Y(n3921) );
  AND2X1 U1774 ( .A(n7446), .B(n10500), .Y(n1237) );
  INVX1 U1776 ( .A(n1237), .Y(n3922) );
  INVX1 U1778 ( .A(n3925), .Y(n3923) );
  INVX1 U1780 ( .A(n3923), .Y(n3924) );
  AND2X1 U1782 ( .A(n7449), .B(n10500), .Y(n1236) );
  INVX1 U1784 ( .A(n1236), .Y(n3925) );
  INVX1 U1786 ( .A(n3928), .Y(n3926) );
  INVX1 U1788 ( .A(n3926), .Y(n3927) );
  AND2X1 U1790 ( .A(n7452), .B(n10500), .Y(n1235) );
  INVX1 U1792 ( .A(n1235), .Y(n3928) );
  INVX1 U1794 ( .A(n3931), .Y(n3929) );
  INVX1 U1796 ( .A(n3929), .Y(n3930) );
  AND2X1 U1798 ( .A(n7455), .B(n10500), .Y(n1234) );
  INVX1 U1800 ( .A(n1234), .Y(n3931) );
  INVX1 U1802 ( .A(n3934), .Y(n3932) );
  INVX1 U1804 ( .A(n3932), .Y(n3933) );
  AND2X1 U1806 ( .A(n7458), .B(n10500), .Y(n1233) );
  INVX1 U1808 ( .A(n1233), .Y(n3934) );
  INVX1 U1810 ( .A(n3937), .Y(n3935) );
  INVX1 U1812 ( .A(n3935), .Y(n3936) );
  AND2X1 U1814 ( .A(n7461), .B(n10500), .Y(n1232) );
  INVX1 U1816 ( .A(n1232), .Y(n3937) );
  INVX1 U1818 ( .A(n3940), .Y(n3938) );
  INVX1 U1820 ( .A(n3938), .Y(n3939) );
  AND2X1 U1822 ( .A(n7464), .B(n10500), .Y(n1231) );
  INVX1 U1824 ( .A(n1231), .Y(n3940) );
  INVX1 U1826 ( .A(n3943), .Y(n3941) );
  INVX1 U1828 ( .A(n3941), .Y(n3942) );
  AND2X1 U1830 ( .A(n7467), .B(n10500), .Y(n1230) );
  INVX1 U1832 ( .A(n1230), .Y(n3943) );
  INVX1 U1834 ( .A(n3946), .Y(n3944) );
  INVX1 U1836 ( .A(n3944), .Y(n3945) );
  AND2X1 U1838 ( .A(n7470), .B(n10500), .Y(n1229) );
  INVX1 U1839 ( .A(n1229), .Y(n3946) );
  INVX1 U1842 ( .A(n3949), .Y(n3947) );
  INVX1 U1844 ( .A(n3947), .Y(n3948) );
  AND2X1 U1846 ( .A(n7473), .B(n10500), .Y(n1228) );
  INVX1 U1848 ( .A(n1228), .Y(n3949) );
  INVX1 U1850 ( .A(n3952), .Y(n3950) );
  INVX1 U1852 ( .A(n3950), .Y(n3951) );
  AND2X1 U1854 ( .A(n7476), .B(n10500), .Y(n1227) );
  INVX1 U1856 ( .A(n1227), .Y(n3952) );
  INVX1 U1858 ( .A(n3955), .Y(n3953) );
  INVX1 U1860 ( .A(n3953), .Y(n3954) );
  AND2X1 U1862 ( .A(n7479), .B(n10500), .Y(n1226) );
  INVX1 U1864 ( .A(n1226), .Y(n3955) );
  INVX1 U1866 ( .A(n3958), .Y(n3956) );
  INVX1 U1868 ( .A(n3956), .Y(n3957) );
  AND2X1 U1870 ( .A(n7482), .B(n10500), .Y(n1225) );
  INVX1 U1872 ( .A(n1225), .Y(n3958) );
  INVX1 U1874 ( .A(n3961), .Y(n3959) );
  INVX1 U1876 ( .A(n3959), .Y(n3960) );
  AND2X1 U1878 ( .A(n7485), .B(n10500), .Y(n1224) );
  INVX1 U1880 ( .A(n1224), .Y(n3961) );
  INVX1 U1882 ( .A(n3964), .Y(n3962) );
  INVX1 U1884 ( .A(n3962), .Y(n3963) );
  AND2X1 U1886 ( .A(n7488), .B(n10500), .Y(n1223) );
  INVX1 U1888 ( .A(n1223), .Y(n3964) );
  INVX1 U1890 ( .A(n3967), .Y(n3965) );
  INVX1 U1892 ( .A(n3965), .Y(n3966) );
  AND2X1 U1894 ( .A(n7491), .B(n10500), .Y(n1222) );
  INVX1 U1896 ( .A(n1222), .Y(n3967) );
  INVX1 U1898 ( .A(n3970), .Y(n3968) );
  INVX1 U1900 ( .A(n3968), .Y(n3969) );
  AND2X1 U1902 ( .A(n7494), .B(n10500), .Y(n1221) );
  INVX1 U1904 ( .A(n1221), .Y(n3970) );
  INVX1 U1906 ( .A(n3973), .Y(n3971) );
  INVX1 U1908 ( .A(n3971), .Y(n3972) );
  AND2X1 U1909 ( .A(n7497), .B(n10500), .Y(n1220) );
  INVX1 U1912 ( .A(n1220), .Y(n3973) );
  INVX1 U1914 ( .A(n3976), .Y(n3974) );
  INVX1 U1916 ( .A(n3974), .Y(n3975) );
  AND2X1 U1918 ( .A(n7500), .B(n10500), .Y(n1219) );
  INVX1 U1920 ( .A(n1219), .Y(n3976) );
  INVX1 U1922 ( .A(n3979), .Y(n3977) );
  INVX1 U1924 ( .A(n3977), .Y(n3978) );
  AND2X1 U1926 ( .A(n7503), .B(n10500), .Y(n1218) );
  INVX1 U1928 ( .A(n1218), .Y(n3979) );
  INVX1 U1930 ( .A(n3982), .Y(n3980) );
  INVX1 U1932 ( .A(n3980), .Y(n3981) );
  AND2X1 U1934 ( .A(n7506), .B(n10500), .Y(n1217) );
  INVX1 U1936 ( .A(n1217), .Y(n3982) );
  INVX1 U1938 ( .A(n3985), .Y(n3983) );
  INVX1 U1940 ( .A(n3983), .Y(n3984) );
  AND2X1 U1942 ( .A(n7509), .B(n10500), .Y(n1216) );
  INVX1 U1944 ( .A(n1216), .Y(n3985) );
  INVX1 U1946 ( .A(n3988), .Y(n3986) );
  INVX1 U1948 ( .A(n3986), .Y(n3987) );
  AND2X1 U1950 ( .A(n7512), .B(n10500), .Y(n1215) );
  INVX1 U1952 ( .A(n1215), .Y(n3988) );
  INVX1 U1954 ( .A(n3991), .Y(n3989) );
  INVX1 U1956 ( .A(n3989), .Y(n3990) );
  AND2X1 U1958 ( .A(n7515), .B(n10500), .Y(n1214) );
  INVX1 U1960 ( .A(n1214), .Y(n3991) );
  INVX1 U1962 ( .A(n3994), .Y(n3992) );
  INVX1 U1964 ( .A(n3992), .Y(n3993) );
  AND2X1 U1966 ( .A(n9048), .B(n1178), .Y(n1212) );
  INVX1 U1968 ( .A(n1212), .Y(n3994) );
  INVX1 U1970 ( .A(n3997), .Y(n3995) );
  INVX1 U1972 ( .A(n3995), .Y(n3996) );
  AND2X1 U1974 ( .A(n9051), .B(n1178), .Y(n1211) );
  INVX1 U1976 ( .A(n1211), .Y(n3997) );
  INVX1 U1978 ( .A(n4000), .Y(n3998) );
  INVX1 U1979 ( .A(n3998), .Y(n3999) );
  AND2X1 U1980 ( .A(n9054), .B(n1178), .Y(n1210) );
  INVX1 U1982 ( .A(n1210), .Y(n4000) );
  INVX1 U1984 ( .A(n4003), .Y(n4001) );
  INVX1 U1986 ( .A(n4001), .Y(n4002) );
  AND2X1 U1988 ( .A(n9057), .B(n1178), .Y(n1209) );
  INVX1 U1990 ( .A(n1209), .Y(n4003) );
  INVX1 U1992 ( .A(n4006), .Y(n4004) );
  INVX1 U1994 ( .A(n4004), .Y(n4005) );
  AND2X1 U1996 ( .A(n9060), .B(n1178), .Y(n1208) );
  INVX1 U1998 ( .A(n1208), .Y(n4006) );
  INVX1 U2000 ( .A(n4009), .Y(n4007) );
  INVX1 U2002 ( .A(n4007), .Y(n4008) );
  AND2X1 U2004 ( .A(n9063), .B(n1178), .Y(n1207) );
  INVX1 U2006 ( .A(n1207), .Y(n4009) );
  INVX1 U2008 ( .A(n4012), .Y(n4010) );
  INVX1 U2010 ( .A(n4010), .Y(n4011) );
  AND2X1 U2012 ( .A(n9066), .B(n1178), .Y(n1206) );
  INVX1 U2014 ( .A(n1206), .Y(n4012) );
  INVX1 U2016 ( .A(n4015), .Y(n4013) );
  INVX1 U2018 ( .A(n4013), .Y(n4014) );
  AND2X1 U2020 ( .A(n9069), .B(n1178), .Y(n1205) );
  INVX1 U2022 ( .A(n1205), .Y(n4015) );
  INVX1 U2024 ( .A(n4018), .Y(n4016) );
  INVX1 U2026 ( .A(n4016), .Y(n4017) );
  AND2X1 U2028 ( .A(n9072), .B(n1178), .Y(n1204) );
  INVX1 U2030 ( .A(n1204), .Y(n4018) );
  INVX1 U2032 ( .A(n4021), .Y(n4019) );
  INVX1 U2034 ( .A(n4019), .Y(n4020) );
  AND2X1 U2036 ( .A(n9075), .B(n1178), .Y(n1203) );
  INVX1 U2038 ( .A(n1203), .Y(n4021) );
  INVX1 U2040 ( .A(n4024), .Y(n4022) );
  INVX1 U2042 ( .A(n4022), .Y(n4023) );
  AND2X1 U2044 ( .A(n9078), .B(n1178), .Y(n1202) );
  INVX1 U2046 ( .A(n1202), .Y(n4024) );
  INVX1 U2048 ( .A(n4027), .Y(n4025) );
  INVX1 U2049 ( .A(n4025), .Y(n4026) );
  AND2X1 U2050 ( .A(n9081), .B(n1178), .Y(n1201) );
  INVX1 U2052 ( .A(n1201), .Y(n4027) );
  INVX1 U2054 ( .A(n4030), .Y(n4028) );
  INVX1 U2056 ( .A(n4028), .Y(n4029) );
  AND2X1 U2058 ( .A(n9084), .B(n1178), .Y(n1200) );
  INVX1 U2060 ( .A(n1200), .Y(n4030) );
  INVX1 U2062 ( .A(n4033), .Y(n4031) );
  INVX1 U2064 ( .A(n4031), .Y(n4032) );
  AND2X1 U2066 ( .A(n9087), .B(n1178), .Y(n1199) );
  INVX1 U2068 ( .A(n1199), .Y(n4033) );
  INVX1 U2070 ( .A(n4036), .Y(n4034) );
  INVX1 U2072 ( .A(n4034), .Y(n4035) );
  AND2X1 U2074 ( .A(n9090), .B(n1178), .Y(n1198) );
  INVX1 U2076 ( .A(n1198), .Y(n4036) );
  INVX1 U2078 ( .A(n4039), .Y(n4037) );
  INVX1 U2080 ( .A(n4037), .Y(n4038) );
  AND2X1 U2082 ( .A(n9093), .B(n1178), .Y(n1197) );
  INVX1 U2084 ( .A(n1197), .Y(n4039) );
  INVX1 U2086 ( .A(n4042), .Y(n4040) );
  INVX1 U2088 ( .A(n4040), .Y(n4041) );
  AND2X1 U2090 ( .A(n9096), .B(n1178), .Y(n1196) );
  INVX1 U2092 ( .A(n1196), .Y(n4042) );
  INVX1 U2094 ( .A(n4045), .Y(n4043) );
  INVX1 U2096 ( .A(n4043), .Y(n4044) );
  AND2X1 U2098 ( .A(n9099), .B(n1178), .Y(n1195) );
  INVX1 U2100 ( .A(n1195), .Y(n4045) );
  INVX1 U2102 ( .A(n4048), .Y(n4046) );
  INVX1 U2104 ( .A(n4046), .Y(n4047) );
  AND2X1 U2106 ( .A(n9102), .B(n1178), .Y(n1194) );
  INVX1 U2108 ( .A(n1194), .Y(n4048) );
  INVX1 U2110 ( .A(n4051), .Y(n4049) );
  INVX1 U2112 ( .A(n4049), .Y(n4050) );
  AND2X1 U2114 ( .A(n9105), .B(n1178), .Y(n1193) );
  INVX1 U2116 ( .A(n1193), .Y(n4051) );
  INVX1 U2118 ( .A(n4054), .Y(n4052) );
  INVX1 U2119 ( .A(n4052), .Y(n4053) );
  AND2X1 U2120 ( .A(n9108), .B(n1178), .Y(n1192) );
  INVX1 U2122 ( .A(n1192), .Y(n4054) );
  INVX1 U2124 ( .A(n4057), .Y(n4055) );
  INVX1 U2126 ( .A(n4055), .Y(n4056) );
  AND2X1 U2128 ( .A(n9111), .B(n1178), .Y(n1191) );
  INVX1 U2130 ( .A(n1191), .Y(n4057) );
  INVX1 U2132 ( .A(n4060), .Y(n4058) );
  INVX1 U2134 ( .A(n4058), .Y(n4059) );
  AND2X1 U2136 ( .A(n9114), .B(n1178), .Y(n1190) );
  INVX1 U2138 ( .A(n1190), .Y(n4060) );
  INVX1 U2140 ( .A(n4063), .Y(n4061) );
  INVX1 U2142 ( .A(n4061), .Y(n4062) );
  AND2X1 U2144 ( .A(n9117), .B(n1178), .Y(n1189) );
  INVX1 U2146 ( .A(n1189), .Y(n4063) );
  INVX1 U2148 ( .A(n4066), .Y(n4064) );
  INVX1 U2150 ( .A(n4064), .Y(n4065) );
  AND2X1 U2152 ( .A(n9120), .B(n1178), .Y(n1188) );
  INVX1 U2154 ( .A(n1188), .Y(n4066) );
  INVX1 U2156 ( .A(n4069), .Y(n4067) );
  INVX1 U2158 ( .A(n4067), .Y(n4068) );
  AND2X1 U2160 ( .A(n9123), .B(n1178), .Y(n1187) );
  INVX1 U2162 ( .A(n1187), .Y(n4069) );
  INVX1 U2164 ( .A(n4072), .Y(n4070) );
  INVX1 U2166 ( .A(n4070), .Y(n4071) );
  AND2X1 U2168 ( .A(n9126), .B(n1178), .Y(n1186) );
  INVX1 U2170 ( .A(n1186), .Y(n4072) );
  INVX1 U2172 ( .A(n4075), .Y(n4073) );
  INVX1 U2174 ( .A(n4073), .Y(n4074) );
  AND2X1 U2176 ( .A(n9129), .B(n1178), .Y(n1185) );
  INVX1 U2178 ( .A(n1185), .Y(n4075) );
  INVX1 U2180 ( .A(n4078), .Y(n4076) );
  INVX1 U2182 ( .A(n4076), .Y(n4077) );
  AND2X1 U2184 ( .A(n9132), .B(n1178), .Y(n1184) );
  INVX1 U2186 ( .A(n1184), .Y(n4078) );
  INVX1 U2188 ( .A(n4081), .Y(n4079) );
  INVX1 U2189 ( .A(n4079), .Y(n4080) );
  AND2X1 U2190 ( .A(n9135), .B(n1178), .Y(n1183) );
  INVX1 U2192 ( .A(n1183), .Y(n4081) );
  INVX1 U2194 ( .A(n4084), .Y(n4082) );
  INVX1 U2196 ( .A(n4082), .Y(n4083) );
  AND2X1 U2198 ( .A(n9138), .B(n1178), .Y(n1182) );
  INVX1 U2200 ( .A(n1182), .Y(n4084) );
  INVX1 U2202 ( .A(n4087), .Y(n4085) );
  INVX1 U2204 ( .A(n4085), .Y(n4086) );
  AND2X1 U2206 ( .A(n9141), .B(n1178), .Y(n1181) );
  INVX1 U2208 ( .A(n1181), .Y(n4087) );
  INVX1 U2210 ( .A(n4090), .Y(n4088) );
  INVX1 U2212 ( .A(n4088), .Y(n4089) );
  AND2X1 U2214 ( .A(n9144), .B(n1178), .Y(n1180) );
  INVX1 U2216 ( .A(n1180), .Y(n4090) );
  INVX1 U2218 ( .A(n4093), .Y(n4091) );
  INVX1 U2220 ( .A(n4091), .Y(n4092) );
  AND2X1 U2222 ( .A(n9147), .B(n1178), .Y(n1179) );
  INVX1 U2224 ( .A(n1179), .Y(n4093) );
  INVX1 U2226 ( .A(n4096), .Y(n4094) );
  INVX1 U2228 ( .A(n4094), .Y(n4095) );
  AND2X1 U2230 ( .A(n7518), .B(n1142), .Y(n1176) );
  INVX1 U2232 ( .A(n1176), .Y(n4096) );
  INVX1 U2234 ( .A(n4099), .Y(n4097) );
  INVX1 U2236 ( .A(n4097), .Y(n4098) );
  AND2X1 U2238 ( .A(n7521), .B(n1142), .Y(n1175) );
  INVX1 U2240 ( .A(n1175), .Y(n4099) );
  INVX1 U2242 ( .A(n4102), .Y(n4100) );
  INVX1 U2244 ( .A(n4100), .Y(n4101) );
  AND2X1 U2246 ( .A(n7524), .B(n1142), .Y(n1174) );
  INVX1 U2248 ( .A(n1174), .Y(n4102) );
  INVX1 U2250 ( .A(n4105), .Y(n4103) );
  INVX1 U2252 ( .A(n4103), .Y(n4104) );
  AND2X1 U2254 ( .A(n7527), .B(n1142), .Y(n1173) );
  INVX1 U2256 ( .A(n1173), .Y(n4105) );
  INVX1 U2258 ( .A(n4108), .Y(n4106) );
  INVX1 U2259 ( .A(n4106), .Y(n4107) );
  AND2X1 U2262 ( .A(n7530), .B(n1142), .Y(n1172) );
  INVX1 U2265 ( .A(n1172), .Y(n4108) );
  INVX1 U2268 ( .A(n4111), .Y(n4109) );
  INVX1 U2271 ( .A(n4109), .Y(n4110) );
  AND2X1 U2274 ( .A(n7533), .B(n1142), .Y(n1171) );
  INVX1 U2277 ( .A(n1171), .Y(n4111) );
  INVX1 U2280 ( .A(n4114), .Y(n4112) );
  INVX1 U2283 ( .A(n4112), .Y(n4113) );
  AND2X1 U2286 ( .A(n7536), .B(n1142), .Y(n1170) );
  INVX1 U2289 ( .A(n1170), .Y(n4114) );
  INVX1 U2292 ( .A(n4117), .Y(n4115) );
  INVX1 U2295 ( .A(n4115), .Y(n4116) );
  AND2X1 U2298 ( .A(n7539), .B(n1142), .Y(n1169) );
  INVX1 U2301 ( .A(n1169), .Y(n4117) );
  INVX1 U2304 ( .A(n4120), .Y(n4118) );
  INVX1 U2307 ( .A(n4118), .Y(n4119) );
  AND2X1 U2310 ( .A(n7542), .B(n1142), .Y(n1168) );
  INVX1 U2313 ( .A(n1168), .Y(n4120) );
  INVX1 U2316 ( .A(n4123), .Y(n4121) );
  INVX1 U2319 ( .A(n4121), .Y(n4122) );
  AND2X1 U2322 ( .A(n7545), .B(n1142), .Y(n1167) );
  INVX1 U2325 ( .A(n1167), .Y(n4123) );
  INVX1 U2328 ( .A(n4126), .Y(n4124) );
  INVX1 U2331 ( .A(n4124), .Y(n4125) );
  AND2X1 U2334 ( .A(n7548), .B(n1142), .Y(n1166) );
  INVX1 U2337 ( .A(n1166), .Y(n4126) );
  INVX1 U2340 ( .A(n4129), .Y(n4127) );
  INVX1 U2343 ( .A(n4127), .Y(n4128) );
  AND2X1 U2346 ( .A(n7551), .B(n1142), .Y(n1165) );
  INVX1 U2349 ( .A(n1165), .Y(n4129) );
  INVX1 U2352 ( .A(n4132), .Y(n4130) );
  INVX1 U2355 ( .A(n4130), .Y(n4131) );
  AND2X1 U2358 ( .A(n7554), .B(n1142), .Y(n1164) );
  INVX1 U2361 ( .A(n1164), .Y(n4132) );
  INVX1 U2362 ( .A(n4135), .Y(n4133) );
  INVX1 U2365 ( .A(n4133), .Y(n4134) );
  AND2X1 U2367 ( .A(n7557), .B(n1142), .Y(n1163) );
  INVX1 U2370 ( .A(n1163), .Y(n4135) );
  INVX1 U2371 ( .A(n4138), .Y(n4136) );
  INVX1 U2373 ( .A(n4136), .Y(n4137) );
  AND2X1 U2385 ( .A(n7560), .B(n1142), .Y(n1162) );
  INVX1 U2387 ( .A(n1162), .Y(n4138) );
  INVX1 U2388 ( .A(n4141), .Y(n4139) );
  INVX1 U2389 ( .A(n4139), .Y(n4140) );
  AND2X1 U2395 ( .A(n7563), .B(n1142), .Y(n1161) );
  INVX1 U2396 ( .A(n1161), .Y(n4141) );
  INVX1 U2398 ( .A(n4144), .Y(n4142) );
  INVX1 U2403 ( .A(n4142), .Y(n4143) );
  AND2X1 U2679 ( .A(n7566), .B(n1142), .Y(n1160) );
  INVX1 U2680 ( .A(n1160), .Y(n4144) );
  INVX1 U2681 ( .A(n4147), .Y(n4145) );
  INVX1 U2682 ( .A(n4145), .Y(n4146) );
  AND2X1 U2683 ( .A(n7569), .B(n1142), .Y(n1159) );
  INVX1 U2684 ( .A(n1159), .Y(n4147) );
  INVX1 U2685 ( .A(n4150), .Y(n4148) );
  INVX1 U2686 ( .A(n4148), .Y(n4149) );
  AND2X1 U2687 ( .A(n7572), .B(n1142), .Y(n1158) );
  INVX1 U2688 ( .A(n1158), .Y(n4150) );
  INVX1 U2689 ( .A(n4153), .Y(n4151) );
  INVX1 U2690 ( .A(n4151), .Y(n4152) );
  AND2X1 U2691 ( .A(n7575), .B(n1142), .Y(n1157) );
  INVX1 U2692 ( .A(n1157), .Y(n4153) );
  INVX1 U2693 ( .A(n4156), .Y(n4154) );
  INVX1 U2694 ( .A(n4154), .Y(n4155) );
  AND2X1 U2695 ( .A(n7578), .B(n1142), .Y(n1156) );
  INVX1 U2696 ( .A(n1156), .Y(n4156) );
  INVX1 U2697 ( .A(n4159), .Y(n4157) );
  INVX1 U2698 ( .A(n4157), .Y(n4158) );
  AND2X1 U2699 ( .A(n7581), .B(n1142), .Y(n1155) );
  INVX1 U2700 ( .A(n1155), .Y(n4159) );
  INVX1 U2701 ( .A(n4162), .Y(n4160) );
  INVX1 U2702 ( .A(n4160), .Y(n4161) );
  AND2X1 U2703 ( .A(n7584), .B(n1142), .Y(n1154) );
  INVX1 U2704 ( .A(n1154), .Y(n4162) );
  INVX1 U2705 ( .A(n4165), .Y(n4163) );
  INVX1 U2706 ( .A(n4163), .Y(n4164) );
  AND2X1 U2707 ( .A(n7587), .B(n1142), .Y(n1153) );
  INVX1 U2708 ( .A(n1153), .Y(n4165) );
  INVX1 U2709 ( .A(n4168), .Y(n4166) );
  INVX1 U2710 ( .A(n4166), .Y(n4167) );
  AND2X1 U2711 ( .A(n7590), .B(n1142), .Y(n1152) );
  INVX1 U2712 ( .A(n1152), .Y(n4168) );
  INVX1 U2713 ( .A(n4171), .Y(n4169) );
  INVX1 U2714 ( .A(n4169), .Y(n4170) );
  AND2X1 U2715 ( .A(n7593), .B(n1142), .Y(n1151) );
  INVX1 U2716 ( .A(n1151), .Y(n4171) );
  INVX1 U2717 ( .A(n4174), .Y(n4172) );
  INVX1 U2718 ( .A(n4172), .Y(n4173) );
  AND2X1 U2719 ( .A(n7596), .B(n1142), .Y(n1150) );
  INVX1 U2720 ( .A(n1150), .Y(n4174) );
  INVX1 U2721 ( .A(n4177), .Y(n4175) );
  INVX1 U2722 ( .A(n4175), .Y(n4176) );
  AND2X1 U2723 ( .A(n7599), .B(n1142), .Y(n1149) );
  INVX1 U2724 ( .A(n1149), .Y(n4177) );
  INVX1 U2725 ( .A(n4180), .Y(n4178) );
  INVX1 U2726 ( .A(n4178), .Y(n4179) );
  AND2X1 U2727 ( .A(n7602), .B(n1142), .Y(n1148) );
  INVX1 U2728 ( .A(n1148), .Y(n4180) );
  INVX1 U2729 ( .A(n4183), .Y(n4181) );
  INVX1 U2730 ( .A(n4181), .Y(n4182) );
  AND2X1 U2731 ( .A(n7605), .B(n1142), .Y(n1147) );
  INVX1 U2732 ( .A(n1147), .Y(n4183) );
  INVX1 U2733 ( .A(n4186), .Y(n4184) );
  INVX1 U2734 ( .A(n4184), .Y(n4185) );
  AND2X1 U2735 ( .A(n7608), .B(n1142), .Y(n1146) );
  INVX1 U2736 ( .A(n1146), .Y(n4186) );
  INVX1 U2737 ( .A(n4189), .Y(n4187) );
  INVX1 U2738 ( .A(n4187), .Y(n4188) );
  AND2X1 U2739 ( .A(n7611), .B(n1142), .Y(n1145) );
  INVX1 U2740 ( .A(n1145), .Y(n4189) );
  INVX1 U2741 ( .A(n4192), .Y(n4190) );
  INVX1 U2742 ( .A(n4190), .Y(n4191) );
  AND2X1 U2743 ( .A(n7614), .B(n1142), .Y(n1144) );
  INVX1 U2744 ( .A(n1144), .Y(n4192) );
  INVX1 U2745 ( .A(n4195), .Y(n4193) );
  INVX1 U2746 ( .A(n4193), .Y(n4194) );
  AND2X1 U2747 ( .A(n7617), .B(n1142), .Y(n1143) );
  INVX1 U2748 ( .A(n1143), .Y(n4195) );
  INVX1 U2749 ( .A(n4198), .Y(n4196) );
  INVX1 U2750 ( .A(n4196), .Y(n4197) );
  AND2X1 U2751 ( .A(n8538), .B(n10116), .Y(n1140) );
  INVX1 U2752 ( .A(n1140), .Y(n4198) );
  INVX1 U2753 ( .A(n4201), .Y(n4199) );
  INVX1 U2754 ( .A(n4199), .Y(n4200) );
  AND2X1 U2755 ( .A(n8541), .B(n10116), .Y(n1139) );
  INVX1 U2756 ( .A(n1139), .Y(n4201) );
  INVX1 U2757 ( .A(n4204), .Y(n4202) );
  INVX1 U2758 ( .A(n4202), .Y(n4203) );
  AND2X1 U2759 ( .A(n8544), .B(n10116), .Y(n1138) );
  INVX1 U2760 ( .A(n1138), .Y(n4204) );
  INVX1 U2761 ( .A(n4207), .Y(n4205) );
  INVX1 U2762 ( .A(n4205), .Y(n4206) );
  AND2X1 U2763 ( .A(n8547), .B(n10116), .Y(n1137) );
  INVX1 U2764 ( .A(n1137), .Y(n4207) );
  INVX1 U2765 ( .A(n4210), .Y(n4208) );
  INVX1 U2766 ( .A(n4208), .Y(n4209) );
  AND2X1 U2767 ( .A(n8550), .B(n10116), .Y(n1136) );
  INVX1 U2768 ( .A(n1136), .Y(n4210) );
  INVX1 U2769 ( .A(n4213), .Y(n4211) );
  INVX1 U2770 ( .A(n4211), .Y(n4212) );
  AND2X1 U2771 ( .A(n8553), .B(n10116), .Y(n1135) );
  INVX1 U2772 ( .A(n1135), .Y(n4213) );
  INVX1 U2773 ( .A(n4216), .Y(n4214) );
  INVX1 U2774 ( .A(n4214), .Y(n4215) );
  AND2X1 U2775 ( .A(n8556), .B(n10116), .Y(n1134) );
  INVX1 U2776 ( .A(n1134), .Y(n4216) );
  INVX1 U2777 ( .A(n4219), .Y(n4217) );
  INVX1 U2778 ( .A(n4217), .Y(n4218) );
  AND2X1 U2779 ( .A(n8559), .B(n10116), .Y(n1133) );
  INVX1 U2780 ( .A(n1133), .Y(n4219) );
  INVX1 U2781 ( .A(n4222), .Y(n4220) );
  INVX1 U2782 ( .A(n4220), .Y(n4221) );
  AND2X1 U2783 ( .A(n8562), .B(n10116), .Y(n1132) );
  INVX1 U2784 ( .A(n1132), .Y(n4222) );
  INVX1 U2785 ( .A(n4225), .Y(n4223) );
  INVX1 U2786 ( .A(n4223), .Y(n4224) );
  AND2X1 U2787 ( .A(n8565), .B(n10116), .Y(n1131) );
  INVX1 U2788 ( .A(n1131), .Y(n4225) );
  INVX1 U2789 ( .A(n4228), .Y(n4226) );
  INVX1 U2790 ( .A(n4226), .Y(n4227) );
  AND2X1 U2791 ( .A(n8568), .B(n10116), .Y(n1130) );
  INVX1 U2792 ( .A(n1130), .Y(n4228) );
  INVX1 U2793 ( .A(n4231), .Y(n4229) );
  INVX1 U2794 ( .A(n4229), .Y(n4230) );
  AND2X1 U2795 ( .A(n8571), .B(n10116), .Y(n1129) );
  INVX1 U2796 ( .A(n1129), .Y(n4231) );
  INVX1 U2797 ( .A(n4234), .Y(n4232) );
  INVX1 U2798 ( .A(n4232), .Y(n4233) );
  AND2X1 U2799 ( .A(n8574), .B(n10116), .Y(n1128) );
  INVX1 U2800 ( .A(n1128), .Y(n4234) );
  INVX1 U2801 ( .A(n4237), .Y(n4235) );
  INVX1 U2802 ( .A(n4235), .Y(n4236) );
  AND2X1 U2803 ( .A(n8577), .B(n10116), .Y(n1127) );
  INVX1 U2804 ( .A(n1127), .Y(n4237) );
  INVX1 U2805 ( .A(n4240), .Y(n4238) );
  INVX1 U2806 ( .A(n4238), .Y(n4239) );
  AND2X1 U2807 ( .A(n8580), .B(n10116), .Y(n1126) );
  INVX1 U2808 ( .A(n1126), .Y(n4240) );
  INVX1 U2809 ( .A(n4243), .Y(n4241) );
  INVX1 U2810 ( .A(n4241), .Y(n4242) );
  AND2X1 U2811 ( .A(n8583), .B(n10116), .Y(n1125) );
  INVX1 U2812 ( .A(n1125), .Y(n4243) );
  INVX1 U2813 ( .A(n4246), .Y(n4244) );
  INVX1 U2814 ( .A(n4244), .Y(n4245) );
  AND2X1 U2815 ( .A(n8586), .B(n10116), .Y(n1124) );
  INVX1 U2816 ( .A(n1124), .Y(n4246) );
  INVX1 U2817 ( .A(n4249), .Y(n4247) );
  INVX1 U2818 ( .A(n4247), .Y(n4248) );
  AND2X1 U2819 ( .A(n8589), .B(n10116), .Y(n1123) );
  INVX1 U2820 ( .A(n1123), .Y(n4249) );
  INVX1 U2821 ( .A(n4252), .Y(n4250) );
  INVX1 U2822 ( .A(n4250), .Y(n4251) );
  AND2X1 U2823 ( .A(n8592), .B(n10116), .Y(n1122) );
  INVX1 U2824 ( .A(n1122), .Y(n4252) );
  INVX1 U2825 ( .A(n4255), .Y(n4253) );
  INVX1 U2826 ( .A(n4253), .Y(n4254) );
  AND2X1 U2827 ( .A(n8595), .B(n10116), .Y(n1121) );
  INVX1 U2828 ( .A(n1121), .Y(n4255) );
  INVX1 U2829 ( .A(n4258), .Y(n4256) );
  INVX1 U2830 ( .A(n4256), .Y(n4257) );
  AND2X1 U2831 ( .A(n8598), .B(n10116), .Y(n1120) );
  INVX1 U2832 ( .A(n1120), .Y(n4258) );
  INVX1 U2833 ( .A(n4261), .Y(n4259) );
  INVX1 U2834 ( .A(n4259), .Y(n4260) );
  AND2X1 U2835 ( .A(n8601), .B(n10116), .Y(n1119) );
  INVX1 U2836 ( .A(n1119), .Y(n4261) );
  INVX1 U2837 ( .A(n4264), .Y(n4262) );
  INVX1 U2838 ( .A(n4262), .Y(n4263) );
  AND2X1 U2839 ( .A(n8604), .B(n10116), .Y(n1118) );
  INVX1 U2840 ( .A(n1118), .Y(n4264) );
  INVX1 U2841 ( .A(n4267), .Y(n4265) );
  INVX1 U2842 ( .A(n4265), .Y(n4266) );
  AND2X1 U2843 ( .A(n8607), .B(n10116), .Y(n1117) );
  INVX1 U2844 ( .A(n1117), .Y(n4267) );
  INVX1 U2845 ( .A(n4270), .Y(n4268) );
  INVX1 U2846 ( .A(n4268), .Y(n4269) );
  AND2X1 U2847 ( .A(n8610), .B(n10116), .Y(n1116) );
  INVX1 U2848 ( .A(n1116), .Y(n4270) );
  INVX1 U2849 ( .A(n4273), .Y(n4271) );
  INVX1 U2850 ( .A(n4271), .Y(n4272) );
  AND2X1 U2851 ( .A(n8613), .B(n10116), .Y(n1115) );
  INVX1 U2852 ( .A(n1115), .Y(n4273) );
  INVX1 U2853 ( .A(n4276), .Y(n4274) );
  INVX1 U2854 ( .A(n4274), .Y(n4275) );
  AND2X1 U2855 ( .A(n8616), .B(n10116), .Y(n1114) );
  INVX1 U2856 ( .A(n1114), .Y(n4276) );
  INVX1 U2857 ( .A(n4279), .Y(n4277) );
  INVX1 U2858 ( .A(n4277), .Y(n4278) );
  AND2X1 U2859 ( .A(n8619), .B(n10116), .Y(n1113) );
  INVX1 U2860 ( .A(n1113), .Y(n4279) );
  INVX1 U2861 ( .A(n4282), .Y(n4280) );
  INVX1 U2862 ( .A(n4280), .Y(n4281) );
  AND2X1 U2863 ( .A(n8622), .B(n10116), .Y(n1112) );
  INVX1 U2864 ( .A(n1112), .Y(n4282) );
  INVX1 U2865 ( .A(n4285), .Y(n4283) );
  INVX1 U2866 ( .A(n4283), .Y(n4284) );
  AND2X1 U2867 ( .A(n8625), .B(n10116), .Y(n1111) );
  INVX1 U2868 ( .A(n1111), .Y(n4285) );
  INVX1 U2869 ( .A(n4288), .Y(n4286) );
  INVX1 U2870 ( .A(n4286), .Y(n4287) );
  AND2X1 U2871 ( .A(n8628), .B(n10116), .Y(n1110) );
  INVX1 U2872 ( .A(n1110), .Y(n4288) );
  INVX1 U2873 ( .A(n4291), .Y(n4289) );
  INVX1 U2874 ( .A(n4289), .Y(n4290) );
  AND2X1 U2875 ( .A(n8631), .B(n10116), .Y(n1109) );
  INVX1 U2876 ( .A(n1109), .Y(n4291) );
  INVX1 U2877 ( .A(n4294), .Y(n4292) );
  INVX1 U2878 ( .A(n4292), .Y(n4293) );
  AND2X1 U2879 ( .A(n8634), .B(n10116), .Y(n1108) );
  INVX1 U2880 ( .A(n1108), .Y(n4294) );
  INVX1 U2881 ( .A(n4297), .Y(n4295) );
  INVX1 U2882 ( .A(n4295), .Y(n4296) );
  AND2X1 U2883 ( .A(n8637), .B(n10116), .Y(n1107) );
  INVX1 U2884 ( .A(n1107), .Y(n4297) );
  INVX1 U2885 ( .A(n4300), .Y(n4298) );
  INVX1 U2886 ( .A(n4298), .Y(n4299) );
  AND2X1 U2887 ( .A(n6906), .B(n10119), .Y(n1105) );
  INVX1 U2888 ( .A(n1105), .Y(n4300) );
  INVX1 U2889 ( .A(n4303), .Y(n4301) );
  INVX1 U2890 ( .A(n4301), .Y(n4302) );
  AND2X1 U2891 ( .A(n6909), .B(n10119), .Y(n1104) );
  INVX1 U2892 ( .A(n1104), .Y(n4303) );
  INVX1 U2893 ( .A(n4306), .Y(n4304) );
  INVX1 U2894 ( .A(n4304), .Y(n4305) );
  AND2X1 U2895 ( .A(n6912), .B(n10119), .Y(n1103) );
  INVX1 U2896 ( .A(n1103), .Y(n4306) );
  INVX1 U2897 ( .A(n4309), .Y(n4307) );
  INVX1 U2898 ( .A(n4307), .Y(n4308) );
  AND2X1 U2899 ( .A(n6915), .B(n10119), .Y(n1102) );
  INVX1 U2900 ( .A(n1102), .Y(n4309) );
  INVX1 U2901 ( .A(n4312), .Y(n4310) );
  INVX1 U2902 ( .A(n4310), .Y(n4311) );
  AND2X1 U2903 ( .A(n6918), .B(n10119), .Y(n1101) );
  INVX1 U2904 ( .A(n1101), .Y(n4312) );
  INVX1 U2905 ( .A(n4315), .Y(n4313) );
  INVX1 U2906 ( .A(n4313), .Y(n4314) );
  AND2X1 U2907 ( .A(n6921), .B(n10119), .Y(n1100) );
  INVX1 U2908 ( .A(n1100), .Y(n4315) );
  INVX1 U2909 ( .A(n4318), .Y(n4316) );
  INVX1 U2910 ( .A(n4316), .Y(n4317) );
  AND2X1 U2911 ( .A(n6924), .B(n10119), .Y(n1099) );
  INVX1 U2912 ( .A(n1099), .Y(n4318) );
  INVX1 U2913 ( .A(n4321), .Y(n4319) );
  INVX1 U2914 ( .A(n4319), .Y(n4320) );
  AND2X1 U2915 ( .A(n6927), .B(n10119), .Y(n1098) );
  INVX1 U2916 ( .A(n1098), .Y(n4321) );
  INVX1 U2917 ( .A(n4324), .Y(n4322) );
  INVX1 U2918 ( .A(n4322), .Y(n4323) );
  AND2X1 U2919 ( .A(n6930), .B(n10119), .Y(n1097) );
  INVX1 U2920 ( .A(n1097), .Y(n4324) );
  INVX1 U2921 ( .A(n4327), .Y(n4325) );
  INVX1 U2922 ( .A(n4325), .Y(n4326) );
  AND2X1 U2923 ( .A(n6933), .B(n10119), .Y(n1096) );
  INVX1 U2924 ( .A(n1096), .Y(n4327) );
  INVX1 U2925 ( .A(n4330), .Y(n4328) );
  INVX1 U2926 ( .A(n4328), .Y(n4329) );
  AND2X1 U2927 ( .A(n6936), .B(n10119), .Y(n1095) );
  INVX1 U2928 ( .A(n1095), .Y(n4330) );
  INVX1 U2929 ( .A(n4333), .Y(n4331) );
  INVX1 U2930 ( .A(n4331), .Y(n4332) );
  AND2X1 U2931 ( .A(n6939), .B(n10119), .Y(n1094) );
  INVX1 U2932 ( .A(n1094), .Y(n4333) );
  INVX1 U2933 ( .A(n4336), .Y(n4334) );
  INVX1 U2934 ( .A(n4334), .Y(n4335) );
  AND2X1 U2935 ( .A(n6942), .B(n10119), .Y(n1093) );
  INVX1 U2936 ( .A(n1093), .Y(n4336) );
  INVX1 U2937 ( .A(n4339), .Y(n4337) );
  INVX1 U2938 ( .A(n4337), .Y(n4338) );
  AND2X1 U2939 ( .A(n6945), .B(n10119), .Y(n1092) );
  INVX1 U2940 ( .A(n1092), .Y(n4339) );
  INVX1 U2941 ( .A(n4342), .Y(n4340) );
  INVX1 U2942 ( .A(n4340), .Y(n4341) );
  AND2X1 U2943 ( .A(n6948), .B(n10119), .Y(n1091) );
  INVX1 U2944 ( .A(n1091), .Y(n4342) );
  INVX1 U2945 ( .A(n4345), .Y(n4343) );
  INVX1 U2946 ( .A(n4343), .Y(n4344) );
  AND2X1 U2947 ( .A(n6951), .B(n10119), .Y(n1090) );
  INVX1 U2948 ( .A(n1090), .Y(n4345) );
  INVX1 U2949 ( .A(n4348), .Y(n4346) );
  INVX1 U2950 ( .A(n4346), .Y(n4347) );
  AND2X1 U3461 ( .A(n6954), .B(n10119), .Y(n1089) );
  INVX1 U3462 ( .A(n1089), .Y(n4348) );
  INVX1 U3463 ( .A(n4351), .Y(n4349) );
  INVX1 U3464 ( .A(n4349), .Y(n4350) );
  AND2X1 U3465 ( .A(n6957), .B(n10119), .Y(n1088) );
  INVX1 U3466 ( .A(n1088), .Y(n4351) );
  INVX1 U3467 ( .A(n4354), .Y(n4352) );
  INVX1 U3468 ( .A(n4352), .Y(n4353) );
  AND2X1 U3469 ( .A(n6960), .B(n10119), .Y(n1087) );
  INVX1 U3470 ( .A(n1087), .Y(n4354) );
  INVX1 U3471 ( .A(n4357), .Y(n4355) );
  INVX1 U3472 ( .A(n4355), .Y(n4356) );
  AND2X1 U3473 ( .A(n6963), .B(n10119), .Y(n1086) );
  INVX1 U3474 ( .A(n1086), .Y(n4357) );
  INVX1 U3475 ( .A(n4360), .Y(n4358) );
  INVX1 U3476 ( .A(n4358), .Y(n4359) );
  AND2X1 U3477 ( .A(n6966), .B(n10119), .Y(n1085) );
  INVX1 U3478 ( .A(n1085), .Y(n4360) );
  INVX1 U3479 ( .A(n4363), .Y(n4361) );
  INVX1 U3480 ( .A(n4361), .Y(n4362) );
  AND2X1 U3481 ( .A(n6969), .B(n10119), .Y(n1084) );
  INVX1 U3482 ( .A(n1084), .Y(n4363) );
  INVX1 U3483 ( .A(n4366), .Y(n4364) );
  INVX1 U3484 ( .A(n4364), .Y(n4365) );
  AND2X1 U3485 ( .A(n6972), .B(n10119), .Y(n1083) );
  INVX1 U3486 ( .A(n1083), .Y(n4366) );
  INVX1 U3487 ( .A(n4369), .Y(n4367) );
  INVX1 U3488 ( .A(n4367), .Y(n4368) );
  AND2X1 U3489 ( .A(n6975), .B(n10119), .Y(n1082) );
  INVX1 U3490 ( .A(n1082), .Y(n4369) );
  INVX1 U3491 ( .A(n4372), .Y(n4370) );
  INVX1 U3492 ( .A(n4370), .Y(n4371) );
  AND2X1 U3493 ( .A(n6978), .B(n10119), .Y(n1081) );
  INVX1 U3494 ( .A(n1081), .Y(n4372) );
  INVX1 U3498 ( .A(n4375), .Y(n4373) );
  INVX1 U3502 ( .A(n4373), .Y(n4374) );
  AND2X1 U3506 ( .A(n6981), .B(n10119), .Y(n1080) );
  INVX1 U3510 ( .A(n1080), .Y(n4375) );
  INVX1 U3511 ( .A(n4378), .Y(n4376) );
  INVX1 U3514 ( .A(n4376), .Y(n4377) );
  AND2X1 U3515 ( .A(n6984), .B(n10119), .Y(n1079) );
  INVX1 U3516 ( .A(n1079), .Y(n4378) );
  INVX1 U3517 ( .A(n4381), .Y(n4379) );
  INVX1 U3518 ( .A(n4379), .Y(n4380) );
  AND2X1 U3519 ( .A(n6987), .B(n10119), .Y(n1078) );
  INVX1 U3520 ( .A(n1078), .Y(n4381) );
  INVX1 U3521 ( .A(n4384), .Y(n4382) );
  INVX1 U3522 ( .A(n4382), .Y(n4383) );
  AND2X1 U3523 ( .A(n6990), .B(n10119), .Y(n1077) );
  INVX1 U3524 ( .A(n1077), .Y(n4384) );
  INVX1 U3525 ( .A(n4387), .Y(n4385) );
  INVX1 U3526 ( .A(n4385), .Y(n4386) );
  AND2X1 U3527 ( .A(n6993), .B(n10119), .Y(n1076) );
  INVX1 U3528 ( .A(n1076), .Y(n4387) );
  INVX1 U3529 ( .A(n4390), .Y(n4388) );
  INVX1 U3530 ( .A(n4388), .Y(n4389) );
  AND2X1 U3531 ( .A(n6996), .B(n10119), .Y(n1075) );
  INVX1 U3532 ( .A(n1075), .Y(n4390) );
  INVX1 U3533 ( .A(n4393), .Y(n4391) );
  INVX1 U3534 ( .A(n4391), .Y(n4392) );
  AND2X1 U3535 ( .A(n6999), .B(n10119), .Y(n1074) );
  INVX1 U3536 ( .A(n1074), .Y(n4393) );
  INVX1 U3537 ( .A(n4396), .Y(n4394) );
  INVX1 U3538 ( .A(n4394), .Y(n4395) );
  AND2X1 U3539 ( .A(n7002), .B(n10119), .Y(n1073) );
  INVX1 U3540 ( .A(n1073), .Y(n4396) );
  INVX1 U3541 ( .A(n4399), .Y(n4397) );
  INVX1 U3542 ( .A(n4397), .Y(n4398) );
  AND2X1 U3543 ( .A(n7005), .B(n10119), .Y(n1072) );
  INVX1 U3544 ( .A(n1072), .Y(n4399) );
  INVX1 U3545 ( .A(n4402), .Y(n4400) );
  INVX1 U3565 ( .A(n4400), .Y(n4401) );
  AND2X1 U3575 ( .A(n8436), .B(n10122), .Y(n1070) );
  INVX1 U3576 ( .A(n1070), .Y(n4402) );
  INVX1 U3577 ( .A(n4405), .Y(n4403) );
  INVX1 U3578 ( .A(n4403), .Y(n4404) );
  AND2X1 U3579 ( .A(n8439), .B(n10122), .Y(n1069) );
  INVX1 U3580 ( .A(n1069), .Y(n4405) );
  INVX1 U3581 ( .A(n4408), .Y(n4406) );
  INVX1 U3582 ( .A(n4406), .Y(n4407) );
  AND2X1 U3583 ( .A(n8442), .B(n10122), .Y(n1068) );
  INVX1 U3584 ( .A(n1068), .Y(n4408) );
  INVX1 U3585 ( .A(n4411), .Y(n4409) );
  INVX1 U3586 ( .A(n4409), .Y(n4410) );
  AND2X1 U3587 ( .A(n8445), .B(n10122), .Y(n1067) );
  INVX1 U3588 ( .A(n1067), .Y(n4411) );
  INVX1 U3589 ( .A(n4414), .Y(n4412) );
  INVX1 U3590 ( .A(n4412), .Y(n4413) );
  AND2X1 U3591 ( .A(n8448), .B(n10122), .Y(n1066) );
  INVX1 U3592 ( .A(n1066), .Y(n4414) );
  INVX1 U3593 ( .A(n4417), .Y(n4415) );
  INVX1 U3594 ( .A(n4415), .Y(n4416) );
  AND2X1 U3595 ( .A(n8451), .B(n10122), .Y(n1065) );
  INVX1 U3596 ( .A(n1065), .Y(n4417) );
  INVX1 U3597 ( .A(n4420), .Y(n4418) );
  INVX1 U3598 ( .A(n4418), .Y(n4419) );
  AND2X1 U3599 ( .A(n8454), .B(n10122), .Y(n1064) );
  INVX1 U3600 ( .A(n1064), .Y(n4420) );
  INVX1 U3601 ( .A(n4423), .Y(n4421) );
  INVX1 U3602 ( .A(n4421), .Y(n4422) );
  AND2X1 U3603 ( .A(n8457), .B(n10122), .Y(n1063) );
  INVX1 U3604 ( .A(n1063), .Y(n4423) );
  INVX1 U3605 ( .A(n4426), .Y(n4424) );
  INVX1 U3606 ( .A(n4424), .Y(n4425) );
  AND2X1 U3607 ( .A(n8460), .B(n10122), .Y(n1062) );
  INVX1 U3608 ( .A(n1062), .Y(n4426) );
  INVX1 U3609 ( .A(n4429), .Y(n4427) );
  INVX1 U3610 ( .A(n4427), .Y(n4428) );
  AND2X1 U3611 ( .A(n8463), .B(n10122), .Y(n1061) );
  INVX1 U3612 ( .A(n1061), .Y(n4429) );
  INVX1 U3613 ( .A(n4432), .Y(n4430) );
  INVX1 U3614 ( .A(n4430), .Y(n4431) );
  AND2X1 U3615 ( .A(n8466), .B(n10122), .Y(n1060) );
  INVX1 U3616 ( .A(n1060), .Y(n4432) );
  INVX1 U3617 ( .A(n4435), .Y(n4433) );
  INVX1 U3618 ( .A(n4433), .Y(n4434) );
  AND2X1 U3619 ( .A(n8469), .B(n10122), .Y(n1059) );
  INVX1 U3620 ( .A(n1059), .Y(n4435) );
  INVX1 U3621 ( .A(n4438), .Y(n4436) );
  INVX1 U3622 ( .A(n4436), .Y(n4437) );
  AND2X1 U3623 ( .A(n8472), .B(n10122), .Y(n1058) );
  INVX1 U3624 ( .A(n1058), .Y(n4438) );
  INVX1 U3625 ( .A(n4441), .Y(n4439) );
  INVX1 U3626 ( .A(n4439), .Y(n4440) );
  AND2X1 U3627 ( .A(n8475), .B(n10122), .Y(n1057) );
  INVX1 U3628 ( .A(n1057), .Y(n4441) );
  INVX1 U3629 ( .A(n4444), .Y(n4442) );
  INVX1 U3630 ( .A(n4442), .Y(n4443) );
  AND2X1 U3631 ( .A(n8478), .B(n10122), .Y(n1056) );
  INVX1 U3632 ( .A(n1056), .Y(n4444) );
  INVX1 U3633 ( .A(n4447), .Y(n4445) );
  INVX1 U3634 ( .A(n4445), .Y(n4446) );
  AND2X1 U3635 ( .A(n8481), .B(n10122), .Y(n1055) );
  INVX1 U3636 ( .A(n1055), .Y(n4447) );
  INVX1 U3637 ( .A(n4450), .Y(n4448) );
  INVX1 U3638 ( .A(n4448), .Y(n4449) );
  AND2X1 U3639 ( .A(n8484), .B(n10122), .Y(n1054) );
  INVX1 U3640 ( .A(n1054), .Y(n4450) );
  INVX1 U3641 ( .A(n4453), .Y(n4451) );
  INVX1 U3642 ( .A(n4451), .Y(n4452) );
  AND2X1 U3643 ( .A(n8487), .B(n10122), .Y(n1053) );
  INVX1 U3644 ( .A(n1053), .Y(n4453) );
  INVX1 U3645 ( .A(n4456), .Y(n4454) );
  INVX1 U3646 ( .A(n4454), .Y(n4455) );
  AND2X1 U3647 ( .A(n8490), .B(n10122), .Y(n1052) );
  INVX1 U3648 ( .A(n1052), .Y(n4456) );
  INVX1 U3649 ( .A(n4459), .Y(n4457) );
  INVX1 U3650 ( .A(n4457), .Y(n4458) );
  AND2X1 U3651 ( .A(n8493), .B(n10122), .Y(n1051) );
  INVX1 U3652 ( .A(n1051), .Y(n4459) );
  INVX1 U3653 ( .A(n4462), .Y(n4460) );
  INVX1 U3654 ( .A(n4460), .Y(n4461) );
  AND2X1 U3655 ( .A(n8496), .B(n10122), .Y(n1050) );
  INVX1 U3656 ( .A(n1050), .Y(n4462) );
  INVX1 U3657 ( .A(n4465), .Y(n4463) );
  INVX1 U3658 ( .A(n4463), .Y(n4464) );
  AND2X1 U3659 ( .A(n8499), .B(n10122), .Y(n1049) );
  INVX1 U3660 ( .A(n1049), .Y(n4465) );
  INVX1 U3661 ( .A(n4468), .Y(n4466) );
  INVX1 U3662 ( .A(n4466), .Y(n4467) );
  AND2X1 U3663 ( .A(n8502), .B(n10122), .Y(n1048) );
  INVX1 U3664 ( .A(n1048), .Y(n4468) );
  INVX1 U3665 ( .A(n4471), .Y(n4469) );
  INVX1 U3666 ( .A(n4469), .Y(n4470) );
  AND2X1 U3667 ( .A(n8505), .B(n10122), .Y(n1047) );
  INVX1 U3668 ( .A(n1047), .Y(n4471) );
  INVX1 U3669 ( .A(n4474), .Y(n4472) );
  INVX1 U3670 ( .A(n4472), .Y(n4473) );
  AND2X1 U3671 ( .A(n8508), .B(n10122), .Y(n1046) );
  INVX1 U3672 ( .A(n1046), .Y(n4474) );
  INVX1 U3673 ( .A(n4477), .Y(n4475) );
  INVX1 U3674 ( .A(n4475), .Y(n4476) );
  AND2X1 U3675 ( .A(n8511), .B(n10122), .Y(n1045) );
  INVX1 U3676 ( .A(n1045), .Y(n4477) );
  INVX1 U3677 ( .A(n4480), .Y(n4478) );
  INVX1 U3678 ( .A(n4478), .Y(n4479) );
  AND2X1 U3679 ( .A(n8514), .B(n10122), .Y(n1044) );
  INVX1 U3680 ( .A(n1044), .Y(n4480) );
  INVX1 U3681 ( .A(n4483), .Y(n4481) );
  INVX1 U3682 ( .A(n4481), .Y(n4482) );
  AND2X1 U3683 ( .A(n8517), .B(n10122), .Y(n1043) );
  INVX1 U3684 ( .A(n1043), .Y(n4483) );
  INVX1 U3685 ( .A(n4486), .Y(n4484) );
  INVX1 U3686 ( .A(n4484), .Y(n4485) );
  AND2X1 U3687 ( .A(n8520), .B(n10122), .Y(n1042) );
  INVX1 U3688 ( .A(n1042), .Y(n4486) );
  INVX1 U3689 ( .A(n4489), .Y(n4487) );
  INVX1 U3690 ( .A(n4487), .Y(n4488) );
  AND2X1 U3691 ( .A(n8523), .B(n10122), .Y(n1041) );
  INVX1 U3692 ( .A(n1041), .Y(n4489) );
  INVX1 U3693 ( .A(n4492), .Y(n4490) );
  INVX1 U3694 ( .A(n4490), .Y(n4491) );
  AND2X1 U3695 ( .A(n8526), .B(n10122), .Y(n1040) );
  INVX1 U3696 ( .A(n1040), .Y(n4492) );
  INVX1 U3697 ( .A(n4495), .Y(n4493) );
  INVX1 U3698 ( .A(n4493), .Y(n4494) );
  AND2X1 U3699 ( .A(n8529), .B(n10122), .Y(n1039) );
  INVX1 U3700 ( .A(n1039), .Y(n4495) );
  INVX1 U3701 ( .A(n4498), .Y(n4496) );
  INVX1 U3702 ( .A(n4496), .Y(n4497) );
  AND2X1 U3703 ( .A(n8532), .B(n10122), .Y(n1038) );
  INVX1 U3704 ( .A(n1038), .Y(n4498) );
  INVX1 U3705 ( .A(n4501), .Y(n4499) );
  INVX1 U3706 ( .A(n4499), .Y(n4500) );
  AND2X1 U3707 ( .A(n8535), .B(n10122), .Y(n1037) );
  INVX1 U3708 ( .A(n1037), .Y(n4501) );
  INVX1 U3709 ( .A(n4504), .Y(n4502) );
  INVX1 U3710 ( .A(n4502), .Y(n4503) );
  AND2X1 U3711 ( .A(n6702), .B(n10125), .Y(n1035) );
  INVX1 U3712 ( .A(n1035), .Y(n4504) );
  INVX1 U3713 ( .A(n4507), .Y(n4505) );
  INVX1 U3714 ( .A(n4505), .Y(n4506) );
  AND2X1 U3715 ( .A(n6705), .B(n10125), .Y(n1034) );
  INVX1 U3716 ( .A(n1034), .Y(n4507) );
  INVX1 U3717 ( .A(n4510), .Y(n4508) );
  INVX1 U3718 ( .A(n4508), .Y(n4509) );
  AND2X1 U3719 ( .A(n6708), .B(n10125), .Y(n1033) );
  INVX1 U3720 ( .A(n1033), .Y(n4510) );
  INVX1 U3721 ( .A(n4513), .Y(n4511) );
  INVX1 U3722 ( .A(n4511), .Y(n4512) );
  AND2X1 U3723 ( .A(n6711), .B(n10125), .Y(n1032) );
  INVX1 U3724 ( .A(n1032), .Y(n4513) );
  INVX1 U3725 ( .A(n4516), .Y(n4514) );
  INVX1 U3726 ( .A(n4514), .Y(n4515) );
  AND2X1 U3727 ( .A(n6714), .B(n10125), .Y(n1031) );
  INVX1 U3728 ( .A(n1031), .Y(n4516) );
  INVX1 U3729 ( .A(n4519), .Y(n4517) );
  INVX1 U3730 ( .A(n4517), .Y(n4518) );
  AND2X1 U3731 ( .A(n6717), .B(n10125), .Y(n1030) );
  INVX1 U3732 ( .A(n1030), .Y(n4519) );
  INVX1 U3733 ( .A(n4522), .Y(n4520) );
  INVX1 U3734 ( .A(n4520), .Y(n4521) );
  AND2X1 U3735 ( .A(n6720), .B(n10125), .Y(n1029) );
  INVX1 U3736 ( .A(n1029), .Y(n4522) );
  INVX1 U3737 ( .A(n4525), .Y(n4523) );
  INVX1 U3738 ( .A(n4523), .Y(n4524) );
  AND2X1 U3739 ( .A(n6723), .B(n10125), .Y(n1028) );
  INVX1 U3740 ( .A(n1028), .Y(n4525) );
  INVX1 U3741 ( .A(n4528), .Y(n4526) );
  INVX1 U3742 ( .A(n4526), .Y(n4527) );
  AND2X1 U3743 ( .A(n6726), .B(n10125), .Y(n1027) );
  INVX1 U3744 ( .A(n1027), .Y(n4528) );
  INVX1 U3745 ( .A(n4531), .Y(n4529) );
  INVX1 U3746 ( .A(n4529), .Y(n4530) );
  AND2X1 U3747 ( .A(n6729), .B(n10125), .Y(n1026) );
  INVX1 U3748 ( .A(n1026), .Y(n4531) );
  INVX1 U3749 ( .A(n4534), .Y(n4532) );
  INVX1 U3750 ( .A(n4532), .Y(n4533) );
  AND2X1 U3751 ( .A(n6732), .B(n10125), .Y(n1025) );
  INVX1 U3752 ( .A(n1025), .Y(n4534) );
  INVX1 U3753 ( .A(n4537), .Y(n4535) );
  INVX1 U3754 ( .A(n4535), .Y(n4536) );
  AND2X1 U3755 ( .A(n6735), .B(n10125), .Y(n1024) );
  INVX1 U3756 ( .A(n1024), .Y(n4537) );
  INVX1 U3757 ( .A(n4540), .Y(n4538) );
  INVX1 U3758 ( .A(n4538), .Y(n4539) );
  AND2X1 U3759 ( .A(n6738), .B(n10125), .Y(n1023) );
  INVX1 U3760 ( .A(n1023), .Y(n4540) );
  INVX1 U3761 ( .A(n4543), .Y(n4541) );
  INVX1 U3762 ( .A(n4541), .Y(n4542) );
  AND2X1 U3763 ( .A(n6741), .B(n10125), .Y(n1022) );
  INVX1 U3764 ( .A(n1022), .Y(n4543) );
  INVX1 U3765 ( .A(n4546), .Y(n4544) );
  INVX1 U3766 ( .A(n4544), .Y(n4545) );
  AND2X1 U3767 ( .A(n6744), .B(n10125), .Y(n1021) );
  INVX1 U3768 ( .A(n1021), .Y(n4546) );
  INVX1 U3769 ( .A(n4549), .Y(n4547) );
  INVX1 U3770 ( .A(n4547), .Y(n4548) );
  AND2X1 U3771 ( .A(n6747), .B(n10125), .Y(n1020) );
  INVX1 U3772 ( .A(n1020), .Y(n4549) );
  INVX1 U3773 ( .A(n4552), .Y(n4550) );
  INVX1 U3774 ( .A(n4550), .Y(n4551) );
  AND2X1 U3775 ( .A(n6750), .B(n10125), .Y(n1019) );
  INVX1 U3776 ( .A(n1019), .Y(n4552) );
  INVX1 U3777 ( .A(n4555), .Y(n4553) );
  INVX1 U3778 ( .A(n4553), .Y(n4554) );
  AND2X1 U3779 ( .A(n6753), .B(n10125), .Y(n1018) );
  INVX1 U3780 ( .A(n1018), .Y(n4555) );
  INVX1 U3781 ( .A(n4558), .Y(n4556) );
  INVX1 U3782 ( .A(n4556), .Y(n4557) );
  AND2X1 U3783 ( .A(n6756), .B(n10125), .Y(n1017) );
  INVX1 U3784 ( .A(n1017), .Y(n4558) );
  INVX1 U3785 ( .A(n4561), .Y(n4559) );
  INVX1 U3786 ( .A(n4559), .Y(n4560) );
  AND2X1 U3787 ( .A(n6759), .B(n10125), .Y(n1016) );
  INVX1 U3788 ( .A(n1016), .Y(n4561) );
  INVX1 U3789 ( .A(n4564), .Y(n4562) );
  INVX1 U3790 ( .A(n4562), .Y(n4563) );
  AND2X1 U3791 ( .A(n6762), .B(n10125), .Y(n1015) );
  INVX1 U3792 ( .A(n1015), .Y(n4564) );
  INVX1 U3793 ( .A(n4567), .Y(n4565) );
  INVX1 U3794 ( .A(n4565), .Y(n4566) );
  AND2X1 U3795 ( .A(n6765), .B(n10125), .Y(n1014) );
  INVX1 U3796 ( .A(n1014), .Y(n4567) );
  INVX1 U3797 ( .A(n4570), .Y(n4568) );
  INVX1 U3798 ( .A(n4568), .Y(n4569) );
  AND2X1 U3799 ( .A(n6768), .B(n10125), .Y(n1013) );
  INVX1 U3800 ( .A(n1013), .Y(n4570) );
  INVX1 U3801 ( .A(n4573), .Y(n4571) );
  INVX1 U3802 ( .A(n4571), .Y(n4572) );
  AND2X1 U3803 ( .A(n6771), .B(n10125), .Y(n1012) );
  INVX1 U3804 ( .A(n1012), .Y(n4573) );
  INVX1 U3805 ( .A(n4576), .Y(n4574) );
  INVX1 U3806 ( .A(n4574), .Y(n4575) );
  AND2X1 U3807 ( .A(n6774), .B(n10125), .Y(n1011) );
  INVX1 U3808 ( .A(n1011), .Y(n4576) );
  INVX1 U3809 ( .A(n4579), .Y(n4577) );
  INVX1 U3810 ( .A(n4577), .Y(n4578) );
  AND2X1 U3811 ( .A(n6777), .B(n10125), .Y(n1010) );
  INVX1 U3812 ( .A(n1010), .Y(n4579) );
  INVX1 U3813 ( .A(n4582), .Y(n4580) );
  INVX1 U3814 ( .A(n4580), .Y(n4581) );
  AND2X1 U3815 ( .A(n6780), .B(n10125), .Y(n1009) );
  INVX1 U3816 ( .A(n1009), .Y(n4582) );
  INVX1 U3817 ( .A(n4585), .Y(n4583) );
  INVX1 U3818 ( .A(n4583), .Y(n4584) );
  AND2X1 U3819 ( .A(n6783), .B(n10125), .Y(n1008) );
  INVX1 U3820 ( .A(n1008), .Y(n4585) );
  INVX1 U3821 ( .A(n4588), .Y(n4586) );
  INVX1 U3822 ( .A(n4586), .Y(n4587) );
  AND2X1 U3823 ( .A(n6786), .B(n10125), .Y(n1007) );
  INVX1 U3824 ( .A(n1007), .Y(n4588) );
  INVX1 U3825 ( .A(n4591), .Y(n4589) );
  INVX1 U3826 ( .A(n4589), .Y(n4590) );
  AND2X1 U3827 ( .A(n6789), .B(n10125), .Y(n1006) );
  INVX1 U3828 ( .A(n1006), .Y(n4591) );
  INVX1 U3829 ( .A(n4594), .Y(n4592) );
  INVX1 U3830 ( .A(n4592), .Y(n4593) );
  AND2X1 U3831 ( .A(n6792), .B(n10125), .Y(n1005) );
  INVX1 U3832 ( .A(n1005), .Y(n4594) );
  INVX1 U3833 ( .A(n4597), .Y(n4595) );
  INVX1 U3834 ( .A(n4595), .Y(n4596) );
  AND2X1 U3835 ( .A(n6795), .B(n10125), .Y(n1004) );
  INVX1 U3836 ( .A(n1004), .Y(n4597) );
  INVX1 U3837 ( .A(n4600), .Y(n4598) );
  INVX1 U3838 ( .A(n4598), .Y(n4599) );
  AND2X1 U3839 ( .A(n6798), .B(n10125), .Y(n1003) );
  INVX1 U3840 ( .A(n1003), .Y(n4600) );
  INVX1 U3841 ( .A(n4603), .Y(n4601) );
  INVX1 U3842 ( .A(n4601), .Y(n4602) );
  AND2X1 U3843 ( .A(n6801), .B(n10125), .Y(n1002) );
  INVX1 U3844 ( .A(n1002), .Y(n4603) );
  INVX1 U3845 ( .A(n4606), .Y(n4604) );
  INVX1 U3846 ( .A(n4604), .Y(n4605) );
  AND2X1 U3847 ( .A(n8334), .B(n10128), .Y(n1000) );
  INVX1 U3848 ( .A(n1000), .Y(n4606) );
  INVX1 U3849 ( .A(n4609), .Y(n4607) );
  INVX1 U3850 ( .A(n4607), .Y(n4608) );
  AND2X1 U3851 ( .A(n8337), .B(n10128), .Y(n999) );
  INVX1 U3852 ( .A(n999), .Y(n4609) );
  INVX1 U3853 ( .A(n4612), .Y(n4610) );
  INVX1 U3854 ( .A(n4610), .Y(n4611) );
  AND2X1 U3855 ( .A(n8340), .B(n10128), .Y(n998) );
  INVX1 U3856 ( .A(n998), .Y(n4612) );
  INVX1 U3857 ( .A(n4615), .Y(n4613) );
  INVX1 U3858 ( .A(n4613), .Y(n4614) );
  AND2X1 U3859 ( .A(n8343), .B(n10128), .Y(n997) );
  INVX1 U3860 ( .A(n997), .Y(n4615) );
  INVX1 U3861 ( .A(n4618), .Y(n4616) );
  INVX1 U3862 ( .A(n4616), .Y(n4617) );
  AND2X1 U3863 ( .A(n8346), .B(n10128), .Y(n996) );
  INVX1 U3864 ( .A(n996), .Y(n4618) );
  INVX1 U3865 ( .A(n4621), .Y(n4619) );
  INVX1 U3866 ( .A(n4619), .Y(n4620) );
  AND2X1 U3867 ( .A(n8349), .B(n10128), .Y(n995) );
  INVX1 U3868 ( .A(n995), .Y(n4621) );
  INVX1 U3869 ( .A(n4624), .Y(n4622) );
  INVX1 U3870 ( .A(n4622), .Y(n4623) );
  AND2X1 U3871 ( .A(n8352), .B(n10128), .Y(n994) );
  INVX1 U3872 ( .A(n994), .Y(n4624) );
  INVX1 U3873 ( .A(n4627), .Y(n4625) );
  INVX1 U3874 ( .A(n4625), .Y(n4626) );
  AND2X1 U3875 ( .A(n8355), .B(n10128), .Y(n993) );
  INVX1 U3876 ( .A(n993), .Y(n4627) );
  INVX1 U3877 ( .A(n4630), .Y(n4628) );
  INVX1 U3878 ( .A(n4628), .Y(n4629) );
  AND2X1 U3879 ( .A(n8358), .B(n10128), .Y(n992) );
  INVX1 U3880 ( .A(n992), .Y(n4630) );
  INVX1 U3881 ( .A(n4633), .Y(n4631) );
  INVX1 U3882 ( .A(n4631), .Y(n4632) );
  AND2X1 U3883 ( .A(n8361), .B(n10128), .Y(n991) );
  INVX1 U3884 ( .A(n991), .Y(n4633) );
  INVX1 U3885 ( .A(n4636), .Y(n4634) );
  INVX1 U3886 ( .A(n4634), .Y(n4635) );
  AND2X1 U3887 ( .A(n8364), .B(n10128), .Y(n990) );
  INVX1 U3888 ( .A(n990), .Y(n4636) );
  INVX1 U3889 ( .A(n4639), .Y(n4637) );
  INVX1 U3890 ( .A(n4637), .Y(n4638) );
  AND2X1 U3891 ( .A(n8367), .B(n10128), .Y(n989) );
  INVX1 U3892 ( .A(n989), .Y(n4639) );
  INVX1 U3893 ( .A(n4642), .Y(n4640) );
  INVX1 U3894 ( .A(n4640), .Y(n4641) );
  AND2X1 U3895 ( .A(n8370), .B(n10128), .Y(n988) );
  INVX1 U3896 ( .A(n988), .Y(n4642) );
  INVX1 U3897 ( .A(n4645), .Y(n4643) );
  INVX1 U3898 ( .A(n4643), .Y(n4644) );
  AND2X1 U3899 ( .A(n8373), .B(n10128), .Y(n987) );
  INVX1 U3900 ( .A(n987), .Y(n4645) );
  INVX1 U3901 ( .A(n4648), .Y(n4646) );
  INVX1 U3902 ( .A(n4646), .Y(n4647) );
  AND2X1 U3903 ( .A(n8376), .B(n10128), .Y(n986) );
  INVX1 U3904 ( .A(n986), .Y(n4648) );
  INVX1 U3905 ( .A(n4651), .Y(n4649) );
  INVX1 U3906 ( .A(n4649), .Y(n4650) );
  AND2X1 U3907 ( .A(n8379), .B(n10128), .Y(n985) );
  INVX1 U3908 ( .A(n985), .Y(n4651) );
  INVX1 U3909 ( .A(n4654), .Y(n4652) );
  INVX1 U3910 ( .A(n4652), .Y(n4653) );
  AND2X1 U3911 ( .A(n8382), .B(n10128), .Y(n984) );
  INVX1 U3912 ( .A(n984), .Y(n4654) );
  INVX1 U3913 ( .A(n4657), .Y(n4655) );
  INVX1 U3914 ( .A(n4655), .Y(n4656) );
  AND2X1 U3915 ( .A(n8385), .B(n10128), .Y(n983) );
  INVX1 U3916 ( .A(n983), .Y(n4657) );
  INVX1 U3917 ( .A(n4660), .Y(n4658) );
  INVX1 U3918 ( .A(n4658), .Y(n4659) );
  AND2X1 U3919 ( .A(n8388), .B(n10128), .Y(n982) );
  INVX1 U3920 ( .A(n982), .Y(n4660) );
  INVX1 U3921 ( .A(n4663), .Y(n4661) );
  INVX1 U3922 ( .A(n4661), .Y(n4662) );
  AND2X1 U3923 ( .A(n8391), .B(n10128), .Y(n981) );
  INVX1 U3924 ( .A(n981), .Y(n4663) );
  INVX1 U3925 ( .A(n4666), .Y(n4664) );
  INVX1 U3926 ( .A(n4664), .Y(n4665) );
  AND2X1 U3927 ( .A(n8394), .B(n10128), .Y(n980) );
  INVX1 U3928 ( .A(n980), .Y(n4666) );
  INVX1 U3929 ( .A(n4669), .Y(n4667) );
  INVX1 U3930 ( .A(n4667), .Y(n4668) );
  AND2X1 U3931 ( .A(n8397), .B(n10128), .Y(n979) );
  INVX1 U3932 ( .A(n979), .Y(n4669) );
  INVX1 U3933 ( .A(n4672), .Y(n4670) );
  INVX1 U3934 ( .A(n4670), .Y(n4671) );
  AND2X1 U3935 ( .A(n8400), .B(n10128), .Y(n978) );
  INVX1 U3936 ( .A(n978), .Y(n4672) );
  INVX1 U3937 ( .A(n4675), .Y(n4673) );
  INVX1 U3938 ( .A(n4673), .Y(n4674) );
  AND2X1 U3939 ( .A(n8403), .B(n10128), .Y(n977) );
  INVX1 U3940 ( .A(n977), .Y(n4675) );
  INVX1 U3941 ( .A(n4678), .Y(n4676) );
  INVX1 U3942 ( .A(n4676), .Y(n4677) );
  AND2X1 U3943 ( .A(n8406), .B(n10128), .Y(n976) );
  INVX1 U3944 ( .A(n976), .Y(n4678) );
  INVX1 U3945 ( .A(n4681), .Y(n4679) );
  INVX1 U3946 ( .A(n4679), .Y(n4680) );
  AND2X1 U3947 ( .A(n8409), .B(n10128), .Y(n975) );
  INVX1 U3948 ( .A(n975), .Y(n4681) );
  INVX1 U3949 ( .A(n4684), .Y(n4682) );
  INVX1 U3950 ( .A(n4682), .Y(n4683) );
  AND2X1 U3951 ( .A(n8412), .B(n10128), .Y(n974) );
  INVX1 U3952 ( .A(n974), .Y(n4684) );
  INVX1 U3953 ( .A(n4687), .Y(n4685) );
  INVX1 U3954 ( .A(n4685), .Y(n4686) );
  AND2X1 U3955 ( .A(n8415), .B(n10128), .Y(n973) );
  INVX1 U3956 ( .A(n973), .Y(n4687) );
  INVX1 U3957 ( .A(n4690), .Y(n4688) );
  INVX1 U3958 ( .A(n4688), .Y(n4689) );
  AND2X1 U3959 ( .A(n8418), .B(n10128), .Y(n972) );
  INVX1 U3960 ( .A(n972), .Y(n4690) );
  INVX1 U3961 ( .A(n4693), .Y(n4691) );
  INVX1 U3962 ( .A(n4691), .Y(n4692) );
  AND2X1 U3963 ( .A(n8421), .B(n10128), .Y(n971) );
  INVX1 U3964 ( .A(n971), .Y(n4693) );
  INVX1 U3965 ( .A(n4696), .Y(n4694) );
  INVX1 U3966 ( .A(n4694), .Y(n4695) );
  AND2X1 U3967 ( .A(n8424), .B(n10128), .Y(n970) );
  INVX1 U3968 ( .A(n970), .Y(n4696) );
  INVX1 U3969 ( .A(n4699), .Y(n4697) );
  INVX1 U3970 ( .A(n4697), .Y(n4698) );
  AND2X1 U3971 ( .A(n8427), .B(n10128), .Y(n969) );
  INVX1 U3972 ( .A(n969), .Y(n4699) );
  INVX1 U3973 ( .A(n4702), .Y(n4700) );
  INVX1 U3974 ( .A(n4700), .Y(n4701) );
  AND2X1 U3975 ( .A(n8430), .B(n10128), .Y(n968) );
  INVX1 U3976 ( .A(n968), .Y(n4702) );
  INVX1 U3977 ( .A(n4705), .Y(n4703) );
  INVX1 U3978 ( .A(n4703), .Y(n4704) );
  AND2X1 U3979 ( .A(n8433), .B(n10128), .Y(n967) );
  INVX1 U3980 ( .A(n967), .Y(n4705) );
  INVX1 U3981 ( .A(n4708), .Y(n4706) );
  INVX1 U3982 ( .A(n4706), .Y(n4707) );
  AND2X1 U3983 ( .A(n6804), .B(n10131), .Y(n965) );
  INVX1 U3984 ( .A(n965), .Y(n4708) );
  INVX1 U3985 ( .A(n4711), .Y(n4709) );
  INVX1 U3986 ( .A(n4709), .Y(n4710) );
  AND2X1 U3987 ( .A(n6807), .B(n10131), .Y(n964) );
  INVX1 U3988 ( .A(n964), .Y(n4711) );
  INVX1 U3989 ( .A(n4714), .Y(n4712) );
  INVX1 U3990 ( .A(n4712), .Y(n4713) );
  AND2X1 U3991 ( .A(n6810), .B(n10131), .Y(n963) );
  INVX1 U3992 ( .A(n963), .Y(n4714) );
  INVX1 U3993 ( .A(n4717), .Y(n4715) );
  INVX1 U3994 ( .A(n4715), .Y(n4716) );
  AND2X1 U3995 ( .A(n6813), .B(n10131), .Y(n962) );
  INVX1 U3996 ( .A(n962), .Y(n4717) );
  INVX1 U3997 ( .A(n4720), .Y(n4718) );
  INVX1 U3998 ( .A(n4718), .Y(n4719) );
  AND2X1 U3999 ( .A(n6816), .B(n10131), .Y(n961) );
  INVX1 U4000 ( .A(n961), .Y(n4720) );
  INVX1 U4001 ( .A(n4723), .Y(n4721) );
  INVX1 U4002 ( .A(n4721), .Y(n4722) );
  AND2X1 U4003 ( .A(n6819), .B(n10131), .Y(n960) );
  INVX1 U4004 ( .A(n960), .Y(n4723) );
  INVX1 U4005 ( .A(n4726), .Y(n4724) );
  INVX1 U4006 ( .A(n4724), .Y(n4725) );
  AND2X1 U4007 ( .A(n6822), .B(n10131), .Y(n959) );
  INVX1 U4008 ( .A(n959), .Y(n4726) );
  INVX1 U4009 ( .A(n4729), .Y(n4727) );
  INVX1 U4010 ( .A(n4727), .Y(n4728) );
  AND2X1 U4011 ( .A(n6825), .B(n10131), .Y(n958) );
  INVX1 U4012 ( .A(n958), .Y(n4729) );
  INVX1 U4013 ( .A(n4732), .Y(n4730) );
  INVX1 U4014 ( .A(n4730), .Y(n4731) );
  AND2X1 U4015 ( .A(n6828), .B(n10131), .Y(n957) );
  INVX1 U4016 ( .A(n957), .Y(n4732) );
  INVX1 U4017 ( .A(n4735), .Y(n4733) );
  INVX1 U4018 ( .A(n4733), .Y(n4734) );
  AND2X1 U4019 ( .A(n6831), .B(n10131), .Y(n956) );
  INVX1 U4020 ( .A(n956), .Y(n4735) );
  INVX1 U4021 ( .A(n4738), .Y(n4736) );
  INVX1 U4022 ( .A(n4736), .Y(n4737) );
  AND2X1 U4023 ( .A(n6834), .B(n10131), .Y(n955) );
  INVX1 U4024 ( .A(n955), .Y(n4738) );
  INVX1 U4025 ( .A(n4741), .Y(n4739) );
  INVX1 U4026 ( .A(n4739), .Y(n4740) );
  AND2X1 U4027 ( .A(n6837), .B(n10131), .Y(n954) );
  INVX1 U4028 ( .A(n954), .Y(n4741) );
  INVX1 U4029 ( .A(n4744), .Y(n4742) );
  INVX1 U4030 ( .A(n4742), .Y(n4743) );
  AND2X1 U4031 ( .A(n6840), .B(n10131), .Y(n953) );
  INVX1 U4032 ( .A(n953), .Y(n4744) );
  INVX1 U4033 ( .A(n4747), .Y(n4745) );
  INVX1 U4034 ( .A(n4745), .Y(n4746) );
  AND2X1 U4035 ( .A(n6843), .B(n10131), .Y(n952) );
  INVX1 U4036 ( .A(n952), .Y(n4747) );
  INVX1 U4037 ( .A(n4750), .Y(n4748) );
  INVX1 U4038 ( .A(n4748), .Y(n4749) );
  AND2X1 U4039 ( .A(n6846), .B(n10131), .Y(n951) );
  INVX1 U4040 ( .A(n951), .Y(n4750) );
  INVX1 U4041 ( .A(n4753), .Y(n4751) );
  INVX1 U4042 ( .A(n4751), .Y(n4752) );
  AND2X1 U4043 ( .A(n6849), .B(n10131), .Y(n950) );
  INVX1 U4044 ( .A(n950), .Y(n4753) );
  INVX1 U4045 ( .A(n4756), .Y(n4754) );
  INVX1 U4046 ( .A(n4754), .Y(n4755) );
  AND2X1 U4047 ( .A(n6852), .B(n10131), .Y(n949) );
  INVX1 U4048 ( .A(n949), .Y(n4756) );
  INVX1 U4049 ( .A(n4759), .Y(n4757) );
  INVX1 U4050 ( .A(n4757), .Y(n4758) );
  AND2X1 U4051 ( .A(n6855), .B(n10131), .Y(n948) );
  INVX1 U4052 ( .A(n948), .Y(n4759) );
  INVX1 U4053 ( .A(n4762), .Y(n4760) );
  INVX1 U4054 ( .A(n4760), .Y(n4761) );
  AND2X1 U4055 ( .A(n6858), .B(n10131), .Y(n947) );
  INVX1 U4056 ( .A(n947), .Y(n4762) );
  INVX1 U4057 ( .A(n4765), .Y(n4763) );
  INVX1 U4058 ( .A(n4763), .Y(n4764) );
  AND2X1 U4059 ( .A(n6861), .B(n10131), .Y(n946) );
  INVX1 U4060 ( .A(n946), .Y(n4765) );
  INVX1 U4061 ( .A(n4768), .Y(n4766) );
  INVX1 U4062 ( .A(n4766), .Y(n4767) );
  AND2X1 U4063 ( .A(n6864), .B(n10131), .Y(n945) );
  INVX1 U4064 ( .A(n945), .Y(n4768) );
  INVX1 U4065 ( .A(n4771), .Y(n4769) );
  INVX1 U4066 ( .A(n4769), .Y(n4770) );
  AND2X1 U4067 ( .A(n6867), .B(n10131), .Y(n944) );
  INVX1 U4068 ( .A(n944), .Y(n4771) );
  INVX1 U4069 ( .A(n4774), .Y(n4772) );
  INVX1 U4070 ( .A(n4772), .Y(n4773) );
  AND2X1 U4071 ( .A(n6870), .B(n10131), .Y(n943) );
  INVX1 U4072 ( .A(n943), .Y(n4774) );
  INVX1 U4073 ( .A(n4777), .Y(n4775) );
  INVX1 U4074 ( .A(n4775), .Y(n4776) );
  AND2X1 U4075 ( .A(n6873), .B(n10131), .Y(n942) );
  INVX1 U4076 ( .A(n942), .Y(n4777) );
  INVX1 U4077 ( .A(n4780), .Y(n4778) );
  INVX1 U4078 ( .A(n4778), .Y(n4779) );
  AND2X1 U4079 ( .A(n6876), .B(n10131), .Y(n941) );
  INVX1 U4080 ( .A(n941), .Y(n4780) );
  INVX1 U4081 ( .A(n4783), .Y(n4781) );
  INVX1 U4082 ( .A(n4781), .Y(n4782) );
  AND2X1 U4083 ( .A(n6879), .B(n10131), .Y(n940) );
  INVX1 U4084 ( .A(n940), .Y(n4783) );
  INVX1 U4085 ( .A(n4786), .Y(n4784) );
  INVX1 U4086 ( .A(n4784), .Y(n4785) );
  AND2X1 U4087 ( .A(n6882), .B(n10131), .Y(n939) );
  INVX1 U4088 ( .A(n939), .Y(n4786) );
  INVX1 U4089 ( .A(n4789), .Y(n4787) );
  INVX1 U4090 ( .A(n4787), .Y(n4788) );
  AND2X1 U4091 ( .A(n6885), .B(n10131), .Y(n938) );
  INVX1 U4092 ( .A(n938), .Y(n4789) );
  INVX1 U4093 ( .A(n4792), .Y(n4790) );
  INVX1 U4094 ( .A(n4790), .Y(n4791) );
  AND2X1 U4095 ( .A(n6888), .B(n10131), .Y(n937) );
  INVX1 U4096 ( .A(n937), .Y(n4792) );
  INVX1 U4097 ( .A(n4795), .Y(n4793) );
  INVX1 U4098 ( .A(n4793), .Y(n4794) );
  AND2X1 U4099 ( .A(n6891), .B(n10131), .Y(n936) );
  INVX1 U4100 ( .A(n936), .Y(n4795) );
  INVX1 U4101 ( .A(n4798), .Y(n4796) );
  INVX1 U4102 ( .A(n4796), .Y(n4797) );
  AND2X1 U4103 ( .A(n6894), .B(n10131), .Y(n935) );
  INVX1 U4104 ( .A(n935), .Y(n4798) );
  INVX1 U4105 ( .A(n4801), .Y(n4799) );
  INVX1 U4106 ( .A(n4799), .Y(n4800) );
  AND2X1 U4107 ( .A(n6897), .B(n10131), .Y(n934) );
  INVX1 U4108 ( .A(n934), .Y(n4801) );
  INVX1 U4109 ( .A(n4804), .Y(n4802) );
  INVX1 U4110 ( .A(n4802), .Y(n4803) );
  AND2X1 U4111 ( .A(n6900), .B(n10131), .Y(n933) );
  INVX1 U4112 ( .A(n933), .Y(n4804) );
  INVX1 U4113 ( .A(n4807), .Y(n4805) );
  INVX1 U4114 ( .A(n4805), .Y(n4806) );
  AND2X1 U4115 ( .A(n6903), .B(n10131), .Y(n932) );
  INVX1 U4116 ( .A(n932), .Y(n4807) );
  INVX1 U4117 ( .A(n4810), .Y(n4808) );
  INVX1 U4118 ( .A(n4808), .Y(n4809) );
  AND2X1 U4119 ( .A(n8640), .B(n10134), .Y(n930) );
  INVX1 U4120 ( .A(n930), .Y(n4810) );
  INVX1 U4121 ( .A(n4813), .Y(n4811) );
  INVX1 U4122 ( .A(n4811), .Y(n4812) );
  AND2X1 U4123 ( .A(n8643), .B(n10134), .Y(n929) );
  INVX1 U4124 ( .A(n929), .Y(n4813) );
  INVX1 U4125 ( .A(n4816), .Y(n4814) );
  INVX1 U4126 ( .A(n4814), .Y(n4815) );
  AND2X1 U4127 ( .A(n8646), .B(n10134), .Y(n928) );
  INVX1 U4128 ( .A(n928), .Y(n4816) );
  INVX1 U4129 ( .A(n4819), .Y(n4817) );
  INVX1 U4130 ( .A(n4817), .Y(n4818) );
  AND2X1 U4131 ( .A(n8649), .B(n10134), .Y(n927) );
  INVX1 U4132 ( .A(n927), .Y(n4819) );
  INVX1 U4133 ( .A(n4822), .Y(n4820) );
  INVX1 U4134 ( .A(n4820), .Y(n4821) );
  AND2X1 U4135 ( .A(n8652), .B(n10134), .Y(n926) );
  INVX1 U4136 ( .A(n926), .Y(n4822) );
  INVX1 U4137 ( .A(n4825), .Y(n4823) );
  INVX1 U4138 ( .A(n4823), .Y(n4824) );
  AND2X1 U4139 ( .A(n8655), .B(n10134), .Y(n925) );
  INVX1 U4140 ( .A(n925), .Y(n4825) );
  INVX1 U4141 ( .A(n4828), .Y(n4826) );
  INVX1 U4142 ( .A(n4826), .Y(n4827) );
  AND2X1 U4143 ( .A(n8658), .B(n10134), .Y(n924) );
  INVX1 U4144 ( .A(n924), .Y(n4828) );
  INVX1 U4145 ( .A(n4831), .Y(n4829) );
  INVX1 U4146 ( .A(n4829), .Y(n4830) );
  AND2X1 U4147 ( .A(n8661), .B(n10134), .Y(n923) );
  INVX1 U4148 ( .A(n923), .Y(n4831) );
  INVX1 U4149 ( .A(n4834), .Y(n4832) );
  INVX1 U4150 ( .A(n4832), .Y(n4833) );
  AND2X1 U4151 ( .A(n8664), .B(n10134), .Y(n922) );
  INVX1 U4152 ( .A(n922), .Y(n4834) );
  INVX1 U4153 ( .A(n4837), .Y(n4835) );
  INVX1 U4154 ( .A(n4835), .Y(n4836) );
  AND2X1 U4155 ( .A(n8667), .B(n10134), .Y(n921) );
  INVX1 U4156 ( .A(n921), .Y(n4837) );
  INVX1 U4157 ( .A(n4840), .Y(n4838) );
  INVX1 U4158 ( .A(n4838), .Y(n4839) );
  AND2X1 U4159 ( .A(n8670), .B(n10134), .Y(n920) );
  INVX1 U4160 ( .A(n920), .Y(n4840) );
  INVX1 U4161 ( .A(n4843), .Y(n4841) );
  INVX1 U4162 ( .A(n4841), .Y(n4842) );
  AND2X1 U4163 ( .A(n8673), .B(n10134), .Y(n919) );
  INVX1 U4164 ( .A(n919), .Y(n4843) );
  INVX1 U4165 ( .A(n4846), .Y(n4844) );
  INVX1 U4166 ( .A(n4844), .Y(n4845) );
  AND2X1 U4167 ( .A(n8676), .B(n10134), .Y(n918) );
  INVX1 U4168 ( .A(n918), .Y(n4846) );
  INVX1 U4169 ( .A(n4849), .Y(n4847) );
  INVX1 U4170 ( .A(n4847), .Y(n4848) );
  AND2X1 U4171 ( .A(n8679), .B(n10134), .Y(n917) );
  INVX1 U4172 ( .A(n917), .Y(n4849) );
  INVX1 U4173 ( .A(n4852), .Y(n4850) );
  INVX1 U4174 ( .A(n4850), .Y(n4851) );
  AND2X1 U4175 ( .A(n8682), .B(n10134), .Y(n916) );
  INVX1 U4176 ( .A(n916), .Y(n4852) );
  INVX1 U4177 ( .A(n4855), .Y(n4853) );
  INVX1 U4178 ( .A(n4853), .Y(n4854) );
  AND2X1 U4179 ( .A(n8685), .B(n10134), .Y(n915) );
  INVX1 U4180 ( .A(n915), .Y(n4855) );
  INVX1 U4181 ( .A(n4858), .Y(n4856) );
  INVX1 U4182 ( .A(n4856), .Y(n4857) );
  AND2X1 U4183 ( .A(n8688), .B(n10134), .Y(n914) );
  INVX1 U4184 ( .A(n914), .Y(n4858) );
  INVX1 U4185 ( .A(n4861), .Y(n4859) );
  INVX1 U4186 ( .A(n4859), .Y(n4860) );
  AND2X1 U4187 ( .A(n8691), .B(n10134), .Y(n913) );
  INVX1 U4188 ( .A(n913), .Y(n4861) );
  INVX1 U4189 ( .A(n4864), .Y(n4862) );
  INVX1 U4190 ( .A(n4862), .Y(n4863) );
  AND2X1 U4191 ( .A(n8694), .B(n10134), .Y(n912) );
  INVX1 U4192 ( .A(n912), .Y(n4864) );
  INVX1 U4193 ( .A(n4867), .Y(n4865) );
  INVX1 U4194 ( .A(n4865), .Y(n4866) );
  AND2X1 U4195 ( .A(n8697), .B(n10134), .Y(n911) );
  INVX1 U4196 ( .A(n911), .Y(n4867) );
  INVX1 U4197 ( .A(n4870), .Y(n4868) );
  INVX1 U4198 ( .A(n4868), .Y(n4869) );
  AND2X1 U4199 ( .A(n8700), .B(n10134), .Y(n910) );
  INVX1 U4200 ( .A(n910), .Y(n4870) );
  INVX1 U4201 ( .A(n4873), .Y(n4871) );
  INVX1 U4202 ( .A(n4871), .Y(n4872) );
  AND2X1 U4203 ( .A(n8703), .B(n10134), .Y(n909) );
  INVX1 U4204 ( .A(n909), .Y(n4873) );
  INVX1 U4205 ( .A(n4876), .Y(n4874) );
  INVX1 U4206 ( .A(n4874), .Y(n4875) );
  AND2X1 U4207 ( .A(n8706), .B(n10134), .Y(n908) );
  INVX1 U4208 ( .A(n908), .Y(n4876) );
  INVX1 U4209 ( .A(n4879), .Y(n4877) );
  INVX1 U4210 ( .A(n4877), .Y(n4878) );
  AND2X1 U4211 ( .A(n8709), .B(n10134), .Y(n907) );
  INVX1 U4212 ( .A(n907), .Y(n4879) );
  INVX1 U4213 ( .A(n4882), .Y(n4880) );
  INVX1 U4214 ( .A(n4880), .Y(n4881) );
  AND2X1 U4215 ( .A(n8712), .B(n10134), .Y(n906) );
  INVX1 U4216 ( .A(n906), .Y(n4882) );
  INVX1 U4217 ( .A(n4885), .Y(n4883) );
  INVX1 U4218 ( .A(n4883), .Y(n4884) );
  AND2X1 U4219 ( .A(n8715), .B(n10134), .Y(n905) );
  INVX1 U4220 ( .A(n905), .Y(n4885) );
  INVX1 U4221 ( .A(n4888), .Y(n4886) );
  INVX1 U4222 ( .A(n4886), .Y(n4887) );
  AND2X1 U4223 ( .A(n8718), .B(n10134), .Y(n904) );
  INVX1 U4224 ( .A(n904), .Y(n4888) );
  INVX1 U4225 ( .A(n4891), .Y(n4889) );
  INVX1 U4226 ( .A(n4889), .Y(n4890) );
  AND2X1 U4227 ( .A(n8721), .B(n10134), .Y(n903) );
  INVX1 U4228 ( .A(n903), .Y(n4891) );
  INVX1 U4229 ( .A(n4894), .Y(n4892) );
  INVX1 U4230 ( .A(n4892), .Y(n4893) );
  AND2X1 U4231 ( .A(n8724), .B(n10134), .Y(n902) );
  INVX1 U4232 ( .A(n902), .Y(n4894) );
  INVX1 U4233 ( .A(n4897), .Y(n4895) );
  INVX1 U4234 ( .A(n4895), .Y(n4896) );
  AND2X1 U4235 ( .A(n8727), .B(n10134), .Y(n901) );
  INVX1 U4236 ( .A(n901), .Y(n4897) );
  INVX1 U4237 ( .A(n4900), .Y(n4898) );
  INVX1 U4238 ( .A(n4898), .Y(n4899) );
  AND2X1 U4239 ( .A(n8730), .B(n10134), .Y(n900) );
  INVX1 U4240 ( .A(n900), .Y(n4900) );
  INVX1 U4241 ( .A(n4903), .Y(n4901) );
  INVX1 U4242 ( .A(n4901), .Y(n4902) );
  AND2X1 U4243 ( .A(n8733), .B(n10134), .Y(n899) );
  INVX1 U4244 ( .A(n899), .Y(n4903) );
  INVX1 U4245 ( .A(n4906), .Y(n4904) );
  INVX1 U4246 ( .A(n4904), .Y(n4905) );
  AND2X1 U4247 ( .A(n8736), .B(n10134), .Y(n898) );
  INVX1 U4248 ( .A(n898), .Y(n4906) );
  INVX1 U4249 ( .A(n4909), .Y(n4907) );
  INVX1 U4250 ( .A(n4907), .Y(n4908) );
  AND2X1 U4251 ( .A(n8739), .B(n10134), .Y(n897) );
  INVX1 U4252 ( .A(n897), .Y(n4909) );
  INVX1 U4253 ( .A(n4912), .Y(n4910) );
  INVX1 U4254 ( .A(n4910), .Y(n4911) );
  AND2X1 U4255 ( .A(n7008), .B(n10137), .Y(n894) );
  INVX1 U4256 ( .A(n894), .Y(n4912) );
  INVX1 U4257 ( .A(n4915), .Y(n4913) );
  INVX1 U4258 ( .A(n4913), .Y(n4914) );
  AND2X1 U4259 ( .A(n7011), .B(n10137), .Y(n893) );
  INVX1 U4260 ( .A(n893), .Y(n4915) );
  INVX1 U4261 ( .A(n4918), .Y(n4916) );
  INVX1 U4262 ( .A(n4916), .Y(n4917) );
  AND2X1 U4263 ( .A(n7014), .B(n10137), .Y(n892) );
  INVX1 U4264 ( .A(n892), .Y(n4918) );
  INVX1 U4265 ( .A(n4921), .Y(n4919) );
  INVX1 U4266 ( .A(n4919), .Y(n4920) );
  AND2X1 U4267 ( .A(n7017), .B(n10137), .Y(n891) );
  INVX1 U4268 ( .A(n891), .Y(n4921) );
  INVX1 U4269 ( .A(n4924), .Y(n4922) );
  INVX1 U4270 ( .A(n4922), .Y(n4923) );
  AND2X1 U4271 ( .A(n7020), .B(n10137), .Y(n890) );
  INVX1 U4272 ( .A(n890), .Y(n4924) );
  INVX1 U4273 ( .A(n4927), .Y(n4925) );
  INVX1 U4274 ( .A(n4925), .Y(n4926) );
  AND2X1 U4275 ( .A(n7023), .B(n10137), .Y(n889) );
  INVX1 U4276 ( .A(n889), .Y(n4927) );
  INVX1 U4277 ( .A(n4930), .Y(n4928) );
  INVX1 U4278 ( .A(n4928), .Y(n4929) );
  AND2X1 U4279 ( .A(n7026), .B(n10137), .Y(n888) );
  INVX1 U4280 ( .A(n888), .Y(n4930) );
  INVX1 U4281 ( .A(n4933), .Y(n4931) );
  INVX1 U4282 ( .A(n4931), .Y(n4932) );
  AND2X1 U4283 ( .A(n7029), .B(n10137), .Y(n887) );
  INVX1 U4284 ( .A(n887), .Y(n4933) );
  INVX1 U4285 ( .A(n4936), .Y(n4934) );
  INVX1 U4286 ( .A(n4934), .Y(n4935) );
  AND2X1 U4287 ( .A(n7032), .B(n10137), .Y(n886) );
  INVX1 U4288 ( .A(n886), .Y(n4936) );
  INVX1 U4289 ( .A(n4939), .Y(n4937) );
  INVX1 U4290 ( .A(n4937), .Y(n4938) );
  AND2X1 U4291 ( .A(n7035), .B(n10137), .Y(n885) );
  INVX1 U4292 ( .A(n885), .Y(n4939) );
  INVX1 U4293 ( .A(n4942), .Y(n4940) );
  INVX1 U4294 ( .A(n4940), .Y(n4941) );
  AND2X1 U4295 ( .A(n7038), .B(n10137), .Y(n884) );
  INVX1 U4296 ( .A(n884), .Y(n4942) );
  INVX1 U4297 ( .A(n4945), .Y(n4943) );
  INVX1 U4298 ( .A(n4943), .Y(n4944) );
  AND2X1 U4299 ( .A(n7041), .B(n10137), .Y(n883) );
  INVX1 U4300 ( .A(n883), .Y(n4945) );
  INVX1 U4301 ( .A(n4948), .Y(n4946) );
  INVX1 U4302 ( .A(n4946), .Y(n4947) );
  AND2X1 U4303 ( .A(n7044), .B(n10137), .Y(n882) );
  INVX1 U4304 ( .A(n882), .Y(n4948) );
  INVX1 U4305 ( .A(n4951), .Y(n4949) );
  INVX1 U4306 ( .A(n4949), .Y(n4950) );
  AND2X1 U4307 ( .A(n7047), .B(n10137), .Y(n881) );
  INVX1 U4308 ( .A(n881), .Y(n4951) );
  INVX1 U4309 ( .A(n4954), .Y(n4952) );
  INVX1 U4310 ( .A(n4952), .Y(n4953) );
  AND2X1 U4311 ( .A(n7050), .B(n10137), .Y(n880) );
  INVX1 U4312 ( .A(n880), .Y(n4954) );
  INVX1 U4313 ( .A(n4957), .Y(n4955) );
  INVX1 U4314 ( .A(n4955), .Y(n4956) );
  AND2X1 U4315 ( .A(n7053), .B(n10137), .Y(n879) );
  INVX1 U4316 ( .A(n879), .Y(n4957) );
  INVX1 U4317 ( .A(n4960), .Y(n4958) );
  INVX1 U4318 ( .A(n4958), .Y(n4959) );
  AND2X1 U4319 ( .A(n7056), .B(n10137), .Y(n878) );
  INVX1 U4320 ( .A(n878), .Y(n4960) );
  INVX1 U4321 ( .A(n4963), .Y(n4961) );
  INVX1 U4322 ( .A(n4961), .Y(n4962) );
  AND2X1 U4323 ( .A(n7059), .B(n10137), .Y(n877) );
  INVX1 U4324 ( .A(n877), .Y(n4963) );
  INVX1 U4325 ( .A(n4966), .Y(n4964) );
  INVX1 U4326 ( .A(n4964), .Y(n4965) );
  AND2X1 U4327 ( .A(n7062), .B(n10137), .Y(n876) );
  INVX1 U4328 ( .A(n876), .Y(n4966) );
  INVX1 U4329 ( .A(n4969), .Y(n4967) );
  INVX1 U4330 ( .A(n4967), .Y(n4968) );
  AND2X1 U4331 ( .A(n7065), .B(n10137), .Y(n875) );
  INVX1 U4332 ( .A(n875), .Y(n4969) );
  INVX1 U4333 ( .A(n4972), .Y(n4970) );
  INVX1 U4334 ( .A(n4970), .Y(n4971) );
  AND2X1 U4335 ( .A(n7068), .B(n10137), .Y(n874) );
  INVX1 U4336 ( .A(n874), .Y(n4972) );
  INVX1 U4337 ( .A(n4975), .Y(n4973) );
  INVX1 U4338 ( .A(n4973), .Y(n4974) );
  AND2X1 U4339 ( .A(n7071), .B(n10137), .Y(n873) );
  INVX1 U4340 ( .A(n873), .Y(n4975) );
  INVX1 U4341 ( .A(n4978), .Y(n4976) );
  INVX1 U4342 ( .A(n4976), .Y(n4977) );
  AND2X1 U4343 ( .A(n7074), .B(n10137), .Y(n872) );
  INVX1 U4344 ( .A(n872), .Y(n4978) );
  INVX1 U4345 ( .A(n4981), .Y(n4979) );
  INVX1 U4346 ( .A(n4979), .Y(n4980) );
  AND2X1 U4347 ( .A(n7077), .B(n10137), .Y(n871) );
  INVX1 U4348 ( .A(n871), .Y(n4981) );
  INVX1 U4349 ( .A(n4984), .Y(n4982) );
  INVX1 U4350 ( .A(n4982), .Y(n4983) );
  AND2X1 U4351 ( .A(n7080), .B(n10137), .Y(n870) );
  INVX1 U4352 ( .A(n870), .Y(n4984) );
  INVX1 U4353 ( .A(n4987), .Y(n4985) );
  INVX1 U4354 ( .A(n4985), .Y(n4986) );
  AND2X1 U4355 ( .A(n7083), .B(n10137), .Y(n869) );
  INVX1 U4356 ( .A(n869), .Y(n4987) );
  INVX1 U4357 ( .A(n4990), .Y(n4988) );
  INVX1 U4358 ( .A(n4988), .Y(n4989) );
  AND2X1 U4359 ( .A(n7086), .B(n10137), .Y(n868) );
  INVX1 U4360 ( .A(n868), .Y(n4990) );
  INVX1 U4361 ( .A(n4993), .Y(n4991) );
  INVX1 U4362 ( .A(n4991), .Y(n4992) );
  AND2X1 U4363 ( .A(n7089), .B(n10137), .Y(n867) );
  INVX1 U4364 ( .A(n867), .Y(n4993) );
  INVX1 U4365 ( .A(n4996), .Y(n4994) );
  INVX1 U4366 ( .A(n4994), .Y(n4995) );
  AND2X1 U4367 ( .A(n7092), .B(n10137), .Y(n866) );
  INVX1 U4368 ( .A(n866), .Y(n4996) );
  INVX1 U4369 ( .A(n4999), .Y(n4997) );
  INVX1 U4370 ( .A(n4997), .Y(n4998) );
  AND2X1 U4371 ( .A(n7095), .B(n10137), .Y(n865) );
  INVX1 U4372 ( .A(n865), .Y(n4999) );
  INVX1 U4373 ( .A(n5002), .Y(n5000) );
  INVX1 U4374 ( .A(n5000), .Y(n5001) );
  AND2X1 U4375 ( .A(n7098), .B(n10137), .Y(n864) );
  INVX1 U4376 ( .A(n864), .Y(n5002) );
  INVX1 U4377 ( .A(n5005), .Y(n5003) );
  INVX1 U4378 ( .A(n5003), .Y(n5004) );
  AND2X1 U4379 ( .A(n7101), .B(n10137), .Y(n863) );
  INVX1 U4380 ( .A(n863), .Y(n5005) );
  INVX1 U4381 ( .A(n5008), .Y(n5006) );
  INVX1 U4382 ( .A(n5006), .Y(n5007) );
  AND2X1 U4383 ( .A(n7104), .B(n10137), .Y(n862) );
  INVX1 U4384 ( .A(n862), .Y(n5008) );
  INVX1 U4385 ( .A(n5011), .Y(n5009) );
  INVX1 U4386 ( .A(n5009), .Y(n5010) );
  AND2X1 U4387 ( .A(n7107), .B(n10137), .Y(n861) );
  INVX1 U4388 ( .A(n861), .Y(n5011) );
  INVX1 U4389 ( .A(n5014), .Y(n5012) );
  INVX1 U4390 ( .A(n5012), .Y(n5013) );
  AND2X1 U4391 ( .A(n9150), .B(n824), .Y(n858) );
  INVX1 U4392 ( .A(n858), .Y(n5014) );
  INVX1 U4393 ( .A(n5017), .Y(n5015) );
  INVX1 U4394 ( .A(n5015), .Y(n5016) );
  AND2X1 U4395 ( .A(n9153), .B(n824), .Y(n857) );
  INVX1 U4396 ( .A(n857), .Y(n5017) );
  INVX1 U4397 ( .A(n5020), .Y(n5018) );
  INVX1 U4398 ( .A(n5018), .Y(n5019) );
  AND2X1 U4399 ( .A(n9156), .B(n824), .Y(n856) );
  INVX1 U4400 ( .A(n856), .Y(n5020) );
  INVX1 U4401 ( .A(n5023), .Y(n5021) );
  INVX1 U4402 ( .A(n5021), .Y(n5022) );
  AND2X1 U4403 ( .A(n9159), .B(n824), .Y(n855) );
  INVX1 U4404 ( .A(n855), .Y(n5023) );
  INVX1 U4405 ( .A(n5026), .Y(n5024) );
  INVX1 U4406 ( .A(n5024), .Y(n5025) );
  AND2X1 U4407 ( .A(n9162), .B(n824), .Y(n854) );
  INVX1 U4408 ( .A(n854), .Y(n5026) );
  INVX1 U4409 ( .A(n5029), .Y(n5027) );
  INVX1 U4410 ( .A(n5027), .Y(n5028) );
  AND2X1 U4411 ( .A(n9165), .B(n824), .Y(n853) );
  INVX1 U4412 ( .A(n853), .Y(n5029) );
  INVX1 U4413 ( .A(n5032), .Y(n5030) );
  INVX1 U4414 ( .A(n5030), .Y(n5031) );
  AND2X1 U4415 ( .A(n9168), .B(n824), .Y(n852) );
  INVX1 U4416 ( .A(n852), .Y(n5032) );
  INVX1 U4417 ( .A(n5035), .Y(n5033) );
  INVX1 U4418 ( .A(n5033), .Y(n5034) );
  AND2X1 U4419 ( .A(n9171), .B(n824), .Y(n851) );
  INVX1 U4420 ( .A(n851), .Y(n5035) );
  INVX1 U4421 ( .A(n5038), .Y(n5036) );
  INVX1 U4422 ( .A(n5036), .Y(n5037) );
  AND2X1 U4423 ( .A(n9174), .B(n824), .Y(n850) );
  INVX1 U4424 ( .A(n850), .Y(n5038) );
  INVX1 U4425 ( .A(n5041), .Y(n5039) );
  INVX1 U4426 ( .A(n5039), .Y(n5040) );
  AND2X1 U4427 ( .A(n9177), .B(n824), .Y(n849) );
  INVX1 U4428 ( .A(n849), .Y(n5041) );
  INVX1 U4429 ( .A(n5044), .Y(n5042) );
  INVX1 U4430 ( .A(n5042), .Y(n5043) );
  AND2X1 U4431 ( .A(n9180), .B(n824), .Y(n848) );
  INVX1 U4432 ( .A(n848), .Y(n5044) );
  INVX1 U4433 ( .A(n5047), .Y(n5045) );
  INVX1 U4434 ( .A(n5045), .Y(n5046) );
  AND2X1 U4435 ( .A(n9183), .B(n824), .Y(n847) );
  INVX1 U4436 ( .A(n847), .Y(n5047) );
  INVX1 U4437 ( .A(n5050), .Y(n5048) );
  INVX1 U4438 ( .A(n5048), .Y(n5049) );
  AND2X1 U4439 ( .A(n9186), .B(n824), .Y(n846) );
  INVX1 U4440 ( .A(n846), .Y(n5050) );
  INVX1 U4441 ( .A(n5053), .Y(n5051) );
  INVX1 U4442 ( .A(n5051), .Y(n5052) );
  AND2X1 U4443 ( .A(n9189), .B(n824), .Y(n845) );
  INVX1 U4444 ( .A(n845), .Y(n5053) );
  INVX1 U4445 ( .A(n5056), .Y(n5054) );
  INVX1 U4446 ( .A(n5054), .Y(n5055) );
  AND2X1 U4447 ( .A(n9192), .B(n824), .Y(n844) );
  INVX1 U4448 ( .A(n844), .Y(n5056) );
  INVX1 U4449 ( .A(n5059), .Y(n5057) );
  INVX1 U4450 ( .A(n5057), .Y(n5058) );
  AND2X1 U4451 ( .A(n9195), .B(n824), .Y(n843) );
  INVX1 U4452 ( .A(n843), .Y(n5059) );
  INVX1 U4453 ( .A(n5062), .Y(n5060) );
  INVX1 U4454 ( .A(n5060), .Y(n5061) );
  AND2X1 U4455 ( .A(n9198), .B(n824), .Y(n842) );
  INVX1 U4456 ( .A(n842), .Y(n5062) );
  INVX1 U4457 ( .A(n5065), .Y(n5063) );
  INVX1 U4458 ( .A(n5063), .Y(n5064) );
  AND2X1 U4459 ( .A(n9201), .B(n824), .Y(n841) );
  INVX1 U4460 ( .A(n841), .Y(n5065) );
  INVX1 U4461 ( .A(n5068), .Y(n5066) );
  INVX1 U4462 ( .A(n5066), .Y(n5067) );
  AND2X1 U4463 ( .A(n9204), .B(n824), .Y(n840) );
  INVX1 U4464 ( .A(n840), .Y(n5068) );
  INVX1 U4465 ( .A(n5071), .Y(n5069) );
  INVX1 U4466 ( .A(n5069), .Y(n5070) );
  AND2X1 U4467 ( .A(n9207), .B(n824), .Y(n839) );
  INVX1 U4468 ( .A(n839), .Y(n5071) );
  INVX1 U4469 ( .A(n5074), .Y(n5072) );
  INVX1 U4470 ( .A(n5072), .Y(n5073) );
  AND2X1 U4471 ( .A(n9210), .B(n824), .Y(n838) );
  INVX1 U4472 ( .A(n838), .Y(n5074) );
  INVX1 U4473 ( .A(n5077), .Y(n5075) );
  INVX1 U4474 ( .A(n5075), .Y(n5076) );
  AND2X1 U4475 ( .A(n9213), .B(n824), .Y(n837) );
  INVX1 U4476 ( .A(n837), .Y(n5077) );
  INVX1 U4477 ( .A(n5080), .Y(n5078) );
  INVX1 U4478 ( .A(n5078), .Y(n5079) );
  AND2X1 U4479 ( .A(n9216), .B(n824), .Y(n836) );
  INVX1 U4480 ( .A(n836), .Y(n5080) );
  INVX1 U4481 ( .A(n5083), .Y(n5081) );
  INVX1 U4482 ( .A(n5081), .Y(n5082) );
  AND2X1 U4483 ( .A(n9219), .B(n824), .Y(n835) );
  INVX1 U4484 ( .A(n835), .Y(n5083) );
  INVX1 U4485 ( .A(n5086), .Y(n5084) );
  INVX1 U4486 ( .A(n5084), .Y(n5085) );
  AND2X1 U4487 ( .A(n9222), .B(n824), .Y(n834) );
  INVX1 U4488 ( .A(n834), .Y(n5086) );
  INVX1 U4489 ( .A(n5089), .Y(n5087) );
  INVX1 U4490 ( .A(n5087), .Y(n5088) );
  AND2X1 U4491 ( .A(n9225), .B(n824), .Y(n833) );
  INVX1 U4492 ( .A(n833), .Y(n5089) );
  INVX1 U4493 ( .A(n5092), .Y(n5090) );
  INVX1 U4494 ( .A(n5090), .Y(n5091) );
  AND2X1 U4495 ( .A(n9228), .B(n824), .Y(n832) );
  INVX1 U4496 ( .A(n832), .Y(n5092) );
  INVX1 U4497 ( .A(n5095), .Y(n5093) );
  INVX1 U4498 ( .A(n5093), .Y(n5094) );
  AND2X1 U4499 ( .A(n9231), .B(n824), .Y(n831) );
  INVX1 U4500 ( .A(n831), .Y(n5095) );
  INVX1 U4501 ( .A(n5098), .Y(n5096) );
  INVX1 U4502 ( .A(n5096), .Y(n5097) );
  AND2X1 U4503 ( .A(n9234), .B(n824), .Y(n830) );
  INVX1 U4504 ( .A(n830), .Y(n5098) );
  INVX1 U4505 ( .A(n5101), .Y(n5099) );
  INVX1 U4506 ( .A(n5099), .Y(n5100) );
  AND2X1 U4507 ( .A(n9237), .B(n824), .Y(n829) );
  INVX1 U4508 ( .A(n829), .Y(n5101) );
  INVX1 U4509 ( .A(n5104), .Y(n5102) );
  INVX1 U4510 ( .A(n5102), .Y(n5103) );
  AND2X1 U4511 ( .A(n9240), .B(n824), .Y(n828) );
  INVX1 U4512 ( .A(n828), .Y(n5104) );
  INVX1 U4513 ( .A(n5107), .Y(n5105) );
  INVX1 U4514 ( .A(n5105), .Y(n5106) );
  AND2X1 U4515 ( .A(n9243), .B(n824), .Y(n827) );
  INVX1 U4516 ( .A(n827), .Y(n5107) );
  INVX1 U4517 ( .A(n5110), .Y(n5108) );
  INVX1 U4518 ( .A(n5108), .Y(n5109) );
  AND2X1 U4519 ( .A(n9246), .B(n824), .Y(n826) );
  INVX1 U4520 ( .A(n826), .Y(n5110) );
  INVX1 U4521 ( .A(n5113), .Y(n5111) );
  INVX1 U4522 ( .A(n5111), .Y(n5112) );
  AND2X1 U4523 ( .A(n9249), .B(n824), .Y(n825) );
  INVX1 U4524 ( .A(n825), .Y(n5113) );
  INVX1 U4525 ( .A(n5116), .Y(n5114) );
  INVX1 U4526 ( .A(n5114), .Y(n5115) );
  AND2X1 U4527 ( .A(n7620), .B(n10511), .Y(n823) );
  INVX1 U4528 ( .A(n823), .Y(n5116) );
  INVX1 U4529 ( .A(n5119), .Y(n5117) );
  INVX1 U4530 ( .A(n5117), .Y(n5118) );
  AND2X1 U4531 ( .A(n7623), .B(n10511), .Y(n822) );
  INVX1 U4532 ( .A(n822), .Y(n5119) );
  INVX1 U4533 ( .A(n5122), .Y(n5120) );
  INVX1 U4534 ( .A(n5120), .Y(n5121) );
  AND2X1 U4535 ( .A(n7626), .B(n10511), .Y(n821) );
  INVX1 U4536 ( .A(n821), .Y(n5122) );
  INVX1 U4537 ( .A(n5125), .Y(n5123) );
  INVX1 U4538 ( .A(n5123), .Y(n5124) );
  AND2X1 U4539 ( .A(n7629), .B(n10511), .Y(n820) );
  INVX1 U4540 ( .A(n820), .Y(n5125) );
  INVX1 U4541 ( .A(n5128), .Y(n5126) );
  INVX1 U4542 ( .A(n5126), .Y(n5127) );
  AND2X1 U4543 ( .A(n7632), .B(n10511), .Y(n819) );
  INVX1 U4544 ( .A(n819), .Y(n5128) );
  INVX1 U4545 ( .A(n5131), .Y(n5129) );
  INVX1 U4546 ( .A(n5129), .Y(n5130) );
  AND2X1 U4547 ( .A(n7635), .B(n10511), .Y(n818) );
  INVX1 U4548 ( .A(n818), .Y(n5131) );
  INVX1 U4549 ( .A(n5134), .Y(n5132) );
  INVX1 U4550 ( .A(n5132), .Y(n5133) );
  AND2X1 U4551 ( .A(n7638), .B(n10511), .Y(n817) );
  INVX1 U4552 ( .A(n817), .Y(n5134) );
  INVX1 U4553 ( .A(n5137), .Y(n5135) );
  INVX1 U4554 ( .A(n5135), .Y(n5136) );
  AND2X1 U4555 ( .A(n7641), .B(n10511), .Y(n816) );
  INVX1 U4556 ( .A(n816), .Y(n5137) );
  INVX1 U4557 ( .A(n5140), .Y(n5138) );
  INVX1 U4558 ( .A(n5138), .Y(n5139) );
  AND2X1 U4559 ( .A(n7644), .B(n10511), .Y(n815) );
  INVX1 U4560 ( .A(n815), .Y(n5140) );
  INVX1 U4561 ( .A(n5143), .Y(n5141) );
  INVX1 U4562 ( .A(n5141), .Y(n5142) );
  AND2X1 U4563 ( .A(n7647), .B(n10511), .Y(n814) );
  INVX1 U4564 ( .A(n814), .Y(n5143) );
  INVX1 U4565 ( .A(n5146), .Y(n5144) );
  INVX1 U4566 ( .A(n5144), .Y(n5145) );
  AND2X1 U4567 ( .A(n7650), .B(n10511), .Y(n813) );
  INVX1 U4568 ( .A(n813), .Y(n5146) );
  INVX1 U4569 ( .A(n5149), .Y(n5147) );
  INVX1 U4570 ( .A(n5147), .Y(n5148) );
  AND2X1 U4571 ( .A(n7653), .B(n10511), .Y(n812) );
  INVX1 U4572 ( .A(n812), .Y(n5149) );
  INVX1 U4573 ( .A(n5152), .Y(n5150) );
  INVX1 U4574 ( .A(n5150), .Y(n5151) );
  AND2X1 U4575 ( .A(n7656), .B(n10511), .Y(n811) );
  INVX1 U4576 ( .A(n811), .Y(n5152) );
  INVX1 U4577 ( .A(n5155), .Y(n5153) );
  INVX1 U4578 ( .A(n5153), .Y(n5154) );
  AND2X1 U4579 ( .A(n7659), .B(n10511), .Y(n810) );
  INVX1 U4580 ( .A(n810), .Y(n5155) );
  INVX1 U4581 ( .A(n5158), .Y(n5156) );
  INVX1 U4582 ( .A(n5156), .Y(n5157) );
  AND2X1 U4583 ( .A(n7662), .B(n10511), .Y(n809) );
  INVX1 U4584 ( .A(n809), .Y(n5158) );
  INVX1 U4585 ( .A(n5161), .Y(n5159) );
  INVX1 U4586 ( .A(n5159), .Y(n5160) );
  AND2X1 U4587 ( .A(n7665), .B(n10511), .Y(n808) );
  INVX1 U4588 ( .A(n808), .Y(n5161) );
  INVX1 U4589 ( .A(n5164), .Y(n5162) );
  INVX1 U4590 ( .A(n5162), .Y(n5163) );
  AND2X1 U4591 ( .A(n7668), .B(n10511), .Y(n807) );
  INVX1 U4592 ( .A(n807), .Y(n5164) );
  INVX1 U4593 ( .A(n5167), .Y(n5165) );
  INVX1 U4594 ( .A(n5165), .Y(n5166) );
  AND2X1 U4595 ( .A(n7671), .B(n10511), .Y(n806) );
  INVX1 U4596 ( .A(n806), .Y(n5167) );
  INVX1 U4597 ( .A(n5170), .Y(n5168) );
  INVX1 U4598 ( .A(n5168), .Y(n5169) );
  AND2X1 U4599 ( .A(n7674), .B(n10511), .Y(n805) );
  INVX1 U4600 ( .A(n805), .Y(n5170) );
  INVX1 U4601 ( .A(n5173), .Y(n5171) );
  INVX1 U4602 ( .A(n5171), .Y(n5172) );
  AND2X1 U4603 ( .A(n7677), .B(n10511), .Y(n804) );
  INVX1 U4604 ( .A(n804), .Y(n5173) );
  INVX1 U4605 ( .A(n5176), .Y(n5174) );
  INVX1 U4606 ( .A(n5174), .Y(n5175) );
  AND2X1 U4607 ( .A(n7680), .B(n10511), .Y(n803) );
  INVX1 U4608 ( .A(n803), .Y(n5176) );
  INVX1 U4609 ( .A(n5179), .Y(n5177) );
  INVX1 U4610 ( .A(n5177), .Y(n5178) );
  AND2X1 U4611 ( .A(n7683), .B(n10511), .Y(n802) );
  INVX1 U4612 ( .A(n802), .Y(n5179) );
  INVX1 U4613 ( .A(n5182), .Y(n5180) );
  INVX1 U4614 ( .A(n5180), .Y(n5181) );
  AND2X1 U4615 ( .A(n7686), .B(n10511), .Y(n801) );
  INVX1 U4616 ( .A(n801), .Y(n5182) );
  INVX1 U4617 ( .A(n5185), .Y(n5183) );
  INVX1 U4618 ( .A(n5183), .Y(n5184) );
  AND2X1 U4619 ( .A(n7689), .B(n10511), .Y(n800) );
  INVX1 U4620 ( .A(n800), .Y(n5185) );
  INVX1 U4621 ( .A(n5188), .Y(n5186) );
  INVX1 U4622 ( .A(n5186), .Y(n5187) );
  AND2X1 U4623 ( .A(n7692), .B(n10511), .Y(n799) );
  INVX1 U4624 ( .A(n799), .Y(n5188) );
  INVX1 U4625 ( .A(n5191), .Y(n5189) );
  INVX1 U4626 ( .A(n5189), .Y(n5190) );
  AND2X1 U4627 ( .A(n7695), .B(n10511), .Y(n798) );
  INVX1 U4628 ( .A(n798), .Y(n5191) );
  INVX1 U4629 ( .A(n5194), .Y(n5192) );
  INVX1 U4630 ( .A(n5192), .Y(n5193) );
  AND2X1 U4631 ( .A(n7698), .B(n10511), .Y(n797) );
  INVX1 U4632 ( .A(n797), .Y(n5194) );
  INVX1 U4633 ( .A(n5197), .Y(n5195) );
  INVX1 U4634 ( .A(n5195), .Y(n5196) );
  AND2X1 U4635 ( .A(n7701), .B(n10511), .Y(n796) );
  INVX1 U4636 ( .A(n796), .Y(n5197) );
  INVX1 U4637 ( .A(n5200), .Y(n5198) );
  INVX1 U4638 ( .A(n5198), .Y(n5199) );
  AND2X1 U4639 ( .A(n7704), .B(n10511), .Y(n795) );
  INVX1 U4640 ( .A(n795), .Y(n5200) );
  INVX1 U4641 ( .A(n5203), .Y(n5201) );
  INVX1 U4642 ( .A(n5201), .Y(n5202) );
  AND2X1 U4643 ( .A(n7707), .B(n10511), .Y(n794) );
  INVX1 U4644 ( .A(n794), .Y(n5203) );
  INVX1 U4645 ( .A(n5206), .Y(n5204) );
  INVX1 U4646 ( .A(n5204), .Y(n5205) );
  AND2X1 U4647 ( .A(n7710), .B(n10511), .Y(n793) );
  INVX1 U4648 ( .A(n793), .Y(n5206) );
  INVX1 U4649 ( .A(n5209), .Y(n5207) );
  INVX1 U4650 ( .A(n5207), .Y(n5208) );
  AND2X1 U4651 ( .A(n7713), .B(n10511), .Y(n792) );
  INVX1 U4652 ( .A(n792), .Y(n5209) );
  INVX1 U4653 ( .A(n5212), .Y(n5210) );
  INVX1 U4654 ( .A(n5210), .Y(n5211) );
  AND2X1 U4655 ( .A(n7716), .B(n10511), .Y(n791) );
  INVX1 U4656 ( .A(n791), .Y(n5212) );
  INVX1 U4657 ( .A(n5215), .Y(n5213) );
  INVX1 U4658 ( .A(n5213), .Y(n5214) );
  AND2X1 U4659 ( .A(n7719), .B(n10511), .Y(n790) );
  INVX1 U4660 ( .A(n790), .Y(n5215) );
  INVX1 U4661 ( .A(n5218), .Y(n5216) );
  INVX1 U4662 ( .A(n5216), .Y(n5217) );
  AND2X1 U4663 ( .A(n9252), .B(n10517), .Y(n788) );
  INVX1 U4664 ( .A(n788), .Y(n5218) );
  INVX1 U4665 ( .A(n5221), .Y(n5219) );
  INVX1 U4666 ( .A(n5219), .Y(n5220) );
  AND2X1 U4667 ( .A(n9255), .B(n10517), .Y(n787) );
  INVX1 U4668 ( .A(n787), .Y(n5221) );
  INVX1 U4669 ( .A(n5224), .Y(n5222) );
  INVX1 U4670 ( .A(n5222), .Y(n5223) );
  AND2X1 U4671 ( .A(n9258), .B(n10517), .Y(n786) );
  INVX1 U4672 ( .A(n786), .Y(n5224) );
  INVX1 U4673 ( .A(n5227), .Y(n5225) );
  INVX1 U4674 ( .A(n5225), .Y(n5226) );
  AND2X1 U4675 ( .A(n9261), .B(n10517), .Y(n785) );
  INVX1 U4676 ( .A(n785), .Y(n5227) );
  INVX1 U4677 ( .A(n5230), .Y(n5228) );
  INVX1 U4678 ( .A(n5228), .Y(n5229) );
  AND2X1 U4679 ( .A(n9264), .B(n10517), .Y(n784) );
  INVX1 U4680 ( .A(n784), .Y(n5230) );
  INVX1 U4681 ( .A(n5233), .Y(n5231) );
  INVX1 U4682 ( .A(n5231), .Y(n5232) );
  AND2X1 U4683 ( .A(n9267), .B(n10517), .Y(n783) );
  INVX1 U4684 ( .A(n783), .Y(n5233) );
  INVX1 U4685 ( .A(n5236), .Y(n5234) );
  INVX1 U4686 ( .A(n5234), .Y(n5235) );
  AND2X1 U4687 ( .A(n9270), .B(n10517), .Y(n782) );
  INVX1 U4688 ( .A(n782), .Y(n5236) );
  INVX1 U4689 ( .A(n5239), .Y(n5237) );
  INVX1 U4690 ( .A(n5237), .Y(n5238) );
  AND2X1 U4691 ( .A(n9273), .B(n10517), .Y(n781) );
  INVX1 U4692 ( .A(n781), .Y(n5239) );
  INVX1 U4693 ( .A(n5242), .Y(n5240) );
  INVX1 U4694 ( .A(n5240), .Y(n5241) );
  AND2X1 U4695 ( .A(n9276), .B(n10517), .Y(n780) );
  INVX1 U4696 ( .A(n780), .Y(n5242) );
  INVX1 U4697 ( .A(n5245), .Y(n5243) );
  INVX1 U4698 ( .A(n5243), .Y(n5244) );
  AND2X1 U4699 ( .A(n9279), .B(n10517), .Y(n779) );
  INVX1 U4700 ( .A(n779), .Y(n5245) );
  INVX1 U4701 ( .A(n5248), .Y(n5246) );
  INVX1 U4702 ( .A(n5246), .Y(n5247) );
  AND2X1 U4703 ( .A(n9282), .B(n10517), .Y(n778) );
  INVX1 U4704 ( .A(n778), .Y(n5248) );
  INVX1 U4705 ( .A(n5251), .Y(n5249) );
  INVX1 U4706 ( .A(n5249), .Y(n5250) );
  AND2X1 U4707 ( .A(n9285), .B(n10517), .Y(n777) );
  INVX1 U4708 ( .A(n777), .Y(n5251) );
  INVX1 U4709 ( .A(n5254), .Y(n5252) );
  INVX1 U4710 ( .A(n5252), .Y(n5253) );
  AND2X1 U4711 ( .A(n9288), .B(n10517), .Y(n776) );
  INVX1 U4712 ( .A(n776), .Y(n5254) );
  INVX1 U4713 ( .A(n5257), .Y(n5255) );
  INVX1 U4714 ( .A(n5255), .Y(n5256) );
  AND2X1 U4715 ( .A(n9291), .B(n10517), .Y(n775) );
  INVX1 U4716 ( .A(n775), .Y(n5257) );
  INVX1 U4717 ( .A(n5260), .Y(n5258) );
  INVX1 U4718 ( .A(n5258), .Y(n5259) );
  AND2X1 U4719 ( .A(n9294), .B(n10517), .Y(n774) );
  INVX1 U4720 ( .A(n774), .Y(n5260) );
  INVX1 U4721 ( .A(n5263), .Y(n5261) );
  INVX1 U4722 ( .A(n5261), .Y(n5262) );
  AND2X1 U4723 ( .A(n9297), .B(n10517), .Y(n773) );
  INVX1 U4724 ( .A(n773), .Y(n5263) );
  INVX1 U4725 ( .A(n5266), .Y(n5264) );
  INVX1 U4726 ( .A(n5264), .Y(n5265) );
  AND2X1 U4727 ( .A(n9300), .B(n10517), .Y(n772) );
  INVX1 U4728 ( .A(n772), .Y(n5266) );
  INVX1 U4729 ( .A(n5269), .Y(n5267) );
  INVX1 U4730 ( .A(n5267), .Y(n5268) );
  AND2X1 U4731 ( .A(n9303), .B(n10517), .Y(n771) );
  INVX1 U4732 ( .A(n771), .Y(n5269) );
  INVX1 U4733 ( .A(n5272), .Y(n5270) );
  INVX1 U4734 ( .A(n5270), .Y(n5271) );
  AND2X1 U4735 ( .A(n9306), .B(n10517), .Y(n770) );
  INVX1 U4736 ( .A(n770), .Y(n5272) );
  INVX1 U4737 ( .A(n5275), .Y(n5273) );
  INVX1 U4738 ( .A(n5273), .Y(n5274) );
  AND2X1 U4739 ( .A(n9309), .B(n10517), .Y(n769) );
  INVX1 U4740 ( .A(n769), .Y(n5275) );
  INVX1 U4741 ( .A(n5278), .Y(n5276) );
  INVX1 U4742 ( .A(n5276), .Y(n5277) );
  AND2X1 U4743 ( .A(n9312), .B(n10517), .Y(n768) );
  INVX1 U4744 ( .A(n768), .Y(n5278) );
  INVX1 U4745 ( .A(n5281), .Y(n5279) );
  INVX1 U4746 ( .A(n5279), .Y(n5280) );
  AND2X1 U4747 ( .A(n9315), .B(n10517), .Y(n767) );
  INVX1 U4748 ( .A(n767), .Y(n5281) );
  INVX1 U4749 ( .A(n5284), .Y(n5282) );
  INVX1 U4750 ( .A(n5282), .Y(n5283) );
  AND2X1 U4751 ( .A(n9318), .B(n10517), .Y(n766) );
  INVX1 U4752 ( .A(n766), .Y(n5284) );
  INVX1 U4753 ( .A(n5287), .Y(n5285) );
  INVX1 U4754 ( .A(n5285), .Y(n5286) );
  AND2X1 U4755 ( .A(n9321), .B(n10517), .Y(n765) );
  INVX1 U4756 ( .A(n765), .Y(n5287) );
  INVX1 U4757 ( .A(n5290), .Y(n5288) );
  INVX1 U4758 ( .A(n5288), .Y(n5289) );
  AND2X1 U4759 ( .A(n9324), .B(n10517), .Y(n764) );
  INVX1 U4760 ( .A(n764), .Y(n5290) );
  INVX1 U4761 ( .A(n5293), .Y(n5291) );
  INVX1 U4762 ( .A(n5291), .Y(n5292) );
  AND2X1 U4763 ( .A(n9327), .B(n10517), .Y(n763) );
  INVX1 U4764 ( .A(n763), .Y(n5293) );
  INVX1 U4765 ( .A(n5296), .Y(n5294) );
  INVX1 U4766 ( .A(n5294), .Y(n5295) );
  AND2X1 U4767 ( .A(n9330), .B(n10517), .Y(n762) );
  INVX1 U4768 ( .A(n762), .Y(n5296) );
  INVX1 U4769 ( .A(n5299), .Y(n5297) );
  INVX1 U4770 ( .A(n5297), .Y(n5298) );
  AND2X1 U4771 ( .A(n9333), .B(n10517), .Y(n761) );
  INVX1 U4772 ( .A(n761), .Y(n5299) );
  INVX1 U4773 ( .A(n5302), .Y(n5300) );
  INVX1 U4774 ( .A(n5300), .Y(n5301) );
  AND2X1 U4775 ( .A(n9336), .B(n10517), .Y(n760) );
  INVX1 U4776 ( .A(n760), .Y(n5302) );
  INVX1 U4777 ( .A(n5305), .Y(n5303) );
  INVX1 U4778 ( .A(n5303), .Y(n5304) );
  AND2X1 U4779 ( .A(n9339), .B(n10517), .Y(n759) );
  INVX1 U4780 ( .A(n759), .Y(n5305) );
  INVX1 U4781 ( .A(n5308), .Y(n5306) );
  INVX1 U4782 ( .A(n5306), .Y(n5307) );
  AND2X1 U4783 ( .A(n9342), .B(n10517), .Y(n758) );
  INVX1 U4784 ( .A(n758), .Y(n5308) );
  INVX1 U4785 ( .A(n5311), .Y(n5309) );
  INVX1 U4786 ( .A(n5309), .Y(n5310) );
  AND2X1 U4787 ( .A(n9345), .B(n10517), .Y(n757) );
  INVX1 U4788 ( .A(n757), .Y(n5311) );
  INVX1 U4789 ( .A(n5314), .Y(n5312) );
  INVX1 U4790 ( .A(n5312), .Y(n5313) );
  AND2X1 U4791 ( .A(n9348), .B(n10517), .Y(n756) );
  INVX1 U4792 ( .A(n756), .Y(n5314) );
  INVX1 U4793 ( .A(n5317), .Y(n5315) );
  INVX1 U4794 ( .A(n5315), .Y(n5316) );
  AND2X1 U4795 ( .A(n9351), .B(n10517), .Y(n755) );
  INVX1 U4796 ( .A(n755), .Y(n5317) );
  INVX1 U4797 ( .A(n5320), .Y(n5318) );
  INVX1 U4798 ( .A(n5318), .Y(n5319) );
  AND2X1 U4799 ( .A(n7722), .B(n719), .Y(n753) );
  INVX1 U4800 ( .A(n753), .Y(n5320) );
  INVX1 U4801 ( .A(n5323), .Y(n5321) );
  INVX1 U4802 ( .A(n5321), .Y(n5322) );
  AND2X1 U4803 ( .A(n7725), .B(n719), .Y(n752) );
  INVX1 U4804 ( .A(n752), .Y(n5323) );
  INVX1 U4805 ( .A(n5326), .Y(n5324) );
  INVX1 U4806 ( .A(n5324), .Y(n5325) );
  AND2X1 U4807 ( .A(n7728), .B(n719), .Y(n751) );
  INVX1 U4808 ( .A(n751), .Y(n5326) );
  INVX1 U4809 ( .A(n5329), .Y(n5327) );
  INVX1 U4810 ( .A(n5327), .Y(n5328) );
  AND2X1 U4811 ( .A(n7731), .B(n719), .Y(n750) );
  INVX1 U4812 ( .A(n750), .Y(n5329) );
  INVX1 U4813 ( .A(n5332), .Y(n5330) );
  INVX1 U4814 ( .A(n5330), .Y(n5331) );
  AND2X1 U4815 ( .A(n7734), .B(n719), .Y(n749) );
  INVX1 U4816 ( .A(n749), .Y(n5332) );
  INVX1 U4817 ( .A(n5335), .Y(n5333) );
  INVX1 U4818 ( .A(n5333), .Y(n5334) );
  AND2X1 U4819 ( .A(n7737), .B(n719), .Y(n748) );
  INVX1 U4820 ( .A(n748), .Y(n5335) );
  INVX1 U4821 ( .A(n5338), .Y(n5336) );
  INVX1 U4822 ( .A(n5336), .Y(n5337) );
  AND2X1 U4823 ( .A(n7740), .B(n719), .Y(n747) );
  INVX1 U4824 ( .A(n747), .Y(n5338) );
  INVX1 U4825 ( .A(n5341), .Y(n5339) );
  INVX1 U4826 ( .A(n5339), .Y(n5340) );
  AND2X1 U4827 ( .A(n7743), .B(n719), .Y(n746) );
  INVX1 U4828 ( .A(n746), .Y(n5341) );
  INVX1 U4829 ( .A(n5344), .Y(n5342) );
  INVX1 U4830 ( .A(n5342), .Y(n5343) );
  AND2X1 U4831 ( .A(n7746), .B(n719), .Y(n745) );
  INVX1 U4832 ( .A(n745), .Y(n5344) );
  INVX1 U4833 ( .A(n5347), .Y(n5345) );
  INVX1 U4834 ( .A(n5345), .Y(n5346) );
  AND2X1 U4835 ( .A(n7749), .B(n719), .Y(n744) );
  INVX1 U4836 ( .A(n744), .Y(n5347) );
  INVX1 U4837 ( .A(n5350), .Y(n5348) );
  INVX1 U4838 ( .A(n5348), .Y(n5349) );
  AND2X1 U4839 ( .A(n7752), .B(n719), .Y(n743) );
  INVX1 U4840 ( .A(n743), .Y(n5350) );
  INVX1 U4841 ( .A(n5353), .Y(n5351) );
  INVX1 U4842 ( .A(n5351), .Y(n5352) );
  AND2X1 U4843 ( .A(n7755), .B(n719), .Y(n742) );
  INVX1 U4844 ( .A(n742), .Y(n5353) );
  INVX1 U4845 ( .A(n5356), .Y(n5354) );
  INVX1 U4846 ( .A(n5354), .Y(n5355) );
  AND2X1 U4847 ( .A(n7758), .B(n719), .Y(n741) );
  INVX1 U4848 ( .A(n741), .Y(n5356) );
  INVX1 U4849 ( .A(n5359), .Y(n5357) );
  INVX1 U4850 ( .A(n5357), .Y(n5358) );
  AND2X1 U4851 ( .A(n7761), .B(n719), .Y(n740) );
  INVX1 U4852 ( .A(n740), .Y(n5359) );
  INVX1 U4853 ( .A(n5362), .Y(n5360) );
  INVX1 U4854 ( .A(n5360), .Y(n5361) );
  AND2X1 U4855 ( .A(n7764), .B(n719), .Y(n739) );
  INVX1 U4856 ( .A(n739), .Y(n5362) );
  INVX1 U4857 ( .A(n5365), .Y(n5363) );
  INVX1 U4858 ( .A(n5363), .Y(n5364) );
  AND2X1 U4859 ( .A(n7767), .B(n719), .Y(n738) );
  INVX1 U4860 ( .A(n738), .Y(n5365) );
  INVX1 U4861 ( .A(n5368), .Y(n5366) );
  INVX1 U4862 ( .A(n5366), .Y(n5367) );
  AND2X1 U4863 ( .A(n7770), .B(n719), .Y(n737) );
  INVX1 U4864 ( .A(n737), .Y(n5368) );
  INVX1 U4865 ( .A(n5371), .Y(n5369) );
  INVX1 U4866 ( .A(n5369), .Y(n5370) );
  AND2X1 U4867 ( .A(n7773), .B(n719), .Y(n736) );
  INVX1 U4868 ( .A(n736), .Y(n5371) );
  INVX1 U4869 ( .A(n5374), .Y(n5372) );
  INVX1 U4870 ( .A(n5372), .Y(n5373) );
  AND2X1 U4871 ( .A(n7776), .B(n719), .Y(n735) );
  INVX1 U4872 ( .A(n735), .Y(n5374) );
  INVX1 U4873 ( .A(n5377), .Y(n5375) );
  INVX1 U4874 ( .A(n5375), .Y(n5376) );
  AND2X1 U4875 ( .A(n7779), .B(n719), .Y(n734) );
  INVX1 U4876 ( .A(n734), .Y(n5377) );
  INVX1 U4877 ( .A(n5380), .Y(n5378) );
  INVX1 U4878 ( .A(n5378), .Y(n5379) );
  AND2X1 U4879 ( .A(n7782), .B(n719), .Y(n733) );
  INVX1 U4880 ( .A(n733), .Y(n5380) );
  INVX1 U4881 ( .A(n5383), .Y(n5381) );
  INVX1 U4882 ( .A(n5381), .Y(n5382) );
  AND2X1 U4883 ( .A(n7785), .B(n719), .Y(n732) );
  INVX1 U4884 ( .A(n732), .Y(n5383) );
  INVX1 U4885 ( .A(n5386), .Y(n5384) );
  INVX1 U4886 ( .A(n5384), .Y(n5385) );
  AND2X1 U4887 ( .A(n7788), .B(n719), .Y(n731) );
  INVX1 U4888 ( .A(n731), .Y(n5386) );
  INVX1 U4889 ( .A(n5389), .Y(n5387) );
  INVX1 U4890 ( .A(n5387), .Y(n5388) );
  AND2X1 U4891 ( .A(n7791), .B(n719), .Y(n730) );
  INVX1 U4892 ( .A(n730), .Y(n5389) );
  INVX1 U4893 ( .A(n5392), .Y(n5390) );
  INVX1 U4894 ( .A(n5390), .Y(n5391) );
  AND2X1 U4895 ( .A(n7794), .B(n719), .Y(n729) );
  INVX1 U4896 ( .A(n729), .Y(n5392) );
  INVX1 U4897 ( .A(n5395), .Y(n5393) );
  INVX1 U4898 ( .A(n5393), .Y(n5394) );
  AND2X1 U4899 ( .A(n7797), .B(n719), .Y(n728) );
  INVX1 U4900 ( .A(n728), .Y(n5395) );
  INVX1 U4901 ( .A(n5398), .Y(n5396) );
  INVX1 U4902 ( .A(n5396), .Y(n5397) );
  AND2X1 U4903 ( .A(n7800), .B(n719), .Y(n727) );
  INVX1 U4904 ( .A(n727), .Y(n5398) );
  INVX1 U4905 ( .A(n5401), .Y(n5399) );
  INVX1 U4906 ( .A(n5399), .Y(n5400) );
  AND2X1 U4907 ( .A(n7803), .B(n719), .Y(n726) );
  INVX1 U4908 ( .A(n726), .Y(n5401) );
  INVX1 U4909 ( .A(n5404), .Y(n5402) );
  INVX1 U4910 ( .A(n5402), .Y(n5403) );
  AND2X1 U4911 ( .A(n7806), .B(n719), .Y(n725) );
  INVX1 U4912 ( .A(n725), .Y(n5404) );
  INVX1 U4913 ( .A(n5407), .Y(n5405) );
  INVX1 U4914 ( .A(n5405), .Y(n5406) );
  AND2X1 U4915 ( .A(n7809), .B(n719), .Y(n724) );
  INVX1 U4916 ( .A(n724), .Y(n5407) );
  INVX1 U4917 ( .A(n5410), .Y(n5408) );
  INVX1 U4918 ( .A(n5408), .Y(n5409) );
  AND2X1 U4919 ( .A(n7812), .B(n719), .Y(n723) );
  INVX1 U4920 ( .A(n723), .Y(n5410) );
  INVX1 U4921 ( .A(n5413), .Y(n5411) );
  INVX1 U4922 ( .A(n5411), .Y(n5412) );
  AND2X1 U4923 ( .A(n7815), .B(n719), .Y(n722) );
  INVX1 U4924 ( .A(n722), .Y(n5413) );
  INVX1 U4925 ( .A(n5416), .Y(n5414) );
  INVX1 U4926 ( .A(n5414), .Y(n5415) );
  AND2X1 U4927 ( .A(n7818), .B(n719), .Y(n721) );
  INVX1 U4928 ( .A(n721), .Y(n5416) );
  INVX1 U4929 ( .A(n5419), .Y(n5417) );
  INVX1 U4930 ( .A(n5417), .Y(n5418) );
  AND2X1 U4931 ( .A(n7821), .B(n719), .Y(n720) );
  INVX1 U4932 ( .A(n720), .Y(n5419) );
  INVX1 U4933 ( .A(n5422), .Y(n5420) );
  INVX1 U4934 ( .A(n5420), .Y(n5421) );
  AND2X1 U4935 ( .A(n9354), .B(n10515), .Y(n718) );
  INVX1 U4936 ( .A(n718), .Y(n5422) );
  INVX1 U4937 ( .A(n5425), .Y(n5423) );
  INVX1 U4938 ( .A(n5423), .Y(n5424) );
  AND2X1 U4939 ( .A(n9357), .B(n10515), .Y(n717) );
  INVX1 U4940 ( .A(n717), .Y(n5425) );
  INVX1 U4941 ( .A(n5428), .Y(n5426) );
  INVX1 U4942 ( .A(n5426), .Y(n5427) );
  AND2X1 U4943 ( .A(n9360), .B(n10515), .Y(n716) );
  INVX1 U4944 ( .A(n716), .Y(n5428) );
  INVX1 U4945 ( .A(n5431), .Y(n5429) );
  INVX1 U4946 ( .A(n5429), .Y(n5430) );
  AND2X1 U4947 ( .A(n9363), .B(n10515), .Y(n715) );
  INVX1 U4948 ( .A(n715), .Y(n5431) );
  INVX1 U4949 ( .A(n5434), .Y(n5432) );
  INVX1 U4950 ( .A(n5432), .Y(n5433) );
  AND2X1 U4951 ( .A(n9366), .B(n10515), .Y(n714) );
  INVX1 U4952 ( .A(n714), .Y(n5434) );
  INVX1 U4953 ( .A(n5437), .Y(n5435) );
  INVX1 U4954 ( .A(n5435), .Y(n5436) );
  AND2X1 U4955 ( .A(n9369), .B(n10515), .Y(n713) );
  INVX1 U4956 ( .A(n713), .Y(n5437) );
  INVX1 U4957 ( .A(n5440), .Y(n5438) );
  INVX1 U4958 ( .A(n5438), .Y(n5439) );
  AND2X1 U4959 ( .A(n9372), .B(n10515), .Y(n712) );
  INVX1 U4960 ( .A(n712), .Y(n5440) );
  INVX1 U4961 ( .A(n5443), .Y(n5441) );
  INVX1 U4962 ( .A(n5441), .Y(n5442) );
  AND2X1 U4963 ( .A(n9375), .B(n10515), .Y(n711) );
  INVX1 U4964 ( .A(n711), .Y(n5443) );
  INVX1 U4965 ( .A(n5446), .Y(n5444) );
  INVX1 U4966 ( .A(n5444), .Y(n5445) );
  AND2X1 U4967 ( .A(n9378), .B(n10515), .Y(n710) );
  INVX1 U4968 ( .A(n710), .Y(n5446) );
  INVX1 U4969 ( .A(n5449), .Y(n5447) );
  INVX1 U4970 ( .A(n5447), .Y(n5448) );
  AND2X1 U4971 ( .A(n9381), .B(n10515), .Y(n709) );
  INVX1 U4972 ( .A(n709), .Y(n5449) );
  INVX1 U4973 ( .A(n5452), .Y(n5450) );
  INVX1 U4974 ( .A(n5450), .Y(n5451) );
  AND2X1 U4975 ( .A(n9384), .B(n10515), .Y(n708) );
  INVX1 U4976 ( .A(n708), .Y(n5452) );
  INVX1 U4977 ( .A(n5455), .Y(n5453) );
  INVX1 U4978 ( .A(n5453), .Y(n5454) );
  AND2X1 U4979 ( .A(n9387), .B(n10515), .Y(n707) );
  INVX1 U4980 ( .A(n707), .Y(n5455) );
  INVX1 U4981 ( .A(n5458), .Y(n5456) );
  INVX1 U4982 ( .A(n5456), .Y(n5457) );
  AND2X1 U4983 ( .A(n9390), .B(n10515), .Y(n706) );
  INVX1 U4984 ( .A(n706), .Y(n5458) );
  INVX1 U4985 ( .A(n5461), .Y(n5459) );
  INVX1 U4986 ( .A(n5459), .Y(n5460) );
  AND2X1 U4987 ( .A(n9393), .B(n10515), .Y(n705) );
  INVX1 U4988 ( .A(n705), .Y(n5461) );
  INVX1 U4989 ( .A(n5464), .Y(n5462) );
  INVX1 U4990 ( .A(n5462), .Y(n5463) );
  AND2X1 U4991 ( .A(n9396), .B(n10515), .Y(n704) );
  INVX1 U4992 ( .A(n704), .Y(n5464) );
  INVX1 U4993 ( .A(n5467), .Y(n5465) );
  INVX1 U4994 ( .A(n5465), .Y(n5466) );
  AND2X1 U4995 ( .A(n9399), .B(n10515), .Y(n703) );
  INVX1 U4996 ( .A(n703), .Y(n5467) );
  INVX1 U4997 ( .A(n5470), .Y(n5468) );
  INVX1 U4998 ( .A(n5468), .Y(n5469) );
  AND2X1 U4999 ( .A(n9402), .B(n10515), .Y(n702) );
  INVX1 U5000 ( .A(n702), .Y(n5470) );
  INVX1 U5001 ( .A(n5473), .Y(n5471) );
  INVX1 U5002 ( .A(n5471), .Y(n5472) );
  AND2X1 U5003 ( .A(n9405), .B(n10515), .Y(n701) );
  INVX1 U5004 ( .A(n701), .Y(n5473) );
  INVX1 U5005 ( .A(n5476), .Y(n5474) );
  INVX1 U5006 ( .A(n5474), .Y(n5475) );
  AND2X1 U5007 ( .A(n9408), .B(n10515), .Y(n700) );
  INVX1 U5008 ( .A(n700), .Y(n5476) );
  INVX1 U5009 ( .A(n5479), .Y(n5477) );
  INVX1 U5010 ( .A(n5477), .Y(n5478) );
  AND2X1 U5011 ( .A(n9411), .B(n10515), .Y(n699) );
  INVX1 U5012 ( .A(n699), .Y(n5479) );
  INVX1 U5013 ( .A(n5482), .Y(n5480) );
  INVX1 U5014 ( .A(n5480), .Y(n5481) );
  AND2X1 U5015 ( .A(n9414), .B(n10515), .Y(n698) );
  INVX1 U5016 ( .A(n698), .Y(n5482) );
  INVX1 U5017 ( .A(n5485), .Y(n5483) );
  INVX1 U5018 ( .A(n5483), .Y(n5484) );
  AND2X1 U5019 ( .A(n9417), .B(n10515), .Y(n697) );
  INVX1 U5020 ( .A(n697), .Y(n5485) );
  INVX1 U5021 ( .A(n5488), .Y(n5486) );
  INVX1 U5022 ( .A(n5486), .Y(n5487) );
  AND2X1 U5023 ( .A(n9420), .B(n10515), .Y(n696) );
  INVX1 U5024 ( .A(n696), .Y(n5488) );
  INVX1 U5025 ( .A(n5491), .Y(n5489) );
  INVX1 U5026 ( .A(n5489), .Y(n5490) );
  AND2X1 U5027 ( .A(n9423), .B(n10515), .Y(n695) );
  INVX1 U5028 ( .A(n695), .Y(n5491) );
  INVX1 U5029 ( .A(n5494), .Y(n5492) );
  INVX1 U5030 ( .A(n5492), .Y(n5493) );
  AND2X1 U5031 ( .A(n9426), .B(n10515), .Y(n694) );
  INVX1 U5032 ( .A(n694), .Y(n5494) );
  INVX1 U5033 ( .A(n5497), .Y(n5495) );
  INVX1 U5034 ( .A(n5495), .Y(n5496) );
  AND2X1 U5035 ( .A(n9429), .B(n10515), .Y(n693) );
  INVX1 U5036 ( .A(n693), .Y(n5497) );
  INVX1 U5037 ( .A(n5500), .Y(n5498) );
  INVX1 U5038 ( .A(n5498), .Y(n5499) );
  AND2X1 U5039 ( .A(n9432), .B(n10515), .Y(n692) );
  INVX1 U5040 ( .A(n692), .Y(n5500) );
  INVX1 U5041 ( .A(n5503), .Y(n5501) );
  INVX1 U5042 ( .A(n5501), .Y(n5502) );
  AND2X1 U5043 ( .A(n9435), .B(n10515), .Y(n691) );
  INVX1 U5044 ( .A(n691), .Y(n5503) );
  INVX1 U5045 ( .A(n5506), .Y(n5504) );
  INVX1 U5046 ( .A(n5504), .Y(n5505) );
  AND2X1 U5047 ( .A(n9438), .B(n10515), .Y(n690) );
  INVX1 U5048 ( .A(n690), .Y(n5506) );
  INVX1 U5049 ( .A(n5509), .Y(n5507) );
  INVX1 U5050 ( .A(n5507), .Y(n5508) );
  AND2X1 U5051 ( .A(n9441), .B(n10515), .Y(n689) );
  INVX1 U5052 ( .A(n689), .Y(n5509) );
  INVX1 U5053 ( .A(n5512), .Y(n5510) );
  INVX1 U5054 ( .A(n5510), .Y(n5511) );
  AND2X1 U5055 ( .A(n9444), .B(n10515), .Y(n688) );
  INVX1 U5056 ( .A(n688), .Y(n5512) );
  INVX1 U5057 ( .A(n5515), .Y(n5513) );
  INVX1 U5058 ( .A(n5513), .Y(n5514) );
  AND2X1 U5059 ( .A(n9447), .B(n10515), .Y(n687) );
  INVX1 U5060 ( .A(n687), .Y(n5515) );
  INVX1 U5061 ( .A(n5518), .Y(n5516) );
  INVX1 U5062 ( .A(n5516), .Y(n5517) );
  AND2X1 U5063 ( .A(n9450), .B(n10515), .Y(n686) );
  INVX1 U5064 ( .A(n686), .Y(n5518) );
  INVX1 U5065 ( .A(n5521), .Y(n5519) );
  INVX1 U5066 ( .A(n5519), .Y(n5520) );
  AND2X1 U5067 ( .A(n9453), .B(n10515), .Y(n685) );
  INVX1 U5068 ( .A(n685), .Y(n5521) );
  INVX1 U5069 ( .A(n5524), .Y(n5522) );
  INVX1 U5070 ( .A(n5522), .Y(n5523) );
  AND2X1 U5071 ( .A(n7824), .B(n649), .Y(n683) );
  INVX1 U5072 ( .A(n683), .Y(n5524) );
  INVX1 U5073 ( .A(n5527), .Y(n5525) );
  INVX1 U5074 ( .A(n5525), .Y(n5526) );
  AND2X1 U5075 ( .A(n7827), .B(n649), .Y(n682) );
  INVX1 U5076 ( .A(n682), .Y(n5527) );
  INVX1 U5077 ( .A(n5530), .Y(n5528) );
  INVX1 U5078 ( .A(n5528), .Y(n5529) );
  AND2X1 U5079 ( .A(n7830), .B(n649), .Y(n681) );
  INVX1 U5080 ( .A(n681), .Y(n5530) );
  INVX1 U5081 ( .A(n5533), .Y(n5531) );
  INVX1 U5082 ( .A(n5531), .Y(n5532) );
  AND2X1 U5083 ( .A(n7833), .B(n649), .Y(n680) );
  INVX1 U5084 ( .A(n680), .Y(n5533) );
  INVX1 U5085 ( .A(n5536), .Y(n5534) );
  INVX1 U5086 ( .A(n5534), .Y(n5535) );
  AND2X1 U5087 ( .A(n7836), .B(n649), .Y(n679) );
  INVX1 U5088 ( .A(n679), .Y(n5536) );
  INVX1 U5089 ( .A(n5539), .Y(n5537) );
  INVX1 U5090 ( .A(n5537), .Y(n5538) );
  AND2X1 U5091 ( .A(n7839), .B(n649), .Y(n678) );
  INVX1 U5092 ( .A(n678), .Y(n5539) );
  INVX1 U5093 ( .A(n5542), .Y(n5540) );
  INVX1 U5094 ( .A(n5540), .Y(n5541) );
  AND2X1 U5095 ( .A(n7842), .B(n649), .Y(n677) );
  INVX1 U5096 ( .A(n677), .Y(n5542) );
  INVX1 U5097 ( .A(n5545), .Y(n5543) );
  INVX1 U5098 ( .A(n5543), .Y(n5544) );
  AND2X1 U5099 ( .A(n7845), .B(n649), .Y(n676) );
  INVX1 U5100 ( .A(n676), .Y(n5545) );
  INVX1 U5101 ( .A(n5548), .Y(n5546) );
  INVX1 U5102 ( .A(n5546), .Y(n5547) );
  AND2X1 U5103 ( .A(n7848), .B(n649), .Y(n675) );
  INVX1 U5104 ( .A(n675), .Y(n5548) );
  INVX1 U5105 ( .A(n5551), .Y(n5549) );
  INVX1 U5106 ( .A(n5549), .Y(n5550) );
  AND2X1 U5107 ( .A(n7851), .B(n649), .Y(n674) );
  INVX1 U5108 ( .A(n674), .Y(n5551) );
  INVX1 U5109 ( .A(n5554), .Y(n5552) );
  INVX1 U5110 ( .A(n5552), .Y(n5553) );
  AND2X1 U5111 ( .A(n7854), .B(n649), .Y(n673) );
  INVX1 U5112 ( .A(n673), .Y(n5554) );
  INVX1 U5113 ( .A(n5557), .Y(n5555) );
  INVX1 U5114 ( .A(n5555), .Y(n5556) );
  AND2X1 U5115 ( .A(n7857), .B(n649), .Y(n672) );
  INVX1 U5116 ( .A(n672), .Y(n5557) );
  INVX1 U5117 ( .A(n5560), .Y(n5558) );
  INVX1 U5118 ( .A(n5558), .Y(n5559) );
  AND2X1 U5119 ( .A(n7860), .B(n649), .Y(n671) );
  INVX1 U5120 ( .A(n671), .Y(n5560) );
  INVX1 U5121 ( .A(n5563), .Y(n5561) );
  INVX1 U5122 ( .A(n5561), .Y(n5562) );
  AND2X1 U5123 ( .A(n7863), .B(n649), .Y(n670) );
  INVX1 U5124 ( .A(n670), .Y(n5563) );
  INVX1 U5125 ( .A(n5566), .Y(n5564) );
  INVX1 U5126 ( .A(n5564), .Y(n5565) );
  AND2X1 U5127 ( .A(n7866), .B(n649), .Y(n669) );
  INVX1 U5128 ( .A(n669), .Y(n5566) );
  INVX1 U5129 ( .A(n5569), .Y(n5567) );
  INVX1 U5130 ( .A(n5567), .Y(n5568) );
  AND2X1 U5131 ( .A(n7869), .B(n649), .Y(n668) );
  INVX1 U5132 ( .A(n668), .Y(n5569) );
  INVX1 U5133 ( .A(n5572), .Y(n5570) );
  INVX1 U5134 ( .A(n5570), .Y(n5571) );
  AND2X1 U5135 ( .A(n7872), .B(n649), .Y(n667) );
  INVX1 U5136 ( .A(n667), .Y(n5572) );
  INVX1 U5137 ( .A(n5575), .Y(n5573) );
  INVX1 U5138 ( .A(n5573), .Y(n5574) );
  AND2X1 U5139 ( .A(n7875), .B(n649), .Y(n666) );
  INVX1 U5140 ( .A(n666), .Y(n5575) );
  INVX1 U5141 ( .A(n5578), .Y(n5576) );
  INVX1 U5142 ( .A(n5576), .Y(n5577) );
  AND2X1 U5143 ( .A(n7878), .B(n649), .Y(n665) );
  INVX1 U5144 ( .A(n665), .Y(n5578) );
  INVX1 U5145 ( .A(n5581), .Y(n5579) );
  INVX1 U5146 ( .A(n5579), .Y(n5580) );
  AND2X1 U5147 ( .A(n7881), .B(n649), .Y(n664) );
  INVX1 U5148 ( .A(n664), .Y(n5581) );
  INVX1 U5149 ( .A(n5584), .Y(n5582) );
  INVX1 U5150 ( .A(n5582), .Y(n5583) );
  AND2X1 U5151 ( .A(n7884), .B(n649), .Y(n663) );
  INVX1 U5152 ( .A(n663), .Y(n5584) );
  INVX1 U5153 ( .A(n5587), .Y(n5585) );
  INVX1 U5154 ( .A(n5585), .Y(n5586) );
  AND2X1 U5155 ( .A(n7887), .B(n649), .Y(n662) );
  INVX1 U5156 ( .A(n662), .Y(n5587) );
  INVX1 U5157 ( .A(n5590), .Y(n5588) );
  INVX1 U5158 ( .A(n5588), .Y(n5589) );
  AND2X1 U5159 ( .A(n7890), .B(n649), .Y(n661) );
  INVX1 U5160 ( .A(n661), .Y(n5590) );
  INVX1 U5161 ( .A(n5593), .Y(n5591) );
  INVX1 U5162 ( .A(n5591), .Y(n5592) );
  AND2X1 U5163 ( .A(n7893), .B(n649), .Y(n660) );
  INVX1 U5164 ( .A(n660), .Y(n5593) );
  INVX1 U5165 ( .A(n5596), .Y(n5594) );
  INVX1 U5166 ( .A(n5594), .Y(n5595) );
  AND2X1 U5167 ( .A(n7896), .B(n649), .Y(n659) );
  INVX1 U5168 ( .A(n659), .Y(n5596) );
  INVX1 U5169 ( .A(n5599), .Y(n5597) );
  INVX1 U5170 ( .A(n5597), .Y(n5598) );
  AND2X1 U5171 ( .A(n7899), .B(n649), .Y(n658) );
  INVX1 U5172 ( .A(n658), .Y(n5599) );
  INVX1 U5173 ( .A(n5602), .Y(n5600) );
  INVX1 U5174 ( .A(n5600), .Y(n5601) );
  AND2X1 U5175 ( .A(n7902), .B(n649), .Y(n657) );
  INVX1 U5176 ( .A(n657), .Y(n5602) );
  INVX1 U5177 ( .A(n5605), .Y(n5603) );
  INVX1 U5178 ( .A(n5603), .Y(n5604) );
  AND2X1 U5179 ( .A(n7905), .B(n649), .Y(n656) );
  INVX1 U5180 ( .A(n656), .Y(n5605) );
  INVX1 U5181 ( .A(n5608), .Y(n5606) );
  INVX1 U5182 ( .A(n5606), .Y(n5607) );
  AND2X1 U5183 ( .A(n7908), .B(n649), .Y(n655) );
  INVX1 U5184 ( .A(n655), .Y(n5608) );
  INVX1 U5185 ( .A(n5611), .Y(n5609) );
  INVX1 U5186 ( .A(n5609), .Y(n5610) );
  AND2X1 U5187 ( .A(n7911), .B(n649), .Y(n654) );
  INVX1 U5188 ( .A(n654), .Y(n5611) );
  INVX1 U5189 ( .A(n5614), .Y(n5612) );
  INVX1 U5190 ( .A(n5612), .Y(n5613) );
  AND2X1 U5191 ( .A(n7914), .B(n649), .Y(n653) );
  INVX1 U5192 ( .A(n653), .Y(n5614) );
  INVX1 U5193 ( .A(n5617), .Y(n5615) );
  INVX1 U5194 ( .A(n5615), .Y(n5616) );
  AND2X1 U5195 ( .A(n7917), .B(n649), .Y(n652) );
  INVX1 U5196 ( .A(n652), .Y(n5617) );
  INVX1 U5197 ( .A(n5620), .Y(n5618) );
  INVX1 U5198 ( .A(n5618), .Y(n5619) );
  AND2X1 U5199 ( .A(n7920), .B(n649), .Y(n651) );
  INVX1 U5200 ( .A(n651), .Y(n5620) );
  INVX1 U5201 ( .A(n5623), .Y(n5621) );
  INVX1 U5202 ( .A(n5621), .Y(n5622) );
  AND2X1 U5203 ( .A(n7923), .B(n649), .Y(n650) );
  INVX1 U5204 ( .A(n650), .Y(n5623) );
  INVX1 U5205 ( .A(n5626), .Y(n5624) );
  INVX1 U5206 ( .A(n5624), .Y(n5625) );
  AND2X1 U5207 ( .A(n9456), .B(n10508), .Y(n648) );
  INVX1 U5208 ( .A(n648), .Y(n5626) );
  INVX1 U5209 ( .A(n5629), .Y(n5627) );
  INVX1 U5210 ( .A(n5627), .Y(n5628) );
  AND2X1 U5211 ( .A(n9459), .B(n10508), .Y(n647) );
  INVX1 U5212 ( .A(n647), .Y(n5629) );
  INVX1 U5213 ( .A(n5632), .Y(n5630) );
  INVX1 U5214 ( .A(n5630), .Y(n5631) );
  AND2X1 U5215 ( .A(n9462), .B(n10508), .Y(n646) );
  INVX1 U5216 ( .A(n646), .Y(n5632) );
  INVX1 U5217 ( .A(n5635), .Y(n5633) );
  INVX1 U5218 ( .A(n5633), .Y(n5634) );
  AND2X1 U5219 ( .A(n9465), .B(n10508), .Y(n645) );
  INVX1 U5220 ( .A(n645), .Y(n5635) );
  INVX1 U5221 ( .A(n5638), .Y(n5636) );
  INVX1 U5222 ( .A(n5636), .Y(n5637) );
  AND2X1 U5223 ( .A(n9468), .B(n10508), .Y(n644) );
  INVX1 U5224 ( .A(n644), .Y(n5638) );
  INVX1 U5225 ( .A(n5641), .Y(n5639) );
  INVX1 U5226 ( .A(n5639), .Y(n5640) );
  AND2X1 U5227 ( .A(n9471), .B(n10508), .Y(n643) );
  INVX1 U5228 ( .A(n643), .Y(n5641) );
  INVX1 U5229 ( .A(n5644), .Y(n5642) );
  INVX1 U5230 ( .A(n5642), .Y(n5643) );
  AND2X1 U5231 ( .A(n9474), .B(n10508), .Y(n642) );
  INVX1 U5232 ( .A(n642), .Y(n5644) );
  INVX1 U5233 ( .A(n5647), .Y(n5645) );
  INVX1 U5234 ( .A(n5645), .Y(n5646) );
  AND2X1 U5235 ( .A(n9477), .B(n10508), .Y(n641) );
  INVX1 U5236 ( .A(n641), .Y(n5647) );
  INVX1 U5237 ( .A(n5650), .Y(n5648) );
  INVX1 U5238 ( .A(n5648), .Y(n5649) );
  AND2X1 U5239 ( .A(n9480), .B(n10508), .Y(n640) );
  INVX1 U5240 ( .A(n640), .Y(n5650) );
  INVX1 U5241 ( .A(n5653), .Y(n5651) );
  INVX1 U5242 ( .A(n5651), .Y(n5652) );
  AND2X1 U5243 ( .A(n9483), .B(n10508), .Y(n639) );
  INVX1 U5244 ( .A(n639), .Y(n5653) );
  INVX1 U5245 ( .A(n5656), .Y(n5654) );
  INVX1 U5246 ( .A(n5654), .Y(n5655) );
  AND2X1 U5247 ( .A(n9486), .B(n10508), .Y(n638) );
  INVX1 U5248 ( .A(n638), .Y(n5656) );
  INVX1 U5249 ( .A(n5659), .Y(n5657) );
  INVX1 U5250 ( .A(n5657), .Y(n5658) );
  AND2X1 U5251 ( .A(n9489), .B(n10508), .Y(n637) );
  INVX1 U5252 ( .A(n637), .Y(n5659) );
  INVX1 U5253 ( .A(n5662), .Y(n5660) );
  INVX1 U5254 ( .A(n5660), .Y(n5661) );
  AND2X1 U5255 ( .A(n9492), .B(n10508), .Y(n636) );
  INVX1 U5256 ( .A(n636), .Y(n5662) );
  INVX1 U5257 ( .A(n5665), .Y(n5663) );
  INVX1 U5258 ( .A(n5663), .Y(n5664) );
  AND2X1 U5259 ( .A(n9495), .B(n10508), .Y(n635) );
  INVX1 U5260 ( .A(n635), .Y(n5665) );
  INVX1 U5261 ( .A(n5668), .Y(n5666) );
  INVX1 U5262 ( .A(n5666), .Y(n5667) );
  AND2X1 U5263 ( .A(n9498), .B(n10508), .Y(n634) );
  INVX1 U5264 ( .A(n634), .Y(n5668) );
  INVX1 U5265 ( .A(n5671), .Y(n5669) );
  INVX1 U5266 ( .A(n5669), .Y(n5670) );
  AND2X1 U5267 ( .A(n9501), .B(n10508), .Y(n633) );
  INVX1 U5268 ( .A(n633), .Y(n5671) );
  INVX1 U5269 ( .A(n5674), .Y(n5672) );
  INVX1 U5270 ( .A(n5672), .Y(n5673) );
  AND2X1 U5271 ( .A(n9504), .B(n10508), .Y(n632) );
  INVX1 U5272 ( .A(n632), .Y(n5674) );
  INVX1 U5273 ( .A(n5677), .Y(n5675) );
  INVX1 U5274 ( .A(n5675), .Y(n5676) );
  AND2X1 U5275 ( .A(n9507), .B(n10508), .Y(n631) );
  INVX1 U5276 ( .A(n631), .Y(n5677) );
  INVX1 U5277 ( .A(n5680), .Y(n5678) );
  INVX1 U5278 ( .A(n5678), .Y(n5679) );
  AND2X1 U5279 ( .A(n9510), .B(n10508), .Y(n630) );
  INVX1 U5280 ( .A(n630), .Y(n5680) );
  INVX1 U5281 ( .A(n5683), .Y(n5681) );
  INVX1 U5282 ( .A(n5681), .Y(n5682) );
  AND2X1 U5283 ( .A(n9513), .B(n10508), .Y(n629) );
  INVX1 U5284 ( .A(n629), .Y(n5683) );
  INVX1 U5285 ( .A(n5686), .Y(n5684) );
  INVX1 U5286 ( .A(n5684), .Y(n5685) );
  AND2X1 U5287 ( .A(n9516), .B(n10508), .Y(n628) );
  INVX1 U5288 ( .A(n628), .Y(n5686) );
  INVX1 U5289 ( .A(n5689), .Y(n5687) );
  INVX1 U5290 ( .A(n5687), .Y(n5688) );
  AND2X1 U5291 ( .A(n9519), .B(n10508), .Y(n627) );
  INVX1 U5292 ( .A(n627), .Y(n5689) );
  INVX1 U5293 ( .A(n5692), .Y(n5690) );
  INVX1 U5294 ( .A(n5690), .Y(n5691) );
  AND2X1 U5295 ( .A(n9522), .B(n10508), .Y(n626) );
  INVX1 U5296 ( .A(n626), .Y(n5692) );
  INVX1 U5297 ( .A(n5695), .Y(n5693) );
  INVX1 U5298 ( .A(n5693), .Y(n5694) );
  AND2X1 U5299 ( .A(n9525), .B(n10508), .Y(n625) );
  INVX1 U5300 ( .A(n625), .Y(n5695) );
  INVX1 U5301 ( .A(n5698), .Y(n5696) );
  INVX1 U5302 ( .A(n5696), .Y(n5697) );
  AND2X1 U5303 ( .A(n9528), .B(n10508), .Y(n624) );
  INVX1 U5304 ( .A(n624), .Y(n5698) );
  INVX1 U5305 ( .A(n5701), .Y(n5699) );
  INVX1 U5306 ( .A(n5699), .Y(n5700) );
  AND2X1 U5307 ( .A(n9531), .B(n10508), .Y(n623) );
  INVX1 U5308 ( .A(n623), .Y(n5701) );
  INVX1 U5309 ( .A(n5704), .Y(n5702) );
  INVX1 U5310 ( .A(n5702), .Y(n5703) );
  AND2X1 U5311 ( .A(n9534), .B(n10508), .Y(n622) );
  INVX1 U5312 ( .A(n622), .Y(n5704) );
  INVX1 U5313 ( .A(n5707), .Y(n5705) );
  INVX1 U5314 ( .A(n5705), .Y(n5706) );
  AND2X1 U5315 ( .A(n9537), .B(n10508), .Y(n621) );
  INVX1 U5316 ( .A(n621), .Y(n5707) );
  INVX1 U5317 ( .A(n5710), .Y(n5708) );
  INVX1 U5318 ( .A(n5708), .Y(n5709) );
  AND2X1 U5319 ( .A(n9540), .B(n10508), .Y(n620) );
  INVX1 U5320 ( .A(n620), .Y(n5710) );
  INVX1 U5321 ( .A(n5713), .Y(n5711) );
  INVX1 U5322 ( .A(n5711), .Y(n5712) );
  AND2X1 U5323 ( .A(n9543), .B(n10508), .Y(n619) );
  INVX1 U5324 ( .A(n619), .Y(n5713) );
  INVX1 U5325 ( .A(n5716), .Y(n5714) );
  INVX1 U5326 ( .A(n5714), .Y(n5715) );
  AND2X1 U5327 ( .A(n9546), .B(n10508), .Y(n618) );
  INVX1 U5328 ( .A(n618), .Y(n5716) );
  INVX1 U5329 ( .A(n5719), .Y(n5717) );
  INVX1 U5330 ( .A(n5717), .Y(n5718) );
  AND2X1 U5331 ( .A(n9549), .B(n10508), .Y(n617) );
  INVX1 U5332 ( .A(n617), .Y(n5719) );
  INVX1 U5333 ( .A(n5722), .Y(n5720) );
  INVX1 U5334 ( .A(n5720), .Y(n5721) );
  AND2X1 U5335 ( .A(n9552), .B(n10508), .Y(n616) );
  INVX1 U5336 ( .A(n616), .Y(n5722) );
  INVX1 U5337 ( .A(n5725), .Y(n5723) );
  INVX1 U5338 ( .A(n5723), .Y(n5724) );
  AND2X1 U5339 ( .A(n9555), .B(n10508), .Y(n615) );
  INVX1 U5340 ( .A(n615), .Y(n5725) );
  INVX1 U5341 ( .A(n5728), .Y(n5726) );
  INVX1 U5342 ( .A(n5726), .Y(n5727) );
  AND2X1 U5343 ( .A(n7926), .B(n10506), .Y(n612) );
  INVX1 U5344 ( .A(n612), .Y(n5728) );
  INVX1 U5345 ( .A(n5731), .Y(n5729) );
  INVX1 U5346 ( .A(n5729), .Y(n5730) );
  AND2X1 U5347 ( .A(n7929), .B(n10506), .Y(n611) );
  INVX1 U5348 ( .A(n611), .Y(n5731) );
  INVX1 U5349 ( .A(n5734), .Y(n5732) );
  INVX1 U5350 ( .A(n5732), .Y(n5733) );
  AND2X1 U5351 ( .A(n7932), .B(n10506), .Y(n610) );
  INVX1 U5352 ( .A(n610), .Y(n5734) );
  INVX1 U5353 ( .A(n5737), .Y(n5735) );
  INVX1 U5354 ( .A(n5735), .Y(n5736) );
  AND2X1 U5355 ( .A(n7935), .B(n10506), .Y(n609) );
  INVX1 U5356 ( .A(n609), .Y(n5737) );
  INVX1 U5357 ( .A(n5740), .Y(n5738) );
  INVX1 U5358 ( .A(n5738), .Y(n5739) );
  AND2X1 U5359 ( .A(n7938), .B(n10506), .Y(n608) );
  INVX1 U5360 ( .A(n608), .Y(n5740) );
  INVX1 U5361 ( .A(n5743), .Y(n5741) );
  INVX1 U5362 ( .A(n5741), .Y(n5742) );
  AND2X1 U5363 ( .A(n7941), .B(n10506), .Y(n607) );
  INVX1 U5364 ( .A(n607), .Y(n5743) );
  INVX1 U5365 ( .A(n5746), .Y(n5744) );
  INVX1 U5366 ( .A(n5744), .Y(n5745) );
  AND2X1 U5367 ( .A(n7944), .B(n10506), .Y(n606) );
  INVX1 U5368 ( .A(n606), .Y(n5746) );
  INVX1 U5369 ( .A(n5749), .Y(n5747) );
  INVX1 U5370 ( .A(n5747), .Y(n5748) );
  AND2X1 U5371 ( .A(n7947), .B(n10506), .Y(n605) );
  INVX1 U5372 ( .A(n605), .Y(n5749) );
  INVX1 U5373 ( .A(n5752), .Y(n5750) );
  INVX1 U5374 ( .A(n5750), .Y(n5751) );
  AND2X1 U5375 ( .A(n7950), .B(n10506), .Y(n604) );
  INVX1 U5376 ( .A(n604), .Y(n5752) );
  INVX1 U5377 ( .A(n5755), .Y(n5753) );
  INVX1 U5378 ( .A(n5753), .Y(n5754) );
  AND2X1 U5379 ( .A(n7953), .B(n10506), .Y(n603) );
  INVX1 U5380 ( .A(n603), .Y(n5755) );
  INVX1 U5381 ( .A(n5758), .Y(n5756) );
  INVX1 U5382 ( .A(n5756), .Y(n5757) );
  AND2X1 U5383 ( .A(n7956), .B(n10506), .Y(n602) );
  INVX1 U5384 ( .A(n602), .Y(n5758) );
  INVX1 U5385 ( .A(n5761), .Y(n5759) );
  INVX1 U5386 ( .A(n5759), .Y(n5760) );
  AND2X1 U5387 ( .A(n7959), .B(n10506), .Y(n601) );
  INVX1 U5388 ( .A(n601), .Y(n5761) );
  INVX1 U5389 ( .A(n5764), .Y(n5762) );
  INVX1 U5390 ( .A(n5762), .Y(n5763) );
  AND2X1 U5391 ( .A(n7962), .B(n10506), .Y(n600) );
  INVX1 U5392 ( .A(n600), .Y(n5764) );
  INVX1 U5393 ( .A(n5767), .Y(n5765) );
  INVX1 U5394 ( .A(n5765), .Y(n5766) );
  AND2X1 U5395 ( .A(n7965), .B(n10506), .Y(n599) );
  INVX1 U5396 ( .A(n599), .Y(n5767) );
  INVX1 U5397 ( .A(n5770), .Y(n5768) );
  INVX1 U5398 ( .A(n5768), .Y(n5769) );
  AND2X1 U5399 ( .A(n7968), .B(n10506), .Y(n598) );
  INVX1 U5400 ( .A(n598), .Y(n5770) );
  INVX1 U5401 ( .A(n5773), .Y(n5771) );
  INVX1 U5402 ( .A(n5771), .Y(n5772) );
  AND2X1 U5403 ( .A(n7971), .B(n10506), .Y(n597) );
  INVX1 U5404 ( .A(n597), .Y(n5773) );
  INVX1 U5405 ( .A(n5776), .Y(n5774) );
  INVX1 U5406 ( .A(n5774), .Y(n5775) );
  AND2X1 U5407 ( .A(n7974), .B(n10506), .Y(n596) );
  INVX1 U5408 ( .A(n596), .Y(n5776) );
  INVX1 U5409 ( .A(n5779), .Y(n5777) );
  INVX1 U5410 ( .A(n5777), .Y(n5778) );
  AND2X1 U5411 ( .A(n7977), .B(n10506), .Y(n595) );
  INVX1 U5412 ( .A(n595), .Y(n5779) );
  INVX1 U5413 ( .A(n5782), .Y(n5780) );
  INVX1 U5414 ( .A(n5780), .Y(n5781) );
  AND2X1 U5415 ( .A(n7980), .B(n10506), .Y(n594) );
  INVX1 U5416 ( .A(n594), .Y(n5782) );
  INVX1 U5417 ( .A(n5785), .Y(n5783) );
  INVX1 U5418 ( .A(n5783), .Y(n5784) );
  AND2X1 U5419 ( .A(n7983), .B(n10506), .Y(n593) );
  INVX1 U5420 ( .A(n593), .Y(n5785) );
  INVX1 U5421 ( .A(n5788), .Y(n5786) );
  INVX1 U5422 ( .A(n5786), .Y(n5787) );
  AND2X1 U5423 ( .A(n7986), .B(n10506), .Y(n592) );
  INVX1 U5424 ( .A(n592), .Y(n5788) );
  INVX1 U5425 ( .A(n5791), .Y(n5789) );
  INVX1 U5426 ( .A(n5789), .Y(n5790) );
  AND2X1 U5427 ( .A(n7989), .B(n10506), .Y(n591) );
  INVX1 U5428 ( .A(n591), .Y(n5791) );
  INVX1 U5429 ( .A(n5794), .Y(n5792) );
  INVX1 U5430 ( .A(n5792), .Y(n5793) );
  AND2X1 U5431 ( .A(n7992), .B(n10506), .Y(n590) );
  INVX1 U5432 ( .A(n590), .Y(n5794) );
  INVX1 U5433 ( .A(n5797), .Y(n5795) );
  INVX1 U5434 ( .A(n5795), .Y(n5796) );
  AND2X1 U5435 ( .A(n7995), .B(n10506), .Y(n589) );
  INVX1 U5436 ( .A(n589), .Y(n5797) );
  INVX1 U5437 ( .A(n5800), .Y(n5798) );
  INVX1 U5438 ( .A(n5798), .Y(n5799) );
  AND2X1 U5439 ( .A(n7998), .B(n10506), .Y(n588) );
  INVX1 U5440 ( .A(n588), .Y(n5800) );
  INVX1 U5441 ( .A(n5803), .Y(n5801) );
  INVX1 U5442 ( .A(n5801), .Y(n5802) );
  AND2X1 U5443 ( .A(n8001), .B(n10506), .Y(n587) );
  INVX1 U5444 ( .A(n587), .Y(n5803) );
  INVX1 U5445 ( .A(n5806), .Y(n5804) );
  INVX1 U5446 ( .A(n5804), .Y(n5805) );
  AND2X1 U5447 ( .A(n8004), .B(n10506), .Y(n586) );
  INVX1 U5448 ( .A(n586), .Y(n5806) );
  INVX1 U5449 ( .A(n5809), .Y(n5807) );
  INVX1 U5450 ( .A(n5807), .Y(n5808) );
  AND2X1 U5451 ( .A(n8007), .B(n10506), .Y(n585) );
  INVX1 U5452 ( .A(n585), .Y(n5809) );
  INVX1 U5453 ( .A(n5812), .Y(n5810) );
  INVX1 U5454 ( .A(n5810), .Y(n5811) );
  AND2X1 U5455 ( .A(n8010), .B(n10506), .Y(n584) );
  INVX1 U5456 ( .A(n584), .Y(n5812) );
  INVX1 U5457 ( .A(n5815), .Y(n5813) );
  INVX1 U5458 ( .A(n5813), .Y(n5814) );
  AND2X1 U5459 ( .A(n8013), .B(n10506), .Y(n583) );
  INVX1 U5460 ( .A(n583), .Y(n5815) );
  INVX1 U5461 ( .A(n5818), .Y(n5816) );
  INVX1 U5462 ( .A(n5816), .Y(n5817) );
  AND2X1 U5463 ( .A(n8016), .B(n10506), .Y(n582) );
  INVX1 U5464 ( .A(n582), .Y(n5818) );
  INVX1 U5465 ( .A(n5821), .Y(n5819) );
  INVX1 U5466 ( .A(n5819), .Y(n5820) );
  AND2X1 U5467 ( .A(n8019), .B(n10506), .Y(n581) );
  INVX1 U5468 ( .A(n581), .Y(n5821) );
  INVX1 U5469 ( .A(n5824), .Y(n5822) );
  INVX1 U5470 ( .A(n5822), .Y(n5823) );
  AND2X1 U5471 ( .A(n8022), .B(n10506), .Y(n580) );
  INVX1 U5472 ( .A(n580), .Y(n5824) );
  INVX1 U5473 ( .A(n5827), .Y(n5825) );
  INVX1 U5474 ( .A(n5825), .Y(n5826) );
  AND2X1 U5475 ( .A(n8025), .B(n10506), .Y(n579) );
  INVX1 U5476 ( .A(n579), .Y(n5827) );
  INVX1 U5477 ( .A(n5830), .Y(n5828) );
  INVX1 U5478 ( .A(n5828), .Y(n5829) );
  AND2X1 U5479 ( .A(n9558), .B(n541), .Y(n575) );
  INVX1 U5480 ( .A(n575), .Y(n5830) );
  INVX1 U5481 ( .A(n5833), .Y(n5831) );
  INVX1 U5482 ( .A(n5831), .Y(n5832) );
  AND2X1 U5483 ( .A(n9561), .B(n541), .Y(n574) );
  INVX1 U5484 ( .A(n574), .Y(n5833) );
  INVX1 U5485 ( .A(n5836), .Y(n5834) );
  INVX1 U5486 ( .A(n5834), .Y(n5835) );
  AND2X1 U5487 ( .A(n9564), .B(n541), .Y(n573) );
  INVX1 U5488 ( .A(n573), .Y(n5836) );
  INVX1 U5489 ( .A(n5839), .Y(n5837) );
  INVX1 U5490 ( .A(n5837), .Y(n5838) );
  AND2X1 U5491 ( .A(n9567), .B(n541), .Y(n572) );
  INVX1 U5492 ( .A(n572), .Y(n5839) );
  INVX1 U5493 ( .A(n5842), .Y(n5840) );
  INVX1 U5494 ( .A(n5840), .Y(n5841) );
  AND2X1 U5495 ( .A(n9570), .B(n541), .Y(n571) );
  INVX1 U5496 ( .A(n571), .Y(n5842) );
  INVX1 U5497 ( .A(n5845), .Y(n5843) );
  INVX1 U5498 ( .A(n5843), .Y(n5844) );
  AND2X1 U5499 ( .A(n9573), .B(n541), .Y(n570) );
  INVX1 U5500 ( .A(n570), .Y(n5845) );
  INVX1 U5501 ( .A(n5848), .Y(n5846) );
  INVX1 U5502 ( .A(n5846), .Y(n5847) );
  AND2X1 U5503 ( .A(n9576), .B(n541), .Y(n569) );
  INVX1 U5504 ( .A(n569), .Y(n5848) );
  INVX1 U5505 ( .A(n5851), .Y(n5849) );
  INVX1 U5506 ( .A(n5849), .Y(n5850) );
  AND2X1 U5507 ( .A(n9579), .B(n541), .Y(n568) );
  INVX1 U5508 ( .A(n568), .Y(n5851) );
  INVX1 U5509 ( .A(n5854), .Y(n5852) );
  INVX1 U5510 ( .A(n5852), .Y(n5853) );
  AND2X1 U5511 ( .A(n9582), .B(n541), .Y(n567) );
  INVX1 U5512 ( .A(n567), .Y(n5854) );
  INVX1 U5513 ( .A(n5857), .Y(n5855) );
  INVX1 U5514 ( .A(n5855), .Y(n5856) );
  AND2X1 U5515 ( .A(n9585), .B(n541), .Y(n566) );
  INVX1 U5516 ( .A(n566), .Y(n5857) );
  INVX1 U5517 ( .A(n5860), .Y(n5858) );
  INVX1 U5518 ( .A(n5858), .Y(n5859) );
  AND2X1 U5519 ( .A(n9588), .B(n541), .Y(n565) );
  INVX1 U5520 ( .A(n565), .Y(n5860) );
  INVX1 U5521 ( .A(n5863), .Y(n5861) );
  INVX1 U5522 ( .A(n5861), .Y(n5862) );
  AND2X1 U5523 ( .A(n9591), .B(n541), .Y(n564) );
  INVX1 U5524 ( .A(n564), .Y(n5863) );
  INVX1 U5525 ( .A(n5866), .Y(n5864) );
  INVX1 U5526 ( .A(n5864), .Y(n5865) );
  AND2X1 U5527 ( .A(n9594), .B(n541), .Y(n563) );
  INVX1 U5528 ( .A(n563), .Y(n5866) );
  INVX1 U5529 ( .A(n5869), .Y(n5867) );
  INVX1 U5530 ( .A(n5867), .Y(n5868) );
  AND2X1 U5531 ( .A(n9597), .B(n541), .Y(n562) );
  INVX1 U5532 ( .A(n562), .Y(n5869) );
  INVX1 U5533 ( .A(n5872), .Y(n5870) );
  INVX1 U5534 ( .A(n5870), .Y(n5871) );
  AND2X1 U5535 ( .A(n9600), .B(n541), .Y(n561) );
  INVX1 U5536 ( .A(n561), .Y(n5872) );
  INVX1 U5537 ( .A(n5875), .Y(n5873) );
  INVX1 U5538 ( .A(n5873), .Y(n5874) );
  AND2X1 U5539 ( .A(n9603), .B(n541), .Y(n560) );
  INVX1 U5540 ( .A(n560), .Y(n5875) );
  INVX1 U5541 ( .A(n5878), .Y(n5876) );
  INVX1 U5542 ( .A(n5876), .Y(n5877) );
  AND2X1 U5543 ( .A(n9606), .B(n541), .Y(n559) );
  INVX1 U5544 ( .A(n559), .Y(n5878) );
  INVX1 U5545 ( .A(n5881), .Y(n5879) );
  INVX1 U5546 ( .A(n5879), .Y(n5880) );
  AND2X1 U5547 ( .A(n9609), .B(n541), .Y(n558) );
  INVX1 U5548 ( .A(n558), .Y(n5881) );
  INVX1 U5549 ( .A(n5884), .Y(n5882) );
  INVX1 U5550 ( .A(n5882), .Y(n5883) );
  AND2X1 U5551 ( .A(n9612), .B(n541), .Y(n557) );
  INVX1 U5552 ( .A(n557), .Y(n5884) );
  INVX1 U5553 ( .A(n5887), .Y(n5885) );
  INVX1 U5554 ( .A(n5885), .Y(n5886) );
  AND2X1 U5555 ( .A(n9615), .B(n541), .Y(n556) );
  INVX1 U5556 ( .A(n556), .Y(n5887) );
  INVX1 U5557 ( .A(n5890), .Y(n5888) );
  INVX1 U5558 ( .A(n5888), .Y(n5889) );
  AND2X1 U5559 ( .A(n9618), .B(n541), .Y(n555) );
  INVX1 U5560 ( .A(n555), .Y(n5890) );
  INVX1 U5561 ( .A(n5893), .Y(n5891) );
  INVX1 U5562 ( .A(n5891), .Y(n5892) );
  AND2X1 U5563 ( .A(n9621), .B(n541), .Y(n554) );
  INVX1 U5564 ( .A(n554), .Y(n5893) );
  INVX1 U5565 ( .A(n5896), .Y(n5894) );
  INVX1 U5566 ( .A(n5894), .Y(n5895) );
  AND2X1 U5567 ( .A(n9624), .B(n541), .Y(n553) );
  INVX1 U5568 ( .A(n553), .Y(n5896) );
  INVX1 U5569 ( .A(n5899), .Y(n5897) );
  INVX1 U5570 ( .A(n5897), .Y(n5898) );
  AND2X1 U5571 ( .A(n9627), .B(n541), .Y(n552) );
  INVX1 U5572 ( .A(n552), .Y(n5899) );
  INVX1 U5573 ( .A(n5902), .Y(n5900) );
  INVX1 U5574 ( .A(n5900), .Y(n5901) );
  AND2X1 U5575 ( .A(n9630), .B(n541), .Y(n551) );
  INVX1 U5576 ( .A(n551), .Y(n5902) );
  INVX1 U5577 ( .A(n5905), .Y(n5903) );
  INVX1 U5578 ( .A(n5903), .Y(n5904) );
  AND2X1 U5579 ( .A(n9633), .B(n541), .Y(n550) );
  INVX1 U5580 ( .A(n550), .Y(n5905) );
  INVX1 U5581 ( .A(n5908), .Y(n5906) );
  INVX1 U5582 ( .A(n5906), .Y(n5907) );
  AND2X1 U5583 ( .A(n9636), .B(n541), .Y(n549) );
  INVX1 U5584 ( .A(n549), .Y(n5908) );
  INVX1 U5585 ( .A(n5911), .Y(n5909) );
  INVX1 U5586 ( .A(n5909), .Y(n5910) );
  AND2X1 U5587 ( .A(n9639), .B(n541), .Y(n548) );
  INVX1 U5588 ( .A(n548), .Y(n5911) );
  INVX1 U5589 ( .A(n5914), .Y(n5912) );
  INVX1 U5590 ( .A(n5912), .Y(n5913) );
  AND2X1 U5591 ( .A(n9642), .B(n541), .Y(n547) );
  INVX1 U5592 ( .A(n547), .Y(n5914) );
  INVX1 U5593 ( .A(n5917), .Y(n5915) );
  INVX1 U5594 ( .A(n5915), .Y(n5916) );
  AND2X1 U5595 ( .A(n9645), .B(n541), .Y(n546) );
  INVX1 U5596 ( .A(n546), .Y(n5917) );
  INVX1 U5597 ( .A(n5920), .Y(n5918) );
  INVX1 U5598 ( .A(n5918), .Y(n5919) );
  AND2X1 U5599 ( .A(n9648), .B(n541), .Y(n545) );
  INVX1 U5600 ( .A(n545), .Y(n5920) );
  INVX1 U5601 ( .A(n5923), .Y(n5921) );
  INVX1 U5602 ( .A(n5921), .Y(n5922) );
  AND2X1 U5603 ( .A(n9651), .B(n541), .Y(n544) );
  INVX1 U5604 ( .A(n544), .Y(n5923) );
  INVX1 U5605 ( .A(n5926), .Y(n5924) );
  INVX1 U5606 ( .A(n5924), .Y(n5925) );
  AND2X1 U5607 ( .A(n9654), .B(n541), .Y(n543) );
  INVX1 U5608 ( .A(n543), .Y(n5926) );
  INVX1 U5609 ( .A(n5929), .Y(n5927) );
  INVX1 U5610 ( .A(n5927), .Y(n5928) );
  AND2X1 U5611 ( .A(n9657), .B(n541), .Y(n542) );
  INVX1 U5612 ( .A(n542), .Y(n5929) );
  INVX1 U5613 ( .A(n5932), .Y(n5930) );
  INVX1 U5614 ( .A(n5930), .Y(n5931) );
  AND2X1 U5615 ( .A(n8028), .B(n505), .Y(n539) );
  INVX1 U5616 ( .A(n539), .Y(n5932) );
  INVX1 U5617 ( .A(n5935), .Y(n5933) );
  INVX1 U5618 ( .A(n5933), .Y(n5934) );
  AND2X1 U5619 ( .A(n8031), .B(n505), .Y(n538) );
  INVX1 U5620 ( .A(n538), .Y(n5935) );
  INVX1 U5621 ( .A(n5938), .Y(n5936) );
  INVX1 U5622 ( .A(n5936), .Y(n5937) );
  AND2X1 U5623 ( .A(n8034), .B(n505), .Y(n537) );
  INVX1 U5624 ( .A(n537), .Y(n5938) );
  INVX1 U5625 ( .A(n5941), .Y(n5939) );
  INVX1 U5626 ( .A(n5939), .Y(n5940) );
  AND2X1 U5627 ( .A(n8037), .B(n505), .Y(n536) );
  INVX1 U5628 ( .A(n536), .Y(n5941) );
  INVX1 U5629 ( .A(n5944), .Y(n5942) );
  INVX1 U5630 ( .A(n5942), .Y(n5943) );
  AND2X1 U5631 ( .A(n8040), .B(n505), .Y(n535) );
  INVX1 U5632 ( .A(n535), .Y(n5944) );
  INVX1 U5633 ( .A(n5947), .Y(n5945) );
  INVX1 U5634 ( .A(n5945), .Y(n5946) );
  AND2X1 U5635 ( .A(n8043), .B(n505), .Y(n534) );
  INVX1 U5636 ( .A(n534), .Y(n5947) );
  INVX1 U5637 ( .A(n5950), .Y(n5948) );
  INVX1 U5638 ( .A(n5948), .Y(n5949) );
  AND2X1 U5639 ( .A(n8046), .B(n505), .Y(n533) );
  INVX1 U5640 ( .A(n533), .Y(n5950) );
  INVX1 U5641 ( .A(n5953), .Y(n5951) );
  INVX1 U5642 ( .A(n5951), .Y(n5952) );
  AND2X1 U5643 ( .A(n8049), .B(n505), .Y(n532) );
  INVX1 U5644 ( .A(n532), .Y(n5953) );
  INVX1 U5645 ( .A(n5956), .Y(n5954) );
  INVX1 U5646 ( .A(n5954), .Y(n5955) );
  AND2X1 U5647 ( .A(n8052), .B(n505), .Y(n531) );
  INVX1 U5648 ( .A(n531), .Y(n5956) );
  INVX1 U5649 ( .A(n5959), .Y(n5957) );
  INVX1 U5650 ( .A(n5957), .Y(n5958) );
  AND2X1 U5651 ( .A(n8055), .B(n505), .Y(n530) );
  INVX1 U5652 ( .A(n530), .Y(n5959) );
  INVX1 U5653 ( .A(n5962), .Y(n5960) );
  INVX1 U5654 ( .A(n5960), .Y(n5961) );
  AND2X1 U5655 ( .A(n8058), .B(n505), .Y(n529) );
  INVX1 U5656 ( .A(n529), .Y(n5962) );
  INVX1 U5657 ( .A(n5965), .Y(n5963) );
  INVX1 U5658 ( .A(n5963), .Y(n5964) );
  AND2X1 U5659 ( .A(n8061), .B(n505), .Y(n528) );
  INVX1 U5660 ( .A(n528), .Y(n5965) );
  INVX1 U5661 ( .A(n5968), .Y(n5966) );
  INVX1 U5662 ( .A(n5966), .Y(n5967) );
  AND2X1 U5663 ( .A(n8064), .B(n505), .Y(n527) );
  INVX1 U5664 ( .A(n527), .Y(n5968) );
  INVX1 U5665 ( .A(n5971), .Y(n5969) );
  INVX1 U5666 ( .A(n5969), .Y(n5970) );
  AND2X1 U5667 ( .A(n8067), .B(n505), .Y(n526) );
  INVX1 U5668 ( .A(n526), .Y(n5971) );
  INVX1 U5669 ( .A(n5974), .Y(n5972) );
  INVX1 U5670 ( .A(n5972), .Y(n5973) );
  AND2X1 U5671 ( .A(n8070), .B(n505), .Y(n525) );
  INVX1 U5672 ( .A(n525), .Y(n5974) );
  INVX1 U5673 ( .A(n5977), .Y(n5975) );
  INVX1 U5674 ( .A(n5975), .Y(n5976) );
  AND2X1 U5675 ( .A(n8073), .B(n505), .Y(n524) );
  INVX1 U5676 ( .A(n524), .Y(n5977) );
  INVX1 U5677 ( .A(n5980), .Y(n5978) );
  INVX1 U5678 ( .A(n5978), .Y(n5979) );
  AND2X1 U5679 ( .A(n8076), .B(n505), .Y(n523) );
  INVX1 U5680 ( .A(n523), .Y(n5980) );
  INVX1 U5681 ( .A(n5983), .Y(n5981) );
  INVX1 U5682 ( .A(n5981), .Y(n5982) );
  AND2X1 U5683 ( .A(n8079), .B(n505), .Y(n522) );
  INVX1 U5684 ( .A(n522), .Y(n5983) );
  INVX1 U5685 ( .A(n5986), .Y(n5984) );
  INVX1 U5686 ( .A(n5984), .Y(n5985) );
  AND2X1 U5687 ( .A(n8082), .B(n505), .Y(n521) );
  INVX1 U5688 ( .A(n521), .Y(n5986) );
  INVX1 U5689 ( .A(n5989), .Y(n5987) );
  INVX1 U5690 ( .A(n5987), .Y(n5988) );
  AND2X1 U5691 ( .A(n8085), .B(n505), .Y(n520) );
  INVX1 U5692 ( .A(n520), .Y(n5989) );
  INVX1 U5693 ( .A(n5992), .Y(n5990) );
  INVX1 U5694 ( .A(n5990), .Y(n5991) );
  AND2X1 U5695 ( .A(n8088), .B(n505), .Y(n519) );
  INVX1 U5696 ( .A(n519), .Y(n5992) );
  INVX1 U5697 ( .A(n5995), .Y(n5993) );
  INVX1 U5698 ( .A(n5993), .Y(n5994) );
  AND2X1 U5699 ( .A(n8091), .B(n505), .Y(n518) );
  INVX1 U5700 ( .A(n518), .Y(n5995) );
  INVX1 U5701 ( .A(n5998), .Y(n5996) );
  INVX1 U5702 ( .A(n5996), .Y(n5997) );
  AND2X1 U5703 ( .A(n8094), .B(n505), .Y(n517) );
  INVX1 U5704 ( .A(n517), .Y(n5998) );
  INVX1 U5705 ( .A(n6001), .Y(n5999) );
  INVX1 U5706 ( .A(n5999), .Y(n6000) );
  AND2X1 U5707 ( .A(n8097), .B(n505), .Y(n516) );
  INVX1 U5708 ( .A(n516), .Y(n6001) );
  INVX1 U5709 ( .A(n6004), .Y(n6002) );
  INVX1 U5710 ( .A(n6002), .Y(n6003) );
  AND2X1 U5711 ( .A(n8100), .B(n505), .Y(n515) );
  INVX1 U5712 ( .A(n515), .Y(n6004) );
  INVX1 U5713 ( .A(n6007), .Y(n6005) );
  INVX1 U5714 ( .A(n6005), .Y(n6006) );
  AND2X1 U5715 ( .A(n8103), .B(n505), .Y(n514) );
  INVX1 U5716 ( .A(n514), .Y(n6007) );
  INVX1 U5717 ( .A(n6010), .Y(n6008) );
  INVX1 U5718 ( .A(n6008), .Y(n6009) );
  AND2X1 U5719 ( .A(n8106), .B(n505), .Y(n513) );
  INVX1 U5720 ( .A(n513), .Y(n6010) );
  INVX1 U5721 ( .A(n6013), .Y(n6011) );
  INVX1 U5722 ( .A(n6011), .Y(n6012) );
  AND2X1 U5723 ( .A(n8109), .B(n505), .Y(n512) );
  INVX1 U5724 ( .A(n512), .Y(n6013) );
  INVX1 U5725 ( .A(n6016), .Y(n6014) );
  INVX1 U5726 ( .A(n6014), .Y(n6015) );
  AND2X1 U5727 ( .A(n8112), .B(n505), .Y(n511) );
  INVX1 U5728 ( .A(n511), .Y(n6016) );
  INVX1 U5729 ( .A(n6019), .Y(n6017) );
  INVX1 U5730 ( .A(n6017), .Y(n6018) );
  AND2X1 U5731 ( .A(n8115), .B(n505), .Y(n510) );
  INVX1 U5732 ( .A(n510), .Y(n6019) );
  INVX1 U5733 ( .A(n6022), .Y(n6020) );
  INVX1 U5734 ( .A(n6020), .Y(n6021) );
  AND2X1 U5735 ( .A(n8118), .B(n505), .Y(n509) );
  INVX1 U5736 ( .A(n509), .Y(n6022) );
  INVX1 U5737 ( .A(n6025), .Y(n6023) );
  INVX1 U5738 ( .A(n6023), .Y(n6024) );
  AND2X1 U5739 ( .A(n8121), .B(n505), .Y(n508) );
  INVX1 U5740 ( .A(n508), .Y(n6025) );
  INVX1 U5741 ( .A(n6028), .Y(n6026) );
  INVX1 U5742 ( .A(n6026), .Y(n6027) );
  AND2X1 U5743 ( .A(n8124), .B(n505), .Y(n507) );
  INVX1 U5744 ( .A(n507), .Y(n6028) );
  INVX1 U5745 ( .A(n6031), .Y(n6029) );
  INVX1 U5746 ( .A(n6029), .Y(n6030) );
  AND2X1 U5747 ( .A(n8127), .B(n505), .Y(n506) );
  INVX1 U5748 ( .A(n506), .Y(n6031) );
  INVX1 U5749 ( .A(n6034), .Y(n6032) );
  INVX1 U5750 ( .A(n6032), .Y(n6033) );
  AND2X1 U5751 ( .A(n9660), .B(n469), .Y(n503) );
  INVX1 U5752 ( .A(n503), .Y(n6034) );
  INVX1 U5753 ( .A(n6037), .Y(n6035) );
  INVX1 U5754 ( .A(n6035), .Y(n6036) );
  AND2X1 U5755 ( .A(n9663), .B(n469), .Y(n502) );
  INVX1 U5756 ( .A(n502), .Y(n6037) );
  INVX1 U5757 ( .A(n6040), .Y(n6038) );
  INVX1 U5758 ( .A(n6038), .Y(n6039) );
  AND2X1 U5759 ( .A(n9666), .B(n469), .Y(n501) );
  INVX1 U5760 ( .A(n501), .Y(n6040) );
  INVX1 U5761 ( .A(n6043), .Y(n6041) );
  INVX1 U5762 ( .A(n6041), .Y(n6042) );
  AND2X1 U5763 ( .A(n9669), .B(n469), .Y(n500) );
  INVX1 U5764 ( .A(n500), .Y(n6043) );
  INVX1 U5765 ( .A(n6046), .Y(n6044) );
  INVX1 U5766 ( .A(n6044), .Y(n6045) );
  AND2X1 U5767 ( .A(n9672), .B(n469), .Y(n499) );
  INVX1 U5768 ( .A(n499), .Y(n6046) );
  INVX1 U5769 ( .A(n6049), .Y(n6047) );
  INVX1 U5770 ( .A(n6047), .Y(n6048) );
  AND2X1 U5771 ( .A(n9675), .B(n469), .Y(n498) );
  INVX1 U5772 ( .A(n498), .Y(n6049) );
  INVX1 U5773 ( .A(n6052), .Y(n6050) );
  INVX1 U5774 ( .A(n6050), .Y(n6051) );
  AND2X1 U5775 ( .A(n9678), .B(n469), .Y(n497) );
  INVX1 U5776 ( .A(n497), .Y(n6052) );
  INVX1 U5777 ( .A(n6055), .Y(n6053) );
  INVX1 U5778 ( .A(n6053), .Y(n6054) );
  AND2X1 U5779 ( .A(n9681), .B(n469), .Y(n496) );
  INVX1 U5780 ( .A(n496), .Y(n6055) );
  INVX1 U5781 ( .A(n6058), .Y(n6056) );
  INVX1 U5782 ( .A(n6056), .Y(n6057) );
  AND2X1 U5783 ( .A(n9684), .B(n469), .Y(n495) );
  INVX1 U5784 ( .A(n495), .Y(n6058) );
  INVX1 U5785 ( .A(n6061), .Y(n6059) );
  INVX1 U5786 ( .A(n6059), .Y(n6060) );
  AND2X1 U5787 ( .A(n9687), .B(n469), .Y(n494) );
  INVX1 U5788 ( .A(n494), .Y(n6061) );
  INVX1 U5789 ( .A(n6064), .Y(n6062) );
  INVX1 U5790 ( .A(n6062), .Y(n6063) );
  AND2X1 U5791 ( .A(n9690), .B(n469), .Y(n493) );
  INVX1 U5792 ( .A(n493), .Y(n6064) );
  INVX1 U5793 ( .A(n6067), .Y(n6065) );
  INVX1 U5794 ( .A(n6065), .Y(n6066) );
  AND2X1 U5795 ( .A(n9693), .B(n469), .Y(n492) );
  INVX1 U5796 ( .A(n492), .Y(n6067) );
  INVX1 U5797 ( .A(n6070), .Y(n6068) );
  INVX1 U5798 ( .A(n6068), .Y(n6069) );
  AND2X1 U5799 ( .A(n9696), .B(n469), .Y(n491) );
  INVX1 U5800 ( .A(n491), .Y(n6070) );
  INVX1 U5801 ( .A(n6073), .Y(n6071) );
  INVX1 U5802 ( .A(n6071), .Y(n6072) );
  AND2X1 U5803 ( .A(n9699), .B(n469), .Y(n490) );
  INVX1 U5804 ( .A(n490), .Y(n6073) );
  INVX1 U5805 ( .A(n6076), .Y(n6074) );
  INVX1 U5806 ( .A(n6074), .Y(n6075) );
  AND2X1 U5807 ( .A(n9702), .B(n469), .Y(n489) );
  INVX1 U5808 ( .A(n489), .Y(n6076) );
  INVX1 U5809 ( .A(n6079), .Y(n6077) );
  INVX1 U5810 ( .A(n6077), .Y(n6078) );
  AND2X1 U5811 ( .A(n9705), .B(n469), .Y(n488) );
  INVX1 U5812 ( .A(n488), .Y(n6079) );
  INVX1 U5813 ( .A(n6082), .Y(n6080) );
  INVX1 U5814 ( .A(n6080), .Y(n6081) );
  AND2X1 U5815 ( .A(n9708), .B(n469), .Y(n487) );
  INVX1 U5816 ( .A(n487), .Y(n6082) );
  INVX1 U5817 ( .A(n6085), .Y(n6083) );
  INVX1 U5818 ( .A(n6083), .Y(n6084) );
  AND2X1 U5819 ( .A(n9711), .B(n469), .Y(n486) );
  INVX1 U5820 ( .A(n486), .Y(n6085) );
  INVX1 U5821 ( .A(n6088), .Y(n6086) );
  INVX1 U5822 ( .A(n6086), .Y(n6087) );
  AND2X1 U5823 ( .A(n9714), .B(n469), .Y(n485) );
  INVX1 U5824 ( .A(n485), .Y(n6088) );
  INVX1 U5825 ( .A(n6091), .Y(n6089) );
  INVX1 U5826 ( .A(n6089), .Y(n6090) );
  AND2X1 U5827 ( .A(n9717), .B(n469), .Y(n484) );
  INVX1 U5828 ( .A(n484), .Y(n6091) );
  INVX1 U5829 ( .A(n6094), .Y(n6092) );
  INVX1 U5830 ( .A(n6092), .Y(n6093) );
  AND2X1 U5831 ( .A(n9720), .B(n469), .Y(n483) );
  INVX1 U5832 ( .A(n483), .Y(n6094) );
  INVX1 U5833 ( .A(n6097), .Y(n6095) );
  INVX1 U5834 ( .A(n6095), .Y(n6096) );
  AND2X1 U5835 ( .A(n9723), .B(n469), .Y(n482) );
  INVX1 U5836 ( .A(n482), .Y(n6097) );
  INVX1 U5837 ( .A(n6100), .Y(n6098) );
  INVX1 U5838 ( .A(n6098), .Y(n6099) );
  AND2X1 U5839 ( .A(n9726), .B(n469), .Y(n481) );
  INVX1 U5840 ( .A(n481), .Y(n6100) );
  INVX1 U5841 ( .A(n6103), .Y(n6101) );
  INVX1 U5842 ( .A(n6101), .Y(n6102) );
  AND2X1 U5843 ( .A(n9729), .B(n469), .Y(n480) );
  INVX1 U5844 ( .A(n480), .Y(n6103) );
  INVX1 U5845 ( .A(n6106), .Y(n6104) );
  INVX1 U5846 ( .A(n6104), .Y(n6105) );
  AND2X1 U5847 ( .A(n9732), .B(n469), .Y(n479) );
  INVX1 U5848 ( .A(n479), .Y(n6106) );
  INVX1 U5849 ( .A(n6109), .Y(n6107) );
  INVX1 U5850 ( .A(n6107), .Y(n6108) );
  AND2X1 U5851 ( .A(n9735), .B(n469), .Y(n478) );
  INVX1 U5852 ( .A(n478), .Y(n6109) );
  INVX1 U5853 ( .A(n6112), .Y(n6110) );
  INVX1 U5854 ( .A(n6110), .Y(n6111) );
  AND2X1 U5855 ( .A(n9738), .B(n469), .Y(n477) );
  INVX1 U5856 ( .A(n477), .Y(n6112) );
  INVX1 U5857 ( .A(n6115), .Y(n6113) );
  INVX1 U5858 ( .A(n6113), .Y(n6114) );
  AND2X1 U5859 ( .A(n9741), .B(n469), .Y(n476) );
  INVX1 U5860 ( .A(n476), .Y(n6115) );
  INVX1 U5861 ( .A(n6118), .Y(n6116) );
  INVX1 U5862 ( .A(n6116), .Y(n6117) );
  AND2X1 U5863 ( .A(n9744), .B(n469), .Y(n475) );
  INVX1 U5864 ( .A(n475), .Y(n6118) );
  INVX1 U5865 ( .A(n6121), .Y(n6119) );
  INVX1 U5866 ( .A(n6119), .Y(n6120) );
  AND2X1 U5867 ( .A(n9747), .B(n469), .Y(n474) );
  INVX1 U5868 ( .A(n474), .Y(n6121) );
  INVX1 U5869 ( .A(n6124), .Y(n6122) );
  INVX1 U5870 ( .A(n6122), .Y(n6123) );
  AND2X1 U5871 ( .A(n9750), .B(n469), .Y(n473) );
  INVX1 U5872 ( .A(n473), .Y(n6124) );
  INVX1 U5873 ( .A(n6127), .Y(n6125) );
  INVX1 U5874 ( .A(n6125), .Y(n6126) );
  AND2X1 U5875 ( .A(n9753), .B(n469), .Y(n472) );
  INVX1 U5876 ( .A(n472), .Y(n6127) );
  INVX1 U5877 ( .A(n6130), .Y(n6128) );
  INVX1 U5878 ( .A(n6128), .Y(n6129) );
  AND2X1 U5879 ( .A(n9756), .B(n469), .Y(n471) );
  INVX1 U5880 ( .A(n471), .Y(n6130) );
  INVX1 U5881 ( .A(n6133), .Y(n6131) );
  INVX1 U5882 ( .A(n6131), .Y(n6132) );
  AND2X1 U5883 ( .A(n9759), .B(n469), .Y(n470) );
  INVX1 U5884 ( .A(n470), .Y(n6133) );
  INVX1 U5885 ( .A(n6136), .Y(n6134) );
  INVX1 U5886 ( .A(n6134), .Y(n6135) );
  AND2X1 U5887 ( .A(n8130), .B(n433), .Y(n467) );
  INVX1 U5888 ( .A(n467), .Y(n6136) );
  INVX1 U5889 ( .A(n6139), .Y(n6137) );
  INVX1 U5890 ( .A(n6137), .Y(n6138) );
  AND2X1 U5891 ( .A(n8133), .B(n433), .Y(n466) );
  INVX1 U5892 ( .A(n466), .Y(n6139) );
  INVX1 U5893 ( .A(n6142), .Y(n6140) );
  INVX1 U5894 ( .A(n6140), .Y(n6141) );
  AND2X1 U5895 ( .A(n8136), .B(n433), .Y(n465) );
  INVX1 U5896 ( .A(n465), .Y(n6142) );
  INVX1 U5897 ( .A(n6145), .Y(n6143) );
  INVX1 U5898 ( .A(n6143), .Y(n6144) );
  AND2X1 U5899 ( .A(n8139), .B(n433), .Y(n464) );
  INVX1 U5900 ( .A(n464), .Y(n6145) );
  INVX1 U5901 ( .A(n6148), .Y(n6146) );
  INVX1 U5902 ( .A(n6146), .Y(n6147) );
  AND2X1 U5903 ( .A(n8142), .B(n433), .Y(n463) );
  INVX1 U5904 ( .A(n463), .Y(n6148) );
  INVX1 U5905 ( .A(n6151), .Y(n6149) );
  INVX1 U5906 ( .A(n6149), .Y(n6150) );
  AND2X1 U5907 ( .A(n8145), .B(n433), .Y(n462) );
  INVX1 U5908 ( .A(n462), .Y(n6151) );
  INVX1 U5909 ( .A(n6154), .Y(n6152) );
  INVX1 U5910 ( .A(n6152), .Y(n6153) );
  AND2X1 U5911 ( .A(n8148), .B(n433), .Y(n461) );
  INVX1 U5912 ( .A(n461), .Y(n6154) );
  INVX1 U5913 ( .A(n6157), .Y(n6155) );
  INVX1 U5914 ( .A(n6155), .Y(n6156) );
  AND2X1 U5915 ( .A(n8151), .B(n433), .Y(n460) );
  INVX1 U5916 ( .A(n460), .Y(n6157) );
  INVX1 U5917 ( .A(n6160), .Y(n6158) );
  INVX1 U5918 ( .A(n6158), .Y(n6159) );
  AND2X1 U5919 ( .A(n8154), .B(n433), .Y(n459) );
  INVX1 U5920 ( .A(n459), .Y(n6160) );
  INVX1 U5921 ( .A(n6163), .Y(n6161) );
  INVX1 U5922 ( .A(n6161), .Y(n6162) );
  AND2X1 U5923 ( .A(n8157), .B(n433), .Y(n458) );
  INVX1 U5924 ( .A(n458), .Y(n6163) );
  INVX1 U5925 ( .A(n6166), .Y(n6164) );
  INVX1 U5926 ( .A(n6164), .Y(n6165) );
  AND2X1 U5927 ( .A(n8160), .B(n433), .Y(n457) );
  INVX1 U5928 ( .A(n457), .Y(n6166) );
  INVX1 U5929 ( .A(n6169), .Y(n6167) );
  INVX1 U5930 ( .A(n6167), .Y(n6168) );
  AND2X1 U5931 ( .A(n8163), .B(n433), .Y(n456) );
  INVX1 U5932 ( .A(n456), .Y(n6169) );
  INVX1 U5933 ( .A(n6172), .Y(n6170) );
  INVX1 U5934 ( .A(n6170), .Y(n6171) );
  AND2X1 U5935 ( .A(n8166), .B(n433), .Y(n455) );
  INVX1 U5936 ( .A(n455), .Y(n6172) );
  INVX1 U5937 ( .A(n6175), .Y(n6173) );
  INVX1 U5938 ( .A(n6173), .Y(n6174) );
  AND2X1 U5939 ( .A(n8169), .B(n433), .Y(n454) );
  INVX1 U5940 ( .A(n454), .Y(n6175) );
  INVX1 U5941 ( .A(n6178), .Y(n6176) );
  INVX1 U5942 ( .A(n6176), .Y(n6177) );
  AND2X1 U5943 ( .A(n8172), .B(n433), .Y(n453) );
  INVX1 U5944 ( .A(n453), .Y(n6178) );
  INVX1 U5945 ( .A(n6181), .Y(n6179) );
  INVX1 U5946 ( .A(n6179), .Y(n6180) );
  AND2X1 U5947 ( .A(n8175), .B(n433), .Y(n452) );
  INVX1 U5948 ( .A(n452), .Y(n6181) );
  INVX1 U5949 ( .A(n6184), .Y(n6182) );
  INVX1 U5950 ( .A(n6182), .Y(n6183) );
  AND2X1 U5951 ( .A(n8178), .B(n433), .Y(n451) );
  INVX1 U5952 ( .A(n451), .Y(n6184) );
  INVX1 U5953 ( .A(n6187), .Y(n6185) );
  INVX1 U5954 ( .A(n6185), .Y(n6186) );
  AND2X1 U5955 ( .A(n8181), .B(n433), .Y(n450) );
  INVX1 U5956 ( .A(n450), .Y(n6187) );
  INVX1 U5957 ( .A(n6190), .Y(n6188) );
  INVX1 U5958 ( .A(n6188), .Y(n6189) );
  AND2X1 U5959 ( .A(n8184), .B(n433), .Y(n449) );
  INVX1 U5960 ( .A(n449), .Y(n6190) );
  INVX1 U5961 ( .A(n6193), .Y(n6191) );
  INVX1 U5962 ( .A(n6191), .Y(n6192) );
  AND2X1 U5963 ( .A(n8187), .B(n433), .Y(n448) );
  INVX1 U5964 ( .A(n448), .Y(n6193) );
  INVX1 U5965 ( .A(n6196), .Y(n6194) );
  INVX1 U5966 ( .A(n6194), .Y(n6195) );
  AND2X1 U5967 ( .A(n8190), .B(n433), .Y(n447) );
  INVX1 U5968 ( .A(n447), .Y(n6196) );
  INVX1 U5969 ( .A(n6199), .Y(n6197) );
  INVX1 U5970 ( .A(n6197), .Y(n6198) );
  AND2X1 U5971 ( .A(n8193), .B(n433), .Y(n446) );
  INVX1 U5972 ( .A(n446), .Y(n6199) );
  INVX1 U5973 ( .A(n6202), .Y(n6200) );
  INVX1 U5974 ( .A(n6200), .Y(n6201) );
  AND2X1 U5975 ( .A(n8196), .B(n433), .Y(n445) );
  INVX1 U5976 ( .A(n445), .Y(n6202) );
  INVX1 U5977 ( .A(n6205), .Y(n6203) );
  INVX1 U5978 ( .A(n6203), .Y(n6204) );
  AND2X1 U5979 ( .A(n8199), .B(n433), .Y(n444) );
  INVX1 U5980 ( .A(n444), .Y(n6205) );
  INVX1 U5981 ( .A(n6208), .Y(n6206) );
  INVX1 U5982 ( .A(n6206), .Y(n6207) );
  AND2X1 U5983 ( .A(n8202), .B(n433), .Y(n443) );
  INVX1 U5984 ( .A(n443), .Y(n6208) );
  INVX1 U5985 ( .A(n6211), .Y(n6209) );
  INVX1 U5986 ( .A(n6209), .Y(n6210) );
  AND2X1 U5987 ( .A(n8205), .B(n433), .Y(n442) );
  INVX1 U5988 ( .A(n442), .Y(n6211) );
  INVX1 U5989 ( .A(n6214), .Y(n6212) );
  INVX1 U5990 ( .A(n6212), .Y(n6213) );
  AND2X1 U5991 ( .A(n8208), .B(n433), .Y(n441) );
  INVX1 U5992 ( .A(n441), .Y(n6214) );
  INVX1 U5993 ( .A(n6217), .Y(n6215) );
  INVX1 U5994 ( .A(n6215), .Y(n6216) );
  AND2X1 U5995 ( .A(n8211), .B(n433), .Y(n440) );
  INVX1 U5996 ( .A(n440), .Y(n6217) );
  INVX1 U5997 ( .A(n6220), .Y(n6218) );
  INVX1 U5998 ( .A(n6218), .Y(n6219) );
  AND2X1 U5999 ( .A(n8214), .B(n433), .Y(n439) );
  INVX1 U6000 ( .A(n439), .Y(n6220) );
  INVX1 U6001 ( .A(n6223), .Y(n6221) );
  INVX1 U6002 ( .A(n6221), .Y(n6222) );
  AND2X1 U6003 ( .A(n8217), .B(n433), .Y(n438) );
  INVX1 U6004 ( .A(n438), .Y(n6223) );
  INVX1 U6005 ( .A(n6226), .Y(n6224) );
  INVX1 U6006 ( .A(n6224), .Y(n6225) );
  AND2X1 U6007 ( .A(n8220), .B(n433), .Y(n437) );
  INVX1 U6008 ( .A(n437), .Y(n6226) );
  INVX1 U6009 ( .A(n6229), .Y(n6227) );
  INVX1 U6010 ( .A(n6227), .Y(n6228) );
  AND2X1 U6011 ( .A(n8223), .B(n433), .Y(n436) );
  INVX1 U6012 ( .A(n436), .Y(n6229) );
  INVX1 U6013 ( .A(n6232), .Y(n6230) );
  INVX1 U6014 ( .A(n6230), .Y(n6231) );
  AND2X1 U6015 ( .A(n8226), .B(n433), .Y(n435) );
  INVX1 U6016 ( .A(n435), .Y(n6232) );
  INVX1 U6017 ( .A(n6235), .Y(n6233) );
  INVX1 U6018 ( .A(n6233), .Y(n6234) );
  AND2X1 U6019 ( .A(n8229), .B(n433), .Y(n434) );
  INVX1 U6020 ( .A(n434), .Y(n6235) );
  INVX1 U6021 ( .A(n6238), .Y(n6236) );
  INVX1 U6022 ( .A(n6236), .Y(n6237) );
  AND2X1 U6023 ( .A(n9762), .B(n397), .Y(n431) );
  INVX1 U6024 ( .A(n431), .Y(n6238) );
  INVX1 U6025 ( .A(n6241), .Y(n6239) );
  INVX1 U6026 ( .A(n6239), .Y(n6240) );
  AND2X1 U6027 ( .A(n9765), .B(n397), .Y(n430) );
  INVX1 U6028 ( .A(n430), .Y(n6241) );
  INVX1 U6029 ( .A(n6244), .Y(n6242) );
  INVX1 U6030 ( .A(n6242), .Y(n6243) );
  AND2X1 U6031 ( .A(n9768), .B(n397), .Y(n429) );
  INVX1 U6032 ( .A(n429), .Y(n6244) );
  INVX1 U6033 ( .A(n6247), .Y(n6245) );
  INVX1 U6034 ( .A(n6245), .Y(n6246) );
  AND2X1 U6035 ( .A(n9771), .B(n397), .Y(n428) );
  INVX1 U6036 ( .A(n428), .Y(n6247) );
  INVX1 U6037 ( .A(n6250), .Y(n6248) );
  INVX1 U6038 ( .A(n6248), .Y(n6249) );
  AND2X1 U6039 ( .A(n9774), .B(n397), .Y(n427) );
  INVX1 U6040 ( .A(n427), .Y(n6250) );
  INVX1 U6041 ( .A(n6253), .Y(n6251) );
  INVX1 U6042 ( .A(n6251), .Y(n6252) );
  AND2X1 U6043 ( .A(n9777), .B(n397), .Y(n426) );
  INVX1 U6044 ( .A(n426), .Y(n6253) );
  INVX1 U6045 ( .A(n6256), .Y(n6254) );
  INVX1 U6046 ( .A(n6254), .Y(n6255) );
  AND2X1 U6047 ( .A(n9780), .B(n397), .Y(n425) );
  INVX1 U6048 ( .A(n425), .Y(n6256) );
  INVX1 U6049 ( .A(n6259), .Y(n6257) );
  INVX1 U6050 ( .A(n6257), .Y(n6258) );
  AND2X1 U6051 ( .A(n9783), .B(n397), .Y(n424) );
  INVX1 U6052 ( .A(n424), .Y(n6259) );
  INVX1 U6053 ( .A(n6262), .Y(n6260) );
  INVX1 U6054 ( .A(n6260), .Y(n6261) );
  AND2X1 U6055 ( .A(n9786), .B(n397), .Y(n423) );
  INVX1 U6056 ( .A(n423), .Y(n6262) );
  INVX1 U6057 ( .A(n6265), .Y(n6263) );
  INVX1 U6058 ( .A(n6263), .Y(n6264) );
  AND2X1 U6059 ( .A(n9789), .B(n397), .Y(n422) );
  INVX1 U6060 ( .A(n422), .Y(n6265) );
  INVX1 U6061 ( .A(n6268), .Y(n6266) );
  INVX1 U6062 ( .A(n6266), .Y(n6267) );
  AND2X1 U6063 ( .A(n9792), .B(n397), .Y(n421) );
  INVX1 U6064 ( .A(n421), .Y(n6268) );
  INVX1 U6065 ( .A(n6271), .Y(n6269) );
  INVX1 U6066 ( .A(n6269), .Y(n6270) );
  AND2X1 U6067 ( .A(n9795), .B(n397), .Y(n420) );
  INVX1 U6068 ( .A(n420), .Y(n6271) );
  INVX1 U6069 ( .A(n6274), .Y(n6272) );
  INVX1 U6070 ( .A(n6272), .Y(n6273) );
  AND2X1 U6071 ( .A(n9798), .B(n397), .Y(n419) );
  INVX1 U6072 ( .A(n419), .Y(n6274) );
  INVX1 U6073 ( .A(n6277), .Y(n6275) );
  INVX1 U6074 ( .A(n6275), .Y(n6276) );
  AND2X1 U6075 ( .A(n9801), .B(n397), .Y(n418) );
  INVX1 U6076 ( .A(n418), .Y(n6277) );
  INVX1 U6077 ( .A(n6280), .Y(n6278) );
  INVX1 U6078 ( .A(n6278), .Y(n6279) );
  AND2X1 U6079 ( .A(n9804), .B(n397), .Y(n417) );
  INVX1 U6080 ( .A(n417), .Y(n6280) );
  INVX1 U6081 ( .A(n6283), .Y(n6281) );
  INVX1 U6082 ( .A(n6281), .Y(n6282) );
  AND2X1 U6083 ( .A(n9807), .B(n397), .Y(n416) );
  INVX1 U6084 ( .A(n416), .Y(n6283) );
  INVX1 U6085 ( .A(n6286), .Y(n6284) );
  INVX1 U6086 ( .A(n6284), .Y(n6285) );
  AND2X1 U6087 ( .A(n9810), .B(n397), .Y(n415) );
  INVX1 U6088 ( .A(n415), .Y(n6286) );
  INVX1 U6089 ( .A(n6289), .Y(n6287) );
  INVX1 U6090 ( .A(n6287), .Y(n6288) );
  AND2X1 U6091 ( .A(n9813), .B(n397), .Y(n414) );
  INVX1 U6092 ( .A(n414), .Y(n6289) );
  INVX1 U6093 ( .A(n6292), .Y(n6290) );
  INVX1 U6094 ( .A(n6290), .Y(n6291) );
  AND2X1 U6095 ( .A(n9816), .B(n397), .Y(n413) );
  INVX1 U6096 ( .A(n413), .Y(n6292) );
  INVX1 U6097 ( .A(n6295), .Y(n6293) );
  INVX1 U6098 ( .A(n6293), .Y(n6294) );
  AND2X1 U6099 ( .A(n9819), .B(n397), .Y(n412) );
  INVX1 U6100 ( .A(n412), .Y(n6295) );
  INVX1 U6101 ( .A(n6298), .Y(n6296) );
  INVX1 U6102 ( .A(n6296), .Y(n6297) );
  AND2X1 U6103 ( .A(n9822), .B(n397), .Y(n411) );
  INVX1 U6104 ( .A(n411), .Y(n6298) );
  INVX1 U6105 ( .A(n6301), .Y(n6299) );
  INVX1 U6106 ( .A(n6299), .Y(n6300) );
  AND2X1 U6107 ( .A(n9825), .B(n397), .Y(n410) );
  INVX1 U6108 ( .A(n410), .Y(n6301) );
  INVX1 U6109 ( .A(n6304), .Y(n6302) );
  INVX1 U6110 ( .A(n6302), .Y(n6303) );
  AND2X1 U6111 ( .A(n9828), .B(n397), .Y(n409) );
  INVX1 U6112 ( .A(n409), .Y(n6304) );
  INVX1 U6113 ( .A(n6307), .Y(n6305) );
  INVX1 U6114 ( .A(n6305), .Y(n6306) );
  AND2X1 U6115 ( .A(n9831), .B(n397), .Y(n408) );
  INVX1 U6116 ( .A(n408), .Y(n6307) );
  INVX1 U6117 ( .A(n6310), .Y(n6308) );
  INVX1 U6118 ( .A(n6308), .Y(n6309) );
  AND2X1 U6119 ( .A(n9834), .B(n397), .Y(n407) );
  INVX1 U6120 ( .A(n407), .Y(n6310) );
  INVX1 U6121 ( .A(n6313), .Y(n6311) );
  INVX1 U6122 ( .A(n6311), .Y(n6312) );
  AND2X1 U6123 ( .A(n9837), .B(n397), .Y(n406) );
  INVX1 U6124 ( .A(n406), .Y(n6313) );
  INVX1 U6125 ( .A(n6316), .Y(n6314) );
  INVX1 U6126 ( .A(n6314), .Y(n6315) );
  AND2X1 U6127 ( .A(n9840), .B(n397), .Y(n405) );
  INVX1 U6128 ( .A(n405), .Y(n6316) );
  INVX1 U6129 ( .A(n6319), .Y(n6317) );
  INVX1 U6130 ( .A(n6317), .Y(n6318) );
  AND2X1 U6131 ( .A(n9843), .B(n397), .Y(n404) );
  INVX1 U6132 ( .A(n404), .Y(n6319) );
  INVX1 U6133 ( .A(n6322), .Y(n6320) );
  INVX1 U6134 ( .A(n6320), .Y(n6321) );
  AND2X1 U6135 ( .A(n9846), .B(n397), .Y(n403) );
  INVX1 U6136 ( .A(n403), .Y(n6322) );
  INVX1 U6137 ( .A(n6325), .Y(n6323) );
  INVX1 U6138 ( .A(n6323), .Y(n6324) );
  AND2X1 U6139 ( .A(n9849), .B(n397), .Y(n402) );
  INVX1 U6140 ( .A(n402), .Y(n6325) );
  INVX1 U6141 ( .A(n6328), .Y(n6326) );
  INVX1 U6142 ( .A(n6326), .Y(n6327) );
  AND2X1 U6143 ( .A(n9852), .B(n397), .Y(n401) );
  INVX1 U6144 ( .A(n401), .Y(n6328) );
  INVX1 U6145 ( .A(n6331), .Y(n6329) );
  INVX1 U6146 ( .A(n6329), .Y(n6330) );
  AND2X1 U6147 ( .A(n9855), .B(n397), .Y(n400) );
  INVX1 U6148 ( .A(n400), .Y(n6331) );
  INVX1 U6149 ( .A(n6334), .Y(n6332) );
  INVX1 U6150 ( .A(n6332), .Y(n6333) );
  AND2X1 U6151 ( .A(n9858), .B(n397), .Y(n399) );
  INVX1 U6152 ( .A(n399), .Y(n6334) );
  INVX1 U6153 ( .A(n6337), .Y(n6335) );
  INVX1 U6154 ( .A(n6335), .Y(n6336) );
  AND2X1 U6155 ( .A(n9861), .B(n397), .Y(n398) );
  INVX1 U6156 ( .A(n398), .Y(n6337) );
  INVX1 U6157 ( .A(n6340), .Y(n6338) );
  INVX1 U6158 ( .A(n6338), .Y(n6339) );
  AND2X1 U6159 ( .A(n8232), .B(n361), .Y(n395) );
  INVX1 U6160 ( .A(n395), .Y(n6340) );
  INVX1 U6161 ( .A(n6343), .Y(n6341) );
  INVX1 U6162 ( .A(n6341), .Y(n6342) );
  AND2X1 U6163 ( .A(n8235), .B(n361), .Y(n394) );
  INVX1 U6164 ( .A(n394), .Y(n6343) );
  INVX1 U6165 ( .A(n6346), .Y(n6344) );
  INVX1 U6166 ( .A(n6344), .Y(n6345) );
  AND2X1 U6167 ( .A(n8238), .B(n361), .Y(n393) );
  INVX1 U6168 ( .A(n393), .Y(n6346) );
  INVX1 U6169 ( .A(n6349), .Y(n6347) );
  INVX1 U6170 ( .A(n6347), .Y(n6348) );
  AND2X1 U6171 ( .A(n8241), .B(n361), .Y(n392) );
  INVX1 U6172 ( .A(n392), .Y(n6349) );
  INVX1 U6173 ( .A(n6352), .Y(n6350) );
  INVX1 U6174 ( .A(n6350), .Y(n6351) );
  AND2X1 U6175 ( .A(n8244), .B(n361), .Y(n391) );
  INVX1 U6176 ( .A(n391), .Y(n6352) );
  INVX1 U6177 ( .A(n6355), .Y(n6353) );
  INVX1 U6178 ( .A(n6353), .Y(n6354) );
  AND2X1 U6179 ( .A(n8247), .B(n361), .Y(n390) );
  INVX1 U6180 ( .A(n390), .Y(n6355) );
  INVX1 U6181 ( .A(n6358), .Y(n6356) );
  INVX1 U6182 ( .A(n6356), .Y(n6357) );
  AND2X1 U6183 ( .A(n8250), .B(n361), .Y(n389) );
  INVX1 U6184 ( .A(n389), .Y(n6358) );
  INVX1 U6185 ( .A(n6361), .Y(n6359) );
  INVX1 U6186 ( .A(n6359), .Y(n6360) );
  AND2X1 U6187 ( .A(n8253), .B(n361), .Y(n388) );
  INVX1 U6188 ( .A(n388), .Y(n6361) );
  INVX1 U6189 ( .A(n6364), .Y(n6362) );
  INVX1 U6190 ( .A(n6362), .Y(n6363) );
  AND2X1 U6191 ( .A(n8256), .B(n361), .Y(n387) );
  INVX1 U6192 ( .A(n387), .Y(n6364) );
  INVX1 U6193 ( .A(n6367), .Y(n6365) );
  INVX1 U6194 ( .A(n6365), .Y(n6366) );
  AND2X1 U6195 ( .A(n8259), .B(n361), .Y(n386) );
  INVX1 U6196 ( .A(n386), .Y(n6367) );
  INVX1 U6197 ( .A(n6370), .Y(n6368) );
  INVX1 U6198 ( .A(n6368), .Y(n6369) );
  AND2X1 U6199 ( .A(n8262), .B(n361), .Y(n385) );
  INVX1 U6200 ( .A(n385), .Y(n6370) );
  INVX1 U6201 ( .A(n6373), .Y(n6371) );
  INVX1 U6202 ( .A(n6371), .Y(n6372) );
  AND2X1 U6203 ( .A(n8265), .B(n361), .Y(n384) );
  INVX1 U6204 ( .A(n384), .Y(n6373) );
  INVX1 U6205 ( .A(n6376), .Y(n6374) );
  INVX1 U6206 ( .A(n6374), .Y(n6375) );
  AND2X1 U6207 ( .A(n8268), .B(n361), .Y(n383) );
  INVX1 U6208 ( .A(n383), .Y(n6376) );
  INVX1 U6209 ( .A(n6379), .Y(n6377) );
  INVX1 U6210 ( .A(n6377), .Y(n6378) );
  AND2X1 U6211 ( .A(n8271), .B(n361), .Y(n382) );
  INVX1 U6212 ( .A(n382), .Y(n6379) );
  INVX1 U6213 ( .A(n6382), .Y(n6380) );
  INVX1 U6214 ( .A(n6380), .Y(n6381) );
  AND2X1 U6215 ( .A(n8274), .B(n361), .Y(n381) );
  INVX1 U6216 ( .A(n381), .Y(n6382) );
  INVX1 U6217 ( .A(n6385), .Y(n6383) );
  INVX1 U6218 ( .A(n6383), .Y(n6384) );
  AND2X1 U6219 ( .A(n8277), .B(n361), .Y(n380) );
  INVX1 U6220 ( .A(n380), .Y(n6385) );
  INVX1 U6221 ( .A(n6388), .Y(n6386) );
  INVX1 U6222 ( .A(n6386), .Y(n6387) );
  AND2X1 U6223 ( .A(n8280), .B(n361), .Y(n379) );
  INVX1 U6224 ( .A(n379), .Y(n6388) );
  INVX1 U6225 ( .A(n6391), .Y(n6389) );
  INVX1 U6226 ( .A(n6389), .Y(n6390) );
  AND2X1 U6227 ( .A(n8283), .B(n361), .Y(n378) );
  INVX1 U6228 ( .A(n378), .Y(n6391) );
  INVX1 U6229 ( .A(n6394), .Y(n6392) );
  INVX1 U6230 ( .A(n6392), .Y(n6393) );
  AND2X1 U6231 ( .A(n8286), .B(n361), .Y(n377) );
  INVX1 U6232 ( .A(n377), .Y(n6394) );
  INVX1 U6233 ( .A(n6397), .Y(n6395) );
  INVX1 U6234 ( .A(n6395), .Y(n6396) );
  AND2X1 U6235 ( .A(n8289), .B(n361), .Y(n376) );
  INVX1 U6236 ( .A(n376), .Y(n6397) );
  INVX1 U6237 ( .A(n6400), .Y(n6398) );
  INVX1 U6238 ( .A(n6398), .Y(n6399) );
  AND2X1 U6239 ( .A(n8292), .B(n361), .Y(n375) );
  INVX1 U6240 ( .A(n375), .Y(n6400) );
  INVX1 U6241 ( .A(n6403), .Y(n6401) );
  INVX1 U6242 ( .A(n6401), .Y(n6402) );
  AND2X1 U6243 ( .A(n8295), .B(n361), .Y(n374) );
  INVX1 U6244 ( .A(n374), .Y(n6403) );
  INVX1 U6245 ( .A(n6406), .Y(n6404) );
  INVX1 U6246 ( .A(n6404), .Y(n6405) );
  AND2X1 U6247 ( .A(n8298), .B(n361), .Y(n373) );
  INVX1 U6248 ( .A(n373), .Y(n6406) );
  INVX1 U6249 ( .A(n6409), .Y(n6407) );
  INVX1 U6250 ( .A(n6407), .Y(n6408) );
  AND2X1 U6251 ( .A(n8301), .B(n361), .Y(n372) );
  INVX1 U6252 ( .A(n372), .Y(n6409) );
  INVX1 U6253 ( .A(n6412), .Y(n6410) );
  INVX1 U6254 ( .A(n6410), .Y(n6411) );
  AND2X1 U6255 ( .A(n8304), .B(n361), .Y(n371) );
  INVX1 U6256 ( .A(n371), .Y(n6412) );
  INVX1 U6257 ( .A(n6415), .Y(n6413) );
  INVX1 U6258 ( .A(n6413), .Y(n6414) );
  AND2X1 U6259 ( .A(n8307), .B(n361), .Y(n370) );
  INVX1 U6260 ( .A(n370), .Y(n6415) );
  INVX1 U6261 ( .A(n6418), .Y(n6416) );
  INVX1 U6262 ( .A(n6416), .Y(n6417) );
  AND2X1 U6263 ( .A(n8310), .B(n361), .Y(n369) );
  INVX1 U6264 ( .A(n369), .Y(n6418) );
  INVX1 U6265 ( .A(n6421), .Y(n6419) );
  INVX1 U6266 ( .A(n6419), .Y(n6420) );
  AND2X1 U6267 ( .A(n8313), .B(n361), .Y(n368) );
  INVX1 U6268 ( .A(n368), .Y(n6421) );
  INVX1 U6269 ( .A(n6424), .Y(n6422) );
  INVX1 U6270 ( .A(n6422), .Y(n6423) );
  AND2X1 U6271 ( .A(n8316), .B(n361), .Y(n367) );
  INVX1 U6272 ( .A(n367), .Y(n6424) );
  INVX1 U6273 ( .A(n6427), .Y(n6425) );
  INVX1 U6274 ( .A(n6425), .Y(n6426) );
  AND2X1 U6275 ( .A(n8319), .B(n361), .Y(n366) );
  INVX1 U6276 ( .A(n366), .Y(n6427) );
  INVX1 U6277 ( .A(n6430), .Y(n6428) );
  INVX1 U6278 ( .A(n6428), .Y(n6429) );
  AND2X1 U6279 ( .A(n8322), .B(n361), .Y(n365) );
  INVX1 U6280 ( .A(n365), .Y(n6430) );
  INVX1 U6281 ( .A(n6433), .Y(n6431) );
  INVX1 U6282 ( .A(n6431), .Y(n6432) );
  AND2X1 U6283 ( .A(n8325), .B(n361), .Y(n364) );
  INVX1 U6284 ( .A(n364), .Y(n6433) );
  INVX1 U6285 ( .A(n6436), .Y(n6434) );
  INVX1 U6286 ( .A(n6434), .Y(n6435) );
  AND2X1 U6287 ( .A(n8328), .B(n361), .Y(n363) );
  INVX1 U6288 ( .A(n363), .Y(n6436) );
  INVX1 U6289 ( .A(n6439), .Y(n6437) );
  INVX1 U6290 ( .A(n6437), .Y(n6438) );
  AND2X1 U6291 ( .A(n8331), .B(n361), .Y(n362) );
  INVX1 U6292 ( .A(n362), .Y(n6439) );
  INVX1 U6293 ( .A(n6442), .Y(n6440) );
  INVX1 U6294 ( .A(n6440), .Y(n6441) );
  AND2X1 U6295 ( .A(n9864), .B(n325), .Y(n359) );
  INVX1 U6296 ( .A(n359), .Y(n6442) );
  INVX1 U6297 ( .A(n6445), .Y(n6443) );
  INVX1 U6298 ( .A(n6443), .Y(n6444) );
  AND2X1 U6299 ( .A(n9867), .B(n325), .Y(n358) );
  INVX1 U6300 ( .A(n358), .Y(n6445) );
  INVX1 U6301 ( .A(n6448), .Y(n6446) );
  INVX1 U6302 ( .A(n6446), .Y(n6447) );
  AND2X1 U6303 ( .A(n9870), .B(n325), .Y(n357) );
  INVX1 U6304 ( .A(n357), .Y(n6448) );
  INVX1 U6305 ( .A(n6451), .Y(n6449) );
  INVX1 U6306 ( .A(n6449), .Y(n6450) );
  AND2X1 U6307 ( .A(n9873), .B(n325), .Y(n356) );
  INVX1 U6308 ( .A(n356), .Y(n6451) );
  INVX1 U6309 ( .A(n6454), .Y(n6452) );
  INVX1 U6310 ( .A(n6452), .Y(n6453) );
  AND2X1 U6311 ( .A(n9876), .B(n325), .Y(n355) );
  INVX1 U6312 ( .A(n355), .Y(n6454) );
  INVX1 U6313 ( .A(n6457), .Y(n6455) );
  INVX1 U6314 ( .A(n6455), .Y(n6456) );
  AND2X1 U6315 ( .A(n9879), .B(n325), .Y(n354) );
  INVX1 U6316 ( .A(n354), .Y(n6457) );
  INVX1 U6317 ( .A(n6460), .Y(n6458) );
  INVX1 U6318 ( .A(n6458), .Y(n6459) );
  AND2X1 U6319 ( .A(n9882), .B(n325), .Y(n353) );
  INVX1 U6320 ( .A(n353), .Y(n6460) );
  INVX1 U6321 ( .A(n6463), .Y(n6461) );
  INVX1 U6322 ( .A(n6461), .Y(n6462) );
  AND2X1 U6323 ( .A(n9885), .B(n325), .Y(n352) );
  INVX1 U6324 ( .A(n352), .Y(n6463) );
  INVX1 U6325 ( .A(n6466), .Y(n6464) );
  INVX1 U6326 ( .A(n6464), .Y(n6465) );
  AND2X1 U6327 ( .A(n9888), .B(n325), .Y(n351) );
  INVX1 U6328 ( .A(n351), .Y(n6466) );
  INVX1 U6329 ( .A(n6469), .Y(n6467) );
  INVX1 U6330 ( .A(n6467), .Y(n6468) );
  AND2X1 U6331 ( .A(n9891), .B(n325), .Y(n350) );
  INVX1 U6332 ( .A(n350), .Y(n6469) );
  INVX1 U6333 ( .A(n6472), .Y(n6470) );
  INVX1 U6334 ( .A(n6470), .Y(n6471) );
  AND2X1 U6335 ( .A(n9894), .B(n325), .Y(n349) );
  INVX1 U6336 ( .A(n349), .Y(n6472) );
  INVX1 U6337 ( .A(n6475), .Y(n6473) );
  INVX1 U6338 ( .A(n6473), .Y(n6474) );
  AND2X1 U6339 ( .A(n9897), .B(n325), .Y(n348) );
  INVX1 U6340 ( .A(n348), .Y(n6475) );
  INVX1 U6341 ( .A(n6478), .Y(n6476) );
  INVX1 U6342 ( .A(n6476), .Y(n6477) );
  AND2X1 U6343 ( .A(n9900), .B(n325), .Y(n347) );
  INVX1 U6344 ( .A(n347), .Y(n6478) );
  INVX1 U6345 ( .A(n6481), .Y(n6479) );
  INVX1 U6346 ( .A(n6479), .Y(n6480) );
  AND2X1 U6347 ( .A(n9903), .B(n325), .Y(n346) );
  INVX1 U6348 ( .A(n346), .Y(n6481) );
  INVX1 U6349 ( .A(n6484), .Y(n6482) );
  INVX1 U6350 ( .A(n6482), .Y(n6483) );
  AND2X1 U6351 ( .A(n9906), .B(n325), .Y(n345) );
  INVX1 U6352 ( .A(n345), .Y(n6484) );
  INVX1 U6353 ( .A(n6487), .Y(n6485) );
  INVX1 U6354 ( .A(n6485), .Y(n6486) );
  AND2X1 U6355 ( .A(n9909), .B(n325), .Y(n344) );
  INVX1 U6356 ( .A(n344), .Y(n6487) );
  INVX1 U6357 ( .A(n6490), .Y(n6488) );
  INVX1 U6358 ( .A(n6488), .Y(n6489) );
  AND2X1 U6359 ( .A(n9912), .B(n325), .Y(n343) );
  INVX1 U6360 ( .A(n343), .Y(n6490) );
  INVX1 U6361 ( .A(n6493), .Y(n6491) );
  INVX1 U6362 ( .A(n6491), .Y(n6492) );
  AND2X1 U6363 ( .A(n9915), .B(n325), .Y(n342) );
  INVX1 U6364 ( .A(n342), .Y(n6493) );
  INVX1 U6365 ( .A(n6496), .Y(n6494) );
  INVX1 U6366 ( .A(n6494), .Y(n6495) );
  AND2X1 U6367 ( .A(n9918), .B(n325), .Y(n341) );
  INVX1 U6368 ( .A(n341), .Y(n6496) );
  INVX1 U6369 ( .A(n6499), .Y(n6497) );
  INVX1 U6370 ( .A(n6497), .Y(n6498) );
  AND2X1 U6371 ( .A(n9921), .B(n325), .Y(n340) );
  INVX1 U6372 ( .A(n340), .Y(n6499) );
  INVX1 U6373 ( .A(n6502), .Y(n6500) );
  INVX1 U6374 ( .A(n6500), .Y(n6501) );
  AND2X1 U6375 ( .A(n9924), .B(n325), .Y(n339) );
  INVX1 U6376 ( .A(n339), .Y(n6502) );
  INVX1 U6377 ( .A(n6505), .Y(n6503) );
  INVX1 U6378 ( .A(n6503), .Y(n6504) );
  AND2X1 U6379 ( .A(n9927), .B(n325), .Y(n338) );
  INVX1 U6380 ( .A(n338), .Y(n6505) );
  INVX1 U6381 ( .A(n6508), .Y(n6506) );
  INVX1 U6382 ( .A(n6506), .Y(n6507) );
  AND2X1 U6383 ( .A(n9930), .B(n325), .Y(n337) );
  INVX1 U6384 ( .A(n337), .Y(n6508) );
  INVX1 U6385 ( .A(n6511), .Y(n6509) );
  INVX1 U6386 ( .A(n6509), .Y(n6510) );
  AND2X1 U6387 ( .A(n9933), .B(n325), .Y(n336) );
  INVX1 U6388 ( .A(n336), .Y(n6511) );
  INVX1 U6389 ( .A(n6514), .Y(n6512) );
  INVX1 U6390 ( .A(n6512), .Y(n6513) );
  AND2X1 U6391 ( .A(n9936), .B(n325), .Y(n335) );
  INVX1 U6392 ( .A(n335), .Y(n6514) );
  INVX1 U6393 ( .A(n6517), .Y(n6515) );
  INVX1 U6394 ( .A(n6515), .Y(n6516) );
  AND2X1 U6395 ( .A(n9939), .B(n325), .Y(n334) );
  INVX1 U6396 ( .A(n334), .Y(n6517) );
  INVX1 U6397 ( .A(n6520), .Y(n6518) );
  INVX1 U6398 ( .A(n6518), .Y(n6519) );
  AND2X1 U6399 ( .A(n9942), .B(n325), .Y(n333) );
  INVX1 U6400 ( .A(n333), .Y(n6520) );
  INVX1 U6401 ( .A(n6523), .Y(n6521) );
  INVX1 U6402 ( .A(n6521), .Y(n6522) );
  AND2X1 U6403 ( .A(n9945), .B(n325), .Y(n332) );
  INVX1 U6404 ( .A(n332), .Y(n6523) );
  INVX1 U6405 ( .A(n6526), .Y(n6524) );
  INVX1 U6406 ( .A(n6524), .Y(n6525) );
  AND2X1 U6407 ( .A(n9948), .B(n325), .Y(n331) );
  INVX1 U6408 ( .A(n331), .Y(n6526) );
  INVX1 U6409 ( .A(n6529), .Y(n6527) );
  INVX1 U6410 ( .A(n6527), .Y(n6528) );
  AND2X1 U6411 ( .A(n9951), .B(n325), .Y(n330) );
  INVX1 U6412 ( .A(n330), .Y(n6529) );
  INVX1 U6413 ( .A(n6532), .Y(n6530) );
  INVX1 U6414 ( .A(n6530), .Y(n6531) );
  AND2X1 U6415 ( .A(n9954), .B(n325), .Y(n329) );
  INVX1 U6416 ( .A(n329), .Y(n6532) );
  INVX1 U6417 ( .A(n6535), .Y(n6533) );
  INVX1 U6418 ( .A(n6533), .Y(n6534) );
  AND2X1 U6419 ( .A(n9957), .B(n325), .Y(n328) );
  INVX1 U6420 ( .A(n328), .Y(n6535) );
  INVX1 U6421 ( .A(n6538), .Y(n6536) );
  INVX1 U6422 ( .A(n6536), .Y(n6537) );
  AND2X1 U6423 ( .A(n9960), .B(n325), .Y(n327) );
  INVX1 U6424 ( .A(n327), .Y(n6538) );
  INVX1 U6425 ( .A(n6541), .Y(n6539) );
  INVX1 U6426 ( .A(n6539), .Y(n6540) );
  AND2X1 U6427 ( .A(n9963), .B(n325), .Y(n326) );
  INVX1 U6428 ( .A(n326), .Y(n6541) );
  INVX1 U6429 ( .A(n6544), .Y(n6542) );
  INVX1 U6430 ( .A(n6542), .Y(n6543) );
  AND2X1 U6431 ( .A(n7110), .B(n10113), .Y(n322) );
  INVX1 U6432 ( .A(n322), .Y(n6544) );
  INVX1 U6433 ( .A(n6547), .Y(n6545) );
  INVX1 U6434 ( .A(n6545), .Y(n6546) );
  AND2X1 U6435 ( .A(n7113), .B(n10113), .Y(n320) );
  INVX1 U6436 ( .A(n320), .Y(n6547) );
  INVX1 U6437 ( .A(n6550), .Y(n6548) );
  INVX1 U6438 ( .A(n6548), .Y(n6549) );
  AND2X1 U6439 ( .A(n7116), .B(n10113), .Y(n318) );
  INVX1 U6440 ( .A(n318), .Y(n6550) );
  INVX1 U6441 ( .A(n6553), .Y(n6551) );
  INVX1 U6442 ( .A(n6551), .Y(n6552) );
  AND2X1 U6443 ( .A(n7119), .B(n10113), .Y(n316) );
  INVX1 U6444 ( .A(n316), .Y(n6553) );
  INVX1 U6445 ( .A(n6556), .Y(n6554) );
  INVX1 U6446 ( .A(n6554), .Y(n6555) );
  AND2X1 U6447 ( .A(n7122), .B(n10113), .Y(n314) );
  INVX1 U6448 ( .A(n314), .Y(n6556) );
  INVX1 U6449 ( .A(n6559), .Y(n6557) );
  INVX1 U6450 ( .A(n6557), .Y(n6558) );
  AND2X1 U6451 ( .A(n7125), .B(n10113), .Y(n312) );
  INVX1 U6452 ( .A(n312), .Y(n6559) );
  INVX1 U6453 ( .A(n6562), .Y(n6560) );
  INVX1 U6454 ( .A(n6560), .Y(n6561) );
  AND2X1 U6455 ( .A(n7128), .B(n10113), .Y(n310) );
  INVX1 U6456 ( .A(n310), .Y(n6562) );
  INVX1 U6457 ( .A(n6565), .Y(n6563) );
  INVX1 U6458 ( .A(n6563), .Y(n6564) );
  AND2X1 U6459 ( .A(n7131), .B(n10113), .Y(n308) );
  INVX1 U6460 ( .A(n308), .Y(n6565) );
  INVX1 U6461 ( .A(n6568), .Y(n6566) );
  INVX1 U6462 ( .A(n6566), .Y(n6567) );
  AND2X1 U6463 ( .A(n7134), .B(n10113), .Y(n306) );
  INVX1 U6464 ( .A(n306), .Y(n6568) );
  INVX1 U6465 ( .A(n6571), .Y(n6569) );
  INVX1 U6466 ( .A(n6569), .Y(n6570) );
  AND2X1 U6467 ( .A(n7137), .B(n10113), .Y(n304) );
  INVX1 U6468 ( .A(n304), .Y(n6571) );
  INVX1 U6469 ( .A(n6574), .Y(n6572) );
  INVX1 U6470 ( .A(n6572), .Y(n6573) );
  AND2X1 U6471 ( .A(n7140), .B(n10113), .Y(n302) );
  INVX1 U6472 ( .A(n302), .Y(n6574) );
  INVX1 U6473 ( .A(n6577), .Y(n6575) );
  INVX1 U6474 ( .A(n6575), .Y(n6576) );
  AND2X1 U6475 ( .A(n7143), .B(n10113), .Y(n300) );
  INVX1 U6476 ( .A(n300), .Y(n6577) );
  INVX1 U6477 ( .A(n6580), .Y(n6578) );
  INVX1 U6478 ( .A(n6578), .Y(n6579) );
  AND2X1 U6479 ( .A(n7146), .B(n10113), .Y(n298) );
  INVX1 U6480 ( .A(n298), .Y(n6580) );
  INVX1 U6481 ( .A(n6583), .Y(n6581) );
  INVX1 U6482 ( .A(n6581), .Y(n6582) );
  AND2X1 U6483 ( .A(n7149), .B(n10113), .Y(n296) );
  INVX1 U6484 ( .A(n296), .Y(n6583) );
  INVX1 U6485 ( .A(n6586), .Y(n6584) );
  INVX1 U6486 ( .A(n6584), .Y(n6585) );
  AND2X1 U6487 ( .A(n7152), .B(n10113), .Y(n294) );
  INVX1 U6488 ( .A(n294), .Y(n6586) );
  INVX1 U6489 ( .A(n6589), .Y(n6587) );
  INVX1 U6490 ( .A(n6587), .Y(n6588) );
  AND2X1 U6491 ( .A(n7155), .B(n10113), .Y(n292) );
  INVX1 U6492 ( .A(n292), .Y(n6589) );
  INVX1 U6493 ( .A(n6592), .Y(n6590) );
  INVX1 U6494 ( .A(n6590), .Y(n6591) );
  AND2X1 U6495 ( .A(n7158), .B(n10113), .Y(n290) );
  INVX1 U6496 ( .A(n290), .Y(n6592) );
  INVX1 U6497 ( .A(n6595), .Y(n6593) );
  INVX1 U6498 ( .A(n6593), .Y(n6594) );
  AND2X1 U6499 ( .A(n7161), .B(n10113), .Y(n288) );
  INVX1 U6500 ( .A(n288), .Y(n6595) );
  INVX1 U6501 ( .A(n6598), .Y(n6596) );
  INVX1 U6502 ( .A(n6596), .Y(n6597) );
  AND2X1 U6503 ( .A(n7164), .B(n10113), .Y(n286) );
  INVX1 U6504 ( .A(n286), .Y(n6598) );
  INVX1 U6505 ( .A(n6601), .Y(n6599) );
  INVX1 U6506 ( .A(n6599), .Y(n6600) );
  AND2X1 U6507 ( .A(n7167), .B(n10113), .Y(n284) );
  INVX1 U6508 ( .A(n284), .Y(n6601) );
  INVX1 U6509 ( .A(n6604), .Y(n6602) );
  INVX1 U6510 ( .A(n6602), .Y(n6603) );
  AND2X1 U6511 ( .A(n7170), .B(n10113), .Y(n282) );
  INVX1 U6512 ( .A(n282), .Y(n6604) );
  INVX1 U6513 ( .A(n6607), .Y(n6605) );
  INVX1 U6514 ( .A(n6605), .Y(n6606) );
  AND2X1 U6515 ( .A(n7173), .B(n10113), .Y(n280) );
  INVX1 U6516 ( .A(n280), .Y(n6607) );
  INVX1 U6517 ( .A(n6610), .Y(n6608) );
  INVX1 U6518 ( .A(n6608), .Y(n6609) );
  AND2X1 U6519 ( .A(n7176), .B(n10113), .Y(n278) );
  INVX1 U6520 ( .A(n278), .Y(n6610) );
  INVX1 U6521 ( .A(n6613), .Y(n6611) );
  INVX1 U6522 ( .A(n6611), .Y(n6612) );
  AND2X1 U6523 ( .A(n7179), .B(n10113), .Y(n276) );
  INVX1 U6524 ( .A(n276), .Y(n6613) );
  INVX1 U6525 ( .A(n6616), .Y(n6614) );
  INVX1 U6526 ( .A(n6614), .Y(n6615) );
  AND2X1 U6527 ( .A(n7182), .B(n10113), .Y(n274) );
  INVX1 U6528 ( .A(n274), .Y(n6616) );
  INVX1 U6529 ( .A(n6619), .Y(n6617) );
  INVX1 U6530 ( .A(n6617), .Y(n6618) );
  AND2X1 U6531 ( .A(n7185), .B(n10113), .Y(n272) );
  INVX1 U6532 ( .A(n272), .Y(n6619) );
  INVX1 U6533 ( .A(n6622), .Y(n6620) );
  INVX1 U6534 ( .A(n6620), .Y(n6621) );
  AND2X1 U6535 ( .A(n7188), .B(n10113), .Y(n270) );
  INVX1 U6536 ( .A(n270), .Y(n6622) );
  INVX1 U6537 ( .A(n6625), .Y(n6623) );
  INVX1 U6538 ( .A(n6623), .Y(n6624) );
  AND2X1 U6539 ( .A(n7191), .B(n10113), .Y(n268) );
  INVX1 U6540 ( .A(n268), .Y(n6625) );
  INVX1 U6541 ( .A(n6628), .Y(n6626) );
  INVX1 U6542 ( .A(n6626), .Y(n6627) );
  AND2X1 U6543 ( .A(n7194), .B(n10113), .Y(n266) );
  INVX1 U6544 ( .A(n266), .Y(n6628) );
  INVX1 U6545 ( .A(n6631), .Y(n6629) );
  INVX1 U6546 ( .A(n6629), .Y(n6630) );
  AND2X1 U6547 ( .A(n7197), .B(n10113), .Y(n264) );
  INVX1 U6548 ( .A(n264), .Y(n6631) );
  INVX1 U6549 ( .A(n6634), .Y(n6632) );
  INVX1 U6550 ( .A(n6632), .Y(n6633) );
  AND2X1 U6551 ( .A(n7200), .B(n10113), .Y(n262) );
  INVX1 U6552 ( .A(n262), .Y(n6634) );
  INVX1 U6553 ( .A(n6637), .Y(n6635) );
  INVX1 U6554 ( .A(n6635), .Y(n6636) );
  AND2X1 U6555 ( .A(n7203), .B(n10113), .Y(n260) );
  INVX1 U6556 ( .A(n260), .Y(n6637) );
  INVX1 U6557 ( .A(n6640), .Y(n6638) );
  INVX1 U6558 ( .A(n6638), .Y(n6639) );
  AND2X1 U6559 ( .A(n7206), .B(n10113), .Y(n258) );
  INVX1 U6560 ( .A(n258), .Y(n6640) );
  INVX1 U6561 ( .A(n6643), .Y(n6641) );
  INVX1 U6562 ( .A(n6641), .Y(n6642) );
  AND2X1 U6563 ( .A(n7209), .B(n10113), .Y(n256) );
  INVX1 U6564 ( .A(n256), .Y(n6643) );
  INVX1 U6565 ( .A(n6646), .Y(n6644) );
  INVX1 U6566 ( .A(n6644), .Y(n6645) );
  AND2X1 U6567 ( .A(n10723), .B(n193), .Y(n253) );
  INVX1 U6568 ( .A(n253), .Y(n6646) );
  INVX1 U6569 ( .A(n6649), .Y(n6647) );
  INVX1 U6570 ( .A(n6647), .Y(n6648) );
  AND2X1 U6571 ( .A(n110), .B(n193), .Y(n251) );
  INVX1 U6572 ( .A(n251), .Y(n6649) );
  INVX1 U6573 ( .A(n6652), .Y(n6650) );
  INVX1 U6574 ( .A(n6650), .Y(n6651) );
  AND2X1 U6575 ( .A(n38), .B(n237), .Y(n249) );
  INVX1 U6576 ( .A(n249), .Y(n6652) );
  INVX1 U6577 ( .A(n6655), .Y(n6653) );
  INVX1 U6578 ( .A(n6653), .Y(n6654) );
  AND2X2 U6579 ( .A(n33), .B(n237), .Y(n247) );
  INVX1 U6580 ( .A(n247), .Y(n6655) );
  INVX1 U6581 ( .A(n6658), .Y(n6656) );
  INVX1 U6582 ( .A(n6656), .Y(n6657) );
  AND2X1 U6583 ( .A(n34), .B(n237), .Y(n245) );
  INVX1 U6584 ( .A(n245), .Y(n6658) );
  INVX1 U6585 ( .A(n6661), .Y(n6659) );
  INVX1 U6586 ( .A(n6659), .Y(n6660) );
  AND2X1 U6587 ( .A(n35), .B(n237), .Y(n243) );
  INVX1 U6588 ( .A(n243), .Y(n6661) );
  INVX1 U6589 ( .A(n6664), .Y(n6662) );
  INVX1 U6590 ( .A(n6662), .Y(n6663) );
  AND2X1 U6591 ( .A(n36), .B(n237), .Y(n241) );
  INVX1 U6592 ( .A(n241), .Y(n6664) );
  INVX1 U6593 ( .A(n6667), .Y(n6665) );
  INVX1 U6594 ( .A(n6665), .Y(n6666) );
  AND2X1 U6595 ( .A(n37), .B(n237), .Y(n239) );
  INVX1 U6596 ( .A(n239), .Y(n6667) );
  INVX1 U6597 ( .A(n6670), .Y(n6668) );
  INVX1 U6598 ( .A(n6668), .Y(n6669) );
  AND2X1 U6599 ( .A(n106), .B(n193), .Y(n201) );
  INVX1 U6600 ( .A(n201), .Y(n6670) );
  INVX1 U6601 ( .A(n6673), .Y(n6671) );
  INVX1 U6602 ( .A(n6671), .Y(n6672) );
  AND2X1 U6603 ( .A(n107), .B(n193), .Y(n199) );
  INVX1 U6604 ( .A(n199), .Y(n6673) );
  INVX1 U6605 ( .A(n6676), .Y(n6674) );
  INVX1 U6606 ( .A(n6674), .Y(n6675) );
  AND2X1 U6607 ( .A(n108), .B(n193), .Y(n197) );
  INVX1 U6608 ( .A(n197), .Y(n6676) );
  INVX1 U6609 ( .A(n6679), .Y(n6677) );
  INVX1 U6610 ( .A(n6677), .Y(n6678) );
  AND2X1 U6611 ( .A(n109), .B(n193), .Y(n195) );
  INVX1 U6612 ( .A(n195), .Y(n6679) );
  INVX1 U6613 ( .A(n6682), .Y(n6680) );
  INVX1 U6614 ( .A(n6680), .Y(n6681) );
  OR2X2 U6615 ( .A(fillcount[1]), .B(fillcount[0]), .Y(n1426) );
  INVX1 U6616 ( .A(n1426), .Y(n6682) );
  INVX1 U6617 ( .A(n10683), .Y(n10687) );
  INVX4 U6618 ( .A(n10688), .Y(n10686) );
  INVX1 U6619 ( .A(n11), .Y(n10688) );
  AND2X1 U6620 ( .A(n576), .B(n324), .Y(n10487) );
  AND2X1 U6621 ( .A(n540), .B(n324), .Y(n10486) );
  AND2X1 U6622 ( .A(n360), .B(n324), .Y(n10488) );
  AND2X1 U6623 ( .A(n10031), .B(n324), .Y(n10489) );
  AND2X1 U6624 ( .A(n10022), .B(n324), .Y(n10490) );
  INVX1 U6625 ( .A(n577), .Y(n324) );
  INVX1 U6626 ( .A(n6685), .Y(n6683) );
  INVX1 U6627 ( .A(n6683), .Y(n6684) );
  BUFX2 U6628 ( .A(n1438), .Y(n6685) );
  INVX1 U6629 ( .A(n6688), .Y(n6686) );
  INVX1 U6630 ( .A(n6686), .Y(n6687) );
  AND2X1 U6631 ( .A(n10104), .B(r301_B_not_4_), .Y(n10523) );
  INVX1 U6632 ( .A(n10523), .Y(n6688) );
  INVX1 U6633 ( .A(n6691), .Y(n6689) );
  INVX1 U6634 ( .A(n6689), .Y(n6690) );
  OR2X2 U6635 ( .A(n10530), .B(n10535), .Y(n1430) );
  INVX1 U6636 ( .A(n1430), .Y(n6691) );
  INVX1 U6637 ( .A(n6694), .Y(n6692) );
  INVX1 U6638 ( .A(n6692), .Y(n6693) );
  BUFX2 U6639 ( .A(rd_ptr_gray_ss[0]), .Y(n6694) );
  INVX1 U6640 ( .A(n6697), .Y(n6695) );
  INVX1 U6641 ( .A(n6695), .Y(n6696) );
  BUFX2 U6642 ( .A(wr_ptr_gray_ss[2]), .Y(n6697) );
  INVX1 U6643 ( .A(n6700), .Y(n6698) );
  INVX1 U6644 ( .A(n6698), .Y(n6699) );
  BUFX2 U6645 ( .A(wr_ptr_gray_ss[3]), .Y(n6700) );
  INVX1 U6646 ( .A(n6703), .Y(n6701) );
  INVX1 U6647 ( .A(n6701), .Y(n6702) );
  BUFX2 U6648 ( .A(fifo[374]), .Y(n6703) );
  INVX1 U6649 ( .A(n6706), .Y(n6704) );
  INVX1 U6650 ( .A(n6704), .Y(n6705) );
  BUFX2 U6651 ( .A(fifo[375]), .Y(n6706) );
  INVX1 U6652 ( .A(n6709), .Y(n6707) );
  INVX1 U6653 ( .A(n6707), .Y(n6708) );
  BUFX2 U6654 ( .A(fifo[376]), .Y(n6709) );
  INVX1 U6655 ( .A(n6712), .Y(n6710) );
  INVX1 U6656 ( .A(n6710), .Y(n6711) );
  BUFX2 U6657 ( .A(fifo[377]), .Y(n6712) );
  INVX1 U6658 ( .A(n6715), .Y(n6713) );
  INVX1 U6659 ( .A(n6713), .Y(n6714) );
  BUFX2 U6660 ( .A(fifo[378]), .Y(n6715) );
  INVX1 U6661 ( .A(n6718), .Y(n6716) );
  INVX1 U6662 ( .A(n6716), .Y(n6717) );
  BUFX2 U6663 ( .A(fifo[379]), .Y(n6718) );
  INVX1 U6664 ( .A(n6721), .Y(n6719) );
  INVX1 U6665 ( .A(n6719), .Y(n6720) );
  BUFX2 U6666 ( .A(fifo[380]), .Y(n6721) );
  INVX1 U6667 ( .A(n6724), .Y(n6722) );
  INVX1 U6668 ( .A(n6722), .Y(n6723) );
  BUFX2 U6669 ( .A(fifo[381]), .Y(n6724) );
  INVX1 U6670 ( .A(n6727), .Y(n6725) );
  INVX1 U6671 ( .A(n6725), .Y(n6726) );
  BUFX2 U6672 ( .A(fifo[382]), .Y(n6727) );
  INVX1 U6673 ( .A(n6730), .Y(n6728) );
  INVX1 U6674 ( .A(n6728), .Y(n6729) );
  BUFX2 U6675 ( .A(fifo[383]), .Y(n6730) );
  INVX1 U6676 ( .A(n6733), .Y(n6731) );
  INVX1 U6677 ( .A(n6731), .Y(n6732) );
  BUFX2 U6678 ( .A(fifo[384]), .Y(n6733) );
  INVX1 U6679 ( .A(n6736), .Y(n6734) );
  INVX1 U6680 ( .A(n6734), .Y(n6735) );
  BUFX2 U6681 ( .A(fifo[385]), .Y(n6736) );
  INVX1 U6682 ( .A(n6739), .Y(n6737) );
  INVX1 U6683 ( .A(n6737), .Y(n6738) );
  BUFX2 U6684 ( .A(fifo[386]), .Y(n6739) );
  INVX1 U6685 ( .A(n6742), .Y(n6740) );
  INVX1 U6686 ( .A(n6740), .Y(n6741) );
  BUFX2 U6687 ( .A(fifo[387]), .Y(n6742) );
  INVX1 U6688 ( .A(n6745), .Y(n6743) );
  INVX1 U6689 ( .A(n6743), .Y(n6744) );
  BUFX2 U6690 ( .A(fifo[388]), .Y(n6745) );
  INVX1 U6691 ( .A(n6748), .Y(n6746) );
  INVX1 U6692 ( .A(n6746), .Y(n6747) );
  BUFX2 U6693 ( .A(fifo[389]), .Y(n6748) );
  INVX1 U6694 ( .A(n6751), .Y(n6749) );
  INVX1 U6695 ( .A(n6749), .Y(n6750) );
  BUFX2 U6696 ( .A(fifo[390]), .Y(n6751) );
  INVX1 U6697 ( .A(n6754), .Y(n6752) );
  INVX1 U6698 ( .A(n6752), .Y(n6753) );
  BUFX2 U6699 ( .A(fifo[391]), .Y(n6754) );
  INVX1 U6700 ( .A(n6757), .Y(n6755) );
  INVX1 U6701 ( .A(n6755), .Y(n6756) );
  BUFX2 U6702 ( .A(fifo[392]), .Y(n6757) );
  INVX1 U6703 ( .A(n6760), .Y(n6758) );
  INVX1 U6704 ( .A(n6758), .Y(n6759) );
  BUFX2 U6705 ( .A(fifo[393]), .Y(n6760) );
  INVX1 U6706 ( .A(n6763), .Y(n6761) );
  INVX1 U6707 ( .A(n6761), .Y(n6762) );
  BUFX2 U6708 ( .A(fifo[394]), .Y(n6763) );
  INVX1 U6709 ( .A(n6766), .Y(n6764) );
  INVX1 U6710 ( .A(n6764), .Y(n6765) );
  BUFX2 U6711 ( .A(fifo[395]), .Y(n6766) );
  INVX1 U6712 ( .A(n6769), .Y(n6767) );
  INVX1 U6713 ( .A(n6767), .Y(n6768) );
  BUFX2 U6714 ( .A(fifo[396]), .Y(n6769) );
  INVX1 U6715 ( .A(n6772), .Y(n6770) );
  INVX1 U6716 ( .A(n6770), .Y(n6771) );
  BUFX2 U6717 ( .A(fifo[397]), .Y(n6772) );
  INVX1 U6718 ( .A(n6775), .Y(n6773) );
  INVX1 U6719 ( .A(n6773), .Y(n6774) );
  BUFX2 U6720 ( .A(fifo[398]), .Y(n6775) );
  INVX1 U6721 ( .A(n6778), .Y(n6776) );
  INVX1 U6722 ( .A(n6776), .Y(n6777) );
  BUFX2 U6723 ( .A(fifo[399]), .Y(n6778) );
  INVX1 U6724 ( .A(n6781), .Y(n6779) );
  INVX1 U6725 ( .A(n6779), .Y(n6780) );
  BUFX2 U6726 ( .A(fifo[400]), .Y(n6781) );
  INVX1 U6727 ( .A(n6784), .Y(n6782) );
  INVX1 U6728 ( .A(n6782), .Y(n6783) );
  BUFX2 U6729 ( .A(fifo[401]), .Y(n6784) );
  INVX1 U6730 ( .A(n6787), .Y(n6785) );
  INVX1 U6731 ( .A(n6785), .Y(n6786) );
  BUFX2 U6732 ( .A(fifo[402]), .Y(n6787) );
  INVX1 U6733 ( .A(n6790), .Y(n6788) );
  INVX1 U6734 ( .A(n6788), .Y(n6789) );
  BUFX2 U6735 ( .A(fifo[403]), .Y(n6790) );
  INVX1 U6736 ( .A(n6793), .Y(n6791) );
  INVX1 U6737 ( .A(n6791), .Y(n6792) );
  BUFX2 U6738 ( .A(fifo[404]), .Y(n6793) );
  INVX1 U6739 ( .A(n6796), .Y(n6794) );
  INVX1 U6740 ( .A(n6794), .Y(n6795) );
  BUFX2 U6741 ( .A(fifo[405]), .Y(n6796) );
  INVX1 U6742 ( .A(n6799), .Y(n6797) );
  INVX1 U6743 ( .A(n6797), .Y(n6798) );
  BUFX2 U6744 ( .A(fifo[406]), .Y(n6799) );
  INVX1 U6745 ( .A(n6802), .Y(n6800) );
  INVX1 U6746 ( .A(n6800), .Y(n6801) );
  BUFX2 U6747 ( .A(fifo[407]), .Y(n6802) );
  INVX1 U6748 ( .A(n6805), .Y(n6803) );
  INVX1 U6749 ( .A(n6803), .Y(n6804) );
  BUFX2 U6750 ( .A(fifo[442]), .Y(n6805) );
  INVX1 U6751 ( .A(n6808), .Y(n6806) );
  INVX1 U6752 ( .A(n6806), .Y(n6807) );
  BUFX2 U6753 ( .A(fifo[443]), .Y(n6808) );
  INVX1 U6754 ( .A(n6811), .Y(n6809) );
  INVX1 U6755 ( .A(n6809), .Y(n6810) );
  BUFX2 U6756 ( .A(fifo[444]), .Y(n6811) );
  INVX1 U6757 ( .A(n6814), .Y(n6812) );
  INVX1 U6758 ( .A(n6812), .Y(n6813) );
  BUFX2 U6759 ( .A(fifo[445]), .Y(n6814) );
  INVX1 U6760 ( .A(n6817), .Y(n6815) );
  INVX1 U6761 ( .A(n6815), .Y(n6816) );
  BUFX2 U6762 ( .A(fifo[446]), .Y(n6817) );
  INVX1 U6763 ( .A(n6820), .Y(n6818) );
  INVX1 U6764 ( .A(n6818), .Y(n6819) );
  BUFX2 U6765 ( .A(fifo[447]), .Y(n6820) );
  INVX1 U6766 ( .A(n6823), .Y(n6821) );
  INVX1 U6767 ( .A(n6821), .Y(n6822) );
  BUFX2 U6768 ( .A(fifo[448]), .Y(n6823) );
  INVX1 U6769 ( .A(n6826), .Y(n6824) );
  INVX1 U6770 ( .A(n6824), .Y(n6825) );
  BUFX2 U6771 ( .A(fifo[449]), .Y(n6826) );
  INVX1 U6772 ( .A(n6829), .Y(n6827) );
  INVX1 U6773 ( .A(n6827), .Y(n6828) );
  BUFX2 U6774 ( .A(fifo[450]), .Y(n6829) );
  INVX1 U6775 ( .A(n6832), .Y(n6830) );
  INVX1 U6776 ( .A(n6830), .Y(n6831) );
  BUFX2 U6777 ( .A(fifo[451]), .Y(n6832) );
  INVX1 U6778 ( .A(n6835), .Y(n6833) );
  INVX1 U6779 ( .A(n6833), .Y(n6834) );
  BUFX2 U6780 ( .A(fifo[452]), .Y(n6835) );
  INVX1 U6781 ( .A(n6838), .Y(n6836) );
  INVX1 U6782 ( .A(n6836), .Y(n6837) );
  BUFX2 U6783 ( .A(fifo[453]), .Y(n6838) );
  INVX1 U6784 ( .A(n6841), .Y(n6839) );
  INVX1 U6785 ( .A(n6839), .Y(n6840) );
  BUFX2 U6786 ( .A(fifo[454]), .Y(n6841) );
  INVX1 U6787 ( .A(n6844), .Y(n6842) );
  INVX1 U6788 ( .A(n6842), .Y(n6843) );
  BUFX2 U6789 ( .A(fifo[455]), .Y(n6844) );
  INVX1 U6790 ( .A(n6847), .Y(n6845) );
  INVX1 U6791 ( .A(n6845), .Y(n6846) );
  BUFX2 U6792 ( .A(fifo[456]), .Y(n6847) );
  INVX1 U6793 ( .A(n6850), .Y(n6848) );
  INVX1 U6794 ( .A(n6848), .Y(n6849) );
  BUFX2 U6795 ( .A(fifo[457]), .Y(n6850) );
  INVX1 U6796 ( .A(n6853), .Y(n6851) );
  INVX1 U6797 ( .A(n6851), .Y(n6852) );
  BUFX2 U6798 ( .A(fifo[458]), .Y(n6853) );
  INVX1 U6799 ( .A(n6856), .Y(n6854) );
  INVX1 U6800 ( .A(n6854), .Y(n6855) );
  BUFX2 U6801 ( .A(fifo[459]), .Y(n6856) );
  INVX1 U6802 ( .A(n6859), .Y(n6857) );
  INVX1 U6803 ( .A(n6857), .Y(n6858) );
  BUFX2 U6804 ( .A(fifo[460]), .Y(n6859) );
  INVX1 U6805 ( .A(n6862), .Y(n6860) );
  INVX1 U6806 ( .A(n6860), .Y(n6861) );
  BUFX2 U6807 ( .A(fifo[461]), .Y(n6862) );
  INVX1 U6808 ( .A(n6865), .Y(n6863) );
  INVX1 U6809 ( .A(n6863), .Y(n6864) );
  BUFX2 U6810 ( .A(fifo[462]), .Y(n6865) );
  INVX1 U6811 ( .A(n6868), .Y(n6866) );
  INVX1 U6812 ( .A(n6866), .Y(n6867) );
  BUFX2 U6813 ( .A(fifo[463]), .Y(n6868) );
  INVX1 U6814 ( .A(n6871), .Y(n6869) );
  INVX1 U6815 ( .A(n6869), .Y(n6870) );
  BUFX2 U6816 ( .A(fifo[464]), .Y(n6871) );
  INVX1 U6817 ( .A(n6874), .Y(n6872) );
  INVX1 U6818 ( .A(n6872), .Y(n6873) );
  BUFX2 U6819 ( .A(fifo[465]), .Y(n6874) );
  INVX1 U6820 ( .A(n6877), .Y(n6875) );
  INVX1 U6821 ( .A(n6875), .Y(n6876) );
  BUFX2 U6822 ( .A(fifo[466]), .Y(n6877) );
  INVX1 U6823 ( .A(n6880), .Y(n6878) );
  INVX1 U6824 ( .A(n6878), .Y(n6879) );
  BUFX2 U6825 ( .A(fifo[467]), .Y(n6880) );
  INVX1 U6826 ( .A(n6883), .Y(n6881) );
  INVX1 U6827 ( .A(n6881), .Y(n6882) );
  BUFX2 U6828 ( .A(fifo[468]), .Y(n6883) );
  INVX1 U6829 ( .A(n6886), .Y(n6884) );
  INVX1 U6830 ( .A(n6884), .Y(n6885) );
  BUFX2 U6831 ( .A(fifo[469]), .Y(n6886) );
  INVX1 U6832 ( .A(n6889), .Y(n6887) );
  INVX1 U6833 ( .A(n6887), .Y(n6888) );
  BUFX2 U6834 ( .A(fifo[470]), .Y(n6889) );
  INVX1 U6835 ( .A(n6892), .Y(n6890) );
  INVX1 U6836 ( .A(n6890), .Y(n6891) );
  BUFX2 U6837 ( .A(fifo[471]), .Y(n6892) );
  INVX1 U6838 ( .A(n6895), .Y(n6893) );
  INVX1 U6839 ( .A(n6893), .Y(n6894) );
  BUFX2 U6840 ( .A(fifo[472]), .Y(n6895) );
  INVX1 U6841 ( .A(n6898), .Y(n6896) );
  INVX1 U6842 ( .A(n6896), .Y(n6897) );
  BUFX2 U6843 ( .A(fifo[473]), .Y(n6898) );
  INVX1 U6844 ( .A(n6901), .Y(n6899) );
  INVX1 U6845 ( .A(n6899), .Y(n6900) );
  BUFX2 U6846 ( .A(fifo[474]), .Y(n6901) );
  INVX1 U6847 ( .A(n6904), .Y(n6902) );
  INVX1 U6848 ( .A(n6902), .Y(n6903) );
  BUFX2 U6849 ( .A(fifo[475]), .Y(n6904) );
  INVX1 U6850 ( .A(n6907), .Y(n6905) );
  INVX1 U6851 ( .A(n6905), .Y(n6906) );
  BUFX2 U6852 ( .A(fifo[306]), .Y(n6907) );
  INVX1 U6853 ( .A(n6910), .Y(n6908) );
  INVX1 U6854 ( .A(n6908), .Y(n6909) );
  BUFX2 U6855 ( .A(fifo[307]), .Y(n6910) );
  INVX1 U6856 ( .A(n6913), .Y(n6911) );
  INVX1 U6857 ( .A(n6911), .Y(n6912) );
  BUFX2 U6858 ( .A(fifo[308]), .Y(n6913) );
  INVX1 U6859 ( .A(n6916), .Y(n6914) );
  INVX1 U6860 ( .A(n6914), .Y(n6915) );
  BUFX2 U6861 ( .A(fifo[309]), .Y(n6916) );
  INVX1 U6862 ( .A(n6919), .Y(n6917) );
  INVX1 U6863 ( .A(n6917), .Y(n6918) );
  BUFX2 U6864 ( .A(fifo[310]), .Y(n6919) );
  INVX1 U6865 ( .A(n6922), .Y(n6920) );
  INVX1 U6866 ( .A(n6920), .Y(n6921) );
  BUFX2 U6867 ( .A(fifo[311]), .Y(n6922) );
  INVX1 U6868 ( .A(n6925), .Y(n6923) );
  INVX1 U6869 ( .A(n6923), .Y(n6924) );
  BUFX2 U6870 ( .A(fifo[312]), .Y(n6925) );
  INVX1 U6871 ( .A(n6928), .Y(n6926) );
  INVX1 U6872 ( .A(n6926), .Y(n6927) );
  BUFX2 U6873 ( .A(fifo[313]), .Y(n6928) );
  INVX1 U6874 ( .A(n6931), .Y(n6929) );
  INVX1 U6875 ( .A(n6929), .Y(n6930) );
  BUFX2 U6876 ( .A(fifo[314]), .Y(n6931) );
  INVX1 U6877 ( .A(n6934), .Y(n6932) );
  INVX1 U6878 ( .A(n6932), .Y(n6933) );
  BUFX2 U6879 ( .A(fifo[315]), .Y(n6934) );
  INVX1 U6880 ( .A(n6937), .Y(n6935) );
  INVX1 U6881 ( .A(n6935), .Y(n6936) );
  BUFX2 U6882 ( .A(fifo[316]), .Y(n6937) );
  INVX1 U6883 ( .A(n6940), .Y(n6938) );
  INVX1 U6884 ( .A(n6938), .Y(n6939) );
  BUFX2 U6885 ( .A(fifo[317]), .Y(n6940) );
  INVX1 U6886 ( .A(n6943), .Y(n6941) );
  INVX1 U6887 ( .A(n6941), .Y(n6942) );
  BUFX2 U6888 ( .A(fifo[318]), .Y(n6943) );
  INVX1 U6889 ( .A(n6946), .Y(n6944) );
  INVX1 U6890 ( .A(n6944), .Y(n6945) );
  BUFX2 U6891 ( .A(fifo[319]), .Y(n6946) );
  INVX1 U6892 ( .A(n6949), .Y(n6947) );
  INVX1 U6893 ( .A(n6947), .Y(n6948) );
  BUFX2 U6894 ( .A(fifo[320]), .Y(n6949) );
  INVX1 U6895 ( .A(n6952), .Y(n6950) );
  INVX1 U6896 ( .A(n6950), .Y(n6951) );
  BUFX2 U6897 ( .A(fifo[321]), .Y(n6952) );
  INVX1 U6898 ( .A(n6955), .Y(n6953) );
  INVX1 U6899 ( .A(n6953), .Y(n6954) );
  BUFX2 U6900 ( .A(fifo[322]), .Y(n6955) );
  INVX1 U6901 ( .A(n6958), .Y(n6956) );
  INVX1 U6902 ( .A(n6956), .Y(n6957) );
  BUFX2 U6903 ( .A(fifo[323]), .Y(n6958) );
  INVX1 U6904 ( .A(n6961), .Y(n6959) );
  INVX1 U6905 ( .A(n6959), .Y(n6960) );
  BUFX2 U6906 ( .A(fifo[324]), .Y(n6961) );
  INVX1 U6907 ( .A(n6964), .Y(n6962) );
  INVX1 U6908 ( .A(n6962), .Y(n6963) );
  BUFX2 U6909 ( .A(fifo[325]), .Y(n6964) );
  INVX1 U6910 ( .A(n6967), .Y(n6965) );
  INVX1 U6911 ( .A(n6965), .Y(n6966) );
  BUFX2 U6912 ( .A(fifo[326]), .Y(n6967) );
  INVX1 U6913 ( .A(n6970), .Y(n6968) );
  INVX1 U6914 ( .A(n6968), .Y(n6969) );
  BUFX2 U6915 ( .A(fifo[327]), .Y(n6970) );
  INVX1 U6916 ( .A(n6973), .Y(n6971) );
  INVX1 U6917 ( .A(n6971), .Y(n6972) );
  BUFX2 U6918 ( .A(fifo[328]), .Y(n6973) );
  INVX1 U6919 ( .A(n6976), .Y(n6974) );
  INVX1 U6920 ( .A(n6974), .Y(n6975) );
  BUFX2 U6921 ( .A(fifo[329]), .Y(n6976) );
  INVX1 U6922 ( .A(n6979), .Y(n6977) );
  INVX1 U6923 ( .A(n6977), .Y(n6978) );
  BUFX2 U6924 ( .A(fifo[330]), .Y(n6979) );
  INVX1 U6925 ( .A(n6982), .Y(n6980) );
  INVX1 U6926 ( .A(n6980), .Y(n6981) );
  BUFX2 U6927 ( .A(fifo[331]), .Y(n6982) );
  INVX1 U6928 ( .A(n6985), .Y(n6983) );
  INVX1 U6929 ( .A(n6983), .Y(n6984) );
  BUFX2 U6930 ( .A(fifo[332]), .Y(n6985) );
  INVX1 U6931 ( .A(n6988), .Y(n6986) );
  INVX1 U6932 ( .A(n6986), .Y(n6987) );
  BUFX2 U6933 ( .A(fifo[333]), .Y(n6988) );
  INVX1 U6934 ( .A(n6991), .Y(n6989) );
  INVX1 U6935 ( .A(n6989), .Y(n6990) );
  BUFX2 U6936 ( .A(fifo[334]), .Y(n6991) );
  INVX1 U6937 ( .A(n6994), .Y(n6992) );
  INVX1 U6938 ( .A(n6992), .Y(n6993) );
  BUFX2 U6939 ( .A(fifo[335]), .Y(n6994) );
  INVX1 U6940 ( .A(n6997), .Y(n6995) );
  INVX1 U6941 ( .A(n6995), .Y(n6996) );
  BUFX2 U6942 ( .A(fifo[336]), .Y(n6997) );
  INVX1 U6943 ( .A(n7000), .Y(n6998) );
  INVX1 U6944 ( .A(n6998), .Y(n6999) );
  BUFX2 U6945 ( .A(fifo[337]), .Y(n7000) );
  INVX1 U6946 ( .A(n7003), .Y(n7001) );
  INVX1 U6947 ( .A(n7001), .Y(n7002) );
  BUFX2 U6948 ( .A(fifo[338]), .Y(n7003) );
  INVX1 U6949 ( .A(n7006), .Y(n7004) );
  INVX1 U6950 ( .A(n7004), .Y(n7005) );
  BUFX2 U6951 ( .A(fifo[339]), .Y(n7006) );
  INVX1 U6952 ( .A(n7009), .Y(n7007) );
  INVX1 U6953 ( .A(n7007), .Y(n7008) );
  BUFX2 U6954 ( .A(fifo[510]), .Y(n7009) );
  INVX1 U6955 ( .A(n7012), .Y(n7010) );
  INVX1 U6956 ( .A(n7010), .Y(n7011) );
  BUFX2 U6957 ( .A(fifo[511]), .Y(n7012) );
  INVX1 U6958 ( .A(n7015), .Y(n7013) );
  INVX1 U6959 ( .A(n7013), .Y(n7014) );
  BUFX2 U6960 ( .A(fifo[512]), .Y(n7015) );
  INVX1 U6961 ( .A(n7018), .Y(n7016) );
  INVX1 U6962 ( .A(n7016), .Y(n7017) );
  BUFX2 U6963 ( .A(fifo[513]), .Y(n7018) );
  INVX1 U6964 ( .A(n7021), .Y(n7019) );
  INVX1 U6965 ( .A(n7019), .Y(n7020) );
  BUFX2 U6966 ( .A(fifo[514]), .Y(n7021) );
  INVX1 U6967 ( .A(n7024), .Y(n7022) );
  INVX1 U6968 ( .A(n7022), .Y(n7023) );
  BUFX2 U6969 ( .A(fifo[515]), .Y(n7024) );
  INVX1 U6970 ( .A(n7027), .Y(n7025) );
  INVX1 U6971 ( .A(n7025), .Y(n7026) );
  BUFX2 U6972 ( .A(fifo[516]), .Y(n7027) );
  INVX1 U6973 ( .A(n7030), .Y(n7028) );
  INVX1 U6974 ( .A(n7028), .Y(n7029) );
  BUFX2 U6975 ( .A(fifo[517]), .Y(n7030) );
  INVX1 U6976 ( .A(n7033), .Y(n7031) );
  INVX1 U6977 ( .A(n7031), .Y(n7032) );
  BUFX2 U6978 ( .A(fifo[518]), .Y(n7033) );
  INVX1 U6979 ( .A(n7036), .Y(n7034) );
  INVX1 U6980 ( .A(n7034), .Y(n7035) );
  BUFX2 U6981 ( .A(fifo[519]), .Y(n7036) );
  INVX1 U6982 ( .A(n7039), .Y(n7037) );
  INVX1 U6983 ( .A(n7037), .Y(n7038) );
  BUFX2 U6984 ( .A(fifo[520]), .Y(n7039) );
  INVX1 U6985 ( .A(n7042), .Y(n7040) );
  INVX1 U6986 ( .A(n7040), .Y(n7041) );
  BUFX2 U6987 ( .A(fifo[521]), .Y(n7042) );
  INVX1 U6988 ( .A(n7045), .Y(n7043) );
  INVX1 U6989 ( .A(n7043), .Y(n7044) );
  BUFX2 U6990 ( .A(fifo[522]), .Y(n7045) );
  INVX1 U6991 ( .A(n7048), .Y(n7046) );
  INVX1 U6992 ( .A(n7046), .Y(n7047) );
  BUFX2 U6993 ( .A(fifo[523]), .Y(n7048) );
  INVX1 U6994 ( .A(n7051), .Y(n7049) );
  INVX1 U6995 ( .A(n7049), .Y(n7050) );
  BUFX2 U6996 ( .A(fifo[524]), .Y(n7051) );
  INVX1 U6997 ( .A(n7054), .Y(n7052) );
  INVX1 U6998 ( .A(n7052), .Y(n7053) );
  BUFX2 U6999 ( .A(fifo[525]), .Y(n7054) );
  INVX1 U7000 ( .A(n7057), .Y(n7055) );
  INVX1 U7001 ( .A(n7055), .Y(n7056) );
  BUFX2 U7002 ( .A(fifo[526]), .Y(n7057) );
  INVX1 U7003 ( .A(n7060), .Y(n7058) );
  INVX1 U7004 ( .A(n7058), .Y(n7059) );
  BUFX2 U7005 ( .A(fifo[527]), .Y(n7060) );
  INVX1 U7006 ( .A(n7063), .Y(n7061) );
  INVX1 U7007 ( .A(n7061), .Y(n7062) );
  BUFX2 U7008 ( .A(fifo[528]), .Y(n7063) );
  INVX1 U7009 ( .A(n7066), .Y(n7064) );
  INVX1 U7010 ( .A(n7064), .Y(n7065) );
  BUFX2 U7011 ( .A(fifo[529]), .Y(n7066) );
  INVX1 U7012 ( .A(n7069), .Y(n7067) );
  INVX1 U7013 ( .A(n7067), .Y(n7068) );
  BUFX2 U7014 ( .A(fifo[530]), .Y(n7069) );
  INVX1 U7015 ( .A(n7072), .Y(n7070) );
  INVX1 U7016 ( .A(n7070), .Y(n7071) );
  BUFX2 U7017 ( .A(fifo[531]), .Y(n7072) );
  INVX1 U7018 ( .A(n7075), .Y(n7073) );
  INVX1 U7019 ( .A(n7073), .Y(n7074) );
  BUFX2 U7020 ( .A(fifo[532]), .Y(n7075) );
  INVX1 U7021 ( .A(n7078), .Y(n7076) );
  INVX1 U7022 ( .A(n7076), .Y(n7077) );
  BUFX2 U7023 ( .A(fifo[533]), .Y(n7078) );
  INVX1 U7024 ( .A(n7081), .Y(n7079) );
  INVX1 U7025 ( .A(n7079), .Y(n7080) );
  BUFX2 U7026 ( .A(fifo[534]), .Y(n7081) );
  INVX1 U7027 ( .A(n7084), .Y(n7082) );
  INVX1 U7028 ( .A(n7082), .Y(n7083) );
  BUFX2 U7029 ( .A(fifo[535]), .Y(n7084) );
  INVX1 U7030 ( .A(n7087), .Y(n7085) );
  INVX1 U7031 ( .A(n7085), .Y(n7086) );
  BUFX2 U7032 ( .A(fifo[536]), .Y(n7087) );
  INVX1 U7033 ( .A(n7090), .Y(n7088) );
  INVX1 U7034 ( .A(n7088), .Y(n7089) );
  BUFX2 U7035 ( .A(fifo[537]), .Y(n7090) );
  INVX1 U7036 ( .A(n7093), .Y(n7091) );
  INVX1 U7037 ( .A(n7091), .Y(n7092) );
  BUFX2 U7038 ( .A(fifo[538]), .Y(n7093) );
  INVX1 U7039 ( .A(n7096), .Y(n7094) );
  INVX1 U7040 ( .A(n7094), .Y(n7095) );
  BUFX2 U7041 ( .A(fifo[539]), .Y(n7096) );
  INVX1 U7042 ( .A(n7099), .Y(n7097) );
  INVX1 U7043 ( .A(n7097), .Y(n7098) );
  BUFX2 U7044 ( .A(fifo[540]), .Y(n7099) );
  INVX1 U7045 ( .A(n7102), .Y(n7100) );
  INVX1 U7046 ( .A(n7100), .Y(n7101) );
  BUFX2 U7047 ( .A(fifo[541]), .Y(n7102) );
  INVX1 U7048 ( .A(n7105), .Y(n7103) );
  INVX1 U7049 ( .A(n7103), .Y(n7104) );
  BUFX2 U7050 ( .A(fifo[542]), .Y(n7105) );
  INVX1 U7051 ( .A(n7108), .Y(n7106) );
  INVX1 U7052 ( .A(n7106), .Y(n7107) );
  BUFX2 U7053 ( .A(fifo[543]), .Y(n7108) );
  INVX1 U7054 ( .A(n7111), .Y(n7109) );
  INVX1 U7055 ( .A(n7109), .Y(n7110) );
  BUFX2 U7056 ( .A(fifo[1054]), .Y(n7111) );
  INVX1 U7057 ( .A(n7114), .Y(n7112) );
  INVX1 U7058 ( .A(n7112), .Y(n7113) );
  BUFX2 U7059 ( .A(fifo[1055]), .Y(n7114) );
  INVX1 U7060 ( .A(n7117), .Y(n7115) );
  INVX1 U7061 ( .A(n7115), .Y(n7116) );
  BUFX2 U7062 ( .A(fifo[1056]), .Y(n7117) );
  INVX1 U7063 ( .A(n7120), .Y(n7118) );
  INVX1 U7064 ( .A(n7118), .Y(n7119) );
  BUFX2 U7065 ( .A(fifo[1057]), .Y(n7120) );
  INVX1 U7066 ( .A(n7123), .Y(n7121) );
  INVX1 U7067 ( .A(n7121), .Y(n7122) );
  BUFX2 U7068 ( .A(fifo[1058]), .Y(n7123) );
  INVX1 U7069 ( .A(n7126), .Y(n7124) );
  INVX1 U7070 ( .A(n7124), .Y(n7125) );
  BUFX2 U7071 ( .A(fifo[1059]), .Y(n7126) );
  INVX1 U7072 ( .A(n7129), .Y(n7127) );
  INVX1 U7073 ( .A(n7127), .Y(n7128) );
  BUFX2 U7074 ( .A(fifo[1060]), .Y(n7129) );
  INVX1 U7075 ( .A(n7132), .Y(n7130) );
  INVX1 U7076 ( .A(n7130), .Y(n7131) );
  BUFX2 U7077 ( .A(fifo[1061]), .Y(n7132) );
  INVX1 U7078 ( .A(n7135), .Y(n7133) );
  INVX1 U7079 ( .A(n7133), .Y(n7134) );
  BUFX2 U7080 ( .A(fifo[1062]), .Y(n7135) );
  INVX1 U7081 ( .A(n7138), .Y(n7136) );
  INVX1 U7082 ( .A(n7136), .Y(n7137) );
  BUFX2 U7083 ( .A(fifo[1063]), .Y(n7138) );
  INVX1 U7084 ( .A(n7141), .Y(n7139) );
  INVX1 U7085 ( .A(n7139), .Y(n7140) );
  BUFX2 U7086 ( .A(fifo[1064]), .Y(n7141) );
  INVX1 U7087 ( .A(n7144), .Y(n7142) );
  INVX1 U7088 ( .A(n7142), .Y(n7143) );
  BUFX2 U7089 ( .A(fifo[1065]), .Y(n7144) );
  INVX1 U7090 ( .A(n7147), .Y(n7145) );
  INVX1 U7091 ( .A(n7145), .Y(n7146) );
  BUFX2 U7092 ( .A(fifo[1066]), .Y(n7147) );
  INVX1 U7093 ( .A(n7150), .Y(n7148) );
  INVX1 U7094 ( .A(n7148), .Y(n7149) );
  BUFX2 U7095 ( .A(fifo[1067]), .Y(n7150) );
  INVX1 U7096 ( .A(n7153), .Y(n7151) );
  INVX1 U7097 ( .A(n7151), .Y(n7152) );
  BUFX2 U7098 ( .A(fifo[1068]), .Y(n7153) );
  INVX1 U7099 ( .A(n7156), .Y(n7154) );
  INVX1 U7100 ( .A(n7154), .Y(n7155) );
  BUFX2 U7101 ( .A(fifo[1069]), .Y(n7156) );
  INVX1 U7102 ( .A(n7159), .Y(n7157) );
  INVX1 U7103 ( .A(n7157), .Y(n7158) );
  BUFX2 U7104 ( .A(fifo[1070]), .Y(n7159) );
  INVX1 U7105 ( .A(n7162), .Y(n7160) );
  INVX1 U7106 ( .A(n7160), .Y(n7161) );
  BUFX2 U7107 ( .A(fifo[1071]), .Y(n7162) );
  INVX1 U7108 ( .A(n7165), .Y(n7163) );
  INVX1 U7109 ( .A(n7163), .Y(n7164) );
  BUFX2 U7110 ( .A(fifo[1072]), .Y(n7165) );
  INVX1 U7111 ( .A(n7168), .Y(n7166) );
  INVX1 U7112 ( .A(n7166), .Y(n7167) );
  BUFX2 U7113 ( .A(fifo[1073]), .Y(n7168) );
  INVX1 U7114 ( .A(n7171), .Y(n7169) );
  INVX1 U7115 ( .A(n7169), .Y(n7170) );
  BUFX2 U7116 ( .A(fifo[1074]), .Y(n7171) );
  INVX1 U7117 ( .A(n7174), .Y(n7172) );
  INVX1 U7118 ( .A(n7172), .Y(n7173) );
  BUFX2 U7119 ( .A(fifo[1075]), .Y(n7174) );
  INVX1 U7120 ( .A(n7177), .Y(n7175) );
  INVX1 U7121 ( .A(n7175), .Y(n7176) );
  BUFX2 U7122 ( .A(fifo[1076]), .Y(n7177) );
  INVX1 U7123 ( .A(n7180), .Y(n7178) );
  INVX1 U7124 ( .A(n7178), .Y(n7179) );
  BUFX2 U7125 ( .A(fifo[1077]), .Y(n7180) );
  INVX1 U7126 ( .A(n7183), .Y(n7181) );
  INVX1 U7127 ( .A(n7181), .Y(n7182) );
  BUFX2 U7128 ( .A(fifo[1078]), .Y(n7183) );
  INVX1 U7129 ( .A(n7186), .Y(n7184) );
  INVX1 U7130 ( .A(n7184), .Y(n7185) );
  BUFX2 U7131 ( .A(fifo[1079]), .Y(n7186) );
  INVX1 U7132 ( .A(n7189), .Y(n7187) );
  INVX1 U7133 ( .A(n7187), .Y(n7188) );
  BUFX2 U7134 ( .A(fifo[1080]), .Y(n7189) );
  INVX1 U7135 ( .A(n7192), .Y(n7190) );
  INVX1 U7136 ( .A(n7190), .Y(n7191) );
  BUFX2 U7137 ( .A(fifo[1081]), .Y(n7192) );
  INVX1 U7138 ( .A(n7195), .Y(n7193) );
  INVX1 U7139 ( .A(n7193), .Y(n7194) );
  BUFX2 U7140 ( .A(fifo[1082]), .Y(n7195) );
  INVX1 U7141 ( .A(n7198), .Y(n7196) );
  INVX1 U7142 ( .A(n7196), .Y(n7197) );
  BUFX2 U7143 ( .A(fifo[1083]), .Y(n7198) );
  INVX1 U7144 ( .A(n7201), .Y(n7199) );
  INVX1 U7145 ( .A(n7199), .Y(n7200) );
  BUFX2 U7146 ( .A(fifo[1084]), .Y(n7201) );
  INVX1 U7147 ( .A(n7204), .Y(n7202) );
  INVX1 U7148 ( .A(n7202), .Y(n7203) );
  BUFX2 U7149 ( .A(fifo[1085]), .Y(n7204) );
  INVX1 U7150 ( .A(n7207), .Y(n7205) );
  INVX1 U7151 ( .A(n7205), .Y(n7206) );
  BUFX2 U7152 ( .A(fifo[1086]), .Y(n7207) );
  INVX1 U7153 ( .A(n7210), .Y(n7208) );
  INVX1 U7154 ( .A(n7208), .Y(n7209) );
  BUFX2 U7155 ( .A(fifo[1087]), .Y(n7210) );
  INVX1 U7156 ( .A(n7213), .Y(n7211) );
  INVX1 U7157 ( .A(n7211), .Y(n7212) );
  BUFX2 U7158 ( .A(fifo[34]), .Y(n7213) );
  INVX1 U7159 ( .A(n7216), .Y(n7214) );
  INVX1 U7160 ( .A(n7214), .Y(n7215) );
  BUFX2 U7161 ( .A(fifo[35]), .Y(n7216) );
  INVX1 U7162 ( .A(n7219), .Y(n7217) );
  INVX1 U7163 ( .A(n7217), .Y(n7218) );
  BUFX2 U7164 ( .A(fifo[36]), .Y(n7219) );
  INVX1 U7165 ( .A(n7222), .Y(n7220) );
  INVX1 U7166 ( .A(n7220), .Y(n7221) );
  BUFX2 U7167 ( .A(fifo[37]), .Y(n7222) );
  INVX1 U7168 ( .A(n7225), .Y(n7223) );
  INVX1 U7169 ( .A(n7223), .Y(n7224) );
  BUFX2 U7170 ( .A(fifo[38]), .Y(n7225) );
  INVX1 U7171 ( .A(n7228), .Y(n7226) );
  INVX1 U7172 ( .A(n7226), .Y(n7227) );
  BUFX2 U7173 ( .A(fifo[39]), .Y(n7228) );
  INVX1 U7174 ( .A(n7231), .Y(n7229) );
  INVX1 U7175 ( .A(n7229), .Y(n7230) );
  BUFX2 U7176 ( .A(fifo[40]), .Y(n7231) );
  INVX1 U7177 ( .A(n7234), .Y(n7232) );
  INVX1 U7178 ( .A(n7232), .Y(n7233) );
  BUFX2 U7179 ( .A(fifo[41]), .Y(n7234) );
  INVX1 U7180 ( .A(n7237), .Y(n7235) );
  INVX1 U7181 ( .A(n7235), .Y(n7236) );
  BUFX2 U7182 ( .A(fifo[42]), .Y(n7237) );
  INVX1 U7183 ( .A(n7240), .Y(n7238) );
  INVX1 U7184 ( .A(n7238), .Y(n7239) );
  BUFX2 U7185 ( .A(fifo[43]), .Y(n7240) );
  INVX1 U7186 ( .A(n7243), .Y(n7241) );
  INVX1 U7187 ( .A(n7241), .Y(n7242) );
  BUFX2 U7188 ( .A(fifo[44]), .Y(n7243) );
  INVX1 U7189 ( .A(n7246), .Y(n7244) );
  INVX1 U7190 ( .A(n7244), .Y(n7245) );
  BUFX2 U7191 ( .A(fifo[45]), .Y(n7246) );
  INVX1 U7192 ( .A(n7249), .Y(n7247) );
  INVX1 U7193 ( .A(n7247), .Y(n7248) );
  BUFX2 U7194 ( .A(fifo[46]), .Y(n7249) );
  INVX1 U7195 ( .A(n7252), .Y(n7250) );
  INVX1 U7196 ( .A(n7250), .Y(n7251) );
  BUFX2 U7197 ( .A(fifo[47]), .Y(n7252) );
  INVX1 U7198 ( .A(n7255), .Y(n7253) );
  INVX1 U7199 ( .A(n7253), .Y(n7254) );
  BUFX2 U7200 ( .A(fifo[48]), .Y(n7255) );
  INVX1 U7201 ( .A(n7258), .Y(n7256) );
  INVX1 U7202 ( .A(n7256), .Y(n7257) );
  BUFX2 U7203 ( .A(fifo[49]), .Y(n7258) );
  INVX1 U7204 ( .A(n7261), .Y(n7259) );
  INVX1 U7205 ( .A(n7259), .Y(n7260) );
  BUFX2 U7206 ( .A(fifo[50]), .Y(n7261) );
  INVX1 U7207 ( .A(n7264), .Y(n7262) );
  INVX1 U7208 ( .A(n7262), .Y(n7263) );
  BUFX2 U7209 ( .A(fifo[51]), .Y(n7264) );
  INVX1 U7210 ( .A(n7267), .Y(n7265) );
  INVX1 U7211 ( .A(n7265), .Y(n7266) );
  BUFX2 U7212 ( .A(fifo[52]), .Y(n7267) );
  INVX1 U7213 ( .A(n7270), .Y(n7268) );
  INVX1 U7214 ( .A(n7268), .Y(n7269) );
  BUFX2 U7215 ( .A(fifo[53]), .Y(n7270) );
  INVX1 U7216 ( .A(n7273), .Y(n7271) );
  INVX1 U7217 ( .A(n7271), .Y(n7272) );
  BUFX2 U7218 ( .A(fifo[54]), .Y(n7273) );
  INVX1 U7219 ( .A(n7276), .Y(n7274) );
  INVX1 U7220 ( .A(n7274), .Y(n7275) );
  BUFX2 U7221 ( .A(fifo[55]), .Y(n7276) );
  INVX1 U7222 ( .A(n7279), .Y(n7277) );
  INVX1 U7223 ( .A(n7277), .Y(n7278) );
  BUFX2 U7224 ( .A(fifo[56]), .Y(n7279) );
  INVX1 U7225 ( .A(n7282), .Y(n7280) );
  INVX1 U7226 ( .A(n7280), .Y(n7281) );
  BUFX2 U7227 ( .A(fifo[57]), .Y(n7282) );
  INVX1 U7228 ( .A(n7285), .Y(n7283) );
  INVX1 U7229 ( .A(n7283), .Y(n7284) );
  BUFX2 U7230 ( .A(fifo[58]), .Y(n7285) );
  INVX1 U7231 ( .A(n7288), .Y(n7286) );
  INVX1 U7232 ( .A(n7286), .Y(n7287) );
  BUFX2 U7233 ( .A(fifo[59]), .Y(n7288) );
  INVX1 U7234 ( .A(n7291), .Y(n7289) );
  INVX1 U7235 ( .A(n7289), .Y(n7290) );
  BUFX2 U7236 ( .A(fifo[60]), .Y(n7291) );
  INVX1 U7237 ( .A(n7294), .Y(n7292) );
  INVX1 U7238 ( .A(n7292), .Y(n7293) );
  BUFX2 U7239 ( .A(fifo[61]), .Y(n7294) );
  INVX1 U7240 ( .A(n7297), .Y(n7295) );
  INVX1 U7241 ( .A(n7295), .Y(n7296) );
  BUFX2 U7242 ( .A(fifo[62]), .Y(n7297) );
  INVX1 U7243 ( .A(n7300), .Y(n7298) );
  INVX1 U7244 ( .A(n7298), .Y(n7299) );
  BUFX2 U7245 ( .A(fifo[63]), .Y(n7300) );
  INVX1 U7246 ( .A(n7303), .Y(n7301) );
  INVX1 U7247 ( .A(n7301), .Y(n7302) );
  BUFX2 U7248 ( .A(fifo[64]), .Y(n7303) );
  INVX1 U7249 ( .A(n7306), .Y(n7304) );
  INVX1 U7250 ( .A(n7304), .Y(n7305) );
  BUFX2 U7251 ( .A(fifo[65]), .Y(n7306) );
  INVX1 U7252 ( .A(n7309), .Y(n7307) );
  INVX1 U7253 ( .A(n7307), .Y(n7308) );
  BUFX2 U7254 ( .A(fifo[66]), .Y(n7309) );
  INVX1 U7255 ( .A(n7312), .Y(n7310) );
  INVX1 U7256 ( .A(n7310), .Y(n7311) );
  BUFX2 U7257 ( .A(fifo[67]), .Y(n7312) );
  INVX1 U7258 ( .A(n7315), .Y(n7313) );
  INVX1 U7259 ( .A(n7313), .Y(n7314) );
  BUFX2 U7260 ( .A(fifo[102]), .Y(n7315) );
  INVX1 U7261 ( .A(n7318), .Y(n7316) );
  INVX1 U7262 ( .A(n7316), .Y(n7317) );
  BUFX2 U7263 ( .A(fifo[103]), .Y(n7318) );
  INVX1 U7264 ( .A(n7321), .Y(n7319) );
  INVX1 U7265 ( .A(n7319), .Y(n7320) );
  BUFX2 U7266 ( .A(fifo[104]), .Y(n7321) );
  INVX1 U7267 ( .A(n7324), .Y(n7322) );
  INVX1 U7268 ( .A(n7322), .Y(n7323) );
  BUFX2 U7269 ( .A(fifo[105]), .Y(n7324) );
  INVX1 U7270 ( .A(n7327), .Y(n7325) );
  INVX1 U7271 ( .A(n7325), .Y(n7326) );
  BUFX2 U7272 ( .A(fifo[106]), .Y(n7327) );
  INVX1 U7273 ( .A(n7330), .Y(n7328) );
  INVX1 U7274 ( .A(n7328), .Y(n7329) );
  BUFX2 U7275 ( .A(fifo[107]), .Y(n7330) );
  INVX1 U7276 ( .A(n7333), .Y(n7331) );
  INVX1 U7277 ( .A(n7331), .Y(n7332) );
  BUFX2 U7278 ( .A(fifo[108]), .Y(n7333) );
  INVX1 U7279 ( .A(n7336), .Y(n7334) );
  INVX1 U7280 ( .A(n7334), .Y(n7335) );
  BUFX2 U7281 ( .A(fifo[109]), .Y(n7336) );
  INVX1 U7282 ( .A(n7339), .Y(n7337) );
  INVX1 U7283 ( .A(n7337), .Y(n7338) );
  BUFX2 U7284 ( .A(fifo[110]), .Y(n7339) );
  INVX1 U7285 ( .A(n7342), .Y(n7340) );
  INVX1 U7286 ( .A(n7340), .Y(n7341) );
  BUFX2 U7287 ( .A(fifo[111]), .Y(n7342) );
  INVX1 U7288 ( .A(n7345), .Y(n7343) );
  INVX1 U7289 ( .A(n7343), .Y(n7344) );
  BUFX2 U7290 ( .A(fifo[112]), .Y(n7345) );
  INVX1 U7291 ( .A(n7348), .Y(n7346) );
  INVX1 U7292 ( .A(n7346), .Y(n7347) );
  BUFX2 U7293 ( .A(fifo[113]), .Y(n7348) );
  INVX1 U7294 ( .A(n7351), .Y(n7349) );
  INVX1 U7295 ( .A(n7349), .Y(n7350) );
  BUFX2 U7296 ( .A(fifo[114]), .Y(n7351) );
  INVX1 U7297 ( .A(n7354), .Y(n7352) );
  INVX1 U7298 ( .A(n7352), .Y(n7353) );
  BUFX2 U7299 ( .A(fifo[115]), .Y(n7354) );
  INVX1 U7300 ( .A(n7357), .Y(n7355) );
  INVX1 U7301 ( .A(n7355), .Y(n7356) );
  BUFX2 U7302 ( .A(fifo[116]), .Y(n7357) );
  INVX1 U7303 ( .A(n7360), .Y(n7358) );
  INVX1 U7304 ( .A(n7358), .Y(n7359) );
  BUFX2 U7305 ( .A(fifo[117]), .Y(n7360) );
  INVX1 U7306 ( .A(n7363), .Y(n7361) );
  INVX1 U7307 ( .A(n7361), .Y(n7362) );
  BUFX2 U7308 ( .A(fifo[118]), .Y(n7363) );
  INVX1 U7309 ( .A(n7366), .Y(n7364) );
  INVX1 U7310 ( .A(n7364), .Y(n7365) );
  BUFX2 U7311 ( .A(fifo[119]), .Y(n7366) );
  INVX1 U7312 ( .A(n7369), .Y(n7367) );
  INVX1 U7313 ( .A(n7367), .Y(n7368) );
  BUFX2 U7314 ( .A(fifo[120]), .Y(n7369) );
  INVX1 U7315 ( .A(n7372), .Y(n7370) );
  INVX1 U7316 ( .A(n7370), .Y(n7371) );
  BUFX2 U7317 ( .A(fifo[121]), .Y(n7372) );
  INVX1 U7318 ( .A(n7375), .Y(n7373) );
  INVX1 U7319 ( .A(n7373), .Y(n7374) );
  BUFX2 U7320 ( .A(fifo[122]), .Y(n7375) );
  INVX1 U7321 ( .A(n7378), .Y(n7376) );
  INVX1 U7322 ( .A(n7376), .Y(n7377) );
  BUFX2 U7323 ( .A(fifo[123]), .Y(n7378) );
  INVX1 U7324 ( .A(n7381), .Y(n7379) );
  INVX1 U7325 ( .A(n7379), .Y(n7380) );
  BUFX2 U7326 ( .A(fifo[124]), .Y(n7381) );
  INVX1 U7327 ( .A(n7384), .Y(n7382) );
  INVX1 U7328 ( .A(n7382), .Y(n7383) );
  BUFX2 U7329 ( .A(fifo[125]), .Y(n7384) );
  INVX1 U7330 ( .A(n7387), .Y(n7385) );
  INVX1 U7331 ( .A(n7385), .Y(n7386) );
  BUFX2 U7332 ( .A(fifo[126]), .Y(n7387) );
  INVX1 U7333 ( .A(n7390), .Y(n7388) );
  INVX1 U7334 ( .A(n7388), .Y(n7389) );
  BUFX2 U7335 ( .A(fifo[127]), .Y(n7390) );
  INVX1 U7336 ( .A(n7393), .Y(n7391) );
  INVX1 U7337 ( .A(n7391), .Y(n7392) );
  BUFX2 U7338 ( .A(fifo[128]), .Y(n7393) );
  INVX1 U7339 ( .A(n7396), .Y(n7394) );
  INVX1 U7340 ( .A(n7394), .Y(n7395) );
  BUFX2 U7341 ( .A(fifo[129]), .Y(n7396) );
  INVX1 U7342 ( .A(n7399), .Y(n7397) );
  INVX1 U7343 ( .A(n7397), .Y(n7398) );
  BUFX2 U7344 ( .A(fifo[130]), .Y(n7399) );
  INVX1 U7345 ( .A(n7402), .Y(n7400) );
  INVX1 U7346 ( .A(n7400), .Y(n7401) );
  BUFX2 U7347 ( .A(fifo[131]), .Y(n7402) );
  INVX1 U7348 ( .A(n7405), .Y(n7403) );
  INVX1 U7349 ( .A(n7403), .Y(n7404) );
  BUFX2 U7350 ( .A(fifo[132]), .Y(n7405) );
  INVX1 U7351 ( .A(n7408), .Y(n7406) );
  INVX1 U7352 ( .A(n7406), .Y(n7407) );
  BUFX2 U7353 ( .A(fifo[133]), .Y(n7408) );
  INVX1 U7354 ( .A(n7411), .Y(n7409) );
  INVX1 U7355 ( .A(n7409), .Y(n7410) );
  BUFX2 U7356 ( .A(fifo[134]), .Y(n7411) );
  INVX1 U7357 ( .A(n7414), .Y(n7412) );
  INVX1 U7358 ( .A(n7412), .Y(n7413) );
  BUFX2 U7359 ( .A(fifo[135]), .Y(n7414) );
  INVX1 U7360 ( .A(n7417), .Y(n7415) );
  INVX1 U7361 ( .A(n7415), .Y(n7416) );
  BUFX2 U7362 ( .A(fifo[170]), .Y(n7417) );
  INVX1 U7363 ( .A(n7420), .Y(n7418) );
  INVX1 U7364 ( .A(n7418), .Y(n7419) );
  BUFX2 U7365 ( .A(fifo[171]), .Y(n7420) );
  INVX1 U7366 ( .A(n7423), .Y(n7421) );
  INVX1 U7367 ( .A(n7421), .Y(n7422) );
  BUFX2 U7368 ( .A(fifo[172]), .Y(n7423) );
  INVX1 U7369 ( .A(n7426), .Y(n7424) );
  INVX1 U7370 ( .A(n7424), .Y(n7425) );
  BUFX2 U7371 ( .A(fifo[173]), .Y(n7426) );
  INVX1 U7372 ( .A(n7429), .Y(n7427) );
  INVX1 U7373 ( .A(n7427), .Y(n7428) );
  BUFX2 U7374 ( .A(fifo[174]), .Y(n7429) );
  INVX1 U7375 ( .A(n7432), .Y(n7430) );
  INVX1 U7376 ( .A(n7430), .Y(n7431) );
  BUFX2 U7377 ( .A(fifo[175]), .Y(n7432) );
  INVX1 U7378 ( .A(n7435), .Y(n7433) );
  INVX1 U7379 ( .A(n7433), .Y(n7434) );
  BUFX2 U7380 ( .A(fifo[176]), .Y(n7435) );
  INVX1 U7381 ( .A(n7438), .Y(n7436) );
  INVX1 U7382 ( .A(n7436), .Y(n7437) );
  BUFX2 U7383 ( .A(fifo[177]), .Y(n7438) );
  INVX1 U7384 ( .A(n7441), .Y(n7439) );
  INVX1 U7385 ( .A(n7439), .Y(n7440) );
  BUFX2 U7386 ( .A(fifo[178]), .Y(n7441) );
  INVX1 U7387 ( .A(n7444), .Y(n7442) );
  INVX1 U7388 ( .A(n7442), .Y(n7443) );
  BUFX2 U7389 ( .A(fifo[179]), .Y(n7444) );
  INVX1 U7390 ( .A(n7447), .Y(n7445) );
  INVX1 U7391 ( .A(n7445), .Y(n7446) );
  BUFX2 U7392 ( .A(fifo[180]), .Y(n7447) );
  INVX1 U7393 ( .A(n7450), .Y(n7448) );
  INVX1 U7394 ( .A(n7448), .Y(n7449) );
  BUFX2 U7395 ( .A(fifo[181]), .Y(n7450) );
  INVX1 U7396 ( .A(n7453), .Y(n7451) );
  INVX1 U7397 ( .A(n7451), .Y(n7452) );
  BUFX2 U7398 ( .A(fifo[182]), .Y(n7453) );
  INVX1 U7399 ( .A(n7456), .Y(n7454) );
  INVX1 U7400 ( .A(n7454), .Y(n7455) );
  BUFX2 U7401 ( .A(fifo[183]), .Y(n7456) );
  INVX1 U7402 ( .A(n7459), .Y(n7457) );
  INVX1 U7403 ( .A(n7457), .Y(n7458) );
  BUFX2 U7404 ( .A(fifo[184]), .Y(n7459) );
  INVX1 U7405 ( .A(n7462), .Y(n7460) );
  INVX1 U7406 ( .A(n7460), .Y(n7461) );
  BUFX2 U7407 ( .A(fifo[185]), .Y(n7462) );
  INVX1 U7408 ( .A(n7465), .Y(n7463) );
  INVX1 U7409 ( .A(n7463), .Y(n7464) );
  BUFX2 U7410 ( .A(fifo[186]), .Y(n7465) );
  INVX1 U7411 ( .A(n7468), .Y(n7466) );
  INVX1 U7412 ( .A(n7466), .Y(n7467) );
  BUFX2 U7413 ( .A(fifo[187]), .Y(n7468) );
  INVX1 U7414 ( .A(n7471), .Y(n7469) );
  INVX1 U7415 ( .A(n7469), .Y(n7470) );
  BUFX2 U7416 ( .A(fifo[188]), .Y(n7471) );
  INVX1 U7417 ( .A(n7474), .Y(n7472) );
  INVX1 U7418 ( .A(n7472), .Y(n7473) );
  BUFX2 U7419 ( .A(fifo[189]), .Y(n7474) );
  INVX1 U7420 ( .A(n7477), .Y(n7475) );
  INVX1 U7421 ( .A(n7475), .Y(n7476) );
  BUFX2 U7422 ( .A(fifo[190]), .Y(n7477) );
  INVX1 U7423 ( .A(n7480), .Y(n7478) );
  INVX1 U7424 ( .A(n7478), .Y(n7479) );
  BUFX2 U7425 ( .A(fifo[191]), .Y(n7480) );
  INVX1 U7426 ( .A(n7483), .Y(n7481) );
  INVX1 U7427 ( .A(n7481), .Y(n7482) );
  BUFX2 U7428 ( .A(fifo[192]), .Y(n7483) );
  INVX1 U7429 ( .A(n7486), .Y(n7484) );
  INVX1 U7430 ( .A(n7484), .Y(n7485) );
  BUFX2 U7431 ( .A(fifo[193]), .Y(n7486) );
  INVX1 U7432 ( .A(n7489), .Y(n7487) );
  INVX1 U7433 ( .A(n7487), .Y(n7488) );
  BUFX2 U7434 ( .A(fifo[194]), .Y(n7489) );
  INVX1 U7435 ( .A(n7492), .Y(n7490) );
  INVX1 U7436 ( .A(n7490), .Y(n7491) );
  BUFX2 U7437 ( .A(fifo[195]), .Y(n7492) );
  INVX1 U7438 ( .A(n7495), .Y(n7493) );
  INVX1 U7439 ( .A(n7493), .Y(n7494) );
  BUFX2 U7440 ( .A(fifo[196]), .Y(n7495) );
  INVX1 U7441 ( .A(n7498), .Y(n7496) );
  INVX1 U7442 ( .A(n7496), .Y(n7497) );
  BUFX2 U7443 ( .A(fifo[197]), .Y(n7498) );
  INVX1 U7444 ( .A(n7501), .Y(n7499) );
  INVX1 U7445 ( .A(n7499), .Y(n7500) );
  BUFX2 U7446 ( .A(fifo[198]), .Y(n7501) );
  INVX1 U7447 ( .A(n7504), .Y(n7502) );
  INVX1 U7448 ( .A(n7502), .Y(n7503) );
  BUFX2 U7449 ( .A(fifo[199]), .Y(n7504) );
  INVX1 U7450 ( .A(n7507), .Y(n7505) );
  INVX1 U7451 ( .A(n7505), .Y(n7506) );
  BUFX2 U7452 ( .A(fifo[200]), .Y(n7507) );
  INVX1 U7453 ( .A(n7510), .Y(n7508) );
  INVX1 U7454 ( .A(n7508), .Y(n7509) );
  BUFX2 U7455 ( .A(fifo[201]), .Y(n7510) );
  INVX1 U7456 ( .A(n7513), .Y(n7511) );
  INVX1 U7457 ( .A(n7511), .Y(n7512) );
  BUFX2 U7458 ( .A(fifo[202]), .Y(n7513) );
  INVX1 U7459 ( .A(n7516), .Y(n7514) );
  INVX1 U7460 ( .A(n7514), .Y(n7515) );
  BUFX2 U7461 ( .A(fifo[203]), .Y(n7516) );
  INVX1 U7462 ( .A(n7519), .Y(n7517) );
  INVX1 U7463 ( .A(n7517), .Y(n7518) );
  BUFX2 U7464 ( .A(fifo[238]), .Y(n7519) );
  INVX1 U7465 ( .A(n7522), .Y(n7520) );
  INVX1 U7466 ( .A(n7520), .Y(n7521) );
  BUFX2 U7467 ( .A(fifo[239]), .Y(n7522) );
  INVX1 U7468 ( .A(n7525), .Y(n7523) );
  INVX1 U7469 ( .A(n7523), .Y(n7524) );
  BUFX2 U7470 ( .A(fifo[240]), .Y(n7525) );
  INVX1 U7471 ( .A(n7528), .Y(n7526) );
  INVX1 U7472 ( .A(n7526), .Y(n7527) );
  BUFX2 U7473 ( .A(fifo[241]), .Y(n7528) );
  INVX1 U7474 ( .A(n7531), .Y(n7529) );
  INVX1 U7475 ( .A(n7529), .Y(n7530) );
  BUFX2 U7476 ( .A(fifo[242]), .Y(n7531) );
  INVX1 U7477 ( .A(n7534), .Y(n7532) );
  INVX1 U7478 ( .A(n7532), .Y(n7533) );
  BUFX2 U7479 ( .A(fifo[243]), .Y(n7534) );
  INVX1 U7480 ( .A(n7537), .Y(n7535) );
  INVX1 U7481 ( .A(n7535), .Y(n7536) );
  BUFX2 U7482 ( .A(fifo[244]), .Y(n7537) );
  INVX1 U7483 ( .A(n7540), .Y(n7538) );
  INVX1 U7484 ( .A(n7538), .Y(n7539) );
  BUFX2 U7485 ( .A(fifo[245]), .Y(n7540) );
  INVX1 U7486 ( .A(n7543), .Y(n7541) );
  INVX1 U7487 ( .A(n7541), .Y(n7542) );
  BUFX2 U7488 ( .A(fifo[246]), .Y(n7543) );
  INVX1 U7489 ( .A(n7546), .Y(n7544) );
  INVX1 U7490 ( .A(n7544), .Y(n7545) );
  BUFX2 U7491 ( .A(fifo[247]), .Y(n7546) );
  INVX1 U7492 ( .A(n7549), .Y(n7547) );
  INVX1 U7493 ( .A(n7547), .Y(n7548) );
  BUFX2 U7494 ( .A(fifo[248]), .Y(n7549) );
  INVX1 U7495 ( .A(n7552), .Y(n7550) );
  INVX1 U7496 ( .A(n7550), .Y(n7551) );
  BUFX2 U7497 ( .A(fifo[249]), .Y(n7552) );
  INVX1 U7498 ( .A(n7555), .Y(n7553) );
  INVX1 U7499 ( .A(n7553), .Y(n7554) );
  BUFX2 U7500 ( .A(fifo[250]), .Y(n7555) );
  INVX1 U7501 ( .A(n7558), .Y(n7556) );
  INVX1 U7502 ( .A(n7556), .Y(n7557) );
  BUFX2 U7503 ( .A(fifo[251]), .Y(n7558) );
  INVX1 U7504 ( .A(n7561), .Y(n7559) );
  INVX1 U7505 ( .A(n7559), .Y(n7560) );
  BUFX2 U7506 ( .A(fifo[252]), .Y(n7561) );
  INVX1 U7507 ( .A(n7564), .Y(n7562) );
  INVX1 U7508 ( .A(n7562), .Y(n7563) );
  BUFX2 U7509 ( .A(fifo[253]), .Y(n7564) );
  INVX1 U7510 ( .A(n7567), .Y(n7565) );
  INVX1 U7511 ( .A(n7565), .Y(n7566) );
  BUFX2 U7512 ( .A(fifo[254]), .Y(n7567) );
  INVX1 U7513 ( .A(n7570), .Y(n7568) );
  INVX1 U7514 ( .A(n7568), .Y(n7569) );
  BUFX2 U7515 ( .A(fifo[255]), .Y(n7570) );
  INVX1 U7516 ( .A(n7573), .Y(n7571) );
  INVX1 U7517 ( .A(n7571), .Y(n7572) );
  BUFX2 U7518 ( .A(fifo[256]), .Y(n7573) );
  INVX1 U7519 ( .A(n7576), .Y(n7574) );
  INVX1 U7520 ( .A(n7574), .Y(n7575) );
  BUFX2 U7521 ( .A(fifo[257]), .Y(n7576) );
  INVX1 U7522 ( .A(n7579), .Y(n7577) );
  INVX1 U7523 ( .A(n7577), .Y(n7578) );
  BUFX2 U7524 ( .A(fifo[258]), .Y(n7579) );
  INVX1 U7525 ( .A(n7582), .Y(n7580) );
  INVX1 U7526 ( .A(n7580), .Y(n7581) );
  BUFX2 U7527 ( .A(fifo[259]), .Y(n7582) );
  INVX1 U7528 ( .A(n7585), .Y(n7583) );
  INVX1 U7529 ( .A(n7583), .Y(n7584) );
  BUFX2 U7530 ( .A(fifo[260]), .Y(n7585) );
  INVX1 U7531 ( .A(n7588), .Y(n7586) );
  INVX1 U7532 ( .A(n7586), .Y(n7587) );
  BUFX2 U7533 ( .A(fifo[261]), .Y(n7588) );
  INVX1 U7534 ( .A(n7591), .Y(n7589) );
  INVX1 U7535 ( .A(n7589), .Y(n7590) );
  BUFX2 U7536 ( .A(fifo[262]), .Y(n7591) );
  INVX1 U7537 ( .A(n7594), .Y(n7592) );
  INVX1 U7538 ( .A(n7592), .Y(n7593) );
  BUFX2 U7539 ( .A(fifo[263]), .Y(n7594) );
  INVX1 U7540 ( .A(n7597), .Y(n7595) );
  INVX1 U7541 ( .A(n7595), .Y(n7596) );
  BUFX2 U7542 ( .A(fifo[264]), .Y(n7597) );
  INVX1 U7543 ( .A(n7600), .Y(n7598) );
  INVX1 U7544 ( .A(n7598), .Y(n7599) );
  BUFX2 U7545 ( .A(fifo[265]), .Y(n7600) );
  INVX1 U7546 ( .A(n7603), .Y(n7601) );
  INVX1 U7547 ( .A(n7601), .Y(n7602) );
  BUFX2 U7548 ( .A(fifo[266]), .Y(n7603) );
  INVX1 U7549 ( .A(n7606), .Y(n7604) );
  INVX1 U7550 ( .A(n7604), .Y(n7605) );
  BUFX2 U7551 ( .A(fifo[267]), .Y(n7606) );
  INVX1 U7552 ( .A(n7609), .Y(n7607) );
  INVX1 U7553 ( .A(n7607), .Y(n7608) );
  BUFX2 U7554 ( .A(fifo[268]), .Y(n7609) );
  INVX1 U7555 ( .A(n7612), .Y(n7610) );
  INVX1 U7556 ( .A(n7610), .Y(n7611) );
  BUFX2 U7557 ( .A(fifo[269]), .Y(n7612) );
  INVX1 U7558 ( .A(n7615), .Y(n7613) );
  INVX1 U7559 ( .A(n7613), .Y(n7614) );
  BUFX2 U7560 ( .A(fifo[270]), .Y(n7615) );
  INVX1 U7561 ( .A(n7618), .Y(n7616) );
  INVX1 U7562 ( .A(n7616), .Y(n7617) );
  BUFX2 U7563 ( .A(fifo[271]), .Y(n7618) );
  INVX1 U7564 ( .A(n7621), .Y(n7619) );
  INVX1 U7565 ( .A(n7619), .Y(n7620) );
  BUFX2 U7566 ( .A(fifo[578]), .Y(n7621) );
  INVX1 U7567 ( .A(n7624), .Y(n7622) );
  INVX1 U7568 ( .A(n7622), .Y(n7623) );
  BUFX2 U7569 ( .A(fifo[579]), .Y(n7624) );
  INVX1 U7570 ( .A(n7627), .Y(n7625) );
  INVX1 U7571 ( .A(n7625), .Y(n7626) );
  BUFX2 U7572 ( .A(fifo[580]), .Y(n7627) );
  INVX1 U7573 ( .A(n7630), .Y(n7628) );
  INVX1 U7574 ( .A(n7628), .Y(n7629) );
  BUFX2 U7575 ( .A(fifo[581]), .Y(n7630) );
  INVX1 U7576 ( .A(n7633), .Y(n7631) );
  INVX1 U7577 ( .A(n7631), .Y(n7632) );
  BUFX2 U7578 ( .A(fifo[582]), .Y(n7633) );
  INVX1 U7579 ( .A(n7636), .Y(n7634) );
  INVX1 U7580 ( .A(n7634), .Y(n7635) );
  BUFX2 U7581 ( .A(fifo[583]), .Y(n7636) );
  INVX1 U7582 ( .A(n7639), .Y(n7637) );
  INVX1 U7583 ( .A(n7637), .Y(n7638) );
  BUFX2 U7584 ( .A(fifo[584]), .Y(n7639) );
  INVX1 U7585 ( .A(n7642), .Y(n7640) );
  INVX1 U7586 ( .A(n7640), .Y(n7641) );
  BUFX2 U7587 ( .A(fifo[585]), .Y(n7642) );
  INVX1 U7588 ( .A(n7645), .Y(n7643) );
  INVX1 U7589 ( .A(n7643), .Y(n7644) );
  BUFX2 U7590 ( .A(fifo[586]), .Y(n7645) );
  INVX1 U7591 ( .A(n7648), .Y(n7646) );
  INVX1 U7592 ( .A(n7646), .Y(n7647) );
  BUFX2 U7593 ( .A(fifo[587]), .Y(n7648) );
  INVX1 U7594 ( .A(n7651), .Y(n7649) );
  INVX1 U7595 ( .A(n7649), .Y(n7650) );
  BUFX2 U7596 ( .A(fifo[588]), .Y(n7651) );
  INVX1 U7597 ( .A(n7654), .Y(n7652) );
  INVX1 U7598 ( .A(n7652), .Y(n7653) );
  BUFX2 U7599 ( .A(fifo[589]), .Y(n7654) );
  INVX1 U7600 ( .A(n7657), .Y(n7655) );
  INVX1 U7601 ( .A(n7655), .Y(n7656) );
  BUFX2 U7602 ( .A(fifo[590]), .Y(n7657) );
  INVX1 U7603 ( .A(n7660), .Y(n7658) );
  INVX1 U7604 ( .A(n7658), .Y(n7659) );
  BUFX2 U7605 ( .A(fifo[591]), .Y(n7660) );
  INVX1 U7606 ( .A(n7663), .Y(n7661) );
  INVX1 U7607 ( .A(n7661), .Y(n7662) );
  BUFX2 U7608 ( .A(fifo[592]), .Y(n7663) );
  INVX1 U7609 ( .A(n7666), .Y(n7664) );
  INVX1 U7610 ( .A(n7664), .Y(n7665) );
  BUFX2 U7611 ( .A(fifo[593]), .Y(n7666) );
  INVX1 U7612 ( .A(n7669), .Y(n7667) );
  INVX1 U7613 ( .A(n7667), .Y(n7668) );
  BUFX2 U7614 ( .A(fifo[594]), .Y(n7669) );
  INVX1 U7615 ( .A(n7672), .Y(n7670) );
  INVX1 U7616 ( .A(n7670), .Y(n7671) );
  BUFX2 U7617 ( .A(fifo[595]), .Y(n7672) );
  INVX1 U7618 ( .A(n7675), .Y(n7673) );
  INVX1 U7619 ( .A(n7673), .Y(n7674) );
  BUFX2 U7620 ( .A(fifo[596]), .Y(n7675) );
  INVX1 U7621 ( .A(n7678), .Y(n7676) );
  INVX1 U7622 ( .A(n7676), .Y(n7677) );
  BUFX2 U7623 ( .A(fifo[597]), .Y(n7678) );
  INVX1 U7624 ( .A(n7681), .Y(n7679) );
  INVX1 U7625 ( .A(n7679), .Y(n7680) );
  BUFX2 U7626 ( .A(fifo[598]), .Y(n7681) );
  INVX1 U7627 ( .A(n7684), .Y(n7682) );
  INVX1 U7628 ( .A(n7682), .Y(n7683) );
  BUFX2 U7629 ( .A(fifo[599]), .Y(n7684) );
  INVX1 U7630 ( .A(n7687), .Y(n7685) );
  INVX1 U7631 ( .A(n7685), .Y(n7686) );
  BUFX2 U7632 ( .A(fifo[600]), .Y(n7687) );
  INVX1 U7633 ( .A(n7690), .Y(n7688) );
  INVX1 U7634 ( .A(n7688), .Y(n7689) );
  BUFX2 U7635 ( .A(fifo[601]), .Y(n7690) );
  INVX1 U7636 ( .A(n7693), .Y(n7691) );
  INVX1 U7637 ( .A(n7691), .Y(n7692) );
  BUFX2 U7638 ( .A(fifo[602]), .Y(n7693) );
  INVX1 U7639 ( .A(n7696), .Y(n7694) );
  INVX1 U7640 ( .A(n7694), .Y(n7695) );
  BUFX2 U7641 ( .A(fifo[603]), .Y(n7696) );
  INVX1 U7642 ( .A(n7699), .Y(n7697) );
  INVX1 U7643 ( .A(n7697), .Y(n7698) );
  BUFX2 U7644 ( .A(fifo[604]), .Y(n7699) );
  INVX1 U7645 ( .A(n7702), .Y(n7700) );
  INVX1 U7646 ( .A(n7700), .Y(n7701) );
  BUFX2 U7647 ( .A(fifo[605]), .Y(n7702) );
  INVX1 U7648 ( .A(n7705), .Y(n7703) );
  INVX1 U7649 ( .A(n7703), .Y(n7704) );
  BUFX2 U7650 ( .A(fifo[606]), .Y(n7705) );
  INVX1 U7651 ( .A(n7708), .Y(n7706) );
  INVX1 U7652 ( .A(n7706), .Y(n7707) );
  BUFX2 U7653 ( .A(fifo[607]), .Y(n7708) );
  INVX1 U7654 ( .A(n7711), .Y(n7709) );
  INVX1 U7655 ( .A(n7709), .Y(n7710) );
  BUFX2 U7656 ( .A(fifo[608]), .Y(n7711) );
  INVX1 U7657 ( .A(n7714), .Y(n7712) );
  INVX1 U7658 ( .A(n7712), .Y(n7713) );
  BUFX2 U7659 ( .A(fifo[609]), .Y(n7714) );
  INVX1 U7660 ( .A(n7717), .Y(n7715) );
  INVX1 U7661 ( .A(n7715), .Y(n7716) );
  BUFX2 U7662 ( .A(fifo[610]), .Y(n7717) );
  INVX1 U7663 ( .A(n7720), .Y(n7718) );
  INVX1 U7664 ( .A(n7718), .Y(n7719) );
  BUFX2 U7665 ( .A(fifo[611]), .Y(n7720) );
  INVX1 U7666 ( .A(n7723), .Y(n7721) );
  INVX1 U7667 ( .A(n7721), .Y(n7722) );
  BUFX2 U7668 ( .A(fifo[646]), .Y(n7723) );
  INVX1 U7669 ( .A(n7726), .Y(n7724) );
  INVX1 U7670 ( .A(n7724), .Y(n7725) );
  BUFX2 U7671 ( .A(fifo[647]), .Y(n7726) );
  INVX1 U7672 ( .A(n7729), .Y(n7727) );
  INVX1 U7673 ( .A(n7727), .Y(n7728) );
  BUFX2 U7674 ( .A(fifo[648]), .Y(n7729) );
  INVX1 U7675 ( .A(n7732), .Y(n7730) );
  INVX1 U7676 ( .A(n7730), .Y(n7731) );
  BUFX2 U7677 ( .A(fifo[649]), .Y(n7732) );
  INVX1 U7678 ( .A(n7735), .Y(n7733) );
  INVX1 U7679 ( .A(n7733), .Y(n7734) );
  BUFX2 U7680 ( .A(fifo[650]), .Y(n7735) );
  INVX1 U7681 ( .A(n7738), .Y(n7736) );
  INVX1 U7682 ( .A(n7736), .Y(n7737) );
  BUFX2 U7683 ( .A(fifo[651]), .Y(n7738) );
  INVX1 U7684 ( .A(n7741), .Y(n7739) );
  INVX1 U7685 ( .A(n7739), .Y(n7740) );
  BUFX2 U7686 ( .A(fifo[652]), .Y(n7741) );
  INVX1 U7687 ( .A(n7744), .Y(n7742) );
  INVX1 U7688 ( .A(n7742), .Y(n7743) );
  BUFX2 U7689 ( .A(fifo[653]), .Y(n7744) );
  INVX1 U7690 ( .A(n7747), .Y(n7745) );
  INVX1 U7691 ( .A(n7745), .Y(n7746) );
  BUFX2 U7692 ( .A(fifo[654]), .Y(n7747) );
  INVX1 U7693 ( .A(n7750), .Y(n7748) );
  INVX1 U7694 ( .A(n7748), .Y(n7749) );
  BUFX2 U7695 ( .A(fifo[655]), .Y(n7750) );
  INVX1 U7696 ( .A(n7753), .Y(n7751) );
  INVX1 U7697 ( .A(n7751), .Y(n7752) );
  BUFX2 U7698 ( .A(fifo[656]), .Y(n7753) );
  INVX1 U7699 ( .A(n7756), .Y(n7754) );
  INVX1 U7700 ( .A(n7754), .Y(n7755) );
  BUFX2 U7701 ( .A(fifo[657]), .Y(n7756) );
  INVX1 U7702 ( .A(n7759), .Y(n7757) );
  INVX1 U7703 ( .A(n7757), .Y(n7758) );
  BUFX2 U7704 ( .A(fifo[658]), .Y(n7759) );
  INVX1 U7705 ( .A(n7762), .Y(n7760) );
  INVX1 U7706 ( .A(n7760), .Y(n7761) );
  BUFX2 U7707 ( .A(fifo[659]), .Y(n7762) );
  INVX1 U7708 ( .A(n7765), .Y(n7763) );
  INVX1 U7709 ( .A(n7763), .Y(n7764) );
  BUFX2 U7710 ( .A(fifo[660]), .Y(n7765) );
  INVX1 U7711 ( .A(n7768), .Y(n7766) );
  INVX1 U7712 ( .A(n7766), .Y(n7767) );
  BUFX2 U7713 ( .A(fifo[661]), .Y(n7768) );
  INVX1 U7714 ( .A(n7771), .Y(n7769) );
  INVX1 U7715 ( .A(n7769), .Y(n7770) );
  BUFX2 U7716 ( .A(fifo[662]), .Y(n7771) );
  INVX1 U7717 ( .A(n7774), .Y(n7772) );
  INVX1 U7718 ( .A(n7772), .Y(n7773) );
  BUFX2 U7719 ( .A(fifo[663]), .Y(n7774) );
  INVX1 U7720 ( .A(n7777), .Y(n7775) );
  INVX1 U7721 ( .A(n7775), .Y(n7776) );
  BUFX2 U7722 ( .A(fifo[664]), .Y(n7777) );
  INVX1 U7723 ( .A(n7780), .Y(n7778) );
  INVX1 U7724 ( .A(n7778), .Y(n7779) );
  BUFX2 U7725 ( .A(fifo[665]), .Y(n7780) );
  INVX1 U7726 ( .A(n7783), .Y(n7781) );
  INVX1 U7727 ( .A(n7781), .Y(n7782) );
  BUFX2 U7728 ( .A(fifo[666]), .Y(n7783) );
  INVX1 U7729 ( .A(n7786), .Y(n7784) );
  INVX1 U7730 ( .A(n7784), .Y(n7785) );
  BUFX2 U7731 ( .A(fifo[667]), .Y(n7786) );
  INVX1 U7732 ( .A(n7789), .Y(n7787) );
  INVX1 U7733 ( .A(n7787), .Y(n7788) );
  BUFX2 U7734 ( .A(fifo[668]), .Y(n7789) );
  INVX1 U7735 ( .A(n7792), .Y(n7790) );
  INVX1 U7736 ( .A(n7790), .Y(n7791) );
  BUFX2 U7737 ( .A(fifo[669]), .Y(n7792) );
  INVX1 U7738 ( .A(n7795), .Y(n7793) );
  INVX1 U7739 ( .A(n7793), .Y(n7794) );
  BUFX2 U7740 ( .A(fifo[670]), .Y(n7795) );
  INVX1 U7741 ( .A(n7798), .Y(n7796) );
  INVX1 U7742 ( .A(n7796), .Y(n7797) );
  BUFX2 U7743 ( .A(fifo[671]), .Y(n7798) );
  INVX1 U7744 ( .A(n7801), .Y(n7799) );
  INVX1 U7745 ( .A(n7799), .Y(n7800) );
  BUFX2 U7746 ( .A(fifo[672]), .Y(n7801) );
  INVX1 U7747 ( .A(n7804), .Y(n7802) );
  INVX1 U7748 ( .A(n7802), .Y(n7803) );
  BUFX2 U7749 ( .A(fifo[673]), .Y(n7804) );
  INVX1 U7750 ( .A(n7807), .Y(n7805) );
  INVX1 U7751 ( .A(n7805), .Y(n7806) );
  BUFX2 U7752 ( .A(fifo[674]), .Y(n7807) );
  INVX1 U7753 ( .A(n7810), .Y(n7808) );
  INVX1 U7754 ( .A(n7808), .Y(n7809) );
  BUFX2 U7755 ( .A(fifo[675]), .Y(n7810) );
  INVX1 U7756 ( .A(n7813), .Y(n7811) );
  INVX1 U7757 ( .A(n7811), .Y(n7812) );
  BUFX2 U7758 ( .A(fifo[676]), .Y(n7813) );
  INVX1 U7759 ( .A(n7816), .Y(n7814) );
  INVX1 U7760 ( .A(n7814), .Y(n7815) );
  BUFX2 U7761 ( .A(fifo[677]), .Y(n7816) );
  INVX1 U7762 ( .A(n7819), .Y(n7817) );
  INVX1 U7763 ( .A(n7817), .Y(n7818) );
  BUFX2 U7764 ( .A(fifo[678]), .Y(n7819) );
  INVX1 U7765 ( .A(n7822), .Y(n7820) );
  INVX1 U7766 ( .A(n7820), .Y(n7821) );
  BUFX2 U7767 ( .A(fifo[679]), .Y(n7822) );
  INVX1 U7768 ( .A(n7825), .Y(n7823) );
  INVX1 U7769 ( .A(n7823), .Y(n7824) );
  BUFX2 U7770 ( .A(fifo[714]), .Y(n7825) );
  INVX1 U7771 ( .A(n7828), .Y(n7826) );
  INVX1 U7772 ( .A(n7826), .Y(n7827) );
  BUFX2 U7773 ( .A(fifo[715]), .Y(n7828) );
  INVX1 U7774 ( .A(n7831), .Y(n7829) );
  INVX1 U7775 ( .A(n7829), .Y(n7830) );
  BUFX2 U7776 ( .A(fifo[716]), .Y(n7831) );
  INVX1 U7777 ( .A(n7834), .Y(n7832) );
  INVX1 U7778 ( .A(n7832), .Y(n7833) );
  BUFX2 U7779 ( .A(fifo[717]), .Y(n7834) );
  INVX1 U7780 ( .A(n7837), .Y(n7835) );
  INVX1 U7781 ( .A(n7835), .Y(n7836) );
  BUFX2 U7782 ( .A(fifo[718]), .Y(n7837) );
  INVX1 U7783 ( .A(n7840), .Y(n7838) );
  INVX1 U7784 ( .A(n7838), .Y(n7839) );
  BUFX2 U7785 ( .A(fifo[719]), .Y(n7840) );
  INVX1 U7786 ( .A(n7843), .Y(n7841) );
  INVX1 U7787 ( .A(n7841), .Y(n7842) );
  BUFX2 U7788 ( .A(fifo[720]), .Y(n7843) );
  INVX1 U7789 ( .A(n7846), .Y(n7844) );
  INVX1 U7790 ( .A(n7844), .Y(n7845) );
  BUFX2 U7791 ( .A(fifo[721]), .Y(n7846) );
  INVX1 U7792 ( .A(n7849), .Y(n7847) );
  INVX1 U7793 ( .A(n7847), .Y(n7848) );
  BUFX2 U7794 ( .A(fifo[722]), .Y(n7849) );
  INVX1 U7795 ( .A(n7852), .Y(n7850) );
  INVX1 U7796 ( .A(n7850), .Y(n7851) );
  BUFX2 U7797 ( .A(fifo[723]), .Y(n7852) );
  INVX1 U7798 ( .A(n7855), .Y(n7853) );
  INVX1 U7799 ( .A(n7853), .Y(n7854) );
  BUFX2 U7800 ( .A(fifo[724]), .Y(n7855) );
  INVX1 U7801 ( .A(n7858), .Y(n7856) );
  INVX1 U7802 ( .A(n7856), .Y(n7857) );
  BUFX2 U7803 ( .A(fifo[725]), .Y(n7858) );
  INVX1 U7804 ( .A(n7861), .Y(n7859) );
  INVX1 U7805 ( .A(n7859), .Y(n7860) );
  BUFX2 U7806 ( .A(fifo[726]), .Y(n7861) );
  INVX1 U7807 ( .A(n7864), .Y(n7862) );
  INVX1 U7808 ( .A(n7862), .Y(n7863) );
  BUFX2 U7809 ( .A(fifo[727]), .Y(n7864) );
  INVX1 U7810 ( .A(n7867), .Y(n7865) );
  INVX1 U7811 ( .A(n7865), .Y(n7866) );
  BUFX2 U7812 ( .A(fifo[728]), .Y(n7867) );
  INVX1 U7813 ( .A(n7870), .Y(n7868) );
  INVX1 U7814 ( .A(n7868), .Y(n7869) );
  BUFX2 U7815 ( .A(fifo[729]), .Y(n7870) );
  INVX1 U7816 ( .A(n7873), .Y(n7871) );
  INVX1 U7817 ( .A(n7871), .Y(n7872) );
  BUFX2 U7818 ( .A(fifo[730]), .Y(n7873) );
  INVX1 U7819 ( .A(n7876), .Y(n7874) );
  INVX1 U7820 ( .A(n7874), .Y(n7875) );
  BUFX2 U7821 ( .A(fifo[731]), .Y(n7876) );
  INVX1 U7822 ( .A(n7879), .Y(n7877) );
  INVX1 U7823 ( .A(n7877), .Y(n7878) );
  BUFX2 U7824 ( .A(fifo[732]), .Y(n7879) );
  INVX1 U7825 ( .A(n7882), .Y(n7880) );
  INVX1 U7826 ( .A(n7880), .Y(n7881) );
  BUFX2 U7827 ( .A(fifo[733]), .Y(n7882) );
  INVX1 U7828 ( .A(n7885), .Y(n7883) );
  INVX1 U7829 ( .A(n7883), .Y(n7884) );
  BUFX2 U7830 ( .A(fifo[734]), .Y(n7885) );
  INVX1 U7831 ( .A(n7888), .Y(n7886) );
  INVX1 U7832 ( .A(n7886), .Y(n7887) );
  BUFX2 U7833 ( .A(fifo[735]), .Y(n7888) );
  INVX1 U7834 ( .A(n7891), .Y(n7889) );
  INVX1 U7835 ( .A(n7889), .Y(n7890) );
  BUFX2 U7836 ( .A(fifo[736]), .Y(n7891) );
  INVX1 U7837 ( .A(n7894), .Y(n7892) );
  INVX1 U7838 ( .A(n7892), .Y(n7893) );
  BUFX2 U7839 ( .A(fifo[737]), .Y(n7894) );
  INVX1 U7840 ( .A(n7897), .Y(n7895) );
  INVX1 U7841 ( .A(n7895), .Y(n7896) );
  BUFX2 U7842 ( .A(fifo[738]), .Y(n7897) );
  INVX1 U7843 ( .A(n7900), .Y(n7898) );
  INVX1 U7844 ( .A(n7898), .Y(n7899) );
  BUFX2 U7845 ( .A(fifo[739]), .Y(n7900) );
  INVX1 U7846 ( .A(n7903), .Y(n7901) );
  INVX1 U7847 ( .A(n7901), .Y(n7902) );
  BUFX2 U7848 ( .A(fifo[740]), .Y(n7903) );
  INVX1 U7849 ( .A(n7906), .Y(n7904) );
  INVX1 U7850 ( .A(n7904), .Y(n7905) );
  BUFX2 U7851 ( .A(fifo[741]), .Y(n7906) );
  INVX1 U7852 ( .A(n7909), .Y(n7907) );
  INVX1 U7853 ( .A(n7907), .Y(n7908) );
  BUFX2 U7854 ( .A(fifo[742]), .Y(n7909) );
  INVX1 U7855 ( .A(n7912), .Y(n7910) );
  INVX1 U7856 ( .A(n7910), .Y(n7911) );
  BUFX2 U7857 ( .A(fifo[743]), .Y(n7912) );
  INVX1 U7858 ( .A(n7915), .Y(n7913) );
  INVX1 U7859 ( .A(n7913), .Y(n7914) );
  BUFX2 U7860 ( .A(fifo[744]), .Y(n7915) );
  INVX1 U7861 ( .A(n7918), .Y(n7916) );
  INVX1 U7862 ( .A(n7916), .Y(n7917) );
  BUFX2 U7863 ( .A(fifo[745]), .Y(n7918) );
  INVX1 U7864 ( .A(n7921), .Y(n7919) );
  INVX1 U7865 ( .A(n7919), .Y(n7920) );
  BUFX2 U7866 ( .A(fifo[746]), .Y(n7921) );
  INVX1 U7867 ( .A(n7924), .Y(n7922) );
  INVX1 U7868 ( .A(n7922), .Y(n7923) );
  BUFX2 U7869 ( .A(fifo[747]), .Y(n7924) );
  INVX1 U7870 ( .A(n7927), .Y(n7925) );
  INVX1 U7871 ( .A(n7925), .Y(n7926) );
  BUFX2 U7872 ( .A(fifo[782]), .Y(n7927) );
  INVX1 U7873 ( .A(n7930), .Y(n7928) );
  INVX1 U7874 ( .A(n7928), .Y(n7929) );
  BUFX2 U7875 ( .A(fifo[783]), .Y(n7930) );
  INVX1 U7876 ( .A(n7933), .Y(n7931) );
  INVX1 U7877 ( .A(n7931), .Y(n7932) );
  BUFX2 U7878 ( .A(fifo[784]), .Y(n7933) );
  INVX1 U7879 ( .A(n7936), .Y(n7934) );
  INVX1 U7880 ( .A(n7934), .Y(n7935) );
  BUFX2 U7881 ( .A(fifo[785]), .Y(n7936) );
  INVX1 U7882 ( .A(n7939), .Y(n7937) );
  INVX1 U7883 ( .A(n7937), .Y(n7938) );
  BUFX2 U7884 ( .A(fifo[786]), .Y(n7939) );
  INVX1 U7885 ( .A(n7942), .Y(n7940) );
  INVX1 U7886 ( .A(n7940), .Y(n7941) );
  BUFX2 U7887 ( .A(fifo[787]), .Y(n7942) );
  INVX1 U7888 ( .A(n7945), .Y(n7943) );
  INVX1 U7889 ( .A(n7943), .Y(n7944) );
  BUFX2 U7890 ( .A(fifo[788]), .Y(n7945) );
  INVX1 U7891 ( .A(n7948), .Y(n7946) );
  INVX1 U7892 ( .A(n7946), .Y(n7947) );
  BUFX2 U7893 ( .A(fifo[789]), .Y(n7948) );
  INVX1 U7894 ( .A(n7951), .Y(n7949) );
  INVX1 U7895 ( .A(n7949), .Y(n7950) );
  BUFX2 U7896 ( .A(fifo[790]), .Y(n7951) );
  INVX1 U7897 ( .A(n7954), .Y(n7952) );
  INVX1 U7898 ( .A(n7952), .Y(n7953) );
  BUFX2 U7899 ( .A(fifo[791]), .Y(n7954) );
  INVX1 U7900 ( .A(n7957), .Y(n7955) );
  INVX1 U7901 ( .A(n7955), .Y(n7956) );
  BUFX2 U7902 ( .A(fifo[792]), .Y(n7957) );
  INVX1 U7903 ( .A(n7960), .Y(n7958) );
  INVX1 U7904 ( .A(n7958), .Y(n7959) );
  BUFX2 U7905 ( .A(fifo[793]), .Y(n7960) );
  INVX1 U7906 ( .A(n7963), .Y(n7961) );
  INVX1 U7907 ( .A(n7961), .Y(n7962) );
  BUFX2 U7908 ( .A(fifo[794]), .Y(n7963) );
  INVX1 U7909 ( .A(n7966), .Y(n7964) );
  INVX1 U7910 ( .A(n7964), .Y(n7965) );
  BUFX2 U7911 ( .A(fifo[795]), .Y(n7966) );
  INVX1 U7912 ( .A(n7969), .Y(n7967) );
  INVX1 U7913 ( .A(n7967), .Y(n7968) );
  BUFX2 U7914 ( .A(fifo[796]), .Y(n7969) );
  INVX1 U7915 ( .A(n7972), .Y(n7970) );
  INVX1 U7916 ( .A(n7970), .Y(n7971) );
  BUFX2 U7917 ( .A(fifo[797]), .Y(n7972) );
  INVX1 U7918 ( .A(n7975), .Y(n7973) );
  INVX1 U7919 ( .A(n7973), .Y(n7974) );
  BUFX2 U7920 ( .A(fifo[798]), .Y(n7975) );
  INVX1 U7921 ( .A(n7978), .Y(n7976) );
  INVX1 U7922 ( .A(n7976), .Y(n7977) );
  BUFX2 U7923 ( .A(fifo[799]), .Y(n7978) );
  INVX1 U7924 ( .A(n7981), .Y(n7979) );
  INVX1 U7925 ( .A(n7979), .Y(n7980) );
  BUFX2 U7926 ( .A(fifo[800]), .Y(n7981) );
  INVX1 U7927 ( .A(n7984), .Y(n7982) );
  INVX1 U7928 ( .A(n7982), .Y(n7983) );
  BUFX2 U7929 ( .A(fifo[801]), .Y(n7984) );
  INVX1 U7930 ( .A(n7987), .Y(n7985) );
  INVX1 U7931 ( .A(n7985), .Y(n7986) );
  BUFX2 U7932 ( .A(fifo[802]), .Y(n7987) );
  INVX1 U7933 ( .A(n7990), .Y(n7988) );
  INVX1 U7934 ( .A(n7988), .Y(n7989) );
  BUFX2 U7935 ( .A(fifo[803]), .Y(n7990) );
  INVX1 U7936 ( .A(n7993), .Y(n7991) );
  INVX1 U7937 ( .A(n7991), .Y(n7992) );
  BUFX2 U7938 ( .A(fifo[804]), .Y(n7993) );
  INVX1 U7939 ( .A(n7996), .Y(n7994) );
  INVX1 U7940 ( .A(n7994), .Y(n7995) );
  BUFX2 U7941 ( .A(fifo[805]), .Y(n7996) );
  INVX1 U7942 ( .A(n7999), .Y(n7997) );
  INVX1 U7943 ( .A(n7997), .Y(n7998) );
  BUFX2 U7944 ( .A(fifo[806]), .Y(n7999) );
  INVX1 U7945 ( .A(n8002), .Y(n8000) );
  INVX1 U7946 ( .A(n8000), .Y(n8001) );
  BUFX2 U7947 ( .A(fifo[807]), .Y(n8002) );
  INVX1 U7948 ( .A(n8005), .Y(n8003) );
  INVX1 U7949 ( .A(n8003), .Y(n8004) );
  BUFX2 U7950 ( .A(fifo[808]), .Y(n8005) );
  INVX1 U7951 ( .A(n8008), .Y(n8006) );
  INVX1 U7952 ( .A(n8006), .Y(n8007) );
  BUFX2 U7953 ( .A(fifo[809]), .Y(n8008) );
  INVX1 U7954 ( .A(n8011), .Y(n8009) );
  INVX1 U7955 ( .A(n8009), .Y(n8010) );
  BUFX2 U7956 ( .A(fifo[810]), .Y(n8011) );
  INVX1 U7957 ( .A(n8014), .Y(n8012) );
  INVX1 U7958 ( .A(n8012), .Y(n8013) );
  BUFX2 U7959 ( .A(fifo[811]), .Y(n8014) );
  INVX1 U7960 ( .A(n8017), .Y(n8015) );
  INVX1 U7961 ( .A(n8015), .Y(n8016) );
  BUFX2 U7962 ( .A(fifo[812]), .Y(n8017) );
  INVX1 U7963 ( .A(n8020), .Y(n8018) );
  INVX1 U7964 ( .A(n8018), .Y(n8019) );
  BUFX2 U7965 ( .A(fifo[813]), .Y(n8020) );
  INVX1 U7966 ( .A(n8023), .Y(n8021) );
  INVX1 U7967 ( .A(n8021), .Y(n8022) );
  BUFX2 U7968 ( .A(fifo[814]), .Y(n8023) );
  INVX1 U7969 ( .A(n8026), .Y(n8024) );
  INVX1 U7970 ( .A(n8024), .Y(n8025) );
  BUFX2 U7971 ( .A(fifo[815]), .Y(n8026) );
  INVX1 U7972 ( .A(n8029), .Y(n8027) );
  INVX1 U7973 ( .A(n8027), .Y(n8028) );
  BUFX2 U7974 ( .A(fifo[850]), .Y(n8029) );
  INVX1 U7975 ( .A(n8032), .Y(n8030) );
  INVX1 U7976 ( .A(n8030), .Y(n8031) );
  BUFX2 U7977 ( .A(fifo[851]), .Y(n8032) );
  INVX1 U7978 ( .A(n8035), .Y(n8033) );
  INVX1 U7979 ( .A(n8033), .Y(n8034) );
  BUFX2 U7980 ( .A(fifo[852]), .Y(n8035) );
  INVX1 U7981 ( .A(n8038), .Y(n8036) );
  INVX1 U7982 ( .A(n8036), .Y(n8037) );
  BUFX2 U7983 ( .A(fifo[853]), .Y(n8038) );
  INVX1 U7984 ( .A(n8041), .Y(n8039) );
  INVX1 U7985 ( .A(n8039), .Y(n8040) );
  BUFX2 U7986 ( .A(fifo[854]), .Y(n8041) );
  INVX1 U7987 ( .A(n8044), .Y(n8042) );
  INVX1 U7988 ( .A(n8042), .Y(n8043) );
  BUFX2 U7989 ( .A(fifo[855]), .Y(n8044) );
  INVX1 U7990 ( .A(n8047), .Y(n8045) );
  INVX1 U7991 ( .A(n8045), .Y(n8046) );
  BUFX2 U7992 ( .A(fifo[856]), .Y(n8047) );
  INVX1 U7993 ( .A(n8050), .Y(n8048) );
  INVX1 U7994 ( .A(n8048), .Y(n8049) );
  BUFX2 U7995 ( .A(fifo[857]), .Y(n8050) );
  INVX1 U7996 ( .A(n8053), .Y(n8051) );
  INVX1 U7997 ( .A(n8051), .Y(n8052) );
  BUFX2 U7998 ( .A(fifo[858]), .Y(n8053) );
  INVX1 U7999 ( .A(n8056), .Y(n8054) );
  INVX1 U8000 ( .A(n8054), .Y(n8055) );
  BUFX2 U8001 ( .A(fifo[859]), .Y(n8056) );
  INVX1 U8002 ( .A(n8059), .Y(n8057) );
  INVX1 U8003 ( .A(n8057), .Y(n8058) );
  BUFX2 U8004 ( .A(fifo[860]), .Y(n8059) );
  INVX1 U8005 ( .A(n8062), .Y(n8060) );
  INVX1 U8006 ( .A(n8060), .Y(n8061) );
  BUFX2 U8007 ( .A(fifo[861]), .Y(n8062) );
  INVX1 U8008 ( .A(n8065), .Y(n8063) );
  INVX1 U8009 ( .A(n8063), .Y(n8064) );
  BUFX2 U8010 ( .A(fifo[862]), .Y(n8065) );
  INVX1 U8011 ( .A(n8068), .Y(n8066) );
  INVX1 U8012 ( .A(n8066), .Y(n8067) );
  BUFX2 U8013 ( .A(fifo[863]), .Y(n8068) );
  INVX1 U8014 ( .A(n8071), .Y(n8069) );
  INVX1 U8015 ( .A(n8069), .Y(n8070) );
  BUFX2 U8016 ( .A(fifo[864]), .Y(n8071) );
  INVX1 U8017 ( .A(n8074), .Y(n8072) );
  INVX1 U8018 ( .A(n8072), .Y(n8073) );
  BUFX2 U8019 ( .A(fifo[865]), .Y(n8074) );
  INVX1 U8020 ( .A(n8077), .Y(n8075) );
  INVX1 U8021 ( .A(n8075), .Y(n8076) );
  BUFX2 U8022 ( .A(fifo[866]), .Y(n8077) );
  INVX1 U8023 ( .A(n8080), .Y(n8078) );
  INVX1 U8024 ( .A(n8078), .Y(n8079) );
  BUFX2 U8025 ( .A(fifo[867]), .Y(n8080) );
  INVX1 U8026 ( .A(n8083), .Y(n8081) );
  INVX1 U8027 ( .A(n8081), .Y(n8082) );
  BUFX2 U8028 ( .A(fifo[868]), .Y(n8083) );
  INVX1 U8029 ( .A(n8086), .Y(n8084) );
  INVX1 U8030 ( .A(n8084), .Y(n8085) );
  BUFX2 U8031 ( .A(fifo[869]), .Y(n8086) );
  INVX1 U8032 ( .A(n8089), .Y(n8087) );
  INVX1 U8033 ( .A(n8087), .Y(n8088) );
  BUFX2 U8034 ( .A(fifo[870]), .Y(n8089) );
  INVX1 U8035 ( .A(n8092), .Y(n8090) );
  INVX1 U8036 ( .A(n8090), .Y(n8091) );
  BUFX2 U8037 ( .A(fifo[871]), .Y(n8092) );
  INVX1 U8038 ( .A(n8095), .Y(n8093) );
  INVX1 U8039 ( .A(n8093), .Y(n8094) );
  BUFX2 U8040 ( .A(fifo[872]), .Y(n8095) );
  INVX1 U8041 ( .A(n8098), .Y(n8096) );
  INVX1 U8042 ( .A(n8096), .Y(n8097) );
  BUFX2 U8043 ( .A(fifo[873]), .Y(n8098) );
  INVX1 U8044 ( .A(n8101), .Y(n8099) );
  INVX1 U8045 ( .A(n8099), .Y(n8100) );
  BUFX2 U8046 ( .A(fifo[874]), .Y(n8101) );
  INVX1 U8047 ( .A(n8104), .Y(n8102) );
  INVX1 U8048 ( .A(n8102), .Y(n8103) );
  BUFX2 U8049 ( .A(fifo[875]), .Y(n8104) );
  INVX1 U8050 ( .A(n8107), .Y(n8105) );
  INVX1 U8051 ( .A(n8105), .Y(n8106) );
  BUFX2 U8052 ( .A(fifo[876]), .Y(n8107) );
  INVX1 U8053 ( .A(n8110), .Y(n8108) );
  INVX1 U8054 ( .A(n8108), .Y(n8109) );
  BUFX2 U8055 ( .A(fifo[877]), .Y(n8110) );
  INVX1 U8056 ( .A(n8113), .Y(n8111) );
  INVX1 U8057 ( .A(n8111), .Y(n8112) );
  BUFX2 U8058 ( .A(fifo[878]), .Y(n8113) );
  INVX1 U8059 ( .A(n8116), .Y(n8114) );
  INVX1 U8060 ( .A(n8114), .Y(n8115) );
  BUFX2 U8061 ( .A(fifo[879]), .Y(n8116) );
  INVX1 U8062 ( .A(n8119), .Y(n8117) );
  INVX1 U8063 ( .A(n8117), .Y(n8118) );
  BUFX2 U8064 ( .A(fifo[880]), .Y(n8119) );
  INVX1 U8065 ( .A(n8122), .Y(n8120) );
  INVX1 U8066 ( .A(n8120), .Y(n8121) );
  BUFX2 U8067 ( .A(fifo[881]), .Y(n8122) );
  INVX1 U8068 ( .A(n8125), .Y(n8123) );
  INVX1 U8069 ( .A(n8123), .Y(n8124) );
  BUFX2 U8070 ( .A(fifo[882]), .Y(n8125) );
  INVX1 U8071 ( .A(n8128), .Y(n8126) );
  INVX1 U8072 ( .A(n8126), .Y(n8127) );
  BUFX2 U8073 ( .A(fifo[883]), .Y(n8128) );
  INVX1 U8074 ( .A(n8131), .Y(n8129) );
  INVX1 U8075 ( .A(n8129), .Y(n8130) );
  BUFX2 U8076 ( .A(fifo[918]), .Y(n8131) );
  INVX1 U8077 ( .A(n8134), .Y(n8132) );
  INVX1 U8078 ( .A(n8132), .Y(n8133) );
  BUFX2 U8079 ( .A(fifo[919]), .Y(n8134) );
  INVX1 U8080 ( .A(n8137), .Y(n8135) );
  INVX1 U8081 ( .A(n8135), .Y(n8136) );
  BUFX2 U8082 ( .A(fifo[920]), .Y(n8137) );
  INVX1 U8083 ( .A(n8140), .Y(n8138) );
  INVX1 U8084 ( .A(n8138), .Y(n8139) );
  BUFX2 U8085 ( .A(fifo[921]), .Y(n8140) );
  INVX1 U8086 ( .A(n8143), .Y(n8141) );
  INVX1 U8087 ( .A(n8141), .Y(n8142) );
  BUFX2 U8088 ( .A(fifo[922]), .Y(n8143) );
  INVX1 U8089 ( .A(n8146), .Y(n8144) );
  INVX1 U8090 ( .A(n8144), .Y(n8145) );
  BUFX2 U8091 ( .A(fifo[923]), .Y(n8146) );
  INVX1 U8092 ( .A(n8149), .Y(n8147) );
  INVX1 U8093 ( .A(n8147), .Y(n8148) );
  BUFX2 U8094 ( .A(fifo[924]), .Y(n8149) );
  INVX1 U8095 ( .A(n8152), .Y(n8150) );
  INVX1 U8096 ( .A(n8150), .Y(n8151) );
  BUFX2 U8097 ( .A(fifo[925]), .Y(n8152) );
  INVX1 U8098 ( .A(n8155), .Y(n8153) );
  INVX1 U8099 ( .A(n8153), .Y(n8154) );
  BUFX2 U8100 ( .A(fifo[926]), .Y(n8155) );
  INVX1 U8101 ( .A(n8158), .Y(n8156) );
  INVX1 U8102 ( .A(n8156), .Y(n8157) );
  BUFX2 U8103 ( .A(fifo[927]), .Y(n8158) );
  INVX1 U8104 ( .A(n8161), .Y(n8159) );
  INVX1 U8105 ( .A(n8159), .Y(n8160) );
  BUFX2 U8106 ( .A(fifo[928]), .Y(n8161) );
  INVX1 U8107 ( .A(n8164), .Y(n8162) );
  INVX1 U8108 ( .A(n8162), .Y(n8163) );
  BUFX2 U8109 ( .A(fifo[929]), .Y(n8164) );
  INVX1 U8110 ( .A(n8167), .Y(n8165) );
  INVX1 U8111 ( .A(n8165), .Y(n8166) );
  BUFX2 U8112 ( .A(fifo[930]), .Y(n8167) );
  INVX1 U8113 ( .A(n8170), .Y(n8168) );
  INVX1 U8114 ( .A(n8168), .Y(n8169) );
  BUFX2 U8115 ( .A(fifo[931]), .Y(n8170) );
  INVX1 U8116 ( .A(n8173), .Y(n8171) );
  INVX1 U8117 ( .A(n8171), .Y(n8172) );
  BUFX2 U8118 ( .A(fifo[932]), .Y(n8173) );
  INVX1 U8119 ( .A(n8176), .Y(n8174) );
  INVX1 U8120 ( .A(n8174), .Y(n8175) );
  BUFX2 U8121 ( .A(fifo[933]), .Y(n8176) );
  INVX1 U8122 ( .A(n8179), .Y(n8177) );
  INVX1 U8123 ( .A(n8177), .Y(n8178) );
  BUFX2 U8124 ( .A(fifo[934]), .Y(n8179) );
  INVX1 U8125 ( .A(n8182), .Y(n8180) );
  INVX1 U8126 ( .A(n8180), .Y(n8181) );
  BUFX2 U8127 ( .A(fifo[935]), .Y(n8182) );
  INVX1 U8128 ( .A(n8185), .Y(n8183) );
  INVX1 U8129 ( .A(n8183), .Y(n8184) );
  BUFX2 U8130 ( .A(fifo[936]), .Y(n8185) );
  INVX1 U8131 ( .A(n8188), .Y(n8186) );
  INVX1 U8132 ( .A(n8186), .Y(n8187) );
  BUFX2 U8133 ( .A(fifo[937]), .Y(n8188) );
  INVX1 U8134 ( .A(n8191), .Y(n8189) );
  INVX1 U8135 ( .A(n8189), .Y(n8190) );
  BUFX2 U8136 ( .A(fifo[938]), .Y(n8191) );
  INVX1 U8137 ( .A(n8194), .Y(n8192) );
  INVX1 U8138 ( .A(n8192), .Y(n8193) );
  BUFX2 U8139 ( .A(fifo[939]), .Y(n8194) );
  INVX1 U8140 ( .A(n8197), .Y(n8195) );
  INVX1 U8141 ( .A(n8195), .Y(n8196) );
  BUFX2 U8142 ( .A(fifo[940]), .Y(n8197) );
  INVX1 U8143 ( .A(n8200), .Y(n8198) );
  INVX1 U8144 ( .A(n8198), .Y(n8199) );
  BUFX2 U8145 ( .A(fifo[941]), .Y(n8200) );
  INVX1 U8146 ( .A(n8203), .Y(n8201) );
  INVX1 U8147 ( .A(n8201), .Y(n8202) );
  BUFX2 U8148 ( .A(fifo[942]), .Y(n8203) );
  INVX1 U8149 ( .A(n8206), .Y(n8204) );
  INVX1 U8150 ( .A(n8204), .Y(n8205) );
  BUFX2 U8151 ( .A(fifo[943]), .Y(n8206) );
  INVX1 U8152 ( .A(n8209), .Y(n8207) );
  INVX1 U8153 ( .A(n8207), .Y(n8208) );
  BUFX2 U8154 ( .A(fifo[944]), .Y(n8209) );
  INVX1 U8155 ( .A(n8212), .Y(n8210) );
  INVX1 U8156 ( .A(n8210), .Y(n8211) );
  BUFX2 U8157 ( .A(fifo[945]), .Y(n8212) );
  INVX1 U8158 ( .A(n8215), .Y(n8213) );
  INVX1 U8159 ( .A(n8213), .Y(n8214) );
  BUFX2 U8160 ( .A(fifo[946]), .Y(n8215) );
  INVX1 U8161 ( .A(n8218), .Y(n8216) );
  INVX1 U8162 ( .A(n8216), .Y(n8217) );
  BUFX2 U8163 ( .A(fifo[947]), .Y(n8218) );
  INVX1 U8164 ( .A(n8221), .Y(n8219) );
  INVX1 U8165 ( .A(n8219), .Y(n8220) );
  BUFX2 U8166 ( .A(fifo[948]), .Y(n8221) );
  INVX1 U8167 ( .A(n8224), .Y(n8222) );
  INVX1 U8168 ( .A(n8222), .Y(n8223) );
  BUFX2 U8169 ( .A(fifo[949]), .Y(n8224) );
  INVX1 U8170 ( .A(n8227), .Y(n8225) );
  INVX1 U8171 ( .A(n8225), .Y(n8226) );
  BUFX2 U8172 ( .A(fifo[950]), .Y(n8227) );
  INVX1 U8173 ( .A(n8230), .Y(n8228) );
  INVX1 U8174 ( .A(n8228), .Y(n8229) );
  BUFX2 U8175 ( .A(fifo[951]), .Y(n8230) );
  INVX1 U8176 ( .A(n8233), .Y(n8231) );
  INVX1 U8177 ( .A(n8231), .Y(n8232) );
  BUFX2 U8178 ( .A(fifo[986]), .Y(n8233) );
  INVX1 U8179 ( .A(n8236), .Y(n8234) );
  INVX1 U8180 ( .A(n8234), .Y(n8235) );
  BUFX2 U8181 ( .A(fifo[987]), .Y(n8236) );
  INVX1 U8182 ( .A(n8239), .Y(n8237) );
  INVX1 U8183 ( .A(n8237), .Y(n8238) );
  BUFX2 U8184 ( .A(fifo[988]), .Y(n8239) );
  INVX1 U8185 ( .A(n8242), .Y(n8240) );
  INVX1 U8186 ( .A(n8240), .Y(n8241) );
  BUFX2 U8187 ( .A(fifo[989]), .Y(n8242) );
  INVX1 U8188 ( .A(n8245), .Y(n8243) );
  INVX1 U8189 ( .A(n8243), .Y(n8244) );
  BUFX2 U8190 ( .A(fifo[990]), .Y(n8245) );
  INVX1 U8191 ( .A(n8248), .Y(n8246) );
  INVX1 U8192 ( .A(n8246), .Y(n8247) );
  BUFX2 U8193 ( .A(fifo[991]), .Y(n8248) );
  INVX1 U8194 ( .A(n8251), .Y(n8249) );
  INVX1 U8195 ( .A(n8249), .Y(n8250) );
  BUFX2 U8196 ( .A(fifo[992]), .Y(n8251) );
  INVX1 U8197 ( .A(n8254), .Y(n8252) );
  INVX1 U8198 ( .A(n8252), .Y(n8253) );
  BUFX2 U8199 ( .A(fifo[993]), .Y(n8254) );
  INVX1 U8200 ( .A(n8257), .Y(n8255) );
  INVX1 U8201 ( .A(n8255), .Y(n8256) );
  BUFX2 U8202 ( .A(fifo[994]), .Y(n8257) );
  INVX1 U8203 ( .A(n8260), .Y(n8258) );
  INVX1 U8204 ( .A(n8258), .Y(n8259) );
  BUFX2 U8205 ( .A(fifo[995]), .Y(n8260) );
  INVX1 U8206 ( .A(n8263), .Y(n8261) );
  INVX1 U8207 ( .A(n8261), .Y(n8262) );
  BUFX2 U8208 ( .A(fifo[996]), .Y(n8263) );
  INVX1 U8209 ( .A(n8266), .Y(n8264) );
  INVX1 U8210 ( .A(n8264), .Y(n8265) );
  BUFX2 U8211 ( .A(fifo[997]), .Y(n8266) );
  INVX1 U8212 ( .A(n8269), .Y(n8267) );
  INVX1 U8213 ( .A(n8267), .Y(n8268) );
  BUFX2 U8214 ( .A(fifo[998]), .Y(n8269) );
  INVX1 U8215 ( .A(n8272), .Y(n8270) );
  INVX1 U8216 ( .A(n8270), .Y(n8271) );
  BUFX2 U8217 ( .A(fifo[999]), .Y(n8272) );
  INVX1 U8218 ( .A(n8275), .Y(n8273) );
  INVX1 U8219 ( .A(n8273), .Y(n8274) );
  BUFX2 U8220 ( .A(fifo[1000]), .Y(n8275) );
  INVX1 U8221 ( .A(n8278), .Y(n8276) );
  INVX1 U8222 ( .A(n8276), .Y(n8277) );
  BUFX2 U8223 ( .A(fifo[1001]), .Y(n8278) );
  INVX1 U8224 ( .A(n8281), .Y(n8279) );
  INVX1 U8225 ( .A(n8279), .Y(n8280) );
  BUFX2 U8226 ( .A(fifo[1002]), .Y(n8281) );
  INVX1 U8227 ( .A(n8284), .Y(n8282) );
  INVX1 U8228 ( .A(n8282), .Y(n8283) );
  BUFX2 U8229 ( .A(fifo[1003]), .Y(n8284) );
  INVX1 U8230 ( .A(n8287), .Y(n8285) );
  INVX1 U8231 ( .A(n8285), .Y(n8286) );
  BUFX2 U8232 ( .A(fifo[1004]), .Y(n8287) );
  INVX1 U8233 ( .A(n8290), .Y(n8288) );
  INVX1 U8234 ( .A(n8288), .Y(n8289) );
  BUFX2 U8235 ( .A(fifo[1005]), .Y(n8290) );
  INVX1 U8236 ( .A(n8293), .Y(n8291) );
  INVX1 U8237 ( .A(n8291), .Y(n8292) );
  BUFX2 U8238 ( .A(fifo[1006]), .Y(n8293) );
  INVX1 U8239 ( .A(n8296), .Y(n8294) );
  INVX1 U8240 ( .A(n8294), .Y(n8295) );
  BUFX2 U8241 ( .A(fifo[1007]), .Y(n8296) );
  INVX1 U8242 ( .A(n8299), .Y(n8297) );
  INVX1 U8243 ( .A(n8297), .Y(n8298) );
  BUFX2 U8244 ( .A(fifo[1008]), .Y(n8299) );
  INVX1 U8245 ( .A(n8302), .Y(n8300) );
  INVX1 U8246 ( .A(n8300), .Y(n8301) );
  BUFX2 U8247 ( .A(fifo[1009]), .Y(n8302) );
  INVX1 U8248 ( .A(n8305), .Y(n8303) );
  INVX1 U8249 ( .A(n8303), .Y(n8304) );
  BUFX2 U8250 ( .A(fifo[1010]), .Y(n8305) );
  INVX1 U8251 ( .A(n8308), .Y(n8306) );
  INVX1 U8252 ( .A(n8306), .Y(n8307) );
  BUFX2 U8253 ( .A(fifo[1011]), .Y(n8308) );
  INVX1 U8254 ( .A(n8311), .Y(n8309) );
  INVX1 U8255 ( .A(n8309), .Y(n8310) );
  BUFX2 U8256 ( .A(fifo[1012]), .Y(n8311) );
  INVX1 U8257 ( .A(n8314), .Y(n8312) );
  INVX1 U8258 ( .A(n8312), .Y(n8313) );
  BUFX2 U8259 ( .A(fifo[1013]), .Y(n8314) );
  INVX1 U8260 ( .A(n8317), .Y(n8315) );
  INVX1 U8261 ( .A(n8315), .Y(n8316) );
  BUFX2 U8262 ( .A(fifo[1014]), .Y(n8317) );
  INVX1 U8263 ( .A(n8320), .Y(n8318) );
  INVX1 U8264 ( .A(n8318), .Y(n8319) );
  BUFX2 U8265 ( .A(fifo[1015]), .Y(n8320) );
  INVX1 U8266 ( .A(n8323), .Y(n8321) );
  INVX1 U8267 ( .A(n8321), .Y(n8322) );
  BUFX2 U8268 ( .A(fifo[1016]), .Y(n8323) );
  INVX1 U8269 ( .A(n8326), .Y(n8324) );
  INVX1 U8270 ( .A(n8324), .Y(n8325) );
  BUFX2 U8271 ( .A(fifo[1017]), .Y(n8326) );
  INVX1 U8272 ( .A(n8329), .Y(n8327) );
  INVX1 U8273 ( .A(n8327), .Y(n8328) );
  BUFX2 U8274 ( .A(fifo[1018]), .Y(n8329) );
  INVX1 U8275 ( .A(n8332), .Y(n8330) );
  INVX1 U8276 ( .A(n8330), .Y(n8331) );
  BUFX2 U8277 ( .A(fifo[1019]), .Y(n8332) );
  INVX1 U8278 ( .A(n8335), .Y(n8333) );
  INVX1 U8279 ( .A(n8333), .Y(n8334) );
  BUFX2 U8280 ( .A(fifo[408]), .Y(n8335) );
  INVX1 U8281 ( .A(n8338), .Y(n8336) );
  INVX1 U8282 ( .A(n8336), .Y(n8337) );
  BUFX2 U8283 ( .A(fifo[409]), .Y(n8338) );
  INVX1 U8284 ( .A(n8341), .Y(n8339) );
  INVX1 U8285 ( .A(n8339), .Y(n8340) );
  BUFX2 U8286 ( .A(fifo[410]), .Y(n8341) );
  INVX1 U8287 ( .A(n8344), .Y(n8342) );
  INVX1 U8288 ( .A(n8342), .Y(n8343) );
  BUFX2 U8289 ( .A(fifo[411]), .Y(n8344) );
  INVX1 U8290 ( .A(n8347), .Y(n8345) );
  INVX1 U8291 ( .A(n8345), .Y(n8346) );
  BUFX2 U8292 ( .A(fifo[412]), .Y(n8347) );
  INVX1 U8293 ( .A(n8350), .Y(n8348) );
  INVX1 U8294 ( .A(n8348), .Y(n8349) );
  BUFX2 U8295 ( .A(fifo[413]), .Y(n8350) );
  INVX1 U8296 ( .A(n8353), .Y(n8351) );
  INVX1 U8297 ( .A(n8351), .Y(n8352) );
  BUFX2 U8298 ( .A(fifo[414]), .Y(n8353) );
  INVX1 U8299 ( .A(n8356), .Y(n8354) );
  INVX1 U8300 ( .A(n8354), .Y(n8355) );
  BUFX2 U8301 ( .A(fifo[415]), .Y(n8356) );
  INVX1 U8302 ( .A(n8359), .Y(n8357) );
  INVX1 U8303 ( .A(n8357), .Y(n8358) );
  BUFX2 U8304 ( .A(fifo[416]), .Y(n8359) );
  INVX1 U8305 ( .A(n8362), .Y(n8360) );
  INVX1 U8306 ( .A(n8360), .Y(n8361) );
  BUFX2 U8307 ( .A(fifo[417]), .Y(n8362) );
  INVX1 U8308 ( .A(n8365), .Y(n8363) );
  INVX1 U8309 ( .A(n8363), .Y(n8364) );
  BUFX2 U8310 ( .A(fifo[418]), .Y(n8365) );
  INVX1 U8311 ( .A(n8368), .Y(n8366) );
  INVX1 U8312 ( .A(n8366), .Y(n8367) );
  BUFX2 U8313 ( .A(fifo[419]), .Y(n8368) );
  INVX1 U8314 ( .A(n8371), .Y(n8369) );
  INVX1 U8315 ( .A(n8369), .Y(n8370) );
  BUFX2 U8316 ( .A(fifo[420]), .Y(n8371) );
  INVX1 U8317 ( .A(n8374), .Y(n8372) );
  INVX1 U8318 ( .A(n8372), .Y(n8373) );
  BUFX2 U8319 ( .A(fifo[421]), .Y(n8374) );
  INVX1 U8320 ( .A(n8377), .Y(n8375) );
  INVX1 U8321 ( .A(n8375), .Y(n8376) );
  BUFX2 U8322 ( .A(fifo[422]), .Y(n8377) );
  INVX1 U8323 ( .A(n8380), .Y(n8378) );
  INVX1 U8324 ( .A(n8378), .Y(n8379) );
  BUFX2 U8325 ( .A(fifo[423]), .Y(n8380) );
  INVX1 U8326 ( .A(n8383), .Y(n8381) );
  INVX1 U8327 ( .A(n8381), .Y(n8382) );
  BUFX2 U8328 ( .A(fifo[424]), .Y(n8383) );
  INVX1 U8329 ( .A(n8386), .Y(n8384) );
  INVX1 U8330 ( .A(n8384), .Y(n8385) );
  BUFX2 U8331 ( .A(fifo[425]), .Y(n8386) );
  INVX1 U8332 ( .A(n8389), .Y(n8387) );
  INVX1 U8333 ( .A(n8387), .Y(n8388) );
  BUFX2 U8334 ( .A(fifo[426]), .Y(n8389) );
  INVX1 U8335 ( .A(n8392), .Y(n8390) );
  INVX1 U8336 ( .A(n8390), .Y(n8391) );
  BUFX2 U8337 ( .A(fifo[427]), .Y(n8392) );
  INVX1 U8338 ( .A(n8395), .Y(n8393) );
  INVX1 U8339 ( .A(n8393), .Y(n8394) );
  BUFX2 U8340 ( .A(fifo[428]), .Y(n8395) );
  INVX1 U8341 ( .A(n8398), .Y(n8396) );
  INVX1 U8342 ( .A(n8396), .Y(n8397) );
  BUFX2 U8343 ( .A(fifo[429]), .Y(n8398) );
  INVX1 U8344 ( .A(n8401), .Y(n8399) );
  INVX1 U8345 ( .A(n8399), .Y(n8400) );
  BUFX2 U8346 ( .A(fifo[430]), .Y(n8401) );
  INVX1 U8347 ( .A(n8404), .Y(n8402) );
  INVX1 U8348 ( .A(n8402), .Y(n8403) );
  BUFX2 U8349 ( .A(fifo[431]), .Y(n8404) );
  INVX1 U8350 ( .A(n8407), .Y(n8405) );
  INVX1 U8351 ( .A(n8405), .Y(n8406) );
  BUFX2 U8352 ( .A(fifo[432]), .Y(n8407) );
  INVX1 U8353 ( .A(n8410), .Y(n8408) );
  INVX1 U8354 ( .A(n8408), .Y(n8409) );
  BUFX2 U8355 ( .A(fifo[433]), .Y(n8410) );
  INVX1 U8356 ( .A(n8413), .Y(n8411) );
  INVX1 U8357 ( .A(n8411), .Y(n8412) );
  BUFX2 U8358 ( .A(fifo[434]), .Y(n8413) );
  INVX1 U8359 ( .A(n8416), .Y(n8414) );
  INVX1 U8360 ( .A(n8414), .Y(n8415) );
  BUFX2 U8361 ( .A(fifo[435]), .Y(n8416) );
  INVX1 U8362 ( .A(n8419), .Y(n8417) );
  INVX1 U8363 ( .A(n8417), .Y(n8418) );
  BUFX2 U8364 ( .A(fifo[436]), .Y(n8419) );
  INVX1 U8365 ( .A(n8422), .Y(n8420) );
  INVX1 U8366 ( .A(n8420), .Y(n8421) );
  BUFX2 U8367 ( .A(fifo[437]), .Y(n8422) );
  INVX1 U8368 ( .A(n8425), .Y(n8423) );
  INVX1 U8369 ( .A(n8423), .Y(n8424) );
  BUFX2 U8370 ( .A(fifo[438]), .Y(n8425) );
  INVX1 U8371 ( .A(n8428), .Y(n8426) );
  INVX1 U8372 ( .A(n8426), .Y(n8427) );
  BUFX2 U8373 ( .A(fifo[439]), .Y(n8428) );
  INVX1 U8374 ( .A(n8431), .Y(n8429) );
  INVX1 U8375 ( .A(n8429), .Y(n8430) );
  BUFX2 U8376 ( .A(fifo[440]), .Y(n8431) );
  INVX1 U8377 ( .A(n8434), .Y(n8432) );
  INVX1 U8378 ( .A(n8432), .Y(n8433) );
  BUFX2 U8379 ( .A(fifo[441]), .Y(n8434) );
  INVX1 U8380 ( .A(n8437), .Y(n8435) );
  INVX1 U8381 ( .A(n8435), .Y(n8436) );
  BUFX2 U8382 ( .A(fifo[340]), .Y(n8437) );
  INVX1 U8383 ( .A(n8440), .Y(n8438) );
  INVX1 U8384 ( .A(n8438), .Y(n8439) );
  BUFX2 U8385 ( .A(fifo[341]), .Y(n8440) );
  INVX1 U8386 ( .A(n8443), .Y(n8441) );
  INVX1 U8387 ( .A(n8441), .Y(n8442) );
  BUFX2 U8388 ( .A(fifo[342]), .Y(n8443) );
  INVX1 U8389 ( .A(n8446), .Y(n8444) );
  INVX1 U8390 ( .A(n8444), .Y(n8445) );
  BUFX2 U8391 ( .A(fifo[343]), .Y(n8446) );
  INVX1 U8392 ( .A(n8449), .Y(n8447) );
  INVX1 U8393 ( .A(n8447), .Y(n8448) );
  BUFX2 U8394 ( .A(fifo[344]), .Y(n8449) );
  INVX1 U8395 ( .A(n8452), .Y(n8450) );
  INVX1 U8396 ( .A(n8450), .Y(n8451) );
  BUFX2 U8397 ( .A(fifo[345]), .Y(n8452) );
  INVX1 U8398 ( .A(n8455), .Y(n8453) );
  INVX1 U8399 ( .A(n8453), .Y(n8454) );
  BUFX2 U8400 ( .A(fifo[346]), .Y(n8455) );
  INVX1 U8401 ( .A(n8458), .Y(n8456) );
  INVX1 U8402 ( .A(n8456), .Y(n8457) );
  BUFX2 U8403 ( .A(fifo[347]), .Y(n8458) );
  INVX1 U8404 ( .A(n8461), .Y(n8459) );
  INVX1 U8405 ( .A(n8459), .Y(n8460) );
  BUFX2 U8406 ( .A(fifo[348]), .Y(n8461) );
  INVX1 U8407 ( .A(n8464), .Y(n8462) );
  INVX1 U8408 ( .A(n8462), .Y(n8463) );
  BUFX2 U8409 ( .A(fifo[349]), .Y(n8464) );
  INVX1 U8410 ( .A(n8467), .Y(n8465) );
  INVX1 U8411 ( .A(n8465), .Y(n8466) );
  BUFX2 U8412 ( .A(fifo[350]), .Y(n8467) );
  INVX1 U8413 ( .A(n8470), .Y(n8468) );
  INVX1 U8414 ( .A(n8468), .Y(n8469) );
  BUFX2 U8415 ( .A(fifo[351]), .Y(n8470) );
  INVX1 U8416 ( .A(n8473), .Y(n8471) );
  INVX1 U8417 ( .A(n8471), .Y(n8472) );
  BUFX2 U8418 ( .A(fifo[352]), .Y(n8473) );
  INVX1 U8419 ( .A(n8476), .Y(n8474) );
  INVX1 U8420 ( .A(n8474), .Y(n8475) );
  BUFX2 U8421 ( .A(fifo[353]), .Y(n8476) );
  INVX1 U8422 ( .A(n8479), .Y(n8477) );
  INVX1 U8423 ( .A(n8477), .Y(n8478) );
  BUFX2 U8424 ( .A(fifo[354]), .Y(n8479) );
  INVX1 U8425 ( .A(n8482), .Y(n8480) );
  INVX1 U8426 ( .A(n8480), .Y(n8481) );
  BUFX2 U8427 ( .A(fifo[355]), .Y(n8482) );
  INVX1 U8428 ( .A(n8485), .Y(n8483) );
  INVX1 U8429 ( .A(n8483), .Y(n8484) );
  BUFX2 U8430 ( .A(fifo[356]), .Y(n8485) );
  INVX1 U8431 ( .A(n8488), .Y(n8486) );
  INVX1 U8432 ( .A(n8486), .Y(n8487) );
  BUFX2 U8433 ( .A(fifo[357]), .Y(n8488) );
  INVX1 U8434 ( .A(n8491), .Y(n8489) );
  INVX1 U8435 ( .A(n8489), .Y(n8490) );
  BUFX2 U8436 ( .A(fifo[358]), .Y(n8491) );
  INVX1 U8437 ( .A(n8494), .Y(n8492) );
  INVX1 U8438 ( .A(n8492), .Y(n8493) );
  BUFX2 U8439 ( .A(fifo[359]), .Y(n8494) );
  INVX1 U8440 ( .A(n8497), .Y(n8495) );
  INVX1 U8441 ( .A(n8495), .Y(n8496) );
  BUFX2 U8442 ( .A(fifo[360]), .Y(n8497) );
  INVX1 U8443 ( .A(n8500), .Y(n8498) );
  INVX1 U8444 ( .A(n8498), .Y(n8499) );
  BUFX2 U8445 ( .A(fifo[361]), .Y(n8500) );
  INVX1 U8446 ( .A(n8503), .Y(n8501) );
  INVX1 U8447 ( .A(n8501), .Y(n8502) );
  BUFX2 U8448 ( .A(fifo[362]), .Y(n8503) );
  INVX1 U8449 ( .A(n8506), .Y(n8504) );
  INVX1 U8450 ( .A(n8504), .Y(n8505) );
  BUFX2 U8451 ( .A(fifo[363]), .Y(n8506) );
  INVX1 U8452 ( .A(n8509), .Y(n8507) );
  INVX1 U8453 ( .A(n8507), .Y(n8508) );
  BUFX2 U8454 ( .A(fifo[364]), .Y(n8509) );
  INVX1 U8455 ( .A(n8512), .Y(n8510) );
  INVX1 U8456 ( .A(n8510), .Y(n8511) );
  BUFX2 U8457 ( .A(fifo[365]), .Y(n8512) );
  INVX1 U8458 ( .A(n8515), .Y(n8513) );
  INVX1 U8459 ( .A(n8513), .Y(n8514) );
  BUFX2 U8460 ( .A(fifo[366]), .Y(n8515) );
  INVX1 U8461 ( .A(n8518), .Y(n8516) );
  INVX1 U8462 ( .A(n8516), .Y(n8517) );
  BUFX2 U8463 ( .A(fifo[367]), .Y(n8518) );
  INVX1 U8464 ( .A(n8521), .Y(n8519) );
  INVX1 U8465 ( .A(n8519), .Y(n8520) );
  BUFX2 U8466 ( .A(fifo[368]), .Y(n8521) );
  INVX1 U8467 ( .A(n8524), .Y(n8522) );
  INVX1 U8468 ( .A(n8522), .Y(n8523) );
  BUFX2 U8469 ( .A(fifo[369]), .Y(n8524) );
  INVX1 U8470 ( .A(n8527), .Y(n8525) );
  INVX1 U8471 ( .A(n8525), .Y(n8526) );
  BUFX2 U8472 ( .A(fifo[370]), .Y(n8527) );
  INVX1 U8473 ( .A(n8530), .Y(n8528) );
  INVX1 U8474 ( .A(n8528), .Y(n8529) );
  BUFX2 U8475 ( .A(fifo[371]), .Y(n8530) );
  INVX1 U8476 ( .A(n8533), .Y(n8531) );
  INVX1 U8477 ( .A(n8531), .Y(n8532) );
  BUFX2 U8478 ( .A(fifo[372]), .Y(n8533) );
  INVX1 U8479 ( .A(n8536), .Y(n8534) );
  INVX1 U8480 ( .A(n8534), .Y(n8535) );
  BUFX2 U8481 ( .A(fifo[373]), .Y(n8536) );
  INVX1 U8482 ( .A(n8539), .Y(n8537) );
  INVX1 U8483 ( .A(n8537), .Y(n8538) );
  BUFX2 U8484 ( .A(fifo[272]), .Y(n8539) );
  INVX1 U8485 ( .A(n8542), .Y(n8540) );
  INVX1 U8486 ( .A(n8540), .Y(n8541) );
  BUFX2 U8487 ( .A(fifo[273]), .Y(n8542) );
  INVX1 U8488 ( .A(n8545), .Y(n8543) );
  INVX1 U8489 ( .A(n8543), .Y(n8544) );
  BUFX2 U8490 ( .A(fifo[274]), .Y(n8545) );
  INVX1 U8491 ( .A(n8548), .Y(n8546) );
  INVX1 U8492 ( .A(n8546), .Y(n8547) );
  BUFX2 U8493 ( .A(fifo[275]), .Y(n8548) );
  INVX1 U8494 ( .A(n8551), .Y(n8549) );
  INVX1 U8495 ( .A(n8549), .Y(n8550) );
  BUFX2 U8496 ( .A(fifo[276]), .Y(n8551) );
  INVX1 U8497 ( .A(n8554), .Y(n8552) );
  INVX1 U8498 ( .A(n8552), .Y(n8553) );
  BUFX2 U8499 ( .A(fifo[277]), .Y(n8554) );
  INVX1 U8500 ( .A(n8557), .Y(n8555) );
  INVX1 U8501 ( .A(n8555), .Y(n8556) );
  BUFX2 U8502 ( .A(fifo[278]), .Y(n8557) );
  INVX1 U8503 ( .A(n8560), .Y(n8558) );
  INVX1 U8504 ( .A(n8558), .Y(n8559) );
  BUFX2 U8505 ( .A(fifo[279]), .Y(n8560) );
  INVX1 U8506 ( .A(n8563), .Y(n8561) );
  INVX1 U8507 ( .A(n8561), .Y(n8562) );
  BUFX2 U8508 ( .A(fifo[280]), .Y(n8563) );
  INVX1 U8509 ( .A(n8566), .Y(n8564) );
  INVX1 U8510 ( .A(n8564), .Y(n8565) );
  BUFX2 U8511 ( .A(fifo[281]), .Y(n8566) );
  INVX1 U8512 ( .A(n8569), .Y(n8567) );
  INVX1 U8513 ( .A(n8567), .Y(n8568) );
  BUFX2 U8514 ( .A(fifo[282]), .Y(n8569) );
  INVX1 U8515 ( .A(n8572), .Y(n8570) );
  INVX1 U8516 ( .A(n8570), .Y(n8571) );
  BUFX2 U8517 ( .A(fifo[283]), .Y(n8572) );
  INVX1 U8518 ( .A(n8575), .Y(n8573) );
  INVX1 U8519 ( .A(n8573), .Y(n8574) );
  BUFX2 U8520 ( .A(fifo[284]), .Y(n8575) );
  INVX1 U8521 ( .A(n8578), .Y(n8576) );
  INVX1 U8522 ( .A(n8576), .Y(n8577) );
  BUFX2 U8523 ( .A(fifo[285]), .Y(n8578) );
  INVX1 U8524 ( .A(n8581), .Y(n8579) );
  INVX1 U8525 ( .A(n8579), .Y(n8580) );
  BUFX2 U8526 ( .A(fifo[286]), .Y(n8581) );
  INVX1 U8527 ( .A(n8584), .Y(n8582) );
  INVX1 U8528 ( .A(n8582), .Y(n8583) );
  BUFX2 U8529 ( .A(fifo[287]), .Y(n8584) );
  INVX1 U8530 ( .A(n8587), .Y(n8585) );
  INVX1 U8531 ( .A(n8585), .Y(n8586) );
  BUFX2 U8532 ( .A(fifo[288]), .Y(n8587) );
  INVX1 U8533 ( .A(n8590), .Y(n8588) );
  INVX1 U8534 ( .A(n8588), .Y(n8589) );
  BUFX2 U8535 ( .A(fifo[289]), .Y(n8590) );
  INVX1 U8536 ( .A(n8593), .Y(n8591) );
  INVX1 U8537 ( .A(n8591), .Y(n8592) );
  BUFX2 U8538 ( .A(fifo[290]), .Y(n8593) );
  INVX1 U8539 ( .A(n8596), .Y(n8594) );
  INVX1 U8540 ( .A(n8594), .Y(n8595) );
  BUFX2 U8541 ( .A(fifo[291]), .Y(n8596) );
  INVX1 U8542 ( .A(n8599), .Y(n8597) );
  INVX1 U8543 ( .A(n8597), .Y(n8598) );
  BUFX2 U8544 ( .A(fifo[292]), .Y(n8599) );
  INVX1 U8545 ( .A(n8602), .Y(n8600) );
  INVX1 U8546 ( .A(n8600), .Y(n8601) );
  BUFX2 U8547 ( .A(fifo[293]), .Y(n8602) );
  INVX1 U8548 ( .A(n8605), .Y(n8603) );
  INVX1 U8549 ( .A(n8603), .Y(n8604) );
  BUFX2 U8550 ( .A(fifo[294]), .Y(n8605) );
  INVX1 U8551 ( .A(n8608), .Y(n8606) );
  INVX1 U8552 ( .A(n8606), .Y(n8607) );
  BUFX2 U8553 ( .A(fifo[295]), .Y(n8608) );
  INVX1 U8554 ( .A(n8611), .Y(n8609) );
  INVX1 U8555 ( .A(n8609), .Y(n8610) );
  BUFX2 U8556 ( .A(fifo[296]), .Y(n8611) );
  INVX1 U8557 ( .A(n8614), .Y(n8612) );
  INVX1 U8558 ( .A(n8612), .Y(n8613) );
  BUFX2 U8559 ( .A(fifo[297]), .Y(n8614) );
  INVX1 U8560 ( .A(n8617), .Y(n8615) );
  INVX1 U8561 ( .A(n8615), .Y(n8616) );
  BUFX2 U8562 ( .A(fifo[298]), .Y(n8617) );
  INVX1 U8563 ( .A(n8620), .Y(n8618) );
  INVX1 U8564 ( .A(n8618), .Y(n8619) );
  BUFX2 U8565 ( .A(fifo[299]), .Y(n8620) );
  INVX1 U8566 ( .A(n8623), .Y(n8621) );
  INVX1 U8567 ( .A(n8621), .Y(n8622) );
  BUFX2 U8568 ( .A(fifo[300]), .Y(n8623) );
  INVX1 U8569 ( .A(n8626), .Y(n8624) );
  INVX1 U8570 ( .A(n8624), .Y(n8625) );
  BUFX2 U8571 ( .A(fifo[301]), .Y(n8626) );
  INVX1 U8572 ( .A(n8629), .Y(n8627) );
  INVX1 U8573 ( .A(n8627), .Y(n8628) );
  BUFX2 U8574 ( .A(fifo[302]), .Y(n8629) );
  INVX1 U8575 ( .A(n8632), .Y(n8630) );
  INVX1 U8576 ( .A(n8630), .Y(n8631) );
  BUFX2 U8577 ( .A(fifo[303]), .Y(n8632) );
  INVX1 U8578 ( .A(n8635), .Y(n8633) );
  INVX1 U8579 ( .A(n8633), .Y(n8634) );
  BUFX2 U8580 ( .A(fifo[304]), .Y(n8635) );
  INVX1 U8581 ( .A(n8638), .Y(n8636) );
  INVX1 U8582 ( .A(n8636), .Y(n8637) );
  BUFX2 U8583 ( .A(fifo[305]), .Y(n8638) );
  INVX1 U8584 ( .A(n8641), .Y(n8639) );
  INVX1 U8585 ( .A(n8639), .Y(n8640) );
  BUFX2 U8586 ( .A(fifo[476]), .Y(n8641) );
  INVX1 U8587 ( .A(n8644), .Y(n8642) );
  INVX1 U8588 ( .A(n8642), .Y(n8643) );
  BUFX2 U8589 ( .A(fifo[477]), .Y(n8644) );
  INVX1 U8590 ( .A(n8647), .Y(n8645) );
  INVX1 U8591 ( .A(n8645), .Y(n8646) );
  BUFX2 U8592 ( .A(fifo[478]), .Y(n8647) );
  INVX1 U8593 ( .A(n8650), .Y(n8648) );
  INVX1 U8594 ( .A(n8648), .Y(n8649) );
  BUFX2 U8595 ( .A(fifo[479]), .Y(n8650) );
  INVX1 U8596 ( .A(n8653), .Y(n8651) );
  INVX1 U8597 ( .A(n8651), .Y(n8652) );
  BUFX2 U8598 ( .A(fifo[480]), .Y(n8653) );
  INVX1 U8599 ( .A(n8656), .Y(n8654) );
  INVX1 U8600 ( .A(n8654), .Y(n8655) );
  BUFX2 U8601 ( .A(fifo[481]), .Y(n8656) );
  INVX1 U8602 ( .A(n8659), .Y(n8657) );
  INVX1 U8603 ( .A(n8657), .Y(n8658) );
  BUFX2 U8604 ( .A(fifo[482]), .Y(n8659) );
  INVX1 U8605 ( .A(n8662), .Y(n8660) );
  INVX1 U8606 ( .A(n8660), .Y(n8661) );
  BUFX2 U8607 ( .A(fifo[483]), .Y(n8662) );
  INVX1 U8608 ( .A(n8665), .Y(n8663) );
  INVX1 U8609 ( .A(n8663), .Y(n8664) );
  BUFX2 U8610 ( .A(fifo[484]), .Y(n8665) );
  INVX1 U8611 ( .A(n8668), .Y(n8666) );
  INVX1 U8612 ( .A(n8666), .Y(n8667) );
  BUFX2 U8613 ( .A(fifo[485]), .Y(n8668) );
  INVX1 U8614 ( .A(n8671), .Y(n8669) );
  INVX1 U8615 ( .A(n8669), .Y(n8670) );
  BUFX2 U8616 ( .A(fifo[486]), .Y(n8671) );
  INVX1 U8617 ( .A(n8674), .Y(n8672) );
  INVX1 U8618 ( .A(n8672), .Y(n8673) );
  BUFX2 U8619 ( .A(fifo[487]), .Y(n8674) );
  INVX1 U8620 ( .A(n8677), .Y(n8675) );
  INVX1 U8621 ( .A(n8675), .Y(n8676) );
  BUFX2 U8622 ( .A(fifo[488]), .Y(n8677) );
  INVX1 U8623 ( .A(n8680), .Y(n8678) );
  INVX1 U8624 ( .A(n8678), .Y(n8679) );
  BUFX2 U8625 ( .A(fifo[489]), .Y(n8680) );
  INVX1 U8626 ( .A(n8683), .Y(n8681) );
  INVX1 U8627 ( .A(n8681), .Y(n8682) );
  BUFX2 U8628 ( .A(fifo[490]), .Y(n8683) );
  INVX1 U8629 ( .A(n8686), .Y(n8684) );
  INVX1 U8630 ( .A(n8684), .Y(n8685) );
  BUFX2 U8631 ( .A(fifo[491]), .Y(n8686) );
  INVX1 U8632 ( .A(n8689), .Y(n8687) );
  INVX1 U8633 ( .A(n8687), .Y(n8688) );
  BUFX2 U8634 ( .A(fifo[492]), .Y(n8689) );
  INVX1 U8635 ( .A(n8692), .Y(n8690) );
  INVX1 U8636 ( .A(n8690), .Y(n8691) );
  BUFX2 U8637 ( .A(fifo[493]), .Y(n8692) );
  INVX1 U8638 ( .A(n8695), .Y(n8693) );
  INVX1 U8639 ( .A(n8693), .Y(n8694) );
  BUFX2 U8640 ( .A(fifo[494]), .Y(n8695) );
  INVX1 U8641 ( .A(n8698), .Y(n8696) );
  INVX1 U8642 ( .A(n8696), .Y(n8697) );
  BUFX2 U8643 ( .A(fifo[495]), .Y(n8698) );
  INVX1 U8644 ( .A(n8701), .Y(n8699) );
  INVX1 U8645 ( .A(n8699), .Y(n8700) );
  BUFX2 U8646 ( .A(fifo[496]), .Y(n8701) );
  INVX1 U8647 ( .A(n8704), .Y(n8702) );
  INVX1 U8648 ( .A(n8702), .Y(n8703) );
  BUFX2 U8649 ( .A(fifo[497]), .Y(n8704) );
  INVX1 U8650 ( .A(n8707), .Y(n8705) );
  INVX1 U8651 ( .A(n8705), .Y(n8706) );
  BUFX2 U8652 ( .A(fifo[498]), .Y(n8707) );
  INVX1 U8653 ( .A(n8710), .Y(n8708) );
  INVX1 U8654 ( .A(n8708), .Y(n8709) );
  BUFX2 U8655 ( .A(fifo[499]), .Y(n8710) );
  INVX1 U8656 ( .A(n8713), .Y(n8711) );
  INVX1 U8657 ( .A(n8711), .Y(n8712) );
  BUFX2 U8658 ( .A(fifo[500]), .Y(n8713) );
  INVX1 U8659 ( .A(n8716), .Y(n8714) );
  INVX1 U8660 ( .A(n8714), .Y(n8715) );
  BUFX2 U8661 ( .A(fifo[501]), .Y(n8716) );
  INVX1 U8662 ( .A(n8719), .Y(n8717) );
  INVX1 U8663 ( .A(n8717), .Y(n8718) );
  BUFX2 U8664 ( .A(fifo[502]), .Y(n8719) );
  INVX1 U8665 ( .A(n8722), .Y(n8720) );
  INVX1 U8666 ( .A(n8720), .Y(n8721) );
  BUFX2 U8667 ( .A(fifo[503]), .Y(n8722) );
  INVX1 U8668 ( .A(n8725), .Y(n8723) );
  INVX1 U8669 ( .A(n8723), .Y(n8724) );
  BUFX2 U8670 ( .A(fifo[504]), .Y(n8725) );
  INVX1 U8671 ( .A(n8728), .Y(n8726) );
  INVX1 U8672 ( .A(n8726), .Y(n8727) );
  BUFX2 U8673 ( .A(fifo[505]), .Y(n8728) );
  INVX1 U8674 ( .A(n8731), .Y(n8729) );
  INVX1 U8675 ( .A(n8729), .Y(n8730) );
  BUFX2 U8676 ( .A(fifo[506]), .Y(n8731) );
  INVX1 U8677 ( .A(n8734), .Y(n8732) );
  INVX1 U8678 ( .A(n8732), .Y(n8733) );
  BUFX2 U8679 ( .A(fifo[507]), .Y(n8734) );
  INVX1 U8680 ( .A(n8737), .Y(n8735) );
  INVX1 U8681 ( .A(n8735), .Y(n8736) );
  BUFX2 U8682 ( .A(fifo[508]), .Y(n8737) );
  INVX1 U8683 ( .A(n8740), .Y(n8738) );
  INVX1 U8684 ( .A(n8738), .Y(n8739) );
  BUFX2 U8685 ( .A(fifo[509]), .Y(n8740) );
  INVX1 U8686 ( .A(n8743), .Y(n8741) );
  INVX1 U8687 ( .A(n8741), .Y(n8742) );
  BUFX2 U8688 ( .A(fifo[0]), .Y(n8743) );
  INVX1 U8689 ( .A(n8746), .Y(n8744) );
  INVX1 U8690 ( .A(n8744), .Y(n8745) );
  BUFX2 U8691 ( .A(fifo[1]), .Y(n8746) );
  INVX1 U8692 ( .A(n8749), .Y(n8747) );
  INVX1 U8693 ( .A(n8747), .Y(n8748) );
  BUFX2 U8694 ( .A(fifo[2]), .Y(n8749) );
  INVX1 U8695 ( .A(n8752), .Y(n8750) );
  INVX1 U8696 ( .A(n8750), .Y(n8751) );
  BUFX2 U8697 ( .A(fifo[3]), .Y(n8752) );
  INVX1 U8698 ( .A(n8755), .Y(n8753) );
  INVX1 U8699 ( .A(n8753), .Y(n8754) );
  BUFX2 U8700 ( .A(fifo[4]), .Y(n8755) );
  INVX1 U8701 ( .A(n8758), .Y(n8756) );
  INVX1 U8702 ( .A(n8756), .Y(n8757) );
  BUFX2 U8703 ( .A(fifo[5]), .Y(n8758) );
  INVX1 U8704 ( .A(n8761), .Y(n8759) );
  INVX1 U8705 ( .A(n8759), .Y(n8760) );
  BUFX2 U8706 ( .A(fifo[6]), .Y(n8761) );
  INVX1 U8707 ( .A(n8764), .Y(n8762) );
  INVX1 U8708 ( .A(n8762), .Y(n8763) );
  BUFX2 U8709 ( .A(fifo[7]), .Y(n8764) );
  INVX1 U8710 ( .A(n8767), .Y(n8765) );
  INVX1 U8711 ( .A(n8765), .Y(n8766) );
  BUFX2 U8712 ( .A(fifo[8]), .Y(n8767) );
  INVX1 U8713 ( .A(n8770), .Y(n8768) );
  INVX1 U8714 ( .A(n8768), .Y(n8769) );
  BUFX2 U8715 ( .A(fifo[9]), .Y(n8770) );
  INVX1 U8716 ( .A(n8773), .Y(n8771) );
  INVX1 U8717 ( .A(n8771), .Y(n8772) );
  BUFX2 U8718 ( .A(fifo[10]), .Y(n8773) );
  INVX1 U8719 ( .A(n8776), .Y(n8774) );
  INVX1 U8720 ( .A(n8774), .Y(n8775) );
  BUFX2 U8721 ( .A(fifo[11]), .Y(n8776) );
  INVX1 U8722 ( .A(n8779), .Y(n8777) );
  INVX1 U8723 ( .A(n8777), .Y(n8778) );
  BUFX2 U8724 ( .A(fifo[12]), .Y(n8779) );
  INVX1 U8725 ( .A(n8782), .Y(n8780) );
  INVX1 U8726 ( .A(n8780), .Y(n8781) );
  BUFX2 U8727 ( .A(fifo[13]), .Y(n8782) );
  INVX1 U8728 ( .A(n8785), .Y(n8783) );
  INVX1 U8729 ( .A(n8783), .Y(n8784) );
  BUFX2 U8730 ( .A(fifo[14]), .Y(n8785) );
  INVX1 U8731 ( .A(n8788), .Y(n8786) );
  INVX1 U8732 ( .A(n8786), .Y(n8787) );
  BUFX2 U8733 ( .A(fifo[15]), .Y(n8788) );
  INVX1 U8734 ( .A(n8791), .Y(n8789) );
  INVX1 U8735 ( .A(n8789), .Y(n8790) );
  BUFX2 U8736 ( .A(fifo[16]), .Y(n8791) );
  INVX1 U8737 ( .A(n8794), .Y(n8792) );
  INVX1 U8738 ( .A(n8792), .Y(n8793) );
  BUFX2 U8739 ( .A(fifo[17]), .Y(n8794) );
  INVX1 U8740 ( .A(n8797), .Y(n8795) );
  INVX1 U8741 ( .A(n8795), .Y(n8796) );
  BUFX2 U8742 ( .A(fifo[18]), .Y(n8797) );
  INVX1 U8743 ( .A(n8800), .Y(n8798) );
  INVX1 U8744 ( .A(n8798), .Y(n8799) );
  BUFX2 U8745 ( .A(fifo[19]), .Y(n8800) );
  INVX1 U8746 ( .A(n8803), .Y(n8801) );
  INVX1 U8747 ( .A(n8801), .Y(n8802) );
  BUFX2 U8748 ( .A(fifo[20]), .Y(n8803) );
  INVX1 U8749 ( .A(n8806), .Y(n8804) );
  INVX1 U8750 ( .A(n8804), .Y(n8805) );
  BUFX2 U8751 ( .A(fifo[21]), .Y(n8806) );
  INVX1 U8752 ( .A(n8809), .Y(n8807) );
  INVX1 U8753 ( .A(n8807), .Y(n8808) );
  BUFX2 U8754 ( .A(fifo[22]), .Y(n8809) );
  INVX1 U8755 ( .A(n8812), .Y(n8810) );
  INVX1 U8756 ( .A(n8810), .Y(n8811) );
  BUFX2 U8757 ( .A(fifo[23]), .Y(n8812) );
  INVX1 U8758 ( .A(n8815), .Y(n8813) );
  INVX1 U8759 ( .A(n8813), .Y(n8814) );
  BUFX2 U8760 ( .A(fifo[24]), .Y(n8815) );
  INVX1 U8761 ( .A(n8818), .Y(n8816) );
  INVX1 U8762 ( .A(n8816), .Y(n8817) );
  BUFX2 U8763 ( .A(fifo[25]), .Y(n8818) );
  INVX1 U8764 ( .A(n8821), .Y(n8819) );
  INVX1 U8765 ( .A(n8819), .Y(n8820) );
  BUFX2 U8766 ( .A(fifo[26]), .Y(n8821) );
  INVX1 U8767 ( .A(n8824), .Y(n8822) );
  INVX1 U8768 ( .A(n8822), .Y(n8823) );
  BUFX2 U8769 ( .A(fifo[27]), .Y(n8824) );
  INVX1 U8770 ( .A(n8827), .Y(n8825) );
  INVX1 U8771 ( .A(n8825), .Y(n8826) );
  BUFX2 U8772 ( .A(fifo[28]), .Y(n8827) );
  INVX1 U8773 ( .A(n8830), .Y(n8828) );
  INVX1 U8774 ( .A(n8828), .Y(n8829) );
  BUFX2 U8775 ( .A(fifo[29]), .Y(n8830) );
  INVX1 U8776 ( .A(n8833), .Y(n8831) );
  INVX1 U8777 ( .A(n8831), .Y(n8832) );
  BUFX2 U8778 ( .A(fifo[30]), .Y(n8833) );
  INVX1 U8779 ( .A(n8836), .Y(n8834) );
  INVX1 U8780 ( .A(n8834), .Y(n8835) );
  BUFX2 U8781 ( .A(fifo[31]), .Y(n8836) );
  INVX1 U8782 ( .A(n8839), .Y(n8837) );
  INVX1 U8783 ( .A(n8837), .Y(n8838) );
  BUFX2 U8784 ( .A(fifo[32]), .Y(n8839) );
  INVX1 U8785 ( .A(n8842), .Y(n8840) );
  INVX1 U8786 ( .A(n8840), .Y(n8841) );
  BUFX2 U8787 ( .A(fifo[33]), .Y(n8842) );
  INVX1 U8788 ( .A(n8845), .Y(n8843) );
  INVX1 U8789 ( .A(n8843), .Y(n8844) );
  BUFX2 U8790 ( .A(fifo[68]), .Y(n8845) );
  INVX1 U8791 ( .A(n8848), .Y(n8846) );
  INVX1 U8792 ( .A(n8846), .Y(n8847) );
  BUFX2 U8793 ( .A(fifo[69]), .Y(n8848) );
  INVX1 U8794 ( .A(n8851), .Y(n8849) );
  INVX1 U8795 ( .A(n8849), .Y(n8850) );
  BUFX2 U8796 ( .A(fifo[70]), .Y(n8851) );
  INVX1 U8797 ( .A(n8854), .Y(n8852) );
  INVX1 U8798 ( .A(n8852), .Y(n8853) );
  BUFX2 U8799 ( .A(fifo[71]), .Y(n8854) );
  INVX1 U8800 ( .A(n8857), .Y(n8855) );
  INVX1 U8801 ( .A(n8855), .Y(n8856) );
  BUFX2 U8802 ( .A(fifo[72]), .Y(n8857) );
  INVX1 U8803 ( .A(n8860), .Y(n8858) );
  INVX1 U8804 ( .A(n8858), .Y(n8859) );
  BUFX2 U8805 ( .A(fifo[73]), .Y(n8860) );
  INVX1 U8806 ( .A(n8863), .Y(n8861) );
  INVX1 U8807 ( .A(n8861), .Y(n8862) );
  BUFX2 U8808 ( .A(fifo[74]), .Y(n8863) );
  INVX1 U8809 ( .A(n8866), .Y(n8864) );
  INVX1 U8810 ( .A(n8864), .Y(n8865) );
  BUFX2 U8811 ( .A(fifo[75]), .Y(n8866) );
  INVX1 U8812 ( .A(n8869), .Y(n8867) );
  INVX1 U8813 ( .A(n8867), .Y(n8868) );
  BUFX2 U8814 ( .A(fifo[76]), .Y(n8869) );
  INVX1 U8815 ( .A(n8872), .Y(n8870) );
  INVX1 U8816 ( .A(n8870), .Y(n8871) );
  BUFX2 U8817 ( .A(fifo[77]), .Y(n8872) );
  INVX1 U8818 ( .A(n8875), .Y(n8873) );
  INVX1 U8819 ( .A(n8873), .Y(n8874) );
  BUFX2 U8820 ( .A(fifo[78]), .Y(n8875) );
  INVX1 U8821 ( .A(n8878), .Y(n8876) );
  INVX1 U8822 ( .A(n8876), .Y(n8877) );
  BUFX2 U8823 ( .A(fifo[79]), .Y(n8878) );
  INVX1 U8824 ( .A(n8881), .Y(n8879) );
  INVX1 U8825 ( .A(n8879), .Y(n8880) );
  BUFX2 U8826 ( .A(fifo[80]), .Y(n8881) );
  INVX1 U8827 ( .A(n8884), .Y(n8882) );
  INVX1 U8828 ( .A(n8882), .Y(n8883) );
  BUFX2 U8829 ( .A(fifo[81]), .Y(n8884) );
  INVX1 U8830 ( .A(n8887), .Y(n8885) );
  INVX1 U8831 ( .A(n8885), .Y(n8886) );
  BUFX2 U8832 ( .A(fifo[82]), .Y(n8887) );
  INVX1 U8833 ( .A(n8890), .Y(n8888) );
  INVX1 U8834 ( .A(n8888), .Y(n8889) );
  BUFX2 U8835 ( .A(fifo[83]), .Y(n8890) );
  INVX1 U8836 ( .A(n8893), .Y(n8891) );
  INVX1 U8837 ( .A(n8891), .Y(n8892) );
  BUFX2 U8838 ( .A(fifo[84]), .Y(n8893) );
  INVX1 U8839 ( .A(n8896), .Y(n8894) );
  INVX1 U8840 ( .A(n8894), .Y(n8895) );
  BUFX2 U8841 ( .A(fifo[85]), .Y(n8896) );
  INVX1 U8842 ( .A(n8899), .Y(n8897) );
  INVX1 U8843 ( .A(n8897), .Y(n8898) );
  BUFX2 U8844 ( .A(fifo[86]), .Y(n8899) );
  INVX1 U8845 ( .A(n8902), .Y(n8900) );
  INVX1 U8846 ( .A(n8900), .Y(n8901) );
  BUFX2 U8847 ( .A(fifo[87]), .Y(n8902) );
  INVX1 U8848 ( .A(n8905), .Y(n8903) );
  INVX1 U8849 ( .A(n8903), .Y(n8904) );
  BUFX2 U8850 ( .A(fifo[88]), .Y(n8905) );
  INVX1 U8851 ( .A(n8908), .Y(n8906) );
  INVX1 U8852 ( .A(n8906), .Y(n8907) );
  BUFX2 U8853 ( .A(fifo[89]), .Y(n8908) );
  INVX1 U8854 ( .A(n8911), .Y(n8909) );
  INVX1 U8855 ( .A(n8909), .Y(n8910) );
  BUFX2 U8856 ( .A(fifo[90]), .Y(n8911) );
  INVX1 U8857 ( .A(n8914), .Y(n8912) );
  INVX1 U8858 ( .A(n8912), .Y(n8913) );
  BUFX2 U8859 ( .A(fifo[91]), .Y(n8914) );
  INVX1 U8860 ( .A(n8917), .Y(n8915) );
  INVX1 U8861 ( .A(n8915), .Y(n8916) );
  BUFX2 U8862 ( .A(fifo[92]), .Y(n8917) );
  INVX1 U8863 ( .A(n8920), .Y(n8918) );
  INVX1 U8864 ( .A(n8918), .Y(n8919) );
  BUFX2 U8865 ( .A(fifo[93]), .Y(n8920) );
  INVX1 U8866 ( .A(n8923), .Y(n8921) );
  INVX1 U8867 ( .A(n8921), .Y(n8922) );
  BUFX2 U8868 ( .A(fifo[94]), .Y(n8923) );
  INVX1 U8869 ( .A(n8926), .Y(n8924) );
  INVX1 U8870 ( .A(n8924), .Y(n8925) );
  BUFX2 U8871 ( .A(fifo[95]), .Y(n8926) );
  INVX1 U8872 ( .A(n8929), .Y(n8927) );
  INVX1 U8873 ( .A(n8927), .Y(n8928) );
  BUFX2 U8874 ( .A(fifo[96]), .Y(n8929) );
  INVX1 U8875 ( .A(n8932), .Y(n8930) );
  INVX1 U8876 ( .A(n8930), .Y(n8931) );
  BUFX2 U8877 ( .A(fifo[97]), .Y(n8932) );
  INVX1 U8878 ( .A(n8935), .Y(n8933) );
  INVX1 U8879 ( .A(n8933), .Y(n8934) );
  BUFX2 U8880 ( .A(fifo[98]), .Y(n8935) );
  INVX1 U8881 ( .A(n8938), .Y(n8936) );
  INVX1 U8882 ( .A(n8936), .Y(n8937) );
  BUFX2 U8883 ( .A(fifo[99]), .Y(n8938) );
  INVX1 U8884 ( .A(n8941), .Y(n8939) );
  INVX1 U8885 ( .A(n8939), .Y(n8940) );
  BUFX2 U8886 ( .A(fifo[100]), .Y(n8941) );
  INVX1 U8887 ( .A(n8944), .Y(n8942) );
  INVX1 U8888 ( .A(n8942), .Y(n8943) );
  BUFX2 U8889 ( .A(fifo[101]), .Y(n8944) );
  INVX1 U8890 ( .A(n8947), .Y(n8945) );
  INVX1 U8891 ( .A(n8945), .Y(n8946) );
  BUFX2 U8892 ( .A(fifo[136]), .Y(n8947) );
  INVX1 U8893 ( .A(n8950), .Y(n8948) );
  INVX1 U8894 ( .A(n8948), .Y(n8949) );
  BUFX2 U8895 ( .A(fifo[137]), .Y(n8950) );
  INVX1 U8896 ( .A(n8953), .Y(n8951) );
  INVX1 U8897 ( .A(n8951), .Y(n8952) );
  BUFX2 U8898 ( .A(fifo[138]), .Y(n8953) );
  INVX1 U8899 ( .A(n8956), .Y(n8954) );
  INVX1 U8900 ( .A(n8954), .Y(n8955) );
  BUFX2 U8901 ( .A(fifo[139]), .Y(n8956) );
  INVX1 U8902 ( .A(n8959), .Y(n8957) );
  INVX1 U8903 ( .A(n8957), .Y(n8958) );
  BUFX2 U8904 ( .A(fifo[140]), .Y(n8959) );
  INVX1 U8905 ( .A(n8962), .Y(n8960) );
  INVX1 U8906 ( .A(n8960), .Y(n8961) );
  BUFX2 U8907 ( .A(fifo[141]), .Y(n8962) );
  INVX1 U8908 ( .A(n8965), .Y(n8963) );
  INVX1 U8909 ( .A(n8963), .Y(n8964) );
  BUFX2 U8910 ( .A(fifo[142]), .Y(n8965) );
  INVX1 U8911 ( .A(n8968), .Y(n8966) );
  INVX1 U8912 ( .A(n8966), .Y(n8967) );
  BUFX2 U8913 ( .A(fifo[143]), .Y(n8968) );
  INVX1 U8914 ( .A(n8971), .Y(n8969) );
  INVX1 U8915 ( .A(n8969), .Y(n8970) );
  BUFX2 U8916 ( .A(fifo[144]), .Y(n8971) );
  INVX1 U8917 ( .A(n8974), .Y(n8972) );
  INVX1 U8918 ( .A(n8972), .Y(n8973) );
  BUFX2 U8919 ( .A(fifo[145]), .Y(n8974) );
  INVX1 U8920 ( .A(n8977), .Y(n8975) );
  INVX1 U8921 ( .A(n8975), .Y(n8976) );
  BUFX2 U8922 ( .A(fifo[146]), .Y(n8977) );
  INVX1 U8923 ( .A(n8980), .Y(n8978) );
  INVX1 U8924 ( .A(n8978), .Y(n8979) );
  BUFX2 U8925 ( .A(fifo[147]), .Y(n8980) );
  INVX1 U8926 ( .A(n8983), .Y(n8981) );
  INVX1 U8927 ( .A(n8981), .Y(n8982) );
  BUFX2 U8928 ( .A(fifo[148]), .Y(n8983) );
  INVX1 U8929 ( .A(n8986), .Y(n8984) );
  INVX1 U8930 ( .A(n8984), .Y(n8985) );
  BUFX2 U8931 ( .A(fifo[149]), .Y(n8986) );
  INVX1 U8932 ( .A(n8989), .Y(n8987) );
  INVX1 U8933 ( .A(n8987), .Y(n8988) );
  BUFX2 U8934 ( .A(fifo[150]), .Y(n8989) );
  INVX1 U8935 ( .A(n8992), .Y(n8990) );
  INVX1 U8936 ( .A(n8990), .Y(n8991) );
  BUFX2 U8937 ( .A(fifo[151]), .Y(n8992) );
  INVX1 U8938 ( .A(n8995), .Y(n8993) );
  INVX1 U8939 ( .A(n8993), .Y(n8994) );
  BUFX2 U8940 ( .A(fifo[152]), .Y(n8995) );
  INVX1 U8941 ( .A(n8998), .Y(n8996) );
  INVX1 U8942 ( .A(n8996), .Y(n8997) );
  BUFX2 U8943 ( .A(fifo[153]), .Y(n8998) );
  INVX1 U8944 ( .A(n9001), .Y(n8999) );
  INVX1 U8945 ( .A(n8999), .Y(n9000) );
  BUFX2 U8946 ( .A(fifo[154]), .Y(n9001) );
  INVX1 U8947 ( .A(n9004), .Y(n9002) );
  INVX1 U8948 ( .A(n9002), .Y(n9003) );
  BUFX2 U8949 ( .A(fifo[155]), .Y(n9004) );
  INVX1 U8950 ( .A(n9007), .Y(n9005) );
  INVX1 U8951 ( .A(n9005), .Y(n9006) );
  BUFX2 U8952 ( .A(fifo[156]), .Y(n9007) );
  INVX1 U8953 ( .A(n9010), .Y(n9008) );
  INVX1 U8954 ( .A(n9008), .Y(n9009) );
  BUFX2 U8955 ( .A(fifo[157]), .Y(n9010) );
  INVX1 U8956 ( .A(n9013), .Y(n9011) );
  INVX1 U8957 ( .A(n9011), .Y(n9012) );
  BUFX2 U8958 ( .A(fifo[158]), .Y(n9013) );
  INVX1 U8959 ( .A(n9016), .Y(n9014) );
  INVX1 U8960 ( .A(n9014), .Y(n9015) );
  BUFX2 U8961 ( .A(fifo[159]), .Y(n9016) );
  INVX1 U8962 ( .A(n9019), .Y(n9017) );
  INVX1 U8963 ( .A(n9017), .Y(n9018) );
  BUFX2 U8964 ( .A(fifo[160]), .Y(n9019) );
  INVX1 U8965 ( .A(n9022), .Y(n9020) );
  INVX1 U8966 ( .A(n9020), .Y(n9021) );
  BUFX2 U8967 ( .A(fifo[161]), .Y(n9022) );
  INVX1 U8968 ( .A(n9025), .Y(n9023) );
  INVX1 U8969 ( .A(n9023), .Y(n9024) );
  BUFX2 U8970 ( .A(fifo[162]), .Y(n9025) );
  INVX1 U8971 ( .A(n9028), .Y(n9026) );
  INVX1 U8972 ( .A(n9026), .Y(n9027) );
  BUFX2 U8973 ( .A(fifo[163]), .Y(n9028) );
  INVX1 U8974 ( .A(n9031), .Y(n9029) );
  INVX1 U8975 ( .A(n9029), .Y(n9030) );
  BUFX2 U8976 ( .A(fifo[164]), .Y(n9031) );
  INVX1 U8977 ( .A(n9034), .Y(n9032) );
  INVX1 U8978 ( .A(n9032), .Y(n9033) );
  BUFX2 U8979 ( .A(fifo[165]), .Y(n9034) );
  INVX1 U8980 ( .A(n9037), .Y(n9035) );
  INVX1 U8981 ( .A(n9035), .Y(n9036) );
  BUFX2 U8982 ( .A(fifo[166]), .Y(n9037) );
  INVX1 U8983 ( .A(n9040), .Y(n9038) );
  INVX1 U8984 ( .A(n9038), .Y(n9039) );
  BUFX2 U8985 ( .A(fifo[167]), .Y(n9040) );
  INVX1 U8986 ( .A(n9043), .Y(n9041) );
  INVX1 U8987 ( .A(n9041), .Y(n9042) );
  BUFX2 U8988 ( .A(fifo[168]), .Y(n9043) );
  INVX1 U8989 ( .A(n9046), .Y(n9044) );
  INVX1 U8990 ( .A(n9044), .Y(n9045) );
  BUFX2 U8991 ( .A(fifo[169]), .Y(n9046) );
  INVX1 U8992 ( .A(n9049), .Y(n9047) );
  INVX1 U8993 ( .A(n9047), .Y(n9048) );
  BUFX2 U8994 ( .A(fifo[204]), .Y(n9049) );
  INVX1 U8995 ( .A(n9052), .Y(n9050) );
  INVX1 U8996 ( .A(n9050), .Y(n9051) );
  BUFX2 U8997 ( .A(fifo[205]), .Y(n9052) );
  INVX1 U8998 ( .A(n9055), .Y(n9053) );
  INVX1 U8999 ( .A(n9053), .Y(n9054) );
  BUFX2 U9000 ( .A(fifo[206]), .Y(n9055) );
  INVX1 U9001 ( .A(n9058), .Y(n9056) );
  INVX1 U9002 ( .A(n9056), .Y(n9057) );
  BUFX2 U9003 ( .A(fifo[207]), .Y(n9058) );
  INVX1 U9004 ( .A(n9061), .Y(n9059) );
  INVX1 U9005 ( .A(n9059), .Y(n9060) );
  BUFX2 U9006 ( .A(fifo[208]), .Y(n9061) );
  INVX1 U9007 ( .A(n9064), .Y(n9062) );
  INVX1 U9008 ( .A(n9062), .Y(n9063) );
  BUFX2 U9009 ( .A(fifo[209]), .Y(n9064) );
  INVX1 U9010 ( .A(n9067), .Y(n9065) );
  INVX1 U9011 ( .A(n9065), .Y(n9066) );
  BUFX2 U9012 ( .A(fifo[210]), .Y(n9067) );
  INVX1 U9013 ( .A(n9070), .Y(n9068) );
  INVX1 U9014 ( .A(n9068), .Y(n9069) );
  BUFX2 U9015 ( .A(fifo[211]), .Y(n9070) );
  INVX1 U9016 ( .A(n9073), .Y(n9071) );
  INVX1 U9017 ( .A(n9071), .Y(n9072) );
  BUFX2 U9018 ( .A(fifo[212]), .Y(n9073) );
  INVX1 U9019 ( .A(n9076), .Y(n9074) );
  INVX1 U9020 ( .A(n9074), .Y(n9075) );
  BUFX2 U9021 ( .A(fifo[213]), .Y(n9076) );
  INVX1 U9022 ( .A(n9079), .Y(n9077) );
  INVX1 U9023 ( .A(n9077), .Y(n9078) );
  BUFX2 U9024 ( .A(fifo[214]), .Y(n9079) );
  INVX1 U9025 ( .A(n9082), .Y(n9080) );
  INVX1 U9026 ( .A(n9080), .Y(n9081) );
  BUFX2 U9027 ( .A(fifo[215]), .Y(n9082) );
  INVX1 U9028 ( .A(n9085), .Y(n9083) );
  INVX1 U9029 ( .A(n9083), .Y(n9084) );
  BUFX2 U9030 ( .A(fifo[216]), .Y(n9085) );
  INVX1 U9031 ( .A(n9088), .Y(n9086) );
  INVX1 U9032 ( .A(n9086), .Y(n9087) );
  BUFX2 U9033 ( .A(fifo[217]), .Y(n9088) );
  INVX1 U9034 ( .A(n9091), .Y(n9089) );
  INVX1 U9035 ( .A(n9089), .Y(n9090) );
  BUFX2 U9036 ( .A(fifo[218]), .Y(n9091) );
  INVX1 U9037 ( .A(n9094), .Y(n9092) );
  INVX1 U9038 ( .A(n9092), .Y(n9093) );
  BUFX2 U9039 ( .A(fifo[219]), .Y(n9094) );
  INVX1 U9040 ( .A(n9097), .Y(n9095) );
  INVX1 U9041 ( .A(n9095), .Y(n9096) );
  BUFX2 U9042 ( .A(fifo[220]), .Y(n9097) );
  INVX1 U9043 ( .A(n9100), .Y(n9098) );
  INVX1 U9044 ( .A(n9098), .Y(n9099) );
  BUFX2 U9045 ( .A(fifo[221]), .Y(n9100) );
  INVX1 U9046 ( .A(n9103), .Y(n9101) );
  INVX1 U9047 ( .A(n9101), .Y(n9102) );
  BUFX2 U9048 ( .A(fifo[222]), .Y(n9103) );
  INVX1 U9049 ( .A(n9106), .Y(n9104) );
  INVX1 U9050 ( .A(n9104), .Y(n9105) );
  BUFX2 U9051 ( .A(fifo[223]), .Y(n9106) );
  INVX1 U9052 ( .A(n9109), .Y(n9107) );
  INVX1 U9053 ( .A(n9107), .Y(n9108) );
  BUFX2 U9054 ( .A(fifo[224]), .Y(n9109) );
  INVX1 U9055 ( .A(n9112), .Y(n9110) );
  INVX1 U9056 ( .A(n9110), .Y(n9111) );
  BUFX2 U9057 ( .A(fifo[225]), .Y(n9112) );
  INVX1 U9058 ( .A(n9115), .Y(n9113) );
  INVX1 U9059 ( .A(n9113), .Y(n9114) );
  BUFX2 U9060 ( .A(fifo[226]), .Y(n9115) );
  INVX1 U9061 ( .A(n9118), .Y(n9116) );
  INVX1 U9062 ( .A(n9116), .Y(n9117) );
  BUFX2 U9063 ( .A(fifo[227]), .Y(n9118) );
  INVX1 U9064 ( .A(n9121), .Y(n9119) );
  INVX1 U9065 ( .A(n9119), .Y(n9120) );
  BUFX2 U9066 ( .A(fifo[228]), .Y(n9121) );
  INVX1 U9067 ( .A(n9124), .Y(n9122) );
  INVX1 U9068 ( .A(n9122), .Y(n9123) );
  BUFX2 U9069 ( .A(fifo[229]), .Y(n9124) );
  INVX1 U9070 ( .A(n9127), .Y(n9125) );
  INVX1 U9071 ( .A(n9125), .Y(n9126) );
  BUFX2 U9072 ( .A(fifo[230]), .Y(n9127) );
  INVX1 U9073 ( .A(n9130), .Y(n9128) );
  INVX1 U9074 ( .A(n9128), .Y(n9129) );
  BUFX2 U9075 ( .A(fifo[231]), .Y(n9130) );
  INVX1 U9076 ( .A(n9133), .Y(n9131) );
  INVX1 U9077 ( .A(n9131), .Y(n9132) );
  BUFX2 U9078 ( .A(fifo[232]), .Y(n9133) );
  INVX1 U9079 ( .A(n9136), .Y(n9134) );
  INVX1 U9080 ( .A(n9134), .Y(n9135) );
  BUFX2 U9081 ( .A(fifo[233]), .Y(n9136) );
  INVX1 U9082 ( .A(n9139), .Y(n9137) );
  INVX1 U9083 ( .A(n9137), .Y(n9138) );
  BUFX2 U9084 ( .A(fifo[234]), .Y(n9139) );
  INVX1 U9085 ( .A(n9142), .Y(n9140) );
  INVX1 U9086 ( .A(n9140), .Y(n9141) );
  BUFX2 U9087 ( .A(fifo[235]), .Y(n9142) );
  INVX1 U9088 ( .A(n9145), .Y(n9143) );
  INVX1 U9089 ( .A(n9143), .Y(n9144) );
  BUFX2 U9090 ( .A(fifo[236]), .Y(n9145) );
  INVX1 U9091 ( .A(n9148), .Y(n9146) );
  INVX1 U9092 ( .A(n9146), .Y(n9147) );
  BUFX2 U9093 ( .A(fifo[237]), .Y(n9148) );
  INVX1 U9094 ( .A(n9151), .Y(n9149) );
  INVX1 U9095 ( .A(n9149), .Y(n9150) );
  BUFX2 U9096 ( .A(fifo[544]), .Y(n9151) );
  INVX1 U9097 ( .A(n9154), .Y(n9152) );
  INVX1 U9098 ( .A(n9152), .Y(n9153) );
  BUFX2 U9099 ( .A(fifo[545]), .Y(n9154) );
  INVX1 U9100 ( .A(n9157), .Y(n9155) );
  INVX1 U9101 ( .A(n9155), .Y(n9156) );
  BUFX2 U9102 ( .A(fifo[546]), .Y(n9157) );
  INVX1 U9103 ( .A(n9160), .Y(n9158) );
  INVX1 U9104 ( .A(n9158), .Y(n9159) );
  BUFX2 U9105 ( .A(fifo[547]), .Y(n9160) );
  INVX1 U9106 ( .A(n9163), .Y(n9161) );
  INVX1 U9107 ( .A(n9161), .Y(n9162) );
  BUFX2 U9108 ( .A(fifo[548]), .Y(n9163) );
  INVX1 U9109 ( .A(n9166), .Y(n9164) );
  INVX1 U9110 ( .A(n9164), .Y(n9165) );
  BUFX2 U9111 ( .A(fifo[549]), .Y(n9166) );
  INVX1 U9112 ( .A(n9169), .Y(n9167) );
  INVX1 U9113 ( .A(n9167), .Y(n9168) );
  BUFX2 U9114 ( .A(fifo[550]), .Y(n9169) );
  INVX1 U9115 ( .A(n9172), .Y(n9170) );
  INVX1 U9116 ( .A(n9170), .Y(n9171) );
  BUFX2 U9117 ( .A(fifo[551]), .Y(n9172) );
  INVX1 U9118 ( .A(n9175), .Y(n9173) );
  INVX1 U9119 ( .A(n9173), .Y(n9174) );
  BUFX2 U9120 ( .A(fifo[552]), .Y(n9175) );
  INVX1 U9121 ( .A(n9178), .Y(n9176) );
  INVX1 U9122 ( .A(n9176), .Y(n9177) );
  BUFX2 U9123 ( .A(fifo[553]), .Y(n9178) );
  INVX1 U9124 ( .A(n9181), .Y(n9179) );
  INVX1 U9125 ( .A(n9179), .Y(n9180) );
  BUFX2 U9126 ( .A(fifo[554]), .Y(n9181) );
  INVX1 U9127 ( .A(n9184), .Y(n9182) );
  INVX1 U9128 ( .A(n9182), .Y(n9183) );
  BUFX2 U9129 ( .A(fifo[555]), .Y(n9184) );
  INVX1 U9130 ( .A(n9187), .Y(n9185) );
  INVX1 U9131 ( .A(n9185), .Y(n9186) );
  BUFX2 U9132 ( .A(fifo[556]), .Y(n9187) );
  INVX1 U9133 ( .A(n9190), .Y(n9188) );
  INVX1 U9134 ( .A(n9188), .Y(n9189) );
  BUFX2 U9135 ( .A(fifo[557]), .Y(n9190) );
  INVX1 U9136 ( .A(n9193), .Y(n9191) );
  INVX1 U9137 ( .A(n9191), .Y(n9192) );
  BUFX2 U9138 ( .A(fifo[558]), .Y(n9193) );
  INVX1 U9139 ( .A(n9196), .Y(n9194) );
  INVX1 U9140 ( .A(n9194), .Y(n9195) );
  BUFX2 U9141 ( .A(fifo[559]), .Y(n9196) );
  INVX1 U9142 ( .A(n9199), .Y(n9197) );
  INVX1 U9143 ( .A(n9197), .Y(n9198) );
  BUFX2 U9144 ( .A(fifo[560]), .Y(n9199) );
  INVX1 U9145 ( .A(n9202), .Y(n9200) );
  INVX1 U9146 ( .A(n9200), .Y(n9201) );
  BUFX2 U9147 ( .A(fifo[561]), .Y(n9202) );
  INVX1 U9148 ( .A(n9205), .Y(n9203) );
  INVX1 U9149 ( .A(n9203), .Y(n9204) );
  BUFX2 U9150 ( .A(fifo[562]), .Y(n9205) );
  INVX1 U9151 ( .A(n9208), .Y(n9206) );
  INVX1 U9152 ( .A(n9206), .Y(n9207) );
  BUFX2 U9153 ( .A(fifo[563]), .Y(n9208) );
  INVX1 U9154 ( .A(n9211), .Y(n9209) );
  INVX1 U9155 ( .A(n9209), .Y(n9210) );
  BUFX2 U9156 ( .A(fifo[564]), .Y(n9211) );
  INVX1 U9157 ( .A(n9214), .Y(n9212) );
  INVX1 U9158 ( .A(n9212), .Y(n9213) );
  BUFX2 U9159 ( .A(fifo[565]), .Y(n9214) );
  INVX1 U9160 ( .A(n9217), .Y(n9215) );
  INVX1 U9161 ( .A(n9215), .Y(n9216) );
  BUFX2 U9162 ( .A(fifo[566]), .Y(n9217) );
  INVX1 U9163 ( .A(n9220), .Y(n9218) );
  INVX1 U9164 ( .A(n9218), .Y(n9219) );
  BUFX2 U9165 ( .A(fifo[567]), .Y(n9220) );
  INVX1 U9166 ( .A(n9223), .Y(n9221) );
  INVX1 U9167 ( .A(n9221), .Y(n9222) );
  BUFX2 U9168 ( .A(fifo[568]), .Y(n9223) );
  INVX1 U9169 ( .A(n9226), .Y(n9224) );
  INVX1 U9170 ( .A(n9224), .Y(n9225) );
  BUFX2 U9171 ( .A(fifo[569]), .Y(n9226) );
  INVX1 U9172 ( .A(n9229), .Y(n9227) );
  INVX1 U9173 ( .A(n9227), .Y(n9228) );
  BUFX2 U9174 ( .A(fifo[570]), .Y(n9229) );
  INVX1 U9175 ( .A(n9232), .Y(n9230) );
  INVX1 U9176 ( .A(n9230), .Y(n9231) );
  BUFX2 U9177 ( .A(fifo[571]), .Y(n9232) );
  INVX1 U9178 ( .A(n9235), .Y(n9233) );
  INVX1 U9179 ( .A(n9233), .Y(n9234) );
  BUFX2 U9180 ( .A(fifo[572]), .Y(n9235) );
  INVX1 U9181 ( .A(n9238), .Y(n9236) );
  INVX1 U9182 ( .A(n9236), .Y(n9237) );
  BUFX2 U9183 ( .A(fifo[573]), .Y(n9238) );
  INVX1 U9184 ( .A(n9241), .Y(n9239) );
  INVX1 U9185 ( .A(n9239), .Y(n9240) );
  BUFX2 U9186 ( .A(fifo[574]), .Y(n9241) );
  INVX1 U9187 ( .A(n9244), .Y(n9242) );
  INVX1 U9188 ( .A(n9242), .Y(n9243) );
  BUFX2 U9189 ( .A(fifo[575]), .Y(n9244) );
  INVX1 U9190 ( .A(n9247), .Y(n9245) );
  INVX1 U9191 ( .A(n9245), .Y(n9246) );
  BUFX2 U9192 ( .A(fifo[576]), .Y(n9247) );
  INVX1 U9193 ( .A(n9250), .Y(n9248) );
  INVX1 U9194 ( .A(n9248), .Y(n9249) );
  BUFX2 U9195 ( .A(fifo[577]), .Y(n9250) );
  INVX1 U9196 ( .A(n9253), .Y(n9251) );
  INVX1 U9197 ( .A(n9251), .Y(n9252) );
  BUFX2 U9198 ( .A(fifo[612]), .Y(n9253) );
  INVX1 U9199 ( .A(n9256), .Y(n9254) );
  INVX1 U9200 ( .A(n9254), .Y(n9255) );
  BUFX2 U9201 ( .A(fifo[613]), .Y(n9256) );
  INVX1 U9202 ( .A(n9259), .Y(n9257) );
  INVX1 U9203 ( .A(n9257), .Y(n9258) );
  BUFX2 U9204 ( .A(fifo[614]), .Y(n9259) );
  INVX1 U9205 ( .A(n9262), .Y(n9260) );
  INVX1 U9206 ( .A(n9260), .Y(n9261) );
  BUFX2 U9207 ( .A(fifo[615]), .Y(n9262) );
  INVX1 U9208 ( .A(n9265), .Y(n9263) );
  INVX1 U9209 ( .A(n9263), .Y(n9264) );
  BUFX2 U9210 ( .A(fifo[616]), .Y(n9265) );
  INVX1 U9211 ( .A(n9268), .Y(n9266) );
  INVX1 U9212 ( .A(n9266), .Y(n9267) );
  BUFX2 U9213 ( .A(fifo[617]), .Y(n9268) );
  INVX1 U9214 ( .A(n9271), .Y(n9269) );
  INVX1 U9215 ( .A(n9269), .Y(n9270) );
  BUFX2 U9216 ( .A(fifo[618]), .Y(n9271) );
  INVX1 U9217 ( .A(n9274), .Y(n9272) );
  INVX1 U9218 ( .A(n9272), .Y(n9273) );
  BUFX2 U9219 ( .A(fifo[619]), .Y(n9274) );
  INVX1 U9220 ( .A(n9277), .Y(n9275) );
  INVX1 U9221 ( .A(n9275), .Y(n9276) );
  BUFX2 U9222 ( .A(fifo[620]), .Y(n9277) );
  INVX1 U9223 ( .A(n9280), .Y(n9278) );
  INVX1 U9224 ( .A(n9278), .Y(n9279) );
  BUFX2 U9225 ( .A(fifo[621]), .Y(n9280) );
  INVX1 U9226 ( .A(n9283), .Y(n9281) );
  INVX1 U9227 ( .A(n9281), .Y(n9282) );
  BUFX2 U9228 ( .A(fifo[622]), .Y(n9283) );
  INVX1 U9229 ( .A(n9286), .Y(n9284) );
  INVX1 U9230 ( .A(n9284), .Y(n9285) );
  BUFX2 U9231 ( .A(fifo[623]), .Y(n9286) );
  INVX1 U9232 ( .A(n9289), .Y(n9287) );
  INVX1 U9233 ( .A(n9287), .Y(n9288) );
  BUFX2 U9234 ( .A(fifo[624]), .Y(n9289) );
  INVX1 U9235 ( .A(n9292), .Y(n9290) );
  INVX1 U9236 ( .A(n9290), .Y(n9291) );
  BUFX2 U9237 ( .A(fifo[625]), .Y(n9292) );
  INVX1 U9238 ( .A(n9295), .Y(n9293) );
  INVX1 U9239 ( .A(n9293), .Y(n9294) );
  BUFX2 U9240 ( .A(fifo[626]), .Y(n9295) );
  INVX1 U9241 ( .A(n9298), .Y(n9296) );
  INVX1 U9242 ( .A(n9296), .Y(n9297) );
  BUFX2 U9243 ( .A(fifo[627]), .Y(n9298) );
  INVX1 U9244 ( .A(n9301), .Y(n9299) );
  INVX1 U9245 ( .A(n9299), .Y(n9300) );
  BUFX2 U9246 ( .A(fifo[628]), .Y(n9301) );
  INVX1 U9247 ( .A(n9304), .Y(n9302) );
  INVX1 U9248 ( .A(n9302), .Y(n9303) );
  BUFX2 U9249 ( .A(fifo[629]), .Y(n9304) );
  INVX1 U9250 ( .A(n9307), .Y(n9305) );
  INVX1 U9251 ( .A(n9305), .Y(n9306) );
  BUFX2 U9252 ( .A(fifo[630]), .Y(n9307) );
  INVX1 U9253 ( .A(n9310), .Y(n9308) );
  INVX1 U9254 ( .A(n9308), .Y(n9309) );
  BUFX2 U9255 ( .A(fifo[631]), .Y(n9310) );
  INVX1 U9256 ( .A(n9313), .Y(n9311) );
  INVX1 U9257 ( .A(n9311), .Y(n9312) );
  BUFX2 U9258 ( .A(fifo[632]), .Y(n9313) );
  INVX1 U9259 ( .A(n9316), .Y(n9314) );
  INVX1 U9260 ( .A(n9314), .Y(n9315) );
  BUFX2 U9261 ( .A(fifo[633]), .Y(n9316) );
  INVX1 U9262 ( .A(n9319), .Y(n9317) );
  INVX1 U9263 ( .A(n9317), .Y(n9318) );
  BUFX2 U9264 ( .A(fifo[634]), .Y(n9319) );
  INVX1 U9265 ( .A(n9322), .Y(n9320) );
  INVX1 U9266 ( .A(n9320), .Y(n9321) );
  BUFX2 U9267 ( .A(fifo[635]), .Y(n9322) );
  INVX1 U9268 ( .A(n9325), .Y(n9323) );
  INVX1 U9269 ( .A(n9323), .Y(n9324) );
  BUFX2 U9270 ( .A(fifo[636]), .Y(n9325) );
  INVX1 U9271 ( .A(n9328), .Y(n9326) );
  INVX1 U9272 ( .A(n9326), .Y(n9327) );
  BUFX2 U9273 ( .A(fifo[637]), .Y(n9328) );
  INVX1 U9274 ( .A(n9331), .Y(n9329) );
  INVX1 U9275 ( .A(n9329), .Y(n9330) );
  BUFX2 U9276 ( .A(fifo[638]), .Y(n9331) );
  INVX1 U9277 ( .A(n9334), .Y(n9332) );
  INVX1 U9278 ( .A(n9332), .Y(n9333) );
  BUFX2 U9279 ( .A(fifo[639]), .Y(n9334) );
  INVX1 U9280 ( .A(n9337), .Y(n9335) );
  INVX1 U9281 ( .A(n9335), .Y(n9336) );
  BUFX2 U9282 ( .A(fifo[640]), .Y(n9337) );
  INVX1 U9283 ( .A(n9340), .Y(n9338) );
  INVX1 U9284 ( .A(n9338), .Y(n9339) );
  BUFX2 U9285 ( .A(fifo[641]), .Y(n9340) );
  INVX1 U9286 ( .A(n9343), .Y(n9341) );
  INVX1 U9287 ( .A(n9341), .Y(n9342) );
  BUFX2 U9288 ( .A(fifo[642]), .Y(n9343) );
  INVX1 U9289 ( .A(n9346), .Y(n9344) );
  INVX1 U9290 ( .A(n9344), .Y(n9345) );
  BUFX2 U9291 ( .A(fifo[643]), .Y(n9346) );
  INVX1 U9292 ( .A(n9349), .Y(n9347) );
  INVX1 U9293 ( .A(n9347), .Y(n9348) );
  BUFX2 U9294 ( .A(fifo[644]), .Y(n9349) );
  INVX1 U9295 ( .A(n9352), .Y(n9350) );
  INVX1 U9296 ( .A(n9350), .Y(n9351) );
  BUFX2 U9297 ( .A(fifo[645]), .Y(n9352) );
  INVX1 U9298 ( .A(n9355), .Y(n9353) );
  INVX1 U9299 ( .A(n9353), .Y(n9354) );
  BUFX2 U9300 ( .A(fifo[680]), .Y(n9355) );
  INVX1 U9301 ( .A(n9358), .Y(n9356) );
  INVX1 U9302 ( .A(n9356), .Y(n9357) );
  BUFX2 U9303 ( .A(fifo[681]), .Y(n9358) );
  INVX1 U9304 ( .A(n9361), .Y(n9359) );
  INVX1 U9305 ( .A(n9359), .Y(n9360) );
  BUFX2 U9306 ( .A(fifo[682]), .Y(n9361) );
  INVX1 U9307 ( .A(n9364), .Y(n9362) );
  INVX1 U9308 ( .A(n9362), .Y(n9363) );
  BUFX2 U9309 ( .A(fifo[683]), .Y(n9364) );
  INVX1 U9310 ( .A(n9367), .Y(n9365) );
  INVX1 U9311 ( .A(n9365), .Y(n9366) );
  BUFX2 U9312 ( .A(fifo[684]), .Y(n9367) );
  INVX1 U9313 ( .A(n9370), .Y(n9368) );
  INVX1 U9314 ( .A(n9368), .Y(n9369) );
  BUFX2 U9315 ( .A(fifo[685]), .Y(n9370) );
  INVX1 U9316 ( .A(n9373), .Y(n9371) );
  INVX1 U9317 ( .A(n9371), .Y(n9372) );
  BUFX2 U9318 ( .A(fifo[686]), .Y(n9373) );
  INVX1 U9319 ( .A(n9376), .Y(n9374) );
  INVX1 U9320 ( .A(n9374), .Y(n9375) );
  BUFX2 U9321 ( .A(fifo[687]), .Y(n9376) );
  INVX1 U9322 ( .A(n9379), .Y(n9377) );
  INVX1 U9323 ( .A(n9377), .Y(n9378) );
  BUFX2 U9324 ( .A(fifo[688]), .Y(n9379) );
  INVX1 U9325 ( .A(n9382), .Y(n9380) );
  INVX1 U9326 ( .A(n9380), .Y(n9381) );
  BUFX2 U9327 ( .A(fifo[689]), .Y(n9382) );
  INVX1 U9328 ( .A(n9385), .Y(n9383) );
  INVX1 U9329 ( .A(n9383), .Y(n9384) );
  BUFX2 U9330 ( .A(fifo[690]), .Y(n9385) );
  INVX1 U9331 ( .A(n9388), .Y(n9386) );
  INVX1 U9332 ( .A(n9386), .Y(n9387) );
  BUFX2 U9333 ( .A(fifo[691]), .Y(n9388) );
  INVX1 U9334 ( .A(n9391), .Y(n9389) );
  INVX1 U9335 ( .A(n9389), .Y(n9390) );
  BUFX2 U9336 ( .A(fifo[692]), .Y(n9391) );
  INVX1 U9337 ( .A(n9394), .Y(n9392) );
  INVX1 U9338 ( .A(n9392), .Y(n9393) );
  BUFX2 U9339 ( .A(fifo[693]), .Y(n9394) );
  INVX1 U9340 ( .A(n9397), .Y(n9395) );
  INVX1 U9341 ( .A(n9395), .Y(n9396) );
  BUFX2 U9342 ( .A(fifo[694]), .Y(n9397) );
  INVX1 U9343 ( .A(n9400), .Y(n9398) );
  INVX1 U9344 ( .A(n9398), .Y(n9399) );
  BUFX2 U9345 ( .A(fifo[695]), .Y(n9400) );
  INVX1 U9346 ( .A(n9403), .Y(n9401) );
  INVX1 U9347 ( .A(n9401), .Y(n9402) );
  BUFX2 U9348 ( .A(fifo[696]), .Y(n9403) );
  INVX1 U9349 ( .A(n9406), .Y(n9404) );
  INVX1 U9350 ( .A(n9404), .Y(n9405) );
  BUFX2 U9351 ( .A(fifo[697]), .Y(n9406) );
  INVX1 U9352 ( .A(n9409), .Y(n9407) );
  INVX1 U9353 ( .A(n9407), .Y(n9408) );
  BUFX2 U9354 ( .A(fifo[698]), .Y(n9409) );
  INVX1 U9355 ( .A(n9412), .Y(n9410) );
  INVX1 U9356 ( .A(n9410), .Y(n9411) );
  BUFX2 U9357 ( .A(fifo[699]), .Y(n9412) );
  INVX1 U9358 ( .A(n9415), .Y(n9413) );
  INVX1 U9359 ( .A(n9413), .Y(n9414) );
  BUFX2 U9360 ( .A(fifo[700]), .Y(n9415) );
  INVX1 U9361 ( .A(n9418), .Y(n9416) );
  INVX1 U9362 ( .A(n9416), .Y(n9417) );
  BUFX2 U9363 ( .A(fifo[701]), .Y(n9418) );
  INVX1 U9364 ( .A(n9421), .Y(n9419) );
  INVX1 U9365 ( .A(n9419), .Y(n9420) );
  BUFX2 U9366 ( .A(fifo[702]), .Y(n9421) );
  INVX1 U9367 ( .A(n9424), .Y(n9422) );
  INVX1 U9368 ( .A(n9422), .Y(n9423) );
  BUFX2 U9369 ( .A(fifo[703]), .Y(n9424) );
  INVX1 U9370 ( .A(n9427), .Y(n9425) );
  INVX1 U9371 ( .A(n9425), .Y(n9426) );
  BUFX2 U9372 ( .A(fifo[704]), .Y(n9427) );
  INVX1 U9373 ( .A(n9430), .Y(n9428) );
  INVX1 U9374 ( .A(n9428), .Y(n9429) );
  BUFX2 U9375 ( .A(fifo[705]), .Y(n9430) );
  INVX1 U9376 ( .A(n9433), .Y(n9431) );
  INVX1 U9377 ( .A(n9431), .Y(n9432) );
  BUFX2 U9378 ( .A(fifo[706]), .Y(n9433) );
  INVX1 U9379 ( .A(n9436), .Y(n9434) );
  INVX1 U9380 ( .A(n9434), .Y(n9435) );
  BUFX2 U9381 ( .A(fifo[707]), .Y(n9436) );
  INVX1 U9382 ( .A(n9439), .Y(n9437) );
  INVX1 U9383 ( .A(n9437), .Y(n9438) );
  BUFX2 U9384 ( .A(fifo[708]), .Y(n9439) );
  INVX1 U9385 ( .A(n9442), .Y(n9440) );
  INVX1 U9386 ( .A(n9440), .Y(n9441) );
  BUFX2 U9387 ( .A(fifo[709]), .Y(n9442) );
  INVX1 U9388 ( .A(n9445), .Y(n9443) );
  INVX1 U9389 ( .A(n9443), .Y(n9444) );
  BUFX2 U9390 ( .A(fifo[710]), .Y(n9445) );
  INVX1 U9391 ( .A(n9448), .Y(n9446) );
  INVX1 U9392 ( .A(n9446), .Y(n9447) );
  BUFX2 U9393 ( .A(fifo[711]), .Y(n9448) );
  INVX1 U9394 ( .A(n9451), .Y(n9449) );
  INVX1 U9395 ( .A(n9449), .Y(n9450) );
  BUFX2 U9396 ( .A(fifo[712]), .Y(n9451) );
  INVX1 U9397 ( .A(n9454), .Y(n9452) );
  INVX1 U9398 ( .A(n9452), .Y(n9453) );
  BUFX2 U9399 ( .A(fifo[713]), .Y(n9454) );
  INVX1 U9400 ( .A(n9457), .Y(n9455) );
  INVX1 U9401 ( .A(n9455), .Y(n9456) );
  BUFX2 U9402 ( .A(fifo[748]), .Y(n9457) );
  INVX1 U9403 ( .A(n9460), .Y(n9458) );
  INVX1 U9404 ( .A(n9458), .Y(n9459) );
  BUFX2 U9405 ( .A(fifo[749]), .Y(n9460) );
  INVX1 U9406 ( .A(n9463), .Y(n9461) );
  INVX1 U9407 ( .A(n9461), .Y(n9462) );
  BUFX2 U9408 ( .A(fifo[750]), .Y(n9463) );
  INVX1 U9409 ( .A(n9466), .Y(n9464) );
  INVX1 U9410 ( .A(n9464), .Y(n9465) );
  BUFX2 U9411 ( .A(fifo[751]), .Y(n9466) );
  INVX1 U9412 ( .A(n9469), .Y(n9467) );
  INVX1 U9413 ( .A(n9467), .Y(n9468) );
  BUFX2 U9414 ( .A(fifo[752]), .Y(n9469) );
  INVX1 U9415 ( .A(n9472), .Y(n9470) );
  INVX1 U9416 ( .A(n9470), .Y(n9471) );
  BUFX2 U9417 ( .A(fifo[753]), .Y(n9472) );
  INVX1 U9418 ( .A(n9475), .Y(n9473) );
  INVX1 U9419 ( .A(n9473), .Y(n9474) );
  BUFX2 U9420 ( .A(fifo[754]), .Y(n9475) );
  INVX1 U9421 ( .A(n9478), .Y(n9476) );
  INVX1 U9422 ( .A(n9476), .Y(n9477) );
  BUFX2 U9423 ( .A(fifo[755]), .Y(n9478) );
  INVX1 U9424 ( .A(n9481), .Y(n9479) );
  INVX1 U9425 ( .A(n9479), .Y(n9480) );
  BUFX2 U9426 ( .A(fifo[756]), .Y(n9481) );
  INVX1 U9427 ( .A(n9484), .Y(n9482) );
  INVX1 U9428 ( .A(n9482), .Y(n9483) );
  BUFX2 U9429 ( .A(fifo[757]), .Y(n9484) );
  INVX1 U9430 ( .A(n9487), .Y(n9485) );
  INVX1 U9431 ( .A(n9485), .Y(n9486) );
  BUFX2 U9432 ( .A(fifo[758]), .Y(n9487) );
  INVX1 U9433 ( .A(n9490), .Y(n9488) );
  INVX1 U9434 ( .A(n9488), .Y(n9489) );
  BUFX2 U9435 ( .A(fifo[759]), .Y(n9490) );
  INVX1 U9436 ( .A(n9493), .Y(n9491) );
  INVX1 U9437 ( .A(n9491), .Y(n9492) );
  BUFX2 U9438 ( .A(fifo[760]), .Y(n9493) );
  INVX1 U9439 ( .A(n9496), .Y(n9494) );
  INVX1 U9440 ( .A(n9494), .Y(n9495) );
  BUFX2 U9441 ( .A(fifo[761]), .Y(n9496) );
  INVX1 U9442 ( .A(n9499), .Y(n9497) );
  INVX1 U9443 ( .A(n9497), .Y(n9498) );
  BUFX2 U9444 ( .A(fifo[762]), .Y(n9499) );
  INVX1 U9445 ( .A(n9502), .Y(n9500) );
  INVX1 U9446 ( .A(n9500), .Y(n9501) );
  BUFX2 U9447 ( .A(fifo[763]), .Y(n9502) );
  INVX1 U9448 ( .A(n9505), .Y(n9503) );
  INVX1 U9449 ( .A(n9503), .Y(n9504) );
  BUFX2 U9450 ( .A(fifo[764]), .Y(n9505) );
  INVX1 U9451 ( .A(n9508), .Y(n9506) );
  INVX1 U9452 ( .A(n9506), .Y(n9507) );
  BUFX2 U9453 ( .A(fifo[765]), .Y(n9508) );
  INVX1 U9454 ( .A(n9511), .Y(n9509) );
  INVX1 U9455 ( .A(n9509), .Y(n9510) );
  BUFX2 U9456 ( .A(fifo[766]), .Y(n9511) );
  INVX1 U9457 ( .A(n9514), .Y(n9512) );
  INVX1 U9458 ( .A(n9512), .Y(n9513) );
  BUFX2 U9459 ( .A(fifo[767]), .Y(n9514) );
  INVX1 U9460 ( .A(n9517), .Y(n9515) );
  INVX1 U9461 ( .A(n9515), .Y(n9516) );
  BUFX2 U9462 ( .A(fifo[768]), .Y(n9517) );
  INVX1 U9463 ( .A(n9520), .Y(n9518) );
  INVX1 U9464 ( .A(n9518), .Y(n9519) );
  BUFX2 U9465 ( .A(fifo[769]), .Y(n9520) );
  INVX1 U9466 ( .A(n9523), .Y(n9521) );
  INVX1 U9467 ( .A(n9521), .Y(n9522) );
  BUFX2 U9468 ( .A(fifo[770]), .Y(n9523) );
  INVX1 U9469 ( .A(n9526), .Y(n9524) );
  INVX1 U9470 ( .A(n9524), .Y(n9525) );
  BUFX2 U9471 ( .A(fifo[771]), .Y(n9526) );
  INVX1 U9472 ( .A(n9529), .Y(n9527) );
  INVX1 U9473 ( .A(n9527), .Y(n9528) );
  BUFX2 U9474 ( .A(fifo[772]), .Y(n9529) );
  INVX1 U9475 ( .A(n9532), .Y(n9530) );
  INVX1 U9476 ( .A(n9530), .Y(n9531) );
  BUFX2 U9477 ( .A(fifo[773]), .Y(n9532) );
  INVX1 U9478 ( .A(n9535), .Y(n9533) );
  INVX1 U9479 ( .A(n9533), .Y(n9534) );
  BUFX2 U9480 ( .A(fifo[774]), .Y(n9535) );
  INVX1 U9481 ( .A(n9538), .Y(n9536) );
  INVX1 U9482 ( .A(n9536), .Y(n9537) );
  BUFX2 U9483 ( .A(fifo[775]), .Y(n9538) );
  INVX1 U9484 ( .A(n9541), .Y(n9539) );
  INVX1 U9485 ( .A(n9539), .Y(n9540) );
  BUFX2 U9486 ( .A(fifo[776]), .Y(n9541) );
  INVX1 U9487 ( .A(n9544), .Y(n9542) );
  INVX1 U9488 ( .A(n9542), .Y(n9543) );
  BUFX2 U9489 ( .A(fifo[777]), .Y(n9544) );
  INVX1 U9490 ( .A(n9547), .Y(n9545) );
  INVX1 U9491 ( .A(n9545), .Y(n9546) );
  BUFX2 U9492 ( .A(fifo[778]), .Y(n9547) );
  INVX1 U9493 ( .A(n9550), .Y(n9548) );
  INVX1 U9494 ( .A(n9548), .Y(n9549) );
  BUFX2 U9495 ( .A(fifo[779]), .Y(n9550) );
  INVX1 U9496 ( .A(n9553), .Y(n9551) );
  INVX1 U9497 ( .A(n9551), .Y(n9552) );
  BUFX2 U9498 ( .A(fifo[780]), .Y(n9553) );
  INVX1 U9499 ( .A(n9556), .Y(n9554) );
  INVX1 U9500 ( .A(n9554), .Y(n9555) );
  BUFX2 U9501 ( .A(fifo[781]), .Y(n9556) );
  INVX1 U9502 ( .A(n9559), .Y(n9557) );
  INVX1 U9503 ( .A(n9557), .Y(n9558) );
  BUFX2 U9504 ( .A(fifo[816]), .Y(n9559) );
  INVX1 U9505 ( .A(n9562), .Y(n9560) );
  INVX1 U9506 ( .A(n9560), .Y(n9561) );
  BUFX2 U9507 ( .A(fifo[817]), .Y(n9562) );
  INVX1 U9508 ( .A(n9565), .Y(n9563) );
  INVX1 U9509 ( .A(n9563), .Y(n9564) );
  BUFX2 U9510 ( .A(fifo[818]), .Y(n9565) );
  INVX1 U9511 ( .A(n9568), .Y(n9566) );
  INVX1 U9512 ( .A(n9566), .Y(n9567) );
  BUFX2 U9513 ( .A(fifo[819]), .Y(n9568) );
  INVX1 U9514 ( .A(n9571), .Y(n9569) );
  INVX1 U9515 ( .A(n9569), .Y(n9570) );
  BUFX2 U9516 ( .A(fifo[820]), .Y(n9571) );
  INVX1 U9517 ( .A(n9574), .Y(n9572) );
  INVX1 U9518 ( .A(n9572), .Y(n9573) );
  BUFX2 U9519 ( .A(fifo[821]), .Y(n9574) );
  INVX1 U9520 ( .A(n9577), .Y(n9575) );
  INVX1 U9521 ( .A(n9575), .Y(n9576) );
  BUFX2 U9522 ( .A(fifo[822]), .Y(n9577) );
  INVX1 U9523 ( .A(n9580), .Y(n9578) );
  INVX1 U9524 ( .A(n9578), .Y(n9579) );
  BUFX2 U9525 ( .A(fifo[823]), .Y(n9580) );
  INVX1 U9526 ( .A(n9583), .Y(n9581) );
  INVX1 U9527 ( .A(n9581), .Y(n9582) );
  BUFX2 U9528 ( .A(fifo[824]), .Y(n9583) );
  INVX1 U9529 ( .A(n9586), .Y(n9584) );
  INVX1 U9530 ( .A(n9584), .Y(n9585) );
  BUFX2 U9531 ( .A(fifo[825]), .Y(n9586) );
  INVX1 U9532 ( .A(n9589), .Y(n9587) );
  INVX1 U9533 ( .A(n9587), .Y(n9588) );
  BUFX2 U9534 ( .A(fifo[826]), .Y(n9589) );
  INVX1 U9535 ( .A(n9592), .Y(n9590) );
  INVX1 U9536 ( .A(n9590), .Y(n9591) );
  BUFX2 U9537 ( .A(fifo[827]), .Y(n9592) );
  INVX1 U9538 ( .A(n9595), .Y(n9593) );
  INVX1 U9539 ( .A(n9593), .Y(n9594) );
  BUFX2 U9540 ( .A(fifo[828]), .Y(n9595) );
  INVX1 U9541 ( .A(n9598), .Y(n9596) );
  INVX1 U9542 ( .A(n9596), .Y(n9597) );
  BUFX2 U9543 ( .A(fifo[829]), .Y(n9598) );
  INVX1 U9544 ( .A(n9601), .Y(n9599) );
  INVX1 U9545 ( .A(n9599), .Y(n9600) );
  BUFX2 U9546 ( .A(fifo[830]), .Y(n9601) );
  INVX1 U9547 ( .A(n9604), .Y(n9602) );
  INVX1 U9548 ( .A(n9602), .Y(n9603) );
  BUFX2 U9549 ( .A(fifo[831]), .Y(n9604) );
  INVX1 U9550 ( .A(n9607), .Y(n9605) );
  INVX1 U9551 ( .A(n9605), .Y(n9606) );
  BUFX2 U9552 ( .A(fifo[832]), .Y(n9607) );
  INVX1 U9553 ( .A(n9610), .Y(n9608) );
  INVX1 U9554 ( .A(n9608), .Y(n9609) );
  BUFX2 U9555 ( .A(fifo[833]), .Y(n9610) );
  INVX1 U9556 ( .A(n9613), .Y(n9611) );
  INVX1 U9557 ( .A(n9611), .Y(n9612) );
  BUFX2 U9558 ( .A(fifo[834]), .Y(n9613) );
  INVX1 U9559 ( .A(n9616), .Y(n9614) );
  INVX1 U9560 ( .A(n9614), .Y(n9615) );
  BUFX2 U9561 ( .A(fifo[835]), .Y(n9616) );
  INVX1 U9562 ( .A(n9619), .Y(n9617) );
  INVX1 U9563 ( .A(n9617), .Y(n9618) );
  BUFX2 U9564 ( .A(fifo[836]), .Y(n9619) );
  INVX1 U9565 ( .A(n9622), .Y(n9620) );
  INVX1 U9566 ( .A(n9620), .Y(n9621) );
  BUFX2 U9567 ( .A(fifo[837]), .Y(n9622) );
  INVX1 U9568 ( .A(n9625), .Y(n9623) );
  INVX1 U9569 ( .A(n9623), .Y(n9624) );
  BUFX2 U9570 ( .A(fifo[838]), .Y(n9625) );
  INVX1 U9571 ( .A(n9628), .Y(n9626) );
  INVX1 U9572 ( .A(n9626), .Y(n9627) );
  BUFX2 U9573 ( .A(fifo[839]), .Y(n9628) );
  INVX1 U9574 ( .A(n9631), .Y(n9629) );
  INVX1 U9575 ( .A(n9629), .Y(n9630) );
  BUFX2 U9576 ( .A(fifo[840]), .Y(n9631) );
  INVX1 U9577 ( .A(n9634), .Y(n9632) );
  INVX1 U9578 ( .A(n9632), .Y(n9633) );
  BUFX2 U9579 ( .A(fifo[841]), .Y(n9634) );
  INVX1 U9580 ( .A(n9637), .Y(n9635) );
  INVX1 U9581 ( .A(n9635), .Y(n9636) );
  BUFX2 U9582 ( .A(fifo[842]), .Y(n9637) );
  INVX1 U9583 ( .A(n9640), .Y(n9638) );
  INVX1 U9584 ( .A(n9638), .Y(n9639) );
  BUFX2 U9585 ( .A(fifo[843]), .Y(n9640) );
  INVX1 U9586 ( .A(n9643), .Y(n9641) );
  INVX1 U9587 ( .A(n9641), .Y(n9642) );
  BUFX2 U9588 ( .A(fifo[844]), .Y(n9643) );
  INVX1 U9589 ( .A(n9646), .Y(n9644) );
  INVX1 U9590 ( .A(n9644), .Y(n9645) );
  BUFX2 U9591 ( .A(fifo[845]), .Y(n9646) );
  INVX1 U9592 ( .A(n9649), .Y(n9647) );
  INVX1 U9593 ( .A(n9647), .Y(n9648) );
  BUFX2 U9594 ( .A(fifo[846]), .Y(n9649) );
  INVX1 U9595 ( .A(n9652), .Y(n9650) );
  INVX1 U9596 ( .A(n9650), .Y(n9651) );
  BUFX2 U9597 ( .A(fifo[847]), .Y(n9652) );
  INVX1 U9598 ( .A(n9655), .Y(n9653) );
  INVX1 U9599 ( .A(n9653), .Y(n9654) );
  BUFX2 U9600 ( .A(fifo[848]), .Y(n9655) );
  INVX1 U9601 ( .A(n9658), .Y(n9656) );
  INVX1 U9602 ( .A(n9656), .Y(n9657) );
  BUFX2 U9603 ( .A(fifo[849]), .Y(n9658) );
  INVX1 U9604 ( .A(n9661), .Y(n9659) );
  INVX1 U9605 ( .A(n9659), .Y(n9660) );
  BUFX2 U9606 ( .A(fifo[884]), .Y(n9661) );
  INVX1 U9607 ( .A(n9664), .Y(n9662) );
  INVX1 U9608 ( .A(n9662), .Y(n9663) );
  BUFX2 U9609 ( .A(fifo[885]), .Y(n9664) );
  INVX1 U9610 ( .A(n9667), .Y(n9665) );
  INVX1 U9611 ( .A(n9665), .Y(n9666) );
  BUFX2 U9612 ( .A(fifo[886]), .Y(n9667) );
  INVX1 U9613 ( .A(n9670), .Y(n9668) );
  INVX1 U9614 ( .A(n9668), .Y(n9669) );
  BUFX2 U9615 ( .A(fifo[887]), .Y(n9670) );
  INVX1 U9616 ( .A(n9673), .Y(n9671) );
  INVX1 U9617 ( .A(n9671), .Y(n9672) );
  BUFX2 U9618 ( .A(fifo[888]), .Y(n9673) );
  INVX1 U9619 ( .A(n9676), .Y(n9674) );
  INVX1 U9620 ( .A(n9674), .Y(n9675) );
  BUFX2 U9621 ( .A(fifo[889]), .Y(n9676) );
  INVX1 U9622 ( .A(n9679), .Y(n9677) );
  INVX1 U9623 ( .A(n9677), .Y(n9678) );
  BUFX2 U9624 ( .A(fifo[890]), .Y(n9679) );
  INVX1 U9625 ( .A(n9682), .Y(n9680) );
  INVX1 U9626 ( .A(n9680), .Y(n9681) );
  BUFX2 U9627 ( .A(fifo[891]), .Y(n9682) );
  INVX1 U9628 ( .A(n9685), .Y(n9683) );
  INVX1 U9629 ( .A(n9683), .Y(n9684) );
  BUFX2 U9630 ( .A(fifo[892]), .Y(n9685) );
  INVX1 U9631 ( .A(n9688), .Y(n9686) );
  INVX1 U9632 ( .A(n9686), .Y(n9687) );
  BUFX2 U9633 ( .A(fifo[893]), .Y(n9688) );
  INVX1 U9634 ( .A(n9691), .Y(n9689) );
  INVX1 U9635 ( .A(n9689), .Y(n9690) );
  BUFX2 U9636 ( .A(fifo[894]), .Y(n9691) );
  INVX1 U9637 ( .A(n9694), .Y(n9692) );
  INVX1 U9638 ( .A(n9692), .Y(n9693) );
  BUFX2 U9639 ( .A(fifo[895]), .Y(n9694) );
  INVX1 U9640 ( .A(n9697), .Y(n9695) );
  INVX1 U9641 ( .A(n9695), .Y(n9696) );
  BUFX2 U9642 ( .A(fifo[896]), .Y(n9697) );
  INVX1 U9643 ( .A(n9700), .Y(n9698) );
  INVX1 U9644 ( .A(n9698), .Y(n9699) );
  BUFX2 U9645 ( .A(fifo[897]), .Y(n9700) );
  INVX1 U9646 ( .A(n9703), .Y(n9701) );
  INVX1 U9647 ( .A(n9701), .Y(n9702) );
  BUFX2 U9648 ( .A(fifo[898]), .Y(n9703) );
  INVX1 U9649 ( .A(n9706), .Y(n9704) );
  INVX1 U9650 ( .A(n9704), .Y(n9705) );
  BUFX2 U9651 ( .A(fifo[899]), .Y(n9706) );
  INVX1 U9652 ( .A(n9709), .Y(n9707) );
  INVX1 U9653 ( .A(n9707), .Y(n9708) );
  BUFX2 U9654 ( .A(fifo[900]), .Y(n9709) );
  INVX1 U9655 ( .A(n9712), .Y(n9710) );
  INVX1 U9656 ( .A(n9710), .Y(n9711) );
  BUFX2 U9657 ( .A(fifo[901]), .Y(n9712) );
  INVX1 U9658 ( .A(n9715), .Y(n9713) );
  INVX1 U9659 ( .A(n9713), .Y(n9714) );
  BUFX2 U9660 ( .A(fifo[902]), .Y(n9715) );
  INVX1 U9661 ( .A(n9718), .Y(n9716) );
  INVX1 U9662 ( .A(n9716), .Y(n9717) );
  BUFX2 U9663 ( .A(fifo[903]), .Y(n9718) );
  INVX1 U9664 ( .A(n9721), .Y(n9719) );
  INVX1 U9665 ( .A(n9719), .Y(n9720) );
  BUFX2 U9666 ( .A(fifo[904]), .Y(n9721) );
  INVX1 U9667 ( .A(n9724), .Y(n9722) );
  INVX1 U9668 ( .A(n9722), .Y(n9723) );
  BUFX2 U9669 ( .A(fifo[905]), .Y(n9724) );
  INVX1 U9670 ( .A(n9727), .Y(n9725) );
  INVX1 U9671 ( .A(n9725), .Y(n9726) );
  BUFX2 U9672 ( .A(fifo[906]), .Y(n9727) );
  INVX1 U9673 ( .A(n9730), .Y(n9728) );
  INVX1 U9674 ( .A(n9728), .Y(n9729) );
  BUFX2 U9675 ( .A(fifo[907]), .Y(n9730) );
  INVX1 U9676 ( .A(n9733), .Y(n9731) );
  INVX1 U9677 ( .A(n9731), .Y(n9732) );
  BUFX2 U9678 ( .A(fifo[908]), .Y(n9733) );
  INVX1 U9679 ( .A(n9736), .Y(n9734) );
  INVX1 U9680 ( .A(n9734), .Y(n9735) );
  BUFX2 U9681 ( .A(fifo[909]), .Y(n9736) );
  INVX1 U9682 ( .A(n9739), .Y(n9737) );
  INVX1 U9683 ( .A(n9737), .Y(n9738) );
  BUFX2 U9684 ( .A(fifo[910]), .Y(n9739) );
  INVX1 U9685 ( .A(n9742), .Y(n9740) );
  INVX1 U9686 ( .A(n9740), .Y(n9741) );
  BUFX2 U9687 ( .A(fifo[911]), .Y(n9742) );
  INVX1 U9688 ( .A(n9745), .Y(n9743) );
  INVX1 U9689 ( .A(n9743), .Y(n9744) );
  BUFX2 U9690 ( .A(fifo[912]), .Y(n9745) );
  INVX1 U9691 ( .A(n9748), .Y(n9746) );
  INVX1 U9692 ( .A(n9746), .Y(n9747) );
  BUFX2 U9693 ( .A(fifo[913]), .Y(n9748) );
  INVX1 U9694 ( .A(n9751), .Y(n9749) );
  INVX1 U9695 ( .A(n9749), .Y(n9750) );
  BUFX2 U9696 ( .A(fifo[914]), .Y(n9751) );
  INVX1 U9697 ( .A(n9754), .Y(n9752) );
  INVX1 U9698 ( .A(n9752), .Y(n9753) );
  BUFX2 U9699 ( .A(fifo[915]), .Y(n9754) );
  INVX1 U9700 ( .A(n9757), .Y(n9755) );
  INVX1 U9701 ( .A(n9755), .Y(n9756) );
  BUFX2 U9702 ( .A(fifo[916]), .Y(n9757) );
  INVX1 U9703 ( .A(n9760), .Y(n9758) );
  INVX1 U9704 ( .A(n9758), .Y(n9759) );
  BUFX2 U9705 ( .A(fifo[917]), .Y(n9760) );
  INVX1 U9706 ( .A(n9763), .Y(n9761) );
  INVX1 U9707 ( .A(n9761), .Y(n9762) );
  BUFX2 U9708 ( .A(fifo[952]), .Y(n9763) );
  INVX1 U9709 ( .A(n9766), .Y(n9764) );
  INVX1 U9710 ( .A(n9764), .Y(n9765) );
  BUFX2 U9711 ( .A(fifo[953]), .Y(n9766) );
  INVX1 U9712 ( .A(n9769), .Y(n9767) );
  INVX1 U9713 ( .A(n9767), .Y(n9768) );
  BUFX2 U9714 ( .A(fifo[954]), .Y(n9769) );
  INVX1 U9715 ( .A(n9772), .Y(n9770) );
  INVX1 U9716 ( .A(n9770), .Y(n9771) );
  BUFX2 U9717 ( .A(fifo[955]), .Y(n9772) );
  INVX1 U9718 ( .A(n9775), .Y(n9773) );
  INVX1 U9719 ( .A(n9773), .Y(n9774) );
  BUFX2 U9720 ( .A(fifo[956]), .Y(n9775) );
  INVX1 U9721 ( .A(n9778), .Y(n9776) );
  INVX1 U9722 ( .A(n9776), .Y(n9777) );
  BUFX2 U9723 ( .A(fifo[957]), .Y(n9778) );
  INVX1 U9724 ( .A(n9781), .Y(n9779) );
  INVX1 U9725 ( .A(n9779), .Y(n9780) );
  BUFX2 U9726 ( .A(fifo[958]), .Y(n9781) );
  INVX1 U9727 ( .A(n9784), .Y(n9782) );
  INVX1 U9728 ( .A(n9782), .Y(n9783) );
  BUFX2 U9729 ( .A(fifo[959]), .Y(n9784) );
  INVX1 U9730 ( .A(n9787), .Y(n9785) );
  INVX1 U9731 ( .A(n9785), .Y(n9786) );
  BUFX2 U9732 ( .A(fifo[960]), .Y(n9787) );
  INVX1 U9733 ( .A(n9790), .Y(n9788) );
  INVX1 U9734 ( .A(n9788), .Y(n9789) );
  BUFX2 U9735 ( .A(fifo[961]), .Y(n9790) );
  INVX1 U9736 ( .A(n9793), .Y(n9791) );
  INVX1 U9737 ( .A(n9791), .Y(n9792) );
  BUFX2 U9738 ( .A(fifo[962]), .Y(n9793) );
  INVX1 U9739 ( .A(n9796), .Y(n9794) );
  INVX1 U9740 ( .A(n9794), .Y(n9795) );
  BUFX2 U9741 ( .A(fifo[963]), .Y(n9796) );
  INVX1 U9742 ( .A(n9799), .Y(n9797) );
  INVX1 U9743 ( .A(n9797), .Y(n9798) );
  BUFX2 U9744 ( .A(fifo[964]), .Y(n9799) );
  INVX1 U9745 ( .A(n9802), .Y(n9800) );
  INVX1 U9746 ( .A(n9800), .Y(n9801) );
  BUFX2 U9747 ( .A(fifo[965]), .Y(n9802) );
  INVX1 U9748 ( .A(n9805), .Y(n9803) );
  INVX1 U9749 ( .A(n9803), .Y(n9804) );
  BUFX2 U9750 ( .A(fifo[966]), .Y(n9805) );
  INVX1 U9751 ( .A(n9808), .Y(n9806) );
  INVX1 U9752 ( .A(n9806), .Y(n9807) );
  BUFX2 U9753 ( .A(fifo[967]), .Y(n9808) );
  INVX1 U9754 ( .A(n9811), .Y(n9809) );
  INVX1 U9755 ( .A(n9809), .Y(n9810) );
  BUFX2 U9756 ( .A(fifo[968]), .Y(n9811) );
  INVX1 U9757 ( .A(n9814), .Y(n9812) );
  INVX1 U9758 ( .A(n9812), .Y(n9813) );
  BUFX2 U9759 ( .A(fifo[969]), .Y(n9814) );
  INVX1 U9760 ( .A(n9817), .Y(n9815) );
  INVX1 U9761 ( .A(n9815), .Y(n9816) );
  BUFX2 U9762 ( .A(fifo[970]), .Y(n9817) );
  INVX1 U9763 ( .A(n9820), .Y(n9818) );
  INVX1 U9764 ( .A(n9818), .Y(n9819) );
  BUFX2 U9765 ( .A(fifo[971]), .Y(n9820) );
  INVX1 U9766 ( .A(n9823), .Y(n9821) );
  INVX1 U9767 ( .A(n9821), .Y(n9822) );
  BUFX2 U9768 ( .A(fifo[972]), .Y(n9823) );
  INVX1 U9769 ( .A(n9826), .Y(n9824) );
  INVX1 U9770 ( .A(n9824), .Y(n9825) );
  BUFX2 U9771 ( .A(fifo[973]), .Y(n9826) );
  INVX1 U9772 ( .A(n9829), .Y(n9827) );
  INVX1 U9773 ( .A(n9827), .Y(n9828) );
  BUFX2 U9774 ( .A(fifo[974]), .Y(n9829) );
  INVX1 U9775 ( .A(n9832), .Y(n9830) );
  INVX1 U9776 ( .A(n9830), .Y(n9831) );
  BUFX2 U9777 ( .A(fifo[975]), .Y(n9832) );
  INVX1 U9778 ( .A(n9835), .Y(n9833) );
  INVX1 U9779 ( .A(n9833), .Y(n9834) );
  BUFX2 U9780 ( .A(fifo[976]), .Y(n9835) );
  INVX1 U9781 ( .A(n9838), .Y(n9836) );
  INVX1 U9782 ( .A(n9836), .Y(n9837) );
  BUFX2 U9783 ( .A(fifo[977]), .Y(n9838) );
  INVX1 U9784 ( .A(n9841), .Y(n9839) );
  INVX1 U9785 ( .A(n9839), .Y(n9840) );
  BUFX2 U9786 ( .A(fifo[978]), .Y(n9841) );
  INVX1 U9787 ( .A(n9844), .Y(n9842) );
  INVX1 U9788 ( .A(n9842), .Y(n9843) );
  BUFX2 U9789 ( .A(fifo[979]), .Y(n9844) );
  INVX1 U9790 ( .A(n9847), .Y(n9845) );
  INVX1 U9791 ( .A(n9845), .Y(n9846) );
  BUFX2 U9792 ( .A(fifo[980]), .Y(n9847) );
  INVX1 U9793 ( .A(n9850), .Y(n9848) );
  INVX1 U9794 ( .A(n9848), .Y(n9849) );
  BUFX2 U9795 ( .A(fifo[981]), .Y(n9850) );
  INVX1 U9796 ( .A(n9853), .Y(n9851) );
  INVX1 U9797 ( .A(n9851), .Y(n9852) );
  BUFX2 U9798 ( .A(fifo[982]), .Y(n9853) );
  INVX1 U9799 ( .A(n9856), .Y(n9854) );
  INVX1 U9800 ( .A(n9854), .Y(n9855) );
  BUFX2 U9801 ( .A(fifo[983]), .Y(n9856) );
  INVX1 U9802 ( .A(n9859), .Y(n9857) );
  INVX1 U9803 ( .A(n9857), .Y(n9858) );
  BUFX2 U9804 ( .A(fifo[984]), .Y(n9859) );
  INVX1 U9805 ( .A(n9862), .Y(n9860) );
  INVX1 U9806 ( .A(n9860), .Y(n9861) );
  BUFX2 U9807 ( .A(fifo[985]), .Y(n9862) );
  INVX1 U9808 ( .A(n9865), .Y(n9863) );
  INVX1 U9809 ( .A(n9863), .Y(n9864) );
  BUFX2 U9810 ( .A(fifo[1020]), .Y(n9865) );
  INVX1 U9811 ( .A(n9868), .Y(n9866) );
  INVX1 U9812 ( .A(n9866), .Y(n9867) );
  BUFX2 U9813 ( .A(fifo[1021]), .Y(n9868) );
  INVX1 U9814 ( .A(n9871), .Y(n9869) );
  INVX1 U9815 ( .A(n9869), .Y(n9870) );
  BUFX2 U9816 ( .A(fifo[1022]), .Y(n9871) );
  INVX1 U9817 ( .A(n9874), .Y(n9872) );
  INVX1 U9818 ( .A(n9872), .Y(n9873) );
  BUFX2 U9819 ( .A(fifo[1023]), .Y(n9874) );
  INVX1 U9820 ( .A(n9877), .Y(n9875) );
  INVX1 U9821 ( .A(n9875), .Y(n9876) );
  BUFX2 U9822 ( .A(fifo[1024]), .Y(n9877) );
  INVX1 U9823 ( .A(n9880), .Y(n9878) );
  INVX1 U9824 ( .A(n9878), .Y(n9879) );
  BUFX2 U9825 ( .A(fifo[1025]), .Y(n9880) );
  INVX1 U9826 ( .A(n9883), .Y(n9881) );
  INVX1 U9827 ( .A(n9881), .Y(n9882) );
  BUFX2 U9828 ( .A(fifo[1026]), .Y(n9883) );
  INVX1 U9829 ( .A(n9886), .Y(n9884) );
  INVX1 U9830 ( .A(n9884), .Y(n9885) );
  BUFX2 U9831 ( .A(fifo[1027]), .Y(n9886) );
  INVX1 U9832 ( .A(n9889), .Y(n9887) );
  INVX1 U9833 ( .A(n9887), .Y(n9888) );
  BUFX2 U9834 ( .A(fifo[1028]), .Y(n9889) );
  INVX1 U9835 ( .A(n9892), .Y(n9890) );
  INVX1 U9836 ( .A(n9890), .Y(n9891) );
  BUFX2 U9837 ( .A(fifo[1029]), .Y(n9892) );
  INVX1 U9838 ( .A(n9895), .Y(n9893) );
  INVX1 U9839 ( .A(n9893), .Y(n9894) );
  BUFX2 U9840 ( .A(fifo[1030]), .Y(n9895) );
  INVX1 U9841 ( .A(n9898), .Y(n9896) );
  INVX1 U9842 ( .A(n9896), .Y(n9897) );
  BUFX2 U9843 ( .A(fifo[1031]), .Y(n9898) );
  INVX1 U9844 ( .A(n9901), .Y(n9899) );
  INVX1 U9845 ( .A(n9899), .Y(n9900) );
  BUFX2 U9846 ( .A(fifo[1032]), .Y(n9901) );
  INVX1 U9847 ( .A(n9904), .Y(n9902) );
  INVX1 U9848 ( .A(n9902), .Y(n9903) );
  BUFX2 U9849 ( .A(fifo[1033]), .Y(n9904) );
  INVX1 U9850 ( .A(n9907), .Y(n9905) );
  INVX1 U9851 ( .A(n9905), .Y(n9906) );
  BUFX2 U9852 ( .A(fifo[1034]), .Y(n9907) );
  INVX1 U9853 ( .A(n9910), .Y(n9908) );
  INVX1 U9854 ( .A(n9908), .Y(n9909) );
  BUFX2 U9855 ( .A(fifo[1035]), .Y(n9910) );
  INVX1 U9856 ( .A(n9913), .Y(n9911) );
  INVX1 U9857 ( .A(n9911), .Y(n9912) );
  BUFX2 U9858 ( .A(fifo[1036]), .Y(n9913) );
  INVX1 U9859 ( .A(n9916), .Y(n9914) );
  INVX1 U9860 ( .A(n9914), .Y(n9915) );
  BUFX2 U9861 ( .A(fifo[1037]), .Y(n9916) );
  INVX1 U9862 ( .A(n9919), .Y(n9917) );
  INVX1 U9863 ( .A(n9917), .Y(n9918) );
  BUFX2 U9864 ( .A(fifo[1038]), .Y(n9919) );
  INVX1 U9865 ( .A(n9922), .Y(n9920) );
  INVX1 U9866 ( .A(n9920), .Y(n9921) );
  BUFX2 U9867 ( .A(fifo[1039]), .Y(n9922) );
  INVX1 U9868 ( .A(n9925), .Y(n9923) );
  INVX1 U9869 ( .A(n9923), .Y(n9924) );
  BUFX2 U9870 ( .A(fifo[1040]), .Y(n9925) );
  INVX1 U9871 ( .A(n9928), .Y(n9926) );
  INVX1 U9872 ( .A(n9926), .Y(n9927) );
  BUFX2 U9873 ( .A(fifo[1041]), .Y(n9928) );
  INVX1 U9874 ( .A(n9931), .Y(n9929) );
  INVX1 U9875 ( .A(n9929), .Y(n9930) );
  BUFX2 U9876 ( .A(fifo[1042]), .Y(n9931) );
  INVX1 U9877 ( .A(n9934), .Y(n9932) );
  INVX1 U9878 ( .A(n9932), .Y(n9933) );
  BUFX2 U9879 ( .A(fifo[1043]), .Y(n9934) );
  INVX1 U9880 ( .A(n9937), .Y(n9935) );
  INVX1 U9881 ( .A(n9935), .Y(n9936) );
  BUFX2 U9882 ( .A(fifo[1044]), .Y(n9937) );
  INVX1 U9883 ( .A(n9940), .Y(n9938) );
  INVX1 U9884 ( .A(n9938), .Y(n9939) );
  BUFX2 U9885 ( .A(fifo[1045]), .Y(n9940) );
  INVX1 U9886 ( .A(n9943), .Y(n9941) );
  INVX1 U9887 ( .A(n9941), .Y(n9942) );
  BUFX2 U9888 ( .A(fifo[1046]), .Y(n9943) );
  INVX1 U9889 ( .A(n9946), .Y(n9944) );
  INVX1 U9890 ( .A(n9944), .Y(n9945) );
  BUFX2 U9891 ( .A(fifo[1047]), .Y(n9946) );
  INVX1 U9892 ( .A(n9949), .Y(n9947) );
  INVX1 U9893 ( .A(n9947), .Y(n9948) );
  BUFX2 U9894 ( .A(fifo[1048]), .Y(n9949) );
  INVX1 U9895 ( .A(n9952), .Y(n9950) );
  INVX1 U9896 ( .A(n9950), .Y(n9951) );
  BUFX2 U9897 ( .A(fifo[1049]), .Y(n9952) );
  INVX1 U9898 ( .A(n9955), .Y(n9953) );
  INVX1 U9899 ( .A(n9953), .Y(n9954) );
  BUFX2 U9900 ( .A(fifo[1050]), .Y(n9955) );
  INVX1 U9901 ( .A(n9958), .Y(n9956) );
  INVX1 U9902 ( .A(n9956), .Y(n9957) );
  BUFX2 U9903 ( .A(fifo[1051]), .Y(n9958) );
  INVX1 U9904 ( .A(n9961), .Y(n9959) );
  INVX1 U9905 ( .A(n9959), .Y(n9960) );
  BUFX2 U9906 ( .A(fifo[1052]), .Y(n9961) );
  INVX1 U9907 ( .A(n9964), .Y(n9962) );
  INVX1 U9908 ( .A(n9962), .Y(n9963) );
  BUFX2 U9909 ( .A(fifo[1053]), .Y(n9964) );
  INVX1 U9910 ( .A(n10), .Y(n10741) );
  INVX1 U9911 ( .A(n12), .Y(n10662) );
  INVX1 U9912 ( .A(rd_ptr_gray_ss[3]), .Y(n10526) );
  INVX1 U9913 ( .A(rd_ptr_gray_ss[2]), .Y(n10524) );
  INVX1 U9914 ( .A(rd_ptr_gray_ss[1]), .Y(n10525) );
  INVX1 U9915 ( .A(rd_ptr_gray_ss[5]), .Y(n9965) );
  INVX1 U9916 ( .A(n9965), .Y(n9966) );
  INVX1 U9917 ( .A(n9969), .Y(n9967) );
  INVX1 U9918 ( .A(n9967), .Y(data_out[13]) );
  BUFX2 U9919 ( .A(n11817), .Y(n9969) );
  INVX1 U9920 ( .A(n9972), .Y(n9970) );
  INVX1 U9921 ( .A(n9970), .Y(data_out[14]) );
  BUFX2 U9922 ( .A(n11816), .Y(n9972) );
  INVX1 U9923 ( .A(n9975), .Y(n9973) );
  INVX1 U9924 ( .A(n9973), .Y(data_out[15]) );
  BUFX2 U9925 ( .A(n11815), .Y(n9975) );
  INVX1 U9926 ( .A(n9978), .Y(n9976) );
  INVX1 U9927 ( .A(n9976), .Y(data_out[16]) );
  BUFX2 U9928 ( .A(n11814), .Y(n9978) );
  INVX1 U9929 ( .A(n9981), .Y(n9979) );
  INVX1 U9930 ( .A(n9979), .Y(data_out[17]) );
  BUFX2 U9931 ( .A(n11813), .Y(n9981) );
  INVX1 U9932 ( .A(n9984), .Y(n9982) );
  INVX1 U9933 ( .A(n9982), .Y(data_out[18]) );
  BUFX2 U9934 ( .A(n11812), .Y(n9984) );
  INVX1 U9935 ( .A(n9987), .Y(n9985) );
  INVX1 U9936 ( .A(n9985), .Y(data_out[19]) );
  BUFX2 U9937 ( .A(n11811), .Y(n9987) );
  INVX1 U9938 ( .A(n9990), .Y(n9988) );
  INVX1 U9939 ( .A(n9988), .Y(data_out[20]) );
  BUFX2 U9940 ( .A(n11810), .Y(n9990) );
  INVX1 U9941 ( .A(n9993), .Y(n9991) );
  INVX1 U9942 ( .A(n9991), .Y(data_out[21]) );
  BUFX2 U9943 ( .A(n11809), .Y(n9993) );
  INVX1 U9944 ( .A(n9996), .Y(n9994) );
  INVX1 U9945 ( .A(n9994), .Y(data_out[22]) );
  BUFX2 U9946 ( .A(n11808), .Y(n9996) );
  INVX1 U9947 ( .A(n9999), .Y(n9997) );
  INVX1 U9948 ( .A(n9997), .Y(n9998) );
  AND2X1 U9949 ( .A(n10088), .B(n242), .Y(n1248) );
  INVX1 U9950 ( .A(n1248), .Y(n9999) );
  INVX1 U9951 ( .A(n10002), .Y(n10000) );
  INVX1 U9952 ( .A(n10000), .Y(n10001) );
  AND2X2 U9953 ( .A(n10091), .B(n244), .Y(n1319) );
  INVX1 U9954 ( .A(n1319), .Y(n10002) );
  INVX1 U9955 ( .A(n10005), .Y(n10003) );
  INVX1 U9956 ( .A(n10003), .Y(data_out[29]) );
  BUFX2 U9957 ( .A(n11801), .Y(n10005) );
  INVX1 U9958 ( .A(n10008), .Y(n10006) );
  INVX1 U9959 ( .A(n10006), .Y(data_out[10]) );
  BUFX2 U9960 ( .A(n11820), .Y(n10008) );
  INVX1 U9961 ( .A(n10011), .Y(n10009) );
  INVX1 U9962 ( .A(n10009), .Y(data_out[11]) );
  BUFX2 U9963 ( .A(n11819), .Y(n10011) );
  INVX1 U9964 ( .A(n10014), .Y(n10012) );
  INVX1 U9965 ( .A(n10012), .Y(data_out[12]) );
  BUFX2 U9966 ( .A(n11818), .Y(n10014) );
  INVX1 U9967 ( .A(wr_ptr_gray_ss[5]), .Y(n10015) );
  INVX1 U9968 ( .A(n10015), .Y(n10016) );
  INVX1 U9969 ( .A(n10015), .Y(n10017) );
  INVX1 U9970 ( .A(n10020), .Y(n10018) );
  INVX1 U9971 ( .A(n10018), .Y(n10019) );
  OR2X2 U9972 ( .A(n10001), .B(n10101), .Y(n468) );
  INVX1 U9973 ( .A(n468), .Y(n10020) );
  INVX1 U9974 ( .A(n10023), .Y(n10021) );
  INVX1 U9975 ( .A(n10021), .Y(n10022) );
  OR2X2 U9976 ( .A(n9998), .B(n246), .Y(n432) );
  INVX1 U9977 ( .A(n432), .Y(n10023) );
  INVX1 U9978 ( .A(n10026), .Y(n10024) );
  INVX1 U9979 ( .A(n10024), .Y(n10025) );
  OR2X2 U9980 ( .A(n9998), .B(n10101), .Y(n396) );
  INVX1 U9981 ( .A(n396), .Y(n10026) );
  INVX1 U9982 ( .A(n10029), .Y(n10027) );
  INVX1 U9983 ( .A(n10027), .Y(data_out[30]) );
  BUFX2 U9984 ( .A(n11800), .Y(n10029) );
  INVX1 U9985 ( .A(n10032), .Y(n10030) );
  INVX1 U9986 ( .A(n10030), .Y(n10031) );
  OR2X2 U9987 ( .A(n10001), .B(n246), .Y(n504) );
  INVX1 U9988 ( .A(n504), .Y(n10032) );
  INVX1 U9989 ( .A(n10035), .Y(n10033) );
  INVX1 U9990 ( .A(n10033), .Y(data_out[23]) );
  BUFX2 U9991 ( .A(n11807), .Y(n10035) );
  INVX1 U9992 ( .A(n10038), .Y(n10036) );
  INVX1 U9993 ( .A(n10036), .Y(data_out[24]) );
  BUFX2 U9994 ( .A(n11806), .Y(n10038) );
  INVX1 U9995 ( .A(n10041), .Y(n10039) );
  INVX1 U9996 ( .A(n10039), .Y(data_out[25]) );
  BUFX2 U9997 ( .A(n11805), .Y(n10041) );
  INVX1 U9998 ( .A(wr_ptr_gray_ss[1]), .Y(n10042) );
  INVX1 U9999 ( .A(n10042), .Y(n10043) );
  INVX1 U10000 ( .A(n10042), .Y(n10044) );
  INVX1 U10001 ( .A(n10048), .Y(n10045) );
  INVX1 U10002 ( .A(n10045), .Y(n10046) );
  INVX1 U10003 ( .A(n10045), .Y(n10047) );
  BUFX2 U10004 ( .A(rd_ptr_bin_5_), .Y(n10048) );
  INVX1 U10005 ( .A(n10051), .Y(n10049) );
  INVX1 U10006 ( .A(n10049), .Y(data_out[9]) );
  BUFX2 U10007 ( .A(n11821), .Y(n10051) );
  INVX1 U10008 ( .A(n11798), .Y(n10052) );
  INVX4 U10009 ( .A(n10052), .Y(data_out[32]) );
  INVX1 U10010 ( .A(n11799), .Y(n10054) );
  INVX4 U10011 ( .A(n10054), .Y(data_out[31]) );
  INVX1 U10012 ( .A(n10058), .Y(n10056) );
  INVX1 U10013 ( .A(n10056), .Y(data_out[1]) );
  BUFX2 U10014 ( .A(n11829), .Y(n10058) );
  INVX1 U10015 ( .A(n10061), .Y(n10059) );
  INVX1 U10016 ( .A(n10059), .Y(data_out[2]) );
  BUFX2 U10017 ( .A(n11828), .Y(n10061) );
  INVX1 U10018 ( .A(n10064), .Y(n10062) );
  INVX1 U10019 ( .A(n10062), .Y(data_out[3]) );
  BUFX2 U10020 ( .A(n11827), .Y(n10064) );
  INVX1 U10021 ( .A(n10067), .Y(n10065) );
  INVX1 U10022 ( .A(n10065), .Y(data_out[4]) );
  BUFX2 U10023 ( .A(n11826), .Y(n10067) );
  INVX1 U10024 ( .A(n10070), .Y(n10068) );
  INVX1 U10025 ( .A(n10068), .Y(data_out[5]) );
  BUFX2 U10026 ( .A(n11825), .Y(n10070) );
  INVX1 U10027 ( .A(n10073), .Y(n10071) );
  INVX1 U10028 ( .A(n10071), .Y(data_out[6]) );
  BUFX2 U10029 ( .A(n11824), .Y(n10073) );
  INVX1 U10030 ( .A(n10076), .Y(n10074) );
  INVX1 U10031 ( .A(n10074), .Y(data_out[7]) );
  BUFX2 U10032 ( .A(n11823), .Y(n10076) );
  INVX1 U10033 ( .A(n10079), .Y(n10077) );
  INVX1 U10034 ( .A(n10077), .Y(data_out[8]) );
  BUFX2 U10035 ( .A(n11822), .Y(n10079) );
  INVX1 U10036 ( .A(n10082), .Y(n10080) );
  INVX1 U10037 ( .A(n10080), .Y(n10081) );
  BUFX2 U10038 ( .A(wr_ptr_bin[5]), .Y(n10082) );
  INVX1 U10039 ( .A(n10085), .Y(n10083) );
  INVX1 U10040 ( .A(n10083), .Y(data_out[0]) );
  BUFX2 U10041 ( .A(n11830), .Y(n10085) );
  INVX1 U10042 ( .A(n10089), .Y(n10086) );
  INVX1 U10043 ( .A(n10086), .Y(n10087) );
  INVX1 U10044 ( .A(n10086), .Y(n10088) );
  BUFX2 U10045 ( .A(wr_ptr_bin[1]), .Y(n10089) );
  INVX1 U10046 ( .A(n10092), .Y(n10090) );
  INVX1 U10047 ( .A(n10090), .Y(n10091) );
  BUFX2 U10048 ( .A(wr_ptr_bin[2]), .Y(n10092) );
  INVX1 U10049 ( .A(n10095), .Y(n10093) );
  INVX2 U10050 ( .A(n10093), .Y(data_out[33]) );
  BUFX2 U10051 ( .A(n11797), .Y(n10095) );
  INVX1 U10052 ( .A(n10098), .Y(n10096) );
  INVX1 U10053 ( .A(n10096), .Y(n10097) );
  BUFX2 U10054 ( .A(wr_ptr_bin[3]), .Y(n10098) );
  INVX1 U10055 ( .A(n10102), .Y(n10099) );
  INVX1 U10056 ( .A(n10099), .Y(n10100) );
  INVX1 U10057 ( .A(n10099), .Y(n10101) );
  BUFX2 U10058 ( .A(wr_ptr_bin[0]), .Y(n10102) );
  INVX1 U10059 ( .A(n10105), .Y(n10103) );
  INVX1 U10060 ( .A(n10103), .Y(n10104) );
  BUFX2 U10061 ( .A(wr_ptr_bin[4]), .Y(n10105) );
  INVX1 U10062 ( .A(n10109), .Y(n10106) );
  INVX1 U10063 ( .A(n10106), .Y(n10107) );
  INVX1 U10064 ( .A(n10106), .Y(n10108) );
  AND2X2 U10065 ( .A(n162), .B(re), .Y(n203) );
  INVX1 U10066 ( .A(n203), .Y(n10109) );
  INVX1 U10067 ( .A(n10533), .Y(n10110) );
  INVX2 U10068 ( .A(n10110), .Y(n10111) );
  INVX1 U10069 ( .A(n10114), .Y(n10112) );
  INVX8 U10070 ( .A(n10112), .Y(n10113) );
  AND2X1 U10071 ( .A(n323), .B(n324), .Y(n254) );
  INVX1 U10072 ( .A(n254), .Y(n10114) );
  INVX1 U10073 ( .A(n10117), .Y(n10115) );
  INVX8 U10074 ( .A(n10115), .Y(n10116) );
  AND2X1 U10075 ( .A(n895), .B(n576), .Y(n1106) );
  INVX1 U10076 ( .A(n1106), .Y(n10117) );
  INVX1 U10077 ( .A(n10120), .Y(n10118) );
  INVX8 U10078 ( .A(n10118), .Y(n10119) );
  AND2X2 U10079 ( .A(n895), .B(n540), .Y(n1071) );
  INVX1 U10080 ( .A(n1071), .Y(n10120) );
  INVX1 U10081 ( .A(n10123), .Y(n10121) );
  INVX8 U10082 ( .A(n10121), .Y(n10122) );
  AND2X2 U10083 ( .A(n895), .B(n10031), .Y(n1036) );
  INVX1 U10084 ( .A(n1036), .Y(n10123) );
  INVX1 U10085 ( .A(n10126), .Y(n10124) );
  INVX8 U10086 ( .A(n10124), .Y(n10125) );
  AND2X2 U10087 ( .A(n895), .B(n10019), .Y(n1001) );
  INVX1 U10088 ( .A(n1001), .Y(n10126) );
  INVX1 U10089 ( .A(n10129), .Y(n10127) );
  INVX8 U10090 ( .A(n10127), .Y(n10128) );
  AND2X2 U10091 ( .A(n895), .B(n10022), .Y(n966) );
  INVX1 U10092 ( .A(n966), .Y(n10129) );
  INVX1 U10093 ( .A(n10132), .Y(n10130) );
  INVX8 U10094 ( .A(n10130), .Y(n10131) );
  AND2X2 U10095 ( .A(n895), .B(n10025), .Y(n931) );
  INVX1 U10096 ( .A(n931), .Y(n10132) );
  INVX1 U10097 ( .A(n10135), .Y(n10133) );
  INVX8 U10098 ( .A(n10133), .Y(n10134) );
  AND2X2 U10099 ( .A(n895), .B(n360), .Y(n896) );
  INVX1 U10100 ( .A(n896), .Y(n10135) );
  INVX1 U10101 ( .A(n10138), .Y(n10136) );
  INVX8 U10102 ( .A(n10136), .Y(n10137) );
  AND2X2 U10103 ( .A(n895), .B(n323), .Y(n860) );
  INVX1 U10104 ( .A(n860), .Y(n10138) );
  INVX1 U10105 ( .A(n2658), .Y(n10645) );
  INVX1 U10106 ( .A(n2658), .Y(n10646) );
  INVX1 U10107 ( .A(n2658), .Y(n10647) );
  INVX1 U10108 ( .A(n2658), .Y(n10648) );
  INVX2 U10109 ( .A(reset), .Y(n2658) );
  INVX2 U10456 ( .A(n10100), .Y(n33) );
  INVX1 U10457 ( .A(rd_ptr_bin_ss[0]), .Y(r301_B_not_0_) );
  INVX8 U10458 ( .A(n10486), .Y(n505) );
  INVX8 U10459 ( .A(n10487), .Y(n541) );
  INVX8 U10460 ( .A(n10488), .Y(n325) );
  INVX8 U10461 ( .A(n10489), .Y(n469) );
  INVX8 U10462 ( .A(n10490), .Y(n397) );
  AND2X2 U10463 ( .A(n10025), .B(n324), .Y(n10491) );
  INVX8 U10464 ( .A(n10491), .Y(n361) );
  AND2X2 U10465 ( .A(n10019), .B(n324), .Y(n10492) );
  INVX8 U10466 ( .A(n10492), .Y(n433) );
  AND2X1 U10467 ( .A(n1177), .B(n323), .Y(n10493) );
  INVX8 U10468 ( .A(n10493), .Y(n1142) );
  INVX8 U10469 ( .A(n10494), .Y(n1178) );
  INVX1 U10470 ( .A(n165), .Y(n10495) );
  INVX8 U10471 ( .A(n10495), .Y(n10496) );
  INVX1 U10472 ( .A(n164), .Y(n10497) );
  INVX8 U10473 ( .A(n10497), .Y(n10498) );
  INVX1 U10474 ( .A(n167), .Y(n10499) );
  INVX8 U10475 ( .A(n10499), .Y(n10500) );
  INVX8 U10476 ( .A(n10501), .Y(n1284) );
  INVX8 U10477 ( .A(n10502), .Y(n1249) );
  INVX1 U10478 ( .A(n166), .Y(n10503) );
  INVX8 U10479 ( .A(n10503), .Y(n10504) );
  INVX1 U10480 ( .A(n172), .Y(n10505) );
  INVX8 U10481 ( .A(n10505), .Y(n10506) );
  INVX1 U10482 ( .A(n171), .Y(n10507) );
  INVX8 U10483 ( .A(n10507), .Y(n10508) );
  INVX8 U10484 ( .A(n10509), .Y(n824) );
  INVX1 U10485 ( .A(n168), .Y(n10510) );
  INVX8 U10486 ( .A(n10510), .Y(n10511) );
  INVX8 U10487 ( .A(n10512), .Y(n649) );
  INVX8 U10488 ( .A(n10513), .Y(n719) );
  INVX1 U10489 ( .A(n170), .Y(n10514) );
  INVX8 U10490 ( .A(n10514), .Y(n10515) );
  INVX1 U10491 ( .A(n169), .Y(n10516) );
  INVX8 U10492 ( .A(n10516), .Y(n10517) );
  AND2X2 U10493 ( .A(n237), .B(n10519), .Y(n895) );
  INVX1 U10494 ( .A(n163), .Y(n10519) );
  XOR2X1 U10495 ( .A(r301_B_not_4_), .B(n10104), .Y(n10520) );
  XOR2X1 U10496 ( .A(n2), .B(n10520), .Y(fillcount[4]) );
  XNOR2X1 U10497 ( .A(rd_ptr_bin_ss[3]), .B(n10524), .Y(rd_ptr_bin_ss[2]) );
  XNOR2X1 U10498 ( .A(rd_ptr_bin_ss[2]), .B(n10525), .Y(rd_ptr_bin_ss[1]) );
  AND2X2 U10499 ( .A(n39), .B(we), .Y(n237) );
  XNOR2X1 U10500 ( .A(rd_ptr_bin_ss[4]), .B(n10526), .Y(rd_ptr_bin_ss[3]) );
  INVX1 U10501 ( .A(n14), .Y(n10527) );
  INVX1 U10502 ( .A(n10527), .Y(n10528) );
  INVX1 U10503 ( .A(n10527), .Y(n10529) );
  XNOR2X1 U10504 ( .A(n194), .B(n1433), .Y(n10530) );
  INVX2 U10505 ( .A(n10528), .Y(n194) );
  INVX1 U10506 ( .A(n13), .Y(n10531) );
  INVX1 U10507 ( .A(n10531), .Y(n10532) );
  INVX1 U10508 ( .A(n196), .Y(n10533) );
  XOR2X1 U10509 ( .A(n10534), .B(n196), .Y(n10535) );
  BUFX2 U10510 ( .A(n196), .Y(n10536) );
  INVX8 U10511 ( .A(n10633), .Y(n10537) );
  INVX8 U10512 ( .A(n10632), .Y(n10538) );
  INVX8 U10513 ( .A(n10632), .Y(n10539) );
  INVX8 U10514 ( .A(n10632), .Y(n10540) );
  INVX8 U10515 ( .A(n10631), .Y(n10541) );
  INVX8 U10516 ( .A(n10631), .Y(n10542) );
  INVX8 U10517 ( .A(n10631), .Y(n10543) );
  INVX8 U10518 ( .A(n10630), .Y(n10544) );
  INVX8 U10519 ( .A(n10630), .Y(n10545) );
  INVX8 U10520 ( .A(n10630), .Y(n10546) );
  INVX8 U10521 ( .A(n10629), .Y(n10547) );
  INVX8 U10522 ( .A(n10629), .Y(n10548) );
  INVX8 U10523 ( .A(n10629), .Y(n10549) );
  INVX8 U10524 ( .A(n10628), .Y(n10550) );
  INVX8 U10525 ( .A(n10628), .Y(n10551) );
  INVX8 U10526 ( .A(n10628), .Y(n10552) );
  INVX8 U10527 ( .A(n10627), .Y(n10553) );
  INVX8 U10528 ( .A(n10627), .Y(n10554) );
  INVX8 U10529 ( .A(n10627), .Y(n10555) );
  INVX8 U10530 ( .A(n10626), .Y(n10556) );
  INVX8 U10531 ( .A(n10626), .Y(n10557) );
  INVX8 U10532 ( .A(n10626), .Y(n10558) );
  INVX8 U10533 ( .A(n10625), .Y(n10559) );
  INVX8 U10534 ( .A(n10625), .Y(n10560) );
  INVX8 U10535 ( .A(n10625), .Y(n10561) );
  INVX8 U10536 ( .A(n10624), .Y(n10562) );
  INVX8 U10537 ( .A(n10624), .Y(n10563) );
  INVX8 U10538 ( .A(n10623), .Y(n10564) );
  INVX8 U10539 ( .A(n10623), .Y(n10565) );
  INVX8 U10540 ( .A(n10623), .Y(n10566) );
  INVX8 U10541 ( .A(n10622), .Y(n10567) );
  INVX8 U10542 ( .A(n10622), .Y(n10568) );
  INVX8 U10543 ( .A(n10622), .Y(n10569) );
  INVX8 U10544 ( .A(n10621), .Y(n10570) );
  INVX8 U10545 ( .A(n10621), .Y(n10571) );
  INVX8 U10546 ( .A(n10621), .Y(n10572) );
  INVX8 U10547 ( .A(n10620), .Y(n10573) );
  INVX8 U10548 ( .A(n10620), .Y(n10574) );
  INVX8 U10549 ( .A(n10620), .Y(n10575) );
  INVX8 U10550 ( .A(n10619), .Y(n10576) );
  INVX8 U10551 ( .A(n10619), .Y(n10577) );
  INVX8 U10552 ( .A(n10619), .Y(n10578) );
  INVX8 U10553 ( .A(n10618), .Y(n10579) );
  INVX8 U10554 ( .A(n10618), .Y(n10580) );
  INVX8 U10555 ( .A(n10618), .Y(n10581) );
  INVX8 U10556 ( .A(n10617), .Y(n10582) );
  INVX8 U10557 ( .A(n10617), .Y(n10583) );
  INVX8 U10558 ( .A(n10617), .Y(n10584) );
  INVX8 U10559 ( .A(n10616), .Y(n10585) );
  INVX8 U10560 ( .A(n10616), .Y(n10586) );
  INVX8 U10561 ( .A(n10616), .Y(n10587) );
  INVX8 U10562 ( .A(n10615), .Y(n10588) );
  INVX8 U10563 ( .A(n10615), .Y(n10589) );
  INVX8 U10564 ( .A(n10615), .Y(n10590) );
  INVX8 U10565 ( .A(n10614), .Y(n10591) );
  INVX8 U10566 ( .A(n10614), .Y(n10592) );
  INVX8 U10567 ( .A(n10614), .Y(n10593) );
  INVX8 U10568 ( .A(n10613), .Y(n10594) );
  INVX8 U10569 ( .A(n10613), .Y(n10595) );
  INVX8 U10570 ( .A(n10613), .Y(n10596) );
  INVX8 U10571 ( .A(n10612), .Y(n10597) );
  INVX8 U10572 ( .A(n10612), .Y(n10598) );
  INVX8 U10573 ( .A(n10612), .Y(n10599) );
  INVX8 U10574 ( .A(n10611), .Y(n10600) );
  INVX8 U10575 ( .A(n10611), .Y(n10601) );
  INVX8 U10576 ( .A(n10611), .Y(n10602) );
  INVX8 U10577 ( .A(n10610), .Y(n10603) );
  INVX8 U10578 ( .A(n10610), .Y(n10604) );
  INVX8 U10579 ( .A(n10610), .Y(n10605) );
  INVX8 U10580 ( .A(n10609), .Y(n10606) );
  INVX8 U10581 ( .A(n10609), .Y(n10607) );
  INVX8 U10582 ( .A(n10609), .Y(n10608) );
  INVX8 U10583 ( .A(n10644), .Y(n10609) );
  INVX8 U10584 ( .A(n10644), .Y(n10610) );
  INVX8 U10585 ( .A(n10644), .Y(n10611) );
  INVX8 U10586 ( .A(n10643), .Y(n10612) );
  INVX8 U10587 ( .A(n10643), .Y(n10613) );
  INVX8 U10588 ( .A(n10643), .Y(n10614) );
  INVX8 U10589 ( .A(n10642), .Y(n10615) );
  INVX8 U10590 ( .A(n10642), .Y(n10616) );
  INVX8 U10591 ( .A(n10642), .Y(n10617) );
  INVX8 U10592 ( .A(n10641), .Y(n10618) );
  INVX8 U10593 ( .A(n10641), .Y(n10619) );
  INVX8 U10594 ( .A(n10641), .Y(n10620) );
  INVX8 U10595 ( .A(n10640), .Y(n10621) );
  INVX8 U10596 ( .A(n10640), .Y(n10622) );
  INVX8 U10597 ( .A(n10640), .Y(n10623) );
  INVX8 U10598 ( .A(n10637), .Y(n10624) );
  INVX8 U10599 ( .A(n10636), .Y(n10625) );
  INVX8 U10600 ( .A(n10636), .Y(n10626) );
  INVX8 U10601 ( .A(n10636), .Y(n10627) );
  INVX8 U10602 ( .A(n10635), .Y(n10628) );
  INVX8 U10603 ( .A(n10635), .Y(n10629) );
  INVX8 U10604 ( .A(n10635), .Y(n10630) );
  INVX8 U10605 ( .A(n10634), .Y(n10631) );
  INVX8 U10606 ( .A(n10634), .Y(n10632) );
  INVX8 U10607 ( .A(n10634), .Y(n10633) );
  INVX8 U10608 ( .A(n10648), .Y(n10634) );
  INVX8 U10609 ( .A(n10648), .Y(n10635) );
  INVX8 U10610 ( .A(n10647), .Y(n10636) );
  INVX8 U10611 ( .A(n10647), .Y(n10637) );
  INVX8 U10612 ( .A(n10647), .Y(n10638) );
  INVX8 U10613 ( .A(n10646), .Y(n10639) );
  INVX8 U10614 ( .A(n10646), .Y(n10640) );
  INVX8 U10615 ( .A(n10646), .Y(n10641) );
  INVX8 U10616 ( .A(n10645), .Y(n10642) );
  INVX8 U10617 ( .A(n10645), .Y(n10643) );
  INVX8 U10618 ( .A(n10645), .Y(n10644) );
  INVX8 U10619 ( .A(n10658), .Y(n10649) );
  INVX8 U10620 ( .A(n10658), .Y(n10650) );
  INVX8 U10621 ( .A(n10658), .Y(n10651) );
  INVX8 U10622 ( .A(n10659), .Y(n10652) );
  INVX8 U10623 ( .A(n10659), .Y(n10653) );
  INVX8 U10624 ( .A(n10660), .Y(n10654) );
  INVX8 U10625 ( .A(n10660), .Y(n10655) );
  INVX8 U10626 ( .A(n10660), .Y(n10656) );
  INVX8 U10627 ( .A(n10659), .Y(n10657) );
  INVX8 U10628 ( .A(n10661), .Y(n10658) );
  INVX8 U10629 ( .A(n10661), .Y(n10659) );
  INVX8 U10630 ( .A(n10661), .Y(n10660) );
  INVX8 U10631 ( .A(n10662), .Y(n10661) );
  INVX8 U10632 ( .A(n10685), .Y(n10663) );
  INVX8 U10633 ( .A(n10685), .Y(n10664) );
  INVX8 U10634 ( .A(n10684), .Y(n10665) );
  INVX8 U10635 ( .A(n10684), .Y(n10666) );
  INVX8 U10636 ( .A(n10684), .Y(n10667) );
  INVX8 U10637 ( .A(n10683), .Y(n10668) );
  INVX8 U10638 ( .A(n10683), .Y(n10669) );
  INVX8 U10639 ( .A(n10683), .Y(n10670) );
  INVX8 U10640 ( .A(n10682), .Y(n10671) );
  INVX8 U10641 ( .A(n10682), .Y(n10672) );
  INVX8 U10642 ( .A(n10682), .Y(n10673) );
  INVX8 U10643 ( .A(n10681), .Y(n10674) );
  INVX8 U10644 ( .A(n10681), .Y(n10675) );
  INVX8 U10645 ( .A(n10681), .Y(n10676) );
  INVX8 U10646 ( .A(n10680), .Y(n10677) );
  INVX8 U10647 ( .A(n10680), .Y(n10678) );
  INVX8 U10648 ( .A(n10680), .Y(n10679) );
  INVX8 U10649 ( .A(n10687), .Y(n10680) );
  INVX8 U10650 ( .A(n10687), .Y(n10681) );
  INVX8 U10651 ( .A(n10687), .Y(n10682) );
  INVX8 U10652 ( .A(n10686), .Y(n10684) );
  INVX8 U10653 ( .A(n10686), .Y(n10685) );
  INVX8 U10654 ( .A(n10722), .Y(n10689) );
  INVX8 U10655 ( .A(n10722), .Y(n10690) );
  INVX8 U10656 ( .A(n10723), .Y(n10691) );
  INVX8 U10657 ( .A(n10723), .Y(n10692) );
  INVX8 U10658 ( .A(n10723), .Y(n10693) );
  INVX8 U10659 ( .A(n10727), .Y(n10694) );
  INVX8 U10660 ( .A(n10724), .Y(n10695) );
  INVX8 U10661 ( .A(n10724), .Y(n10696) );
  INVX8 U10662 ( .A(n10724), .Y(n10697) );
  INVX8 U10663 ( .A(n10725), .Y(n10698) );
  INVX8 U10664 ( .A(n10725), .Y(n10699) );
  INVX8 U10665 ( .A(n10725), .Y(n10700) );
  INVX8 U10666 ( .A(n10726), .Y(n10701) );
  INVX8 U10667 ( .A(n10726), .Y(n10702) );
  INVX8 U10668 ( .A(n10726), .Y(n10703) );
  INVX8 U10669 ( .A(n10727), .Y(n10704) );
  INVX8 U10670 ( .A(n10727), .Y(n10705) );
  INVX8 U10671 ( .A(n10728), .Y(n10706) );
  INVX8 U10672 ( .A(n10728), .Y(n10707) );
  INVX8 U10673 ( .A(n10728), .Y(n10708) );
  INVX8 U10674 ( .A(n10729), .Y(n10709) );
  INVX8 U10675 ( .A(n10729), .Y(n10710) );
  INVX8 U10676 ( .A(n10729), .Y(n10711) );
  INVX8 U10677 ( .A(n10730), .Y(n10712) );
  INVX8 U10678 ( .A(n10730), .Y(n10713) );
  INVX8 U10679 ( .A(n10730), .Y(n10714) );
  INVX8 U10680 ( .A(n10731), .Y(n10715) );
  INVX8 U10681 ( .A(n10731), .Y(n10716) );
  INVX8 U10682 ( .A(n10732), .Y(n10717) );
  INVX8 U10683 ( .A(n10732), .Y(n10718) );
  INVX8 U10684 ( .A(n10732), .Y(n10719) );
  INVX8 U10685 ( .A(n10731), .Y(n10720) );
  INVX8 U10686 ( .A(n10722), .Y(n10721) );
  INVX8 U10687 ( .A(n10737), .Y(n10722) );
  INVX8 U10688 ( .A(n10737), .Y(n10723) );
  INVX8 U10689 ( .A(n10737), .Y(n10724) );
  INVX8 U10690 ( .A(n10736), .Y(n10725) );
  INVX8 U10691 ( .A(n10736), .Y(n10726) );
  INVX8 U10692 ( .A(n10736), .Y(n10727) );
  INVX8 U10693 ( .A(n10735), .Y(n10728) );
  INVX8 U10694 ( .A(n10735), .Y(n10729) );
  INVX8 U10695 ( .A(n10735), .Y(n10730) );
  INVX8 U10696 ( .A(n10734), .Y(n10731) );
  INVX8 U10697 ( .A(n10734), .Y(n10732) );
  INVX8 U10698 ( .A(n10734), .Y(n10733) );
  INVX8 U10699 ( .A(n10739), .Y(n10734) );
  INVX8 U10700 ( .A(n10738), .Y(n10735) );
  INVX8 U10701 ( .A(n10738), .Y(n10736) );
  INVX8 U10702 ( .A(n10738), .Y(n10737) );
  INVX8 U10703 ( .A(n10740), .Y(n10738) );
  MUX2X1 U10704 ( .B(n10743), .A(n10744), .S(n10679), .Y(n10742) );
  MUX2X1 U10705 ( .B(n10746), .A(n10747), .S(n10679), .Y(n10745) );
  MUX2X1 U10706 ( .B(n10749), .A(n10750), .S(n10679), .Y(n10748) );
  MUX2X1 U10707 ( .B(n10752), .A(n10753), .S(n10679), .Y(n10751) );
  MUX2X1 U10708 ( .B(n10755), .A(n10756), .S(n10111), .Y(n10754) );
  MUX2X1 U10709 ( .B(n10758), .A(n10759), .S(n10679), .Y(n10757) );
  MUX2X1 U10710 ( .B(n10761), .A(n10762), .S(n10678), .Y(n10760) );
  MUX2X1 U10711 ( .B(n10764), .A(n10765), .S(n10678), .Y(n10763) );
  MUX2X1 U10712 ( .B(n10767), .A(n10768), .S(n10678), .Y(n10766) );
  MUX2X1 U10713 ( .B(n10770), .A(n10771), .S(n10111), .Y(n10769) );
  MUX2X1 U10714 ( .B(n10773), .A(n10774), .S(n10678), .Y(n10772) );
  MUX2X1 U10715 ( .B(n10776), .A(n10777), .S(n10678), .Y(n10775) );
  MUX2X1 U10716 ( .B(n10779), .A(n10780), .S(n10678), .Y(n10778) );
  MUX2X1 U10717 ( .B(n10782), .A(n10783), .S(n10678), .Y(n10781) );
  MUX2X1 U10718 ( .B(n10785), .A(n10786), .S(n10111), .Y(n10784) );
  MUX2X1 U10719 ( .B(n10788), .A(n10789), .S(n10678), .Y(n10787) );
  MUX2X1 U10720 ( .B(n10791), .A(n10792), .S(n10678), .Y(n10790) );
  MUX2X1 U10721 ( .B(n10794), .A(n10795), .S(n10678), .Y(n10793) );
  MUX2X1 U10722 ( .B(n10797), .A(n10798), .S(n10678), .Y(n10796) );
  MUX2X1 U10723 ( .B(n10800), .A(n10801), .S(n10111), .Y(n10799) );
  MUX2X1 U10724 ( .B(n10803), .A(n10804), .S(n10678), .Y(n10802) );
  MUX2X1 U10725 ( .B(n10806), .A(n10807), .S(n10678), .Y(n10805) );
  MUX2X1 U10726 ( .B(n10809), .A(n10810), .S(n10678), .Y(n10808) );
  MUX2X1 U10727 ( .B(n10812), .A(n10813), .S(n10678), .Y(n10811) );
  MUX2X1 U10728 ( .B(n10815), .A(n10816), .S(n10111), .Y(n10814) );
  MUX2X1 U10729 ( .B(n10818), .A(n10819), .S(n10678), .Y(n10817) );
  MUX2X1 U10730 ( .B(n10821), .A(n10822), .S(n10678), .Y(n10820) );
  MUX2X1 U10731 ( .B(n10824), .A(n10825), .S(n10677), .Y(n10823) );
  MUX2X1 U10732 ( .B(n10827), .A(n10828), .S(n10677), .Y(n10826) );
  MUX2X1 U10733 ( .B(n10830), .A(n10831), .S(n10111), .Y(n10829) );
  MUX2X1 U10734 ( .B(n10833), .A(n10834), .S(n10677), .Y(n10832) );
  MUX2X1 U10735 ( .B(n10836), .A(n10837), .S(n10677), .Y(n10835) );
  MUX2X1 U10736 ( .B(n10839), .A(n10840), .S(n10677), .Y(n10838) );
  MUX2X1 U10737 ( .B(n10842), .A(n10843), .S(n10677), .Y(n10841) );
  MUX2X1 U10738 ( .B(n10845), .A(n10846), .S(n10111), .Y(n10844) );
  MUX2X1 U10739 ( .B(n10848), .A(n10849), .S(n10677), .Y(n10847) );
  MUX2X1 U10740 ( .B(n10851), .A(n10852), .S(n10677), .Y(n10850) );
  MUX2X1 U10741 ( .B(n10854), .A(n10855), .S(n10677), .Y(n10853) );
  MUX2X1 U10742 ( .B(n10857), .A(n10858), .S(n10677), .Y(n10856) );
  MUX2X1 U10743 ( .B(n10860), .A(n10861), .S(n10111), .Y(n10859) );
  MUX2X1 U10744 ( .B(n10863), .A(n10864), .S(n10677), .Y(n10862) );
  MUX2X1 U10745 ( .B(n10866), .A(n10867), .S(n10677), .Y(n10865) );
  MUX2X1 U10746 ( .B(n10869), .A(n10870), .S(n10677), .Y(n10868) );
  MUX2X1 U10747 ( .B(n10872), .A(n10873), .S(n10677), .Y(n10871) );
  MUX2X1 U10748 ( .B(n10875), .A(n10876), .S(n10111), .Y(n10874) );
  MUX2X1 U10749 ( .B(n10878), .A(n10879), .S(n10677), .Y(n10877) );
  MUX2X1 U10750 ( .B(n10881), .A(n10882), .S(n10677), .Y(n10880) );
  MUX2X1 U10751 ( .B(n10884), .A(n10885), .S(n10677), .Y(n10883) );
  MUX2X1 U10752 ( .B(n10887), .A(n10888), .S(n10676), .Y(n10886) );
  MUX2X1 U10753 ( .B(n10890), .A(n10891), .S(n10111), .Y(n10889) );
  MUX2X1 U10754 ( .B(n10893), .A(n10894), .S(n10676), .Y(n10892) );
  MUX2X1 U10755 ( .B(n10896), .A(n10897), .S(n10676), .Y(n10895) );
  MUX2X1 U10756 ( .B(n10899), .A(n10900), .S(n10676), .Y(n10898) );
  MUX2X1 U10757 ( .B(n10902), .A(n10903), .S(n10676), .Y(n10901) );
  MUX2X1 U10758 ( .B(n10905), .A(n10906), .S(n10111), .Y(n10904) );
  MUX2X1 U10759 ( .B(n10908), .A(n10909), .S(n10676), .Y(n10907) );
  MUX2X1 U10760 ( .B(n10911), .A(n10912), .S(n10676), .Y(n10910) );
  MUX2X1 U10761 ( .B(n10914), .A(n10915), .S(n10676), .Y(n10913) );
  MUX2X1 U10762 ( .B(n10917), .A(n10918), .S(n10676), .Y(n10916) );
  MUX2X1 U10763 ( .B(n10920), .A(n10921), .S(n10111), .Y(n10919) );
  MUX2X1 U10764 ( .B(n10923), .A(n10924), .S(n10676), .Y(n10922) );
  MUX2X1 U10765 ( .B(n10926), .A(n10927), .S(n10676), .Y(n10925) );
  MUX2X1 U10766 ( .B(n10929), .A(n10930), .S(n10676), .Y(n10928) );
  MUX2X1 U10767 ( .B(n10932), .A(n10933), .S(n10676), .Y(n10931) );
  MUX2X1 U10768 ( .B(n10935), .A(n10936), .S(n10111), .Y(n10934) );
  MUX2X1 U10769 ( .B(n10938), .A(n10939), .S(n10676), .Y(n10937) );
  MUX2X1 U10770 ( .B(n10941), .A(n10942), .S(n10676), .Y(n10940) );
  MUX2X1 U10771 ( .B(n10944), .A(n10945), .S(n10676), .Y(n10943) );
  MUX2X1 U10772 ( .B(n10947), .A(n10948), .S(n10676), .Y(n10946) );
  MUX2X1 U10773 ( .B(n10950), .A(n10951), .S(n10111), .Y(n10949) );
  MUX2X1 U10774 ( .B(n10953), .A(n10954), .S(n10675), .Y(n10952) );
  MUX2X1 U10775 ( .B(n10956), .A(n10957), .S(n10675), .Y(n10955) );
  MUX2X1 U10776 ( .B(n10959), .A(n10960), .S(n10675), .Y(n10958) );
  MUX2X1 U10777 ( .B(n10962), .A(n10963), .S(n10675), .Y(n10961) );
  MUX2X1 U10778 ( .B(n10965), .A(n10966), .S(n10111), .Y(n10964) );
  MUX2X1 U10779 ( .B(n10968), .A(n10969), .S(n10675), .Y(n10967) );
  MUX2X1 U10780 ( .B(n10971), .A(n10972), .S(n10675), .Y(n10970) );
  MUX2X1 U10781 ( .B(n10974), .A(n10975), .S(n10675), .Y(n10973) );
  MUX2X1 U10782 ( .B(n10977), .A(n10978), .S(n10675), .Y(n10976) );
  MUX2X1 U10783 ( .B(n10980), .A(n10981), .S(n10111), .Y(n10979) );
  MUX2X1 U10784 ( .B(n10983), .A(n10984), .S(n10675), .Y(n10982) );
  MUX2X1 U10785 ( .B(n10986), .A(n10987), .S(n10675), .Y(n10985) );
  MUX2X1 U10786 ( .B(n10989), .A(n10990), .S(n10675), .Y(n10988) );
  MUX2X1 U10787 ( .B(n10992), .A(n10993), .S(n10675), .Y(n10991) );
  MUX2X1 U10788 ( .B(n10995), .A(n10996), .S(n10111), .Y(n10994) );
  MUX2X1 U10789 ( .B(n10998), .A(n10999), .S(n10675), .Y(n10997) );
  MUX2X1 U10790 ( .B(n11001), .A(n11002), .S(n10675), .Y(n11000) );
  MUX2X1 U10791 ( .B(n11004), .A(n11005), .S(n10675), .Y(n11003) );
  MUX2X1 U10792 ( .B(n11007), .A(n11008), .S(n10675), .Y(n11006) );
  MUX2X1 U10793 ( .B(n11010), .A(n11011), .S(n10111), .Y(n11009) );
  MUX2X1 U10794 ( .B(n11013), .A(n11014), .S(n10675), .Y(n11012) );
  MUX2X1 U10795 ( .B(n11016), .A(n11017), .S(n10674), .Y(n11015) );
  MUX2X1 U10796 ( .B(n11019), .A(n11020), .S(n10674), .Y(n11018) );
  MUX2X1 U10797 ( .B(n11022), .A(n11023), .S(n10674), .Y(n11021) );
  MUX2X1 U10798 ( .B(n11025), .A(n11026), .S(n10111), .Y(n11024) );
  MUX2X1 U10799 ( .B(n11028), .A(n11029), .S(n10674), .Y(n11027) );
  MUX2X1 U10800 ( .B(n11031), .A(n11032), .S(n10674), .Y(n11030) );
  MUX2X1 U10801 ( .B(n11034), .A(n11035), .S(n10674), .Y(n11033) );
  MUX2X1 U10802 ( .B(n11037), .A(n11038), .S(n10674), .Y(n11036) );
  MUX2X1 U10803 ( .B(n11040), .A(n11041), .S(n10111), .Y(n11039) );
  MUX2X1 U10804 ( .B(n11043), .A(n11044), .S(n10674), .Y(n11042) );
  MUX2X1 U10805 ( .B(n11046), .A(n11047), .S(n10674), .Y(n11045) );
  MUX2X1 U10806 ( .B(n11049), .A(n11050), .S(n10674), .Y(n11048) );
  MUX2X1 U10807 ( .B(n11052), .A(n11053), .S(n10674), .Y(n11051) );
  MUX2X1 U10808 ( .B(n11055), .A(n11056), .S(n10111), .Y(n11054) );
  MUX2X1 U10809 ( .B(n11058), .A(n11059), .S(n10674), .Y(n11057) );
  MUX2X1 U10810 ( .B(n11061), .A(n11062), .S(n10674), .Y(n11060) );
  MUX2X1 U10811 ( .B(n11064), .A(n11065), .S(n10674), .Y(n11063) );
  MUX2X1 U10812 ( .B(n11067), .A(n11068), .S(n10674), .Y(n11066) );
  MUX2X1 U10813 ( .B(n11070), .A(n11071), .S(n10111), .Y(n11069) );
  MUX2X1 U10814 ( .B(n11073), .A(n11074), .S(n10674), .Y(n11072) );
  MUX2X1 U10815 ( .B(n11076), .A(n11077), .S(n10674), .Y(n11075) );
  MUX2X1 U10816 ( .B(n11079), .A(n11080), .S(n10673), .Y(n11078) );
  MUX2X1 U10817 ( .B(n11082), .A(n11083), .S(n10673), .Y(n11081) );
  MUX2X1 U10818 ( .B(n11085), .A(n11086), .S(n10111), .Y(n11084) );
  MUX2X1 U10819 ( .B(n11088), .A(n11089), .S(n10673), .Y(n11087) );
  MUX2X1 U10820 ( .B(n11091), .A(n11092), .S(n10673), .Y(n11090) );
  MUX2X1 U10821 ( .B(n11094), .A(n11095), .S(n10673), .Y(n11093) );
  MUX2X1 U10822 ( .B(n11097), .A(n11098), .S(n10673), .Y(n11096) );
  MUX2X1 U10823 ( .B(n11100), .A(n11101), .S(n10111), .Y(n11099) );
  MUX2X1 U10824 ( .B(n11103), .A(n11104), .S(n10673), .Y(n11102) );
  MUX2X1 U10825 ( .B(n11106), .A(n11107), .S(n10673), .Y(n11105) );
  MUX2X1 U10826 ( .B(n11109), .A(n11110), .S(n10673), .Y(n11108) );
  MUX2X1 U10827 ( .B(n11112), .A(n11113), .S(n10673), .Y(n11111) );
  MUX2X1 U10828 ( .B(n11115), .A(n11116), .S(n10111), .Y(n11114) );
  MUX2X1 U10829 ( .B(n11118), .A(n11119), .S(n10673), .Y(n11117) );
  MUX2X1 U10830 ( .B(n11121), .A(n11122), .S(n10673), .Y(n11120) );
  MUX2X1 U10831 ( .B(n11124), .A(n11125), .S(n10673), .Y(n11123) );
  MUX2X1 U10832 ( .B(n11127), .A(n11128), .S(n10673), .Y(n11126) );
  MUX2X1 U10833 ( .B(n11130), .A(n11131), .S(n10111), .Y(n11129) );
  MUX2X1 U10834 ( .B(n11133), .A(n11134), .S(n10673), .Y(n11132) );
  MUX2X1 U10835 ( .B(n11136), .A(n11137), .S(n10673), .Y(n11135) );
  MUX2X1 U10836 ( .B(n11139), .A(n11140), .S(n10673), .Y(n11138) );
  MUX2X1 U10837 ( .B(n11142), .A(n11143), .S(n10672), .Y(n11141) );
  MUX2X1 U10838 ( .B(n11145), .A(n11146), .S(n10111), .Y(n11144) );
  MUX2X1 U10839 ( .B(n11148), .A(n11149), .S(n10672), .Y(n11147) );
  MUX2X1 U10840 ( .B(n11151), .A(n11152), .S(n10672), .Y(n11150) );
  MUX2X1 U10841 ( .B(n11154), .A(n11155), .S(n10672), .Y(n11153) );
  MUX2X1 U10842 ( .B(n11157), .A(n11158), .S(n10672), .Y(n11156) );
  MUX2X1 U10843 ( .B(n11160), .A(n11161), .S(n10111), .Y(n11159) );
  MUX2X1 U10844 ( .B(n11163), .A(n11164), .S(n10672), .Y(n11162) );
  MUX2X1 U10845 ( .B(n11166), .A(n11167), .S(n10672), .Y(n11165) );
  MUX2X1 U10846 ( .B(n11169), .A(n11170), .S(n10672), .Y(n11168) );
  MUX2X1 U10847 ( .B(n11172), .A(n11173), .S(n10672), .Y(n11171) );
  MUX2X1 U10848 ( .B(n11175), .A(n11176), .S(n10111), .Y(n11174) );
  MUX2X1 U10849 ( .B(n11178), .A(n11179), .S(n10672), .Y(n11177) );
  MUX2X1 U10850 ( .B(n11181), .A(n11182), .S(n10672), .Y(n11180) );
  MUX2X1 U10851 ( .B(n11184), .A(n11185), .S(n10672), .Y(n11183) );
  MUX2X1 U10852 ( .B(n11187), .A(n11188), .S(n10672), .Y(n11186) );
  MUX2X1 U10853 ( .B(n11190), .A(n11191), .S(n10111), .Y(n11189) );
  MUX2X1 U10854 ( .B(n11193), .A(n11194), .S(n10672), .Y(n11192) );
  MUX2X1 U10855 ( .B(n11196), .A(n11197), .S(n10672), .Y(n11195) );
  MUX2X1 U10856 ( .B(n11199), .A(n11200), .S(n10672), .Y(n11198) );
  MUX2X1 U10857 ( .B(n11202), .A(n11203), .S(n10672), .Y(n11201) );
  MUX2X1 U10858 ( .B(n11205), .A(n11206), .S(n10111), .Y(n11204) );
  MUX2X1 U10859 ( .B(n11208), .A(n11209), .S(n10671), .Y(n11207) );
  MUX2X1 U10860 ( .B(n11211), .A(n11212), .S(n10671), .Y(n11210) );
  MUX2X1 U10861 ( .B(n11214), .A(n11215), .S(n10671), .Y(n11213) );
  MUX2X1 U10862 ( .B(n11217), .A(n11218), .S(n10671), .Y(n11216) );
  MUX2X1 U10863 ( .B(n11220), .A(n11221), .S(n10111), .Y(n11219) );
  MUX2X1 U10864 ( .B(n11223), .A(n11224), .S(n10671), .Y(n11222) );
  MUX2X1 U10865 ( .B(n11226), .A(n11227), .S(n10671), .Y(n11225) );
  MUX2X1 U10866 ( .B(n11229), .A(n11230), .S(n10671), .Y(n11228) );
  MUX2X1 U10867 ( .B(n11232), .A(n11233), .S(n10671), .Y(n11231) );
  MUX2X1 U10868 ( .B(n11235), .A(n11236), .S(n10111), .Y(n11234) );
  MUX2X1 U10869 ( .B(n11238), .A(n11239), .S(n10671), .Y(n11237) );
  MUX2X1 U10870 ( .B(n11241), .A(n11242), .S(n10671), .Y(n11240) );
  MUX2X1 U10871 ( .B(n11244), .A(n11245), .S(n10671), .Y(n11243) );
  MUX2X1 U10872 ( .B(n11247), .A(n11248), .S(n10671), .Y(n11246) );
  MUX2X1 U10873 ( .B(n11250), .A(n11251), .S(n10111), .Y(n11249) );
  MUX2X1 U10874 ( .B(n11253), .A(n11254), .S(n10671), .Y(n11252) );
  MUX2X1 U10875 ( .B(n11256), .A(n11257), .S(n10671), .Y(n11255) );
  MUX2X1 U10876 ( .B(n11259), .A(n11260), .S(n10671), .Y(n11258) );
  MUX2X1 U10877 ( .B(n11262), .A(n11263), .S(n10671), .Y(n11261) );
  MUX2X1 U10878 ( .B(n11265), .A(n11266), .S(n10111), .Y(n11264) );
  MUX2X1 U10879 ( .B(n11268), .A(n11269), .S(n10671), .Y(n11267) );
  MUX2X1 U10880 ( .B(n11271), .A(n11272), .S(n10670), .Y(n11270) );
  MUX2X1 U10881 ( .B(n11274), .A(n11275), .S(n10670), .Y(n11273) );
  MUX2X1 U10882 ( .B(n11277), .A(n11278), .S(n10670), .Y(n11276) );
  MUX2X1 U10883 ( .B(n11280), .A(n11281), .S(n10111), .Y(n11279) );
  MUX2X1 U10884 ( .B(n11283), .A(n11284), .S(n10670), .Y(n11282) );
  MUX2X1 U10885 ( .B(n11286), .A(n11287), .S(n10670), .Y(n11285) );
  MUX2X1 U10886 ( .B(n11289), .A(n11290), .S(n10670), .Y(n11288) );
  MUX2X1 U10887 ( .B(n11292), .A(n11293), .S(n10670), .Y(n11291) );
  MUX2X1 U10888 ( .B(n11295), .A(n11296), .S(n10111), .Y(n11294) );
  MUX2X1 U10889 ( .B(n11298), .A(n11299), .S(n10670), .Y(n11297) );
  MUX2X1 U10890 ( .B(n11301), .A(n11302), .S(n10670), .Y(n11300) );
  MUX2X1 U10891 ( .B(n11304), .A(n11305), .S(n10670), .Y(n11303) );
  MUX2X1 U10892 ( .B(n11307), .A(n11308), .S(n10670), .Y(n11306) );
  MUX2X1 U10893 ( .B(n11310), .A(n11311), .S(n10111), .Y(n11309) );
  MUX2X1 U10894 ( .B(n11313), .A(n11314), .S(n10670), .Y(n11312) );
  MUX2X1 U10895 ( .B(n11316), .A(n11317), .S(n10670), .Y(n11315) );
  MUX2X1 U10896 ( .B(n11319), .A(n11320), .S(n10670), .Y(n11318) );
  MUX2X1 U10897 ( .B(n11322), .A(n11323), .S(n10670), .Y(n11321) );
  MUX2X1 U10898 ( .B(n11325), .A(n11326), .S(n10111), .Y(n11324) );
  MUX2X1 U10899 ( .B(n11328), .A(n11329), .S(n10670), .Y(n11327) );
  MUX2X1 U10900 ( .B(n11331), .A(n11332), .S(n10670), .Y(n11330) );
  MUX2X1 U10901 ( .B(n11334), .A(n11335), .S(n10669), .Y(n11333) );
  MUX2X1 U10902 ( .B(n11337), .A(n11338), .S(n10669), .Y(n11336) );
  MUX2X1 U10903 ( .B(n11340), .A(n11341), .S(n10111), .Y(n11339) );
  MUX2X1 U10904 ( .B(n11343), .A(n11344), .S(n10669), .Y(n11342) );
  MUX2X1 U10905 ( .B(n11346), .A(n11347), .S(n10669), .Y(n11345) );
  MUX2X1 U10906 ( .B(n11349), .A(n11350), .S(n10669), .Y(n11348) );
  MUX2X1 U10907 ( .B(n11352), .A(n11353), .S(n10669), .Y(n11351) );
  MUX2X1 U10908 ( .B(n11355), .A(n11356), .S(n10111), .Y(n11354) );
  MUX2X1 U10909 ( .B(n11358), .A(n11359), .S(n10669), .Y(n11357) );
  MUX2X1 U10910 ( .B(n11361), .A(n11362), .S(n10669), .Y(n11360) );
  MUX2X1 U10911 ( .B(n11364), .A(n11365), .S(n10669), .Y(n11363) );
  MUX2X1 U10912 ( .B(n11367), .A(n11368), .S(n10669), .Y(n11366) );
  MUX2X1 U10913 ( .B(n11370), .A(n11371), .S(n10111), .Y(n11369) );
  MUX2X1 U10914 ( .B(n11373), .A(n11374), .S(n10669), .Y(n11372) );
  MUX2X1 U10915 ( .B(n11376), .A(n11377), .S(n10669), .Y(n11375) );
  MUX2X1 U10916 ( .B(n11379), .A(n11380), .S(n10669), .Y(n11378) );
  MUX2X1 U10917 ( .B(n11382), .A(n11383), .S(n10669), .Y(n11381) );
  MUX2X1 U10918 ( .B(n11385), .A(n11386), .S(n10111), .Y(n11384) );
  MUX2X1 U10919 ( .B(n11388), .A(n11389), .S(n10669), .Y(n11387) );
  MUX2X1 U10920 ( .B(n11391), .A(n11392), .S(n10669), .Y(n11390) );
  MUX2X1 U10921 ( .B(n11394), .A(n11395), .S(n10669), .Y(n11393) );
  MUX2X1 U10922 ( .B(n11397), .A(n11398), .S(n10668), .Y(n11396) );
  MUX2X1 U10923 ( .B(n11400), .A(n11401), .S(n10111), .Y(n11399) );
  MUX2X1 U10924 ( .B(n11403), .A(n11404), .S(n10668), .Y(n11402) );
  MUX2X1 U10925 ( .B(n11406), .A(n11407), .S(n10668), .Y(n11405) );
  MUX2X1 U10926 ( .B(n11409), .A(n11410), .S(n10668), .Y(n11408) );
  MUX2X1 U10927 ( .B(n11412), .A(n11413), .S(n10668), .Y(n11411) );
  MUX2X1 U10928 ( .B(n11415), .A(n11416), .S(n10111), .Y(n11414) );
  MUX2X1 U10929 ( .B(n11418), .A(n11419), .S(n10668), .Y(n11417) );
  MUX2X1 U10930 ( .B(n11421), .A(n11422), .S(n10668), .Y(n11420) );
  MUX2X1 U10931 ( .B(n11424), .A(n11425), .S(n10668), .Y(n11423) );
  MUX2X1 U10932 ( .B(n11427), .A(n11428), .S(n10668), .Y(n11426) );
  MUX2X1 U10933 ( .B(n11430), .A(n11431), .S(n10111), .Y(n11429) );
  MUX2X1 U10934 ( .B(n11433), .A(n11434), .S(n10668), .Y(n11432) );
  MUX2X1 U10935 ( .B(n11436), .A(n11437), .S(n10668), .Y(n11435) );
  MUX2X1 U10936 ( .B(n11439), .A(n11440), .S(n10668), .Y(n11438) );
  MUX2X1 U10937 ( .B(n11442), .A(n11443), .S(n10668), .Y(n11441) );
  MUX2X1 U10938 ( .B(n11445), .A(n11446), .S(n10111), .Y(n11444) );
  MUX2X1 U10939 ( .B(n11448), .A(n11449), .S(n10668), .Y(n11447) );
  MUX2X1 U10940 ( .B(n11451), .A(n11452), .S(n10668), .Y(n11450) );
  MUX2X1 U10941 ( .B(n11454), .A(n11455), .S(n10668), .Y(n11453) );
  MUX2X1 U10942 ( .B(n11457), .A(n11458), .S(n10668), .Y(n11456) );
  MUX2X1 U10943 ( .B(n11460), .A(n11461), .S(n10111), .Y(n11459) );
  MUX2X1 U10944 ( .B(n11463), .A(n11464), .S(n10667), .Y(n11462) );
  MUX2X1 U10945 ( .B(n11466), .A(n11467), .S(n10667), .Y(n11465) );
  MUX2X1 U10946 ( .B(n11469), .A(n11470), .S(n10667), .Y(n11468) );
  MUX2X1 U10947 ( .B(n11472), .A(n11473), .S(n10667), .Y(n11471) );
  MUX2X1 U10948 ( .B(n11475), .A(n11476), .S(n10111), .Y(n11474) );
  MUX2X1 U10949 ( .B(n11478), .A(n11479), .S(n10667), .Y(n11477) );
  MUX2X1 U10950 ( .B(n11481), .A(n11482), .S(n10667), .Y(n11480) );
  MUX2X1 U10951 ( .B(n11484), .A(n11485), .S(n10667), .Y(n11483) );
  MUX2X1 U10952 ( .B(n11487), .A(n11488), .S(n10667), .Y(n11486) );
  MUX2X1 U10953 ( .B(n11490), .A(n11491), .S(n10111), .Y(n11489) );
  MUX2X1 U10954 ( .B(n11493), .A(n11494), .S(n10667), .Y(n11492) );
  MUX2X1 U10955 ( .B(n11496), .A(n11497), .S(n10667), .Y(n11495) );
  MUX2X1 U10956 ( .B(n11499), .A(n11500), .S(n10667), .Y(n11498) );
  MUX2X1 U10957 ( .B(n11502), .A(n11503), .S(n10667), .Y(n11501) );
  MUX2X1 U10958 ( .B(n11505), .A(n11506), .S(n10111), .Y(n11504) );
  MUX2X1 U10959 ( .B(n11508), .A(n11509), .S(n10667), .Y(n11507) );
  MUX2X1 U10960 ( .B(n11511), .A(n11512), .S(n10667), .Y(n11510) );
  MUX2X1 U10961 ( .B(n11514), .A(n11515), .S(n10667), .Y(n11513) );
  MUX2X1 U10962 ( .B(n11517), .A(n11518), .S(n10667), .Y(n11516) );
  MUX2X1 U10963 ( .B(n11520), .A(n11521), .S(n10111), .Y(n11519) );
  MUX2X1 U10964 ( .B(n11523), .A(n11524), .S(n10667), .Y(n11522) );
  MUX2X1 U10965 ( .B(n11526), .A(n11527), .S(n10666), .Y(n11525) );
  MUX2X1 U10966 ( .B(n11529), .A(n11530), .S(n10666), .Y(n11528) );
  MUX2X1 U10967 ( .B(n11532), .A(n11533), .S(n10666), .Y(n11531) );
  MUX2X1 U10968 ( .B(n11535), .A(n11536), .S(n10111), .Y(n11534) );
  MUX2X1 U10969 ( .B(n11538), .A(n11539), .S(n10666), .Y(n11537) );
  MUX2X1 U10970 ( .B(n11541), .A(n11542), .S(n10666), .Y(n11540) );
  MUX2X1 U10971 ( .B(n11544), .A(n11545), .S(n10666), .Y(n11543) );
  MUX2X1 U10972 ( .B(n11547), .A(n11548), .S(n10666), .Y(n11546) );
  MUX2X1 U10973 ( .B(n11550), .A(n11551), .S(n10111), .Y(n11549) );
  MUX2X1 U10974 ( .B(n11553), .A(n11554), .S(n10666), .Y(n11552) );
  MUX2X1 U10975 ( .B(n11556), .A(n11557), .S(n10666), .Y(n11555) );
  MUX2X1 U10976 ( .B(n11559), .A(n11560), .S(n10666), .Y(n11558) );
  MUX2X1 U10977 ( .B(n11562), .A(n11563), .S(n10666), .Y(n11561) );
  MUX2X1 U10978 ( .B(n11565), .A(n11566), .S(n10111), .Y(n11564) );
  MUX2X1 U10979 ( .B(n11568), .A(n11569), .S(n10666), .Y(n11567) );
  MUX2X1 U10980 ( .B(n11571), .A(n11572), .S(n10666), .Y(n11570) );
  MUX2X1 U10981 ( .B(n11574), .A(n11575), .S(n10666), .Y(n11573) );
  MUX2X1 U10982 ( .B(n11577), .A(n11578), .S(n10666), .Y(n11576) );
  MUX2X1 U10983 ( .B(n11580), .A(n11581), .S(n10111), .Y(n11579) );
  MUX2X1 U10984 ( .B(n11583), .A(n11584), .S(n10666), .Y(n11582) );
  MUX2X1 U10985 ( .B(n11586), .A(n11587), .S(n10666), .Y(n11585) );
  MUX2X1 U10986 ( .B(n11589), .A(n11590), .S(n10665), .Y(n11588) );
  MUX2X1 U10987 ( .B(n11592), .A(n11593), .S(n10665), .Y(n11591) );
  MUX2X1 U10988 ( .B(n11595), .A(n11596), .S(n10111), .Y(n11594) );
  MUX2X1 U10989 ( .B(n11598), .A(n11599), .S(n10665), .Y(n11597) );
  MUX2X1 U10990 ( .B(n11601), .A(n11602), .S(n10665), .Y(n11600) );
  MUX2X1 U10991 ( .B(n11604), .A(n11605), .S(n10665), .Y(n11603) );
  MUX2X1 U10992 ( .B(n11607), .A(n11608), .S(n10665), .Y(n11606) );
  MUX2X1 U10993 ( .B(n11610), .A(n11611), .S(n10111), .Y(n11609) );
  MUX2X1 U10994 ( .B(n11613), .A(n11614), .S(n10665), .Y(n11612) );
  MUX2X1 U10995 ( .B(n11616), .A(n11617), .S(n10665), .Y(n11615) );
  MUX2X1 U10996 ( .B(n11619), .A(n11620), .S(n10665), .Y(n11618) );
  MUX2X1 U10997 ( .B(n11622), .A(n11623), .S(n10665), .Y(n11621) );
  MUX2X1 U10998 ( .B(n11625), .A(n11626), .S(n10111), .Y(n11624) );
  MUX2X1 U10999 ( .B(n11628), .A(n11629), .S(n10665), .Y(n11627) );
  MUX2X1 U11000 ( .B(n11631), .A(n11632), .S(n10665), .Y(n11630) );
  MUX2X1 U11001 ( .B(n11634), .A(n11635), .S(n10665), .Y(n11633) );
  MUX2X1 U11002 ( .B(n11637), .A(n11638), .S(n10665), .Y(n11636) );
  MUX2X1 U11003 ( .B(n11640), .A(n11641), .S(n10111), .Y(n11639) );
  MUX2X1 U11004 ( .B(n11643), .A(n11644), .S(n10665), .Y(n11642) );
  MUX2X1 U11005 ( .B(n11646), .A(n11647), .S(n10665), .Y(n11645) );
  MUX2X1 U11006 ( .B(n11649), .A(n11650), .S(n10665), .Y(n11648) );
  MUX2X1 U11007 ( .B(n11652), .A(n11653), .S(n10664), .Y(n11651) );
  MUX2X1 U11008 ( .B(n11655), .A(n11656), .S(n10111), .Y(n11654) );
  MUX2X1 U11009 ( .B(n11658), .A(n11659), .S(n10664), .Y(n11657) );
  MUX2X1 U11010 ( .B(n11661), .A(n11662), .S(n10664), .Y(n11660) );
  MUX2X1 U11011 ( .B(n11664), .A(n11665), .S(n10664), .Y(n11663) );
  MUX2X1 U11012 ( .B(n11667), .A(n11668), .S(n10664), .Y(n11666) );
  MUX2X1 U11013 ( .B(n11670), .A(n11671), .S(n10111), .Y(n11669) );
  MUX2X1 U11014 ( .B(n11673), .A(n11674), .S(n10664), .Y(n11672) );
  MUX2X1 U11015 ( .B(n11676), .A(n11677), .S(n10664), .Y(n11675) );
  MUX2X1 U11016 ( .B(n11679), .A(n11680), .S(n10664), .Y(n11678) );
  MUX2X1 U11017 ( .B(n11682), .A(n11683), .S(n10664), .Y(n11681) );
  MUX2X1 U11018 ( .B(n11685), .A(n11686), .S(n10111), .Y(n11684) );
  MUX2X1 U11019 ( .B(n11688), .A(n11689), .S(n10664), .Y(n11687) );
  MUX2X1 U11020 ( .B(n11691), .A(n11692), .S(n10664), .Y(n11690) );
  MUX2X1 U11021 ( .B(n11694), .A(n11695), .S(n10664), .Y(n11693) );
  MUX2X1 U11022 ( .B(n11697), .A(n11698), .S(n10664), .Y(n11696) );
  MUX2X1 U11023 ( .B(n11700), .A(n11701), .S(n10111), .Y(n11699) );
  MUX2X1 U11024 ( .B(n11703), .A(n11704), .S(n10664), .Y(n11702) );
  MUX2X1 U11025 ( .B(n11706), .A(n11707), .S(n10664), .Y(n11705) );
  MUX2X1 U11026 ( .B(n11709), .A(n11710), .S(n10664), .Y(n11708) );
  MUX2X1 U11027 ( .B(n11712), .A(n11713), .S(n10664), .Y(n11711) );
  MUX2X1 U11028 ( .B(n11715), .A(n11716), .S(n10111), .Y(n11714) );
  MUX2X1 U11029 ( .B(n11718), .A(n11719), .S(n10663), .Y(n11717) );
  MUX2X1 U11030 ( .B(n11721), .A(n11722), .S(n10663), .Y(n11720) );
  MUX2X1 U11031 ( .B(n11724), .A(n11725), .S(n10663), .Y(n11723) );
  MUX2X1 U11032 ( .B(n11727), .A(n11728), .S(n10663), .Y(n11726) );
  MUX2X1 U11033 ( .B(n11730), .A(n11731), .S(n10111), .Y(n11729) );
  MUX2X1 U11034 ( .B(n11733), .A(n11734), .S(n10663), .Y(n11732) );
  MUX2X1 U11035 ( .B(n11736), .A(n11737), .S(n10663), .Y(n11735) );
  MUX2X1 U11036 ( .B(n11739), .A(n11740), .S(n10663), .Y(n11738) );
  MUX2X1 U11037 ( .B(n11742), .A(n11743), .S(n10663), .Y(n11741) );
  MUX2X1 U11038 ( .B(n11745), .A(n11746), .S(n10111), .Y(n11744) );
  MUX2X1 U11039 ( .B(n11748), .A(n11749), .S(n10663), .Y(n11747) );
  MUX2X1 U11040 ( .B(n11751), .A(n11752), .S(n10663), .Y(n11750) );
  MUX2X1 U11041 ( .B(n11754), .A(n11755), .S(n10663), .Y(n11753) );
  MUX2X1 U11042 ( .B(n11757), .A(n11758), .S(n10663), .Y(n11756) );
  MUX2X1 U11043 ( .B(n11760), .A(n11761), .S(n10111), .Y(n11759) );
  MUX2X1 U11044 ( .B(n7212), .A(n8742), .S(n10689), .Y(n10744) );
  MUX2X1 U11045 ( .B(n7314), .A(n8844), .S(n10713), .Y(n10743) );
  MUX2X1 U11046 ( .B(n7416), .A(n8946), .S(n10713), .Y(n10747) );
  MUX2X1 U11047 ( .B(n7518), .A(n9048), .S(n10713), .Y(n10746) );
  MUX2X1 U11048 ( .B(n10745), .A(n10742), .S(n10649), .Y(n10756) );
  MUX2X1 U11049 ( .B(n6906), .A(n8538), .S(n10712), .Y(n10750) );
  MUX2X1 U11050 ( .B(n6702), .A(n8436), .S(n10712), .Y(n10749) );
  MUX2X1 U11051 ( .B(n6804), .A(n8334), .S(n10712), .Y(n10753) );
  MUX2X1 U11052 ( .B(n7008), .A(n8640), .S(n10712), .Y(n10752) );
  MUX2X1 U11053 ( .B(n10751), .A(n10748), .S(n10657), .Y(n10755) );
  MUX2X1 U11054 ( .B(n7620), .A(n9150), .S(n10712), .Y(n10759) );
  MUX2X1 U11055 ( .B(n7722), .A(n9252), .S(n10712), .Y(n10758) );
  MUX2X1 U11056 ( .B(n7824), .A(n9354), .S(n10712), .Y(n10762) );
  MUX2X1 U11057 ( .B(n7926), .A(n9456), .S(n10712), .Y(n10761) );
  MUX2X1 U11058 ( .B(n10760), .A(n10757), .S(n10657), .Y(n10771) );
  MUX2X1 U11059 ( .B(n8028), .A(n9558), .S(n10712), .Y(n10765) );
  MUX2X1 U11060 ( .B(n8130), .A(n9660), .S(n10712), .Y(n10764) );
  MUX2X1 U11061 ( .B(n8232), .A(n9762), .S(n10712), .Y(n10768) );
  MUX2X1 U11062 ( .B(n7110), .A(n9864), .S(n10712), .Y(n10767) );
  MUX2X1 U11063 ( .B(n10766), .A(n10763), .S(n10657), .Y(n10770) );
  MUX2X1 U11064 ( .B(n10769), .A(n10754), .S(n10529), .Y(n11762) );
  INVX2 U11065 ( .A(n11762), .Y(n104) );
  MUX2X1 U11066 ( .B(n7215), .A(n8745), .S(n10712), .Y(n10774) );
  MUX2X1 U11067 ( .B(n7317), .A(n8847), .S(n10712), .Y(n10773) );
  MUX2X1 U11068 ( .B(n7419), .A(n8949), .S(n10712), .Y(n10777) );
  MUX2X1 U11069 ( .B(n7521), .A(n9051), .S(n10712), .Y(n10776) );
  MUX2X1 U11070 ( .B(n10775), .A(n10772), .S(n10657), .Y(n10786) );
  MUX2X1 U11071 ( .B(n6909), .A(n8541), .S(n10712), .Y(n10780) );
  MUX2X1 U11072 ( .B(n6705), .A(n8439), .S(n10711), .Y(n10779) );
  MUX2X1 U11073 ( .B(n6807), .A(n8337), .S(n10711), .Y(n10783) );
  MUX2X1 U11074 ( .B(n7011), .A(n8643), .S(n10711), .Y(n10782) );
  MUX2X1 U11075 ( .B(n10781), .A(n10778), .S(n10656), .Y(n10785) );
  MUX2X1 U11076 ( .B(n7623), .A(n9153), .S(n10711), .Y(n10789) );
  MUX2X1 U11077 ( .B(n7725), .A(n9255), .S(n10711), .Y(n10788) );
  MUX2X1 U11078 ( .B(n7827), .A(n9357), .S(n10711), .Y(n10792) );
  MUX2X1 U11079 ( .B(n7929), .A(n9459), .S(n10711), .Y(n10791) );
  MUX2X1 U11080 ( .B(n10790), .A(n10787), .S(n10656), .Y(n10801) );
  MUX2X1 U11081 ( .B(n8031), .A(n9561), .S(n10711), .Y(n10795) );
  MUX2X1 U11082 ( .B(n8133), .A(n9663), .S(n10711), .Y(n10794) );
  MUX2X1 U11083 ( .B(n8235), .A(n9765), .S(n10711), .Y(n10798) );
  MUX2X1 U11084 ( .B(n7113), .A(n9867), .S(n10711), .Y(n10797) );
  MUX2X1 U11085 ( .B(n10796), .A(n10793), .S(n10656), .Y(n10800) );
  MUX2X1 U11086 ( .B(n10799), .A(n10784), .S(n10529), .Y(n11763) );
  INVX2 U11087 ( .A(n11763), .Y(n103) );
  MUX2X1 U11088 ( .B(n7218), .A(n8748), .S(n10711), .Y(n10804) );
  MUX2X1 U11089 ( .B(n7320), .A(n8850), .S(n10711), .Y(n10803) );
  MUX2X1 U11090 ( .B(n7422), .A(n8952), .S(n10711), .Y(n10807) );
  MUX2X1 U11091 ( .B(n7524), .A(n9054), .S(n10711), .Y(n10806) );
  MUX2X1 U11092 ( .B(n10805), .A(n10802), .S(n10656), .Y(n10816) );
  MUX2X1 U11093 ( .B(n6912), .A(n8544), .S(n10711), .Y(n10810) );
  MUX2X1 U11094 ( .B(n6708), .A(n8442), .S(n10711), .Y(n10809) );
  MUX2X1 U11095 ( .B(n6810), .A(n8340), .S(n10710), .Y(n10813) );
  MUX2X1 U11096 ( .B(n7014), .A(n8646), .S(n10710), .Y(n10812) );
  MUX2X1 U11097 ( .B(n10811), .A(n10808), .S(n10656), .Y(n10815) );
  MUX2X1 U11098 ( .B(n7626), .A(n9156), .S(n10710), .Y(n10819) );
  MUX2X1 U11099 ( .B(n7728), .A(n9258), .S(n10710), .Y(n10818) );
  MUX2X1 U11100 ( .B(n7830), .A(n9360), .S(n10710), .Y(n10822) );
  MUX2X1 U11101 ( .B(n7932), .A(n9462), .S(n10710), .Y(n10821) );
  MUX2X1 U11102 ( .B(n10820), .A(n10817), .S(n10656), .Y(n10831) );
  MUX2X1 U11103 ( .B(n8034), .A(n9564), .S(n10710), .Y(n10825) );
  MUX2X1 U11104 ( .B(n8136), .A(n9666), .S(n10710), .Y(n10824) );
  MUX2X1 U11105 ( .B(n8238), .A(n9768), .S(n10710), .Y(n10828) );
  MUX2X1 U11106 ( .B(n7116), .A(n9870), .S(n10710), .Y(n10827) );
  MUX2X1 U11107 ( .B(n10826), .A(n10823), .S(n10656), .Y(n10830) );
  MUX2X1 U11108 ( .B(n10829), .A(n10814), .S(n10529), .Y(n11764) );
  INVX2 U11109 ( .A(n11764), .Y(n102) );
  MUX2X1 U11110 ( .B(n7221), .A(n8751), .S(n10710), .Y(n10834) );
  MUX2X1 U11111 ( .B(n7323), .A(n8853), .S(n10710), .Y(n10833) );
  MUX2X1 U11112 ( .B(n7425), .A(n8955), .S(n10710), .Y(n10837) );
  MUX2X1 U11113 ( .B(n7527), .A(n9057), .S(n10710), .Y(n10836) );
  MUX2X1 U11114 ( .B(n10835), .A(n10832), .S(n10656), .Y(n10846) );
  MUX2X1 U11115 ( .B(n6915), .A(n8547), .S(n10710), .Y(n10840) );
  MUX2X1 U11116 ( .B(n6711), .A(n8445), .S(n10710), .Y(n10839) );
  MUX2X1 U11117 ( .B(n6813), .A(n8343), .S(n10710), .Y(n10843) );
  MUX2X1 U11118 ( .B(n7017), .A(n8649), .S(n10709), .Y(n10842) );
  MUX2X1 U11119 ( .B(n10841), .A(n10838), .S(n10656), .Y(n10845) );
  MUX2X1 U11120 ( .B(n7629), .A(n9159), .S(n10709), .Y(n10849) );
  MUX2X1 U11121 ( .B(n7731), .A(n9261), .S(n10709), .Y(n10848) );
  MUX2X1 U11122 ( .B(n7833), .A(n9363), .S(n10709), .Y(n10852) );
  MUX2X1 U11123 ( .B(n7935), .A(n9465), .S(n10709), .Y(n10851) );
  MUX2X1 U11124 ( .B(n10850), .A(n10847), .S(n10656), .Y(n10861) );
  MUX2X1 U11125 ( .B(n8037), .A(n9567), .S(n10709), .Y(n10855) );
  MUX2X1 U11126 ( .B(n8139), .A(n9669), .S(n10709), .Y(n10854) );
  MUX2X1 U11127 ( .B(n8241), .A(n9771), .S(n10709), .Y(n10858) );
  MUX2X1 U11128 ( .B(n7119), .A(n9873), .S(n10709), .Y(n10857) );
  MUX2X1 U11129 ( .B(n10856), .A(n10853), .S(n10656), .Y(n10860) );
  MUX2X1 U11130 ( .B(n10859), .A(n10844), .S(n10529), .Y(n11765) );
  INVX2 U11131 ( .A(n11765), .Y(n101) );
  MUX2X1 U11132 ( .B(n7224), .A(n8754), .S(n10709), .Y(n10864) );
  MUX2X1 U11133 ( .B(n7326), .A(n8856), .S(n10709), .Y(n10863) );
  MUX2X1 U11134 ( .B(n7428), .A(n8958), .S(n10709), .Y(n10867) );
  MUX2X1 U11135 ( .B(n7530), .A(n9060), .S(n10709), .Y(n10866) );
  MUX2X1 U11136 ( .B(n10865), .A(n10862), .S(n10656), .Y(n10876) );
  MUX2X1 U11137 ( .B(n6918), .A(n8550), .S(n10709), .Y(n10870) );
  MUX2X1 U11138 ( .B(n6714), .A(n8448), .S(n10709), .Y(n10869) );
  MUX2X1 U11139 ( .B(n6816), .A(n8346), .S(n10709), .Y(n10873) );
  MUX2X1 U11140 ( .B(n7020), .A(n8652), .S(n10708), .Y(n10872) );
  MUX2X1 U11141 ( .B(n10871), .A(n10868), .S(n10656), .Y(n10875) );
  MUX2X1 U11142 ( .B(n7632), .A(n9162), .S(n10708), .Y(n10879) );
  MUX2X1 U11143 ( .B(n7734), .A(n9264), .S(n10708), .Y(n10878) );
  MUX2X1 U11144 ( .B(n7836), .A(n9366), .S(n10708), .Y(n10882) );
  MUX2X1 U11145 ( .B(n7938), .A(n9468), .S(n10708), .Y(n10881) );
  MUX2X1 U11146 ( .B(n10880), .A(n10877), .S(n10656), .Y(n10891) );
  MUX2X1 U11147 ( .B(n8040), .A(n9570), .S(n10708), .Y(n10885) );
  MUX2X1 U11148 ( .B(n8142), .A(n9672), .S(n10708), .Y(n10884) );
  MUX2X1 U11149 ( .B(n8244), .A(n9774), .S(n10708), .Y(n10888) );
  MUX2X1 U11150 ( .B(n7122), .A(n9876), .S(n10708), .Y(n10887) );
  MUX2X1 U11151 ( .B(n10886), .A(n10883), .S(n10656), .Y(n10890) );
  MUX2X1 U11152 ( .B(n10889), .A(n10874), .S(n10529), .Y(n11766) );
  INVX2 U11153 ( .A(n11766), .Y(n100) );
  MUX2X1 U11154 ( .B(n7227), .A(n8757), .S(n10708), .Y(n10894) );
  MUX2X1 U11155 ( .B(n7329), .A(n8859), .S(n10708), .Y(n10893) );
  MUX2X1 U11156 ( .B(n7431), .A(n8961), .S(n10708), .Y(n10897) );
  MUX2X1 U11157 ( .B(n7533), .A(n9063), .S(n10708), .Y(n10896) );
  MUX2X1 U11158 ( .B(n10895), .A(n10892), .S(n10656), .Y(n10906) );
  MUX2X1 U11159 ( .B(n6921), .A(n8553), .S(n10708), .Y(n10900) );
  MUX2X1 U11160 ( .B(n6717), .A(n8451), .S(n10708), .Y(n10899) );
  MUX2X1 U11161 ( .B(n6819), .A(n8349), .S(n10708), .Y(n10903) );
  MUX2X1 U11162 ( .B(n7023), .A(n8655), .S(n10708), .Y(n10902) );
  MUX2X1 U11163 ( .B(n10901), .A(n10898), .S(n10655), .Y(n10905) );
  MUX2X1 U11164 ( .B(n7635), .A(n9165), .S(n10707), .Y(n10909) );
  MUX2X1 U11165 ( .B(n7737), .A(n9267), .S(n10707), .Y(n10908) );
  MUX2X1 U11166 ( .B(n7839), .A(n9369), .S(n10707), .Y(n10912) );
  MUX2X1 U11167 ( .B(n7941), .A(n9471), .S(n10707), .Y(n10911) );
  MUX2X1 U11168 ( .B(n10910), .A(n10907), .S(n10656), .Y(n10921) );
  MUX2X1 U11169 ( .B(n8043), .A(n9573), .S(n10707), .Y(n10915) );
  MUX2X1 U11170 ( .B(n8145), .A(n9675), .S(n10707), .Y(n10914) );
  MUX2X1 U11171 ( .B(n8247), .A(n9777), .S(n10707), .Y(n10918) );
  MUX2X1 U11172 ( .B(n7125), .A(n9879), .S(n10707), .Y(n10917) );
  MUX2X1 U11173 ( .B(n10916), .A(n10913), .S(n10655), .Y(n10920) );
  MUX2X1 U11174 ( .B(n10919), .A(n10904), .S(n10529), .Y(n11767) );
  INVX2 U11175 ( .A(n11767), .Y(n99) );
  MUX2X1 U11176 ( .B(n7230), .A(n8760), .S(n10707), .Y(n10924) );
  MUX2X1 U11177 ( .B(n7332), .A(n8862), .S(n10707), .Y(n10923) );
  MUX2X1 U11178 ( .B(n7434), .A(n8964), .S(n10707), .Y(n10927) );
  MUX2X1 U11179 ( .B(n7536), .A(n9066), .S(n10707), .Y(n10926) );
  MUX2X1 U11180 ( .B(n10925), .A(n10922), .S(n10655), .Y(n10936) );
  MUX2X1 U11181 ( .B(n6924), .A(n8556), .S(n10707), .Y(n10930) );
  MUX2X1 U11182 ( .B(n6720), .A(n8454), .S(n10707), .Y(n10929) );
  MUX2X1 U11183 ( .B(n6822), .A(n8352), .S(n10707), .Y(n10933) );
  MUX2X1 U11184 ( .B(n7026), .A(n8658), .S(n10707), .Y(n10932) );
  MUX2X1 U11185 ( .B(n10931), .A(n10928), .S(n10655), .Y(n10935) );
  MUX2X1 U11186 ( .B(n7638), .A(n9168), .S(n10707), .Y(n10939) );
  MUX2X1 U11187 ( .B(n7740), .A(n9270), .S(n10706), .Y(n10938) );
  MUX2X1 U11188 ( .B(n7842), .A(n9372), .S(n10706), .Y(n10942) );
  MUX2X1 U11189 ( .B(n7944), .A(n9474), .S(n10706), .Y(n10941) );
  MUX2X1 U11190 ( .B(n10940), .A(n10937), .S(n10655), .Y(n10951) );
  MUX2X1 U11191 ( .B(n8046), .A(n9576), .S(n10706), .Y(n10945) );
  MUX2X1 U11192 ( .B(n8148), .A(n9678), .S(n10706), .Y(n10944) );
  MUX2X1 U11193 ( .B(n8250), .A(n9780), .S(n10706), .Y(n10948) );
  MUX2X1 U11194 ( .B(n7128), .A(n9882), .S(n10706), .Y(n10947) );
  MUX2X1 U11195 ( .B(n10946), .A(n10943), .S(n10655), .Y(n10950) );
  MUX2X1 U11196 ( .B(n10949), .A(n10934), .S(n10529), .Y(n11768) );
  INVX2 U11197 ( .A(n11768), .Y(n98) );
  MUX2X1 U11198 ( .B(n7233), .A(n8763), .S(n10706), .Y(n10954) );
  MUX2X1 U11199 ( .B(n7335), .A(n8865), .S(n10706), .Y(n10953) );
  MUX2X1 U11200 ( .B(n7437), .A(n8967), .S(n10706), .Y(n10957) );
  MUX2X1 U11201 ( .B(n7539), .A(n9069), .S(n10706), .Y(n10956) );
  MUX2X1 U11202 ( .B(n10955), .A(n10952), .S(n10655), .Y(n10966) );
  MUX2X1 U11203 ( .B(n6927), .A(n8559), .S(n10706), .Y(n10960) );
  MUX2X1 U11204 ( .B(n6723), .A(n8457), .S(n10706), .Y(n10959) );
  MUX2X1 U11205 ( .B(n6825), .A(n8355), .S(n10706), .Y(n10963) );
  MUX2X1 U11206 ( .B(n7029), .A(n8661), .S(n10706), .Y(n10962) );
  MUX2X1 U11207 ( .B(n10961), .A(n10958), .S(n10655), .Y(n10965) );
  MUX2X1 U11208 ( .B(n7641), .A(n9171), .S(n10706), .Y(n10969) );
  MUX2X1 U11209 ( .B(n7743), .A(n9273), .S(n10706), .Y(n10968) );
  MUX2X1 U11210 ( .B(n7845), .A(n9375), .S(n10705), .Y(n10972) );
  MUX2X1 U11211 ( .B(n7947), .A(n9477), .S(n10705), .Y(n10971) );
  MUX2X1 U11212 ( .B(n10970), .A(n10967), .S(n10655), .Y(n10981) );
  MUX2X1 U11213 ( .B(n8049), .A(n9579), .S(n10705), .Y(n10975) );
  MUX2X1 U11214 ( .B(n8151), .A(n9681), .S(n10705), .Y(n10974) );
  MUX2X1 U11215 ( .B(n8253), .A(n9783), .S(n10705), .Y(n10978) );
  MUX2X1 U11216 ( .B(n7131), .A(n9885), .S(n10705), .Y(n10977) );
  MUX2X1 U11217 ( .B(n10976), .A(n10973), .S(n10655), .Y(n10980) );
  MUX2X1 U11218 ( .B(n10979), .A(n10964), .S(n10529), .Y(n11769) );
  INVX2 U11219 ( .A(n11769), .Y(n97) );
  MUX2X1 U11220 ( .B(n7236), .A(n8766), .S(n10705), .Y(n10984) );
  MUX2X1 U11221 ( .B(n7338), .A(n8868), .S(n10705), .Y(n10983) );
  MUX2X1 U11222 ( .B(n7440), .A(n8970), .S(n10705), .Y(n10987) );
  MUX2X1 U11223 ( .B(n7542), .A(n9072), .S(n10705), .Y(n10986) );
  MUX2X1 U11224 ( .B(n10985), .A(n10982), .S(n10655), .Y(n10996) );
  MUX2X1 U11225 ( .B(n6930), .A(n8562), .S(n10705), .Y(n10990) );
  MUX2X1 U11226 ( .B(n6726), .A(n8460), .S(n10705), .Y(n10989) );
  MUX2X1 U11227 ( .B(n6828), .A(n8358), .S(n10705), .Y(n10993) );
  MUX2X1 U11228 ( .B(n7032), .A(n8664), .S(n10705), .Y(n10992) );
  MUX2X1 U11229 ( .B(n10991), .A(n10988), .S(n10655), .Y(n10995) );
  MUX2X1 U11230 ( .B(n7644), .A(n9174), .S(n10709), .Y(n10999) );
  MUX2X1 U11231 ( .B(n7746), .A(n9276), .S(n10721), .Y(n10998) );
  MUX2X1 U11232 ( .B(n7848), .A(n9378), .S(n10721), .Y(n11002) );
  MUX2X1 U11233 ( .B(n7950), .A(n9480), .S(n10721), .Y(n11001) );
  MUX2X1 U11234 ( .B(n11000), .A(n10997), .S(n10655), .Y(n11011) );
  MUX2X1 U11235 ( .B(n8052), .A(n9582), .S(n10720), .Y(n11005) );
  MUX2X1 U11236 ( .B(n8154), .A(n9684), .S(n10720), .Y(n11004) );
  MUX2X1 U11237 ( .B(n8256), .A(n9786), .S(n10720), .Y(n11008) );
  MUX2X1 U11238 ( .B(n7134), .A(n9888), .S(n10720), .Y(n11007) );
  MUX2X1 U11239 ( .B(n11006), .A(n11003), .S(n10655), .Y(n11010) );
  MUX2X1 U11240 ( .B(n11009), .A(n10994), .S(n10529), .Y(n11770) );
  INVX2 U11241 ( .A(n11770), .Y(n96) );
  MUX2X1 U11242 ( .B(n7239), .A(n8769), .S(n10720), .Y(n11014) );
  MUX2X1 U11243 ( .B(n7341), .A(n8871), .S(n10720), .Y(n11013) );
  MUX2X1 U11244 ( .B(n7443), .A(n8973), .S(n10720), .Y(n11017) );
  MUX2X1 U11245 ( .B(n7545), .A(n9075), .S(n10720), .Y(n11016) );
  MUX2X1 U11246 ( .B(n11015), .A(n11012), .S(n10655), .Y(n11026) );
  MUX2X1 U11247 ( .B(n6933), .A(n8565), .S(n10720), .Y(n11020) );
  MUX2X1 U11248 ( .B(n6729), .A(n8463), .S(n10720), .Y(n11019) );
  MUX2X1 U11249 ( .B(n6831), .A(n8361), .S(n10720), .Y(n11023) );
  MUX2X1 U11250 ( .B(n7035), .A(n8667), .S(n10720), .Y(n11022) );
  MUX2X1 U11251 ( .B(n11021), .A(n11018), .S(n10655), .Y(n11025) );
  MUX2X1 U11252 ( .B(n7647), .A(n9177), .S(n10720), .Y(n11029) );
  MUX2X1 U11253 ( .B(n7749), .A(n9279), .S(n10720), .Y(n11028) );
  MUX2X1 U11254 ( .B(n7851), .A(n9381), .S(n10720), .Y(n11032) );
  MUX2X1 U11255 ( .B(n7953), .A(n9483), .S(n10720), .Y(n11031) );
  MUX2X1 U11256 ( .B(n11030), .A(n11027), .S(n10655), .Y(n11041) );
  MUX2X1 U11257 ( .B(n8055), .A(n9585), .S(n10720), .Y(n11035) );
  MUX2X1 U11258 ( .B(n8157), .A(n9687), .S(n10719), .Y(n11034) );
  MUX2X1 U11259 ( .B(n8259), .A(n9789), .S(n10719), .Y(n11038) );
  MUX2X1 U11260 ( .B(n7137), .A(n9891), .S(n10719), .Y(n11037) );
  MUX2X1 U11261 ( .B(n11036), .A(n11033), .S(n10654), .Y(n11040) );
  MUX2X1 U11262 ( .B(n11039), .A(n11024), .S(n10529), .Y(n11771) );
  INVX2 U11263 ( .A(n11771), .Y(n95) );
  MUX2X1 U11264 ( .B(n7242), .A(n8772), .S(n10719), .Y(n11044) );
  MUX2X1 U11265 ( .B(n7344), .A(n8874), .S(n10719), .Y(n11043) );
  MUX2X1 U11266 ( .B(n7446), .A(n8976), .S(n10719), .Y(n11047) );
  MUX2X1 U11267 ( .B(n7548), .A(n9078), .S(n10719), .Y(n11046) );
  MUX2X1 U11268 ( .B(n11045), .A(n11042), .S(n10654), .Y(n11056) );
  MUX2X1 U11269 ( .B(n6936), .A(n8568), .S(n10719), .Y(n11050) );
  MUX2X1 U11270 ( .B(n6732), .A(n8466), .S(n10719), .Y(n11049) );
  MUX2X1 U11271 ( .B(n6834), .A(n8364), .S(n10719), .Y(n11053) );
  MUX2X1 U11272 ( .B(n7038), .A(n8670), .S(n10719), .Y(n11052) );
  MUX2X1 U11273 ( .B(n11051), .A(n11048), .S(n10654), .Y(n11055) );
  MUX2X1 U11274 ( .B(n7650), .A(n9180), .S(n10719), .Y(n11059) );
  MUX2X1 U11275 ( .B(n7752), .A(n9282), .S(n10719), .Y(n11058) );
  MUX2X1 U11276 ( .B(n7854), .A(n9384), .S(n10719), .Y(n11062) );
  MUX2X1 U11277 ( .B(n7956), .A(n9486), .S(n10719), .Y(n11061) );
  MUX2X1 U11278 ( .B(n11060), .A(n11057), .S(n10654), .Y(n11071) );
  MUX2X1 U11279 ( .B(n8058), .A(n9588), .S(n10719), .Y(n11065) );
  MUX2X1 U11280 ( .B(n8160), .A(n9690), .S(n10719), .Y(n11064) );
  MUX2X1 U11281 ( .B(n8262), .A(n9792), .S(n10718), .Y(n11068) );
  MUX2X1 U11282 ( .B(n7140), .A(n9894), .S(n10718), .Y(n11067) );
  MUX2X1 U11283 ( .B(n11066), .A(n11063), .S(n10654), .Y(n11070) );
  MUX2X1 U11284 ( .B(n11069), .A(n11054), .S(n10529), .Y(n11772) );
  INVX2 U11285 ( .A(n11772), .Y(n94) );
  MUX2X1 U11286 ( .B(n7245), .A(n8775), .S(n10718), .Y(n11074) );
  MUX2X1 U11287 ( .B(n7347), .A(n8877), .S(n10718), .Y(n11073) );
  MUX2X1 U11288 ( .B(n7449), .A(n8979), .S(n10718), .Y(n11077) );
  MUX2X1 U11289 ( .B(n7551), .A(n9081), .S(n10718), .Y(n11076) );
  MUX2X1 U11290 ( .B(n11075), .A(n11072), .S(n10654), .Y(n11086) );
  MUX2X1 U11291 ( .B(n6939), .A(n8571), .S(n10718), .Y(n11080) );
  MUX2X1 U11292 ( .B(n6735), .A(n8469), .S(n10718), .Y(n11079) );
  MUX2X1 U11293 ( .B(n6837), .A(n8367), .S(n10718), .Y(n11083) );
  MUX2X1 U11294 ( .B(n7041), .A(n8673), .S(n10718), .Y(n11082) );
  MUX2X1 U11295 ( .B(n11081), .A(n11078), .S(n10654), .Y(n11085) );
  MUX2X1 U11296 ( .B(n7653), .A(n9183), .S(n10718), .Y(n11089) );
  MUX2X1 U11297 ( .B(n7755), .A(n9285), .S(n10718), .Y(n11088) );
  MUX2X1 U11298 ( .B(n7857), .A(n9387), .S(n10718), .Y(n11092) );
  MUX2X1 U11299 ( .B(n7959), .A(n9489), .S(n10718), .Y(n11091) );
  MUX2X1 U11300 ( .B(n11090), .A(n11087), .S(n10654), .Y(n11101) );
  MUX2X1 U11301 ( .B(n8061), .A(n9591), .S(n10718), .Y(n11095) );
  MUX2X1 U11302 ( .B(n8163), .A(n9693), .S(n10718), .Y(n11094) );
  MUX2X1 U11303 ( .B(n8265), .A(n9795), .S(n10718), .Y(n11098) );
  MUX2X1 U11304 ( .B(n7143), .A(n9897), .S(n10717), .Y(n11097) );
  MUX2X1 U11305 ( .B(n11096), .A(n11093), .S(n10654), .Y(n11100) );
  MUX2X1 U11306 ( .B(n11099), .A(n11084), .S(n10529), .Y(n11773) );
  INVX2 U11307 ( .A(n11773), .Y(n93) );
  MUX2X1 U11308 ( .B(n7248), .A(n8778), .S(n10717), .Y(n11104) );
  MUX2X1 U11309 ( .B(n7350), .A(n8880), .S(n10717), .Y(n11103) );
  MUX2X1 U11310 ( .B(n7452), .A(n8982), .S(n10717), .Y(n11107) );
  MUX2X1 U11311 ( .B(n7554), .A(n9084), .S(n10717), .Y(n11106) );
  MUX2X1 U11312 ( .B(n11105), .A(n11102), .S(n10654), .Y(n11116) );
  MUX2X1 U11313 ( .B(n6942), .A(n8574), .S(n10717), .Y(n11110) );
  MUX2X1 U11314 ( .B(n6738), .A(n8472), .S(n10717), .Y(n11109) );
  MUX2X1 U11315 ( .B(n6840), .A(n8370), .S(n10717), .Y(n11113) );
  MUX2X1 U11316 ( .B(n7044), .A(n8676), .S(n10717), .Y(n11112) );
  MUX2X1 U11317 ( .B(n11111), .A(n11108), .S(n10654), .Y(n11115) );
  MUX2X1 U11318 ( .B(n7656), .A(n9186), .S(n10717), .Y(n11119) );
  MUX2X1 U11319 ( .B(n7758), .A(n9288), .S(n10717), .Y(n11118) );
  MUX2X1 U11320 ( .B(n7860), .A(n9390), .S(n10717), .Y(n11122) );
  MUX2X1 U11321 ( .B(n7962), .A(n9492), .S(n10717), .Y(n11121) );
  MUX2X1 U11322 ( .B(n11120), .A(n11117), .S(n10654), .Y(n11131) );
  MUX2X1 U11323 ( .B(n8064), .A(n9594), .S(n10717), .Y(n11125) );
  MUX2X1 U11324 ( .B(n8166), .A(n9696), .S(n10717), .Y(n11124) );
  MUX2X1 U11325 ( .B(n8268), .A(n9798), .S(n10717), .Y(n11128) );
  MUX2X1 U11326 ( .B(n7146), .A(n9900), .S(n10716), .Y(n11127) );
  MUX2X1 U11327 ( .B(n11126), .A(n11123), .S(n10654), .Y(n11130) );
  MUX2X1 U11328 ( .B(n11129), .A(n11114), .S(n10529), .Y(n11774) );
  INVX2 U11329 ( .A(n11774), .Y(n92) );
  MUX2X1 U11330 ( .B(n7251), .A(n8781), .S(n10716), .Y(n11134) );
  MUX2X1 U11331 ( .B(n7353), .A(n8883), .S(n10716), .Y(n11133) );
  MUX2X1 U11332 ( .B(n7455), .A(n8985), .S(n10716), .Y(n11137) );
  MUX2X1 U11333 ( .B(n7557), .A(n9087), .S(n10716), .Y(n11136) );
  MUX2X1 U11334 ( .B(n11135), .A(n11132), .S(n10654), .Y(n11146) );
  MUX2X1 U11335 ( .B(n6945), .A(n8577), .S(n10716), .Y(n11140) );
  MUX2X1 U11336 ( .B(n6741), .A(n8475), .S(n10716), .Y(n11139) );
  MUX2X1 U11337 ( .B(n6843), .A(n8373), .S(n10716), .Y(n11143) );
  MUX2X1 U11338 ( .B(n7047), .A(n8679), .S(n10716), .Y(n11142) );
  MUX2X1 U11339 ( .B(n11141), .A(n11138), .S(n10654), .Y(n11145) );
  MUX2X1 U11340 ( .B(n7659), .A(n9189), .S(n10716), .Y(n11149) );
  MUX2X1 U11341 ( .B(n7761), .A(n9291), .S(n10716), .Y(n11148) );
  MUX2X1 U11342 ( .B(n7863), .A(n9393), .S(n10716), .Y(n11152) );
  MUX2X1 U11343 ( .B(n7965), .A(n9495), .S(n10716), .Y(n11151) );
  MUX2X1 U11344 ( .B(n11150), .A(n11147), .S(n10654), .Y(n11161) );
  MUX2X1 U11345 ( .B(n8067), .A(n9597), .S(n10716), .Y(n11155) );
  MUX2X1 U11346 ( .B(n8169), .A(n9699), .S(n10716), .Y(n11154) );
  MUX2X1 U11347 ( .B(n8271), .A(n9801), .S(n10716), .Y(n11158) );
  MUX2X1 U11348 ( .B(n7149), .A(n9903), .S(n10716), .Y(n11157) );
  MUX2X1 U11349 ( .B(n11156), .A(n11153), .S(n10654), .Y(n11160) );
  MUX2X1 U11350 ( .B(n11159), .A(n11144), .S(n10529), .Y(n11775) );
  INVX2 U11351 ( .A(n11775), .Y(n91) );
  MUX2X1 U11352 ( .B(n7254), .A(n8784), .S(n10715), .Y(n11164) );
  MUX2X1 U11353 ( .B(n7356), .A(n8886), .S(n10715), .Y(n11163) );
  MUX2X1 U11354 ( .B(n7458), .A(n8988), .S(n10715), .Y(n11167) );
  MUX2X1 U11355 ( .B(n7560), .A(n9090), .S(n10715), .Y(n11166) );
  MUX2X1 U11356 ( .B(n11165), .A(n11162), .S(n10653), .Y(n11176) );
  MUX2X1 U11357 ( .B(n6948), .A(n8580), .S(n10715), .Y(n11170) );
  MUX2X1 U11358 ( .B(n6744), .A(n8478), .S(n10715), .Y(n11169) );
  MUX2X1 U11359 ( .B(n6846), .A(n8376), .S(n10715), .Y(n11173) );
  MUX2X1 U11360 ( .B(n7050), .A(n8682), .S(n10715), .Y(n11172) );
  MUX2X1 U11361 ( .B(n11171), .A(n11168), .S(n10653), .Y(n11175) );
  MUX2X1 U11362 ( .B(n7662), .A(n9192), .S(n10715), .Y(n11179) );
  MUX2X1 U11363 ( .B(n7764), .A(n9294), .S(n10715), .Y(n11178) );
  MUX2X1 U11364 ( .B(n7866), .A(n9396), .S(n10715), .Y(n11182) );
  MUX2X1 U11365 ( .B(n7968), .A(n9498), .S(n10715), .Y(n11181) );
  MUX2X1 U11366 ( .B(n11180), .A(n11177), .S(n10653), .Y(n11191) );
  MUX2X1 U11367 ( .B(n8070), .A(n9600), .S(n10715), .Y(n11185) );
  MUX2X1 U11368 ( .B(n8172), .A(n9702), .S(n10715), .Y(n11184) );
  MUX2X1 U11369 ( .B(n8274), .A(n9804), .S(n10715), .Y(n11188) );
  MUX2X1 U11370 ( .B(n7152), .A(n9906), .S(n10715), .Y(n11187) );
  MUX2X1 U11371 ( .B(n11186), .A(n11183), .S(n10653), .Y(n11190) );
  MUX2X1 U11372 ( .B(n11189), .A(n11174), .S(n10529), .Y(n11776) );
  INVX2 U11373 ( .A(n11776), .Y(n90) );
  MUX2X1 U11374 ( .B(n7257), .A(n8787), .S(n10715), .Y(n11194) );
  MUX2X1 U11375 ( .B(n7359), .A(n8889), .S(n10714), .Y(n11193) );
  MUX2X1 U11376 ( .B(n7461), .A(n8991), .S(n10714), .Y(n11197) );
  MUX2X1 U11377 ( .B(n7563), .A(n9093), .S(n10714), .Y(n11196) );
  MUX2X1 U11378 ( .B(n11195), .A(n11192), .S(n10653), .Y(n11206) );
  MUX2X1 U11379 ( .B(n6951), .A(n8583), .S(n10714), .Y(n11200) );
  MUX2X1 U11380 ( .B(n6747), .A(n8481), .S(n10714), .Y(n11199) );
  MUX2X1 U11381 ( .B(n6849), .A(n8379), .S(n10714), .Y(n11203) );
  MUX2X1 U11382 ( .B(n7053), .A(n8685), .S(n10714), .Y(n11202) );
  MUX2X1 U11383 ( .B(n11201), .A(n11198), .S(n10653), .Y(n11205) );
  MUX2X1 U11384 ( .B(n7665), .A(n9195), .S(n10714), .Y(n11209) );
  MUX2X1 U11385 ( .B(n7767), .A(n9297), .S(n10714), .Y(n11208) );
  MUX2X1 U11386 ( .B(n7869), .A(n9399), .S(n10714), .Y(n11212) );
  MUX2X1 U11387 ( .B(n7971), .A(n9501), .S(n10714), .Y(n11211) );
  MUX2X1 U11388 ( .B(n11210), .A(n11207), .S(n10653), .Y(n11221) );
  MUX2X1 U11389 ( .B(n8073), .A(n9603), .S(n10714), .Y(n11215) );
  MUX2X1 U11390 ( .B(n8175), .A(n9705), .S(n10714), .Y(n11214) );
  MUX2X1 U11391 ( .B(n8277), .A(n9807), .S(n10714), .Y(n11218) );
  MUX2X1 U11392 ( .B(n7155), .A(n9909), .S(n10714), .Y(n11217) );
  MUX2X1 U11393 ( .B(n11216), .A(n11213), .S(n10653), .Y(n11220) );
  MUX2X1 U11394 ( .B(n11219), .A(n11204), .S(n10529), .Y(n11777) );
  INVX2 U11395 ( .A(n11777), .Y(n89) );
  MUX2X1 U11396 ( .B(n7260), .A(n8790), .S(n10714), .Y(n11224) );
  MUX2X1 U11397 ( .B(n7362), .A(n8892), .S(n10714), .Y(n11223) );
  MUX2X1 U11398 ( .B(n7464), .A(n8994), .S(n10713), .Y(n11227) );
  MUX2X1 U11399 ( .B(n7566), .A(n9096), .S(n10713), .Y(n11226) );
  MUX2X1 U11400 ( .B(n11225), .A(n11222), .S(n10653), .Y(n11236) );
  MUX2X1 U11401 ( .B(n6954), .A(n8586), .S(n10713), .Y(n11230) );
  MUX2X1 U11402 ( .B(n6750), .A(n8484), .S(n10713), .Y(n11229) );
  MUX2X1 U11403 ( .B(n6852), .A(n8382), .S(n10713), .Y(n11233) );
  MUX2X1 U11404 ( .B(n7056), .A(n8688), .S(n10713), .Y(n11232) );
  MUX2X1 U11405 ( .B(n11231), .A(n11228), .S(n10653), .Y(n11235) );
  MUX2X1 U11406 ( .B(n7668), .A(n9198), .S(n10713), .Y(n11239) );
  MUX2X1 U11407 ( .B(n7770), .A(n9300), .S(n10713), .Y(n11238) );
  MUX2X1 U11408 ( .B(n7872), .A(n9402), .S(n10713), .Y(n11242) );
  MUX2X1 U11409 ( .B(n7974), .A(n9504), .S(n10713), .Y(n11241) );
  MUX2X1 U11410 ( .B(n11240), .A(n11237), .S(n10653), .Y(n11251) );
  MUX2X1 U11411 ( .B(n8076), .A(n9606), .S(n10713), .Y(n11245) );
  MUX2X1 U11412 ( .B(n8178), .A(n9708), .S(n10713), .Y(n11244) );
  MUX2X1 U11413 ( .B(n8280), .A(n9810), .S(n10713), .Y(n11248) );
  MUX2X1 U11414 ( .B(n7158), .A(n9912), .S(n10713), .Y(n11247) );
  MUX2X1 U11415 ( .B(n11246), .A(n11243), .S(n10653), .Y(n11250) );
  MUX2X1 U11416 ( .B(n11249), .A(n11234), .S(n10529), .Y(n11778) );
  INVX2 U11417 ( .A(n11778), .Y(n88) );
  MUX2X1 U11418 ( .B(n7263), .A(n8793), .S(n10717), .Y(n11254) );
  MUX2X1 U11419 ( .B(n7365), .A(n8895), .S(n10697), .Y(n11253) );
  MUX2X1 U11420 ( .B(n7467), .A(n8997), .S(n10697), .Y(n11257) );
  MUX2X1 U11421 ( .B(n7569), .A(n9099), .S(n10697), .Y(n11256) );
  MUX2X1 U11422 ( .B(n11255), .A(n11252), .S(n10653), .Y(n11266) );
  MUX2X1 U11423 ( .B(n6957), .A(n8589), .S(n10696), .Y(n11260) );
  MUX2X1 U11424 ( .B(n6753), .A(n8487), .S(n10696), .Y(n11259) );
  MUX2X1 U11425 ( .B(n6855), .A(n8385), .S(n10696), .Y(n11263) );
  MUX2X1 U11426 ( .B(n7059), .A(n8691), .S(n10696), .Y(n11262) );
  MUX2X1 U11427 ( .B(n11261), .A(n11258), .S(n10653), .Y(n11265) );
  MUX2X1 U11428 ( .B(n7671), .A(n9201), .S(n10696), .Y(n11269) );
  MUX2X1 U11429 ( .B(n7773), .A(n9303), .S(n10696), .Y(n11268) );
  MUX2X1 U11430 ( .B(n7875), .A(n9405), .S(n10696), .Y(n11272) );
  MUX2X1 U11431 ( .B(n7977), .A(n9507), .S(n10696), .Y(n11271) );
  MUX2X1 U11432 ( .B(n11270), .A(n11267), .S(n10653), .Y(n11281) );
  MUX2X1 U11433 ( .B(n8079), .A(n9609), .S(n10696), .Y(n11275) );
  MUX2X1 U11434 ( .B(n8181), .A(n9711), .S(n10696), .Y(n11274) );
  MUX2X1 U11435 ( .B(n8283), .A(n9813), .S(n10696), .Y(n11278) );
  MUX2X1 U11436 ( .B(n7161), .A(n9915), .S(n10696), .Y(n11277) );
  MUX2X1 U11437 ( .B(n11276), .A(n11273), .S(n10653), .Y(n11280) );
  MUX2X1 U11438 ( .B(n11279), .A(n11264), .S(n10529), .Y(n11779) );
  INVX2 U11439 ( .A(n11779), .Y(n87) );
  MUX2X1 U11440 ( .B(n7266), .A(n8796), .S(n10696), .Y(n11284) );
  MUX2X1 U11441 ( .B(n7368), .A(n8898), .S(n10696), .Y(n11283) );
  MUX2X1 U11442 ( .B(n7470), .A(n9000), .S(n10696), .Y(n11287) );
  MUX2X1 U11443 ( .B(n7572), .A(n9102), .S(n10696), .Y(n11286) );
  MUX2X1 U11444 ( .B(n11285), .A(n11282), .S(n10652), .Y(n11296) );
  MUX2X1 U11445 ( .B(n6960), .A(n8592), .S(n10696), .Y(n11290) );
  MUX2X1 U11446 ( .B(n6756), .A(n8490), .S(n10695), .Y(n11289) );
  MUX2X1 U11447 ( .B(n6858), .A(n8388), .S(n10695), .Y(n11293) );
  MUX2X1 U11448 ( .B(n7062), .A(n8694), .S(n10695), .Y(n11292) );
  MUX2X1 U11449 ( .B(n11291), .A(n11288), .S(n10652), .Y(n11295) );
  MUX2X1 U11450 ( .B(n7674), .A(n9204), .S(n10695), .Y(n11299) );
  MUX2X1 U11451 ( .B(n7776), .A(n9306), .S(n10695), .Y(n11298) );
  MUX2X1 U11452 ( .B(n7878), .A(n9408), .S(n10695), .Y(n11302) );
  MUX2X1 U11453 ( .B(n7980), .A(n9510), .S(n10695), .Y(n11301) );
  MUX2X1 U11454 ( .B(n11300), .A(n11297), .S(n10652), .Y(n11311) );
  MUX2X1 U11455 ( .B(n8082), .A(n9612), .S(n10695), .Y(n11305) );
  MUX2X1 U11456 ( .B(n8184), .A(n9714), .S(n10695), .Y(n11304) );
  MUX2X1 U11457 ( .B(n8286), .A(n9816), .S(n10695), .Y(n11308) );
  MUX2X1 U11458 ( .B(n7164), .A(n9918), .S(n10695), .Y(n11307) );
  MUX2X1 U11459 ( .B(n11306), .A(n11303), .S(n10652), .Y(n11310) );
  MUX2X1 U11460 ( .B(n11309), .A(n11294), .S(n10529), .Y(n11780) );
  INVX2 U11461 ( .A(n11780), .Y(n86) );
  MUX2X1 U11462 ( .B(n7269), .A(n8799), .S(n10695), .Y(n11314) );
  MUX2X1 U11463 ( .B(n7371), .A(n8901), .S(n10695), .Y(n11313) );
  MUX2X1 U11464 ( .B(n7473), .A(n9003), .S(n10695), .Y(n11317) );
  MUX2X1 U11465 ( .B(n7575), .A(n9105), .S(n10695), .Y(n11316) );
  MUX2X1 U11466 ( .B(n11315), .A(n11312), .S(n10652), .Y(n11326) );
  MUX2X1 U11467 ( .B(n6963), .A(n8595), .S(n10695), .Y(n11320) );
  MUX2X1 U11468 ( .B(n6759), .A(n8493), .S(n10695), .Y(n11319) );
  MUX2X1 U11469 ( .B(n6861), .A(n8391), .S(n10694), .Y(n11323) );
  MUX2X1 U11470 ( .B(n7065), .A(n8697), .S(n10694), .Y(n11322) );
  MUX2X1 U11471 ( .B(n11321), .A(n11318), .S(n10652), .Y(n11325) );
  MUX2X1 U11472 ( .B(n7677), .A(n9207), .S(n10694), .Y(n11329) );
  MUX2X1 U11473 ( .B(n7779), .A(n9309), .S(n10694), .Y(n11328) );
  MUX2X1 U11474 ( .B(n7881), .A(n9411), .S(n10694), .Y(n11332) );
  MUX2X1 U11475 ( .B(n7983), .A(n9513), .S(n10694), .Y(n11331) );
  MUX2X1 U11476 ( .B(n11330), .A(n11327), .S(n10652), .Y(n11341) );
  MUX2X1 U11477 ( .B(n8085), .A(n9615), .S(n10694), .Y(n11335) );
  MUX2X1 U11478 ( .B(n8187), .A(n9717), .S(n10694), .Y(n11334) );
  MUX2X1 U11479 ( .B(n8289), .A(n9819), .S(n10694), .Y(n11338) );
  MUX2X1 U11480 ( .B(n7167), .A(n9921), .S(n10694), .Y(n11337) );
  MUX2X1 U11481 ( .B(n11336), .A(n11333), .S(n10652), .Y(n11340) );
  MUX2X1 U11482 ( .B(n11339), .A(n11324), .S(n10529), .Y(n11781) );
  INVX2 U11483 ( .A(n11781), .Y(n85) );
  MUX2X1 U11484 ( .B(n7272), .A(n8802), .S(n10694), .Y(n11344) );
  MUX2X1 U11485 ( .B(n7374), .A(n8904), .S(n10694), .Y(n11343) );
  MUX2X1 U11486 ( .B(n7476), .A(n9006), .S(n10694), .Y(n11347) );
  MUX2X1 U11487 ( .B(n7578), .A(n9108), .S(n10694), .Y(n11346) );
  MUX2X1 U11488 ( .B(n11345), .A(n11342), .S(n10652), .Y(n11356) );
  MUX2X1 U11489 ( .B(n6966), .A(n8598), .S(n10694), .Y(n11350) );
  MUX2X1 U11490 ( .B(n6762), .A(n8496), .S(n10694), .Y(n11349) );
  MUX2X1 U11491 ( .B(n6864), .A(n8394), .S(n10694), .Y(n11353) );
  MUX2X1 U11492 ( .B(n7068), .A(n8700), .S(n10693), .Y(n11352) );
  MUX2X1 U11493 ( .B(n11351), .A(n11348), .S(n10652), .Y(n11355) );
  MUX2X1 U11494 ( .B(n7680), .A(n9210), .S(n10693), .Y(n11359) );
  MUX2X1 U11495 ( .B(n7782), .A(n9312), .S(n10693), .Y(n11358) );
  MUX2X1 U11496 ( .B(n7884), .A(n9414), .S(n10693), .Y(n11362) );
  MUX2X1 U11497 ( .B(n7986), .A(n9516), .S(n10693), .Y(n11361) );
  MUX2X1 U11498 ( .B(n11360), .A(n11357), .S(n10652), .Y(n11371) );
  MUX2X1 U11499 ( .B(n8088), .A(n9618), .S(n10693), .Y(n11365) );
  MUX2X1 U11500 ( .B(n8190), .A(n9720), .S(n10693), .Y(n11364) );
  MUX2X1 U11501 ( .B(n8292), .A(n9822), .S(n10693), .Y(n11368) );
  MUX2X1 U11502 ( .B(n7170), .A(n9924), .S(n10693), .Y(n11367) );
  MUX2X1 U11503 ( .B(n11366), .A(n11363), .S(n10652), .Y(n11370) );
  MUX2X1 U11504 ( .B(n11369), .A(n11354), .S(n10529), .Y(n11782) );
  INVX2 U11505 ( .A(n11782), .Y(n84) );
  MUX2X1 U11506 ( .B(n7275), .A(n8805), .S(n10693), .Y(n11374) );
  MUX2X1 U11507 ( .B(n7377), .A(n8907), .S(n10693), .Y(n11373) );
  MUX2X1 U11508 ( .B(n7479), .A(n9009), .S(n10693), .Y(n11377) );
  MUX2X1 U11509 ( .B(n7581), .A(n9111), .S(n10693), .Y(n11376) );
  MUX2X1 U11510 ( .B(n11375), .A(n11372), .S(n10652), .Y(n11386) );
  MUX2X1 U11511 ( .B(n6969), .A(n8601), .S(n10693), .Y(n11380) );
  MUX2X1 U11512 ( .B(n6765), .A(n8499), .S(n10693), .Y(n11379) );
  MUX2X1 U11513 ( .B(n6867), .A(n8397), .S(n10693), .Y(n11383) );
  MUX2X1 U11514 ( .B(n7071), .A(n8703), .S(n10692), .Y(n11382) );
  MUX2X1 U11515 ( .B(n11381), .A(n11378), .S(n10652), .Y(n11385) );
  MUX2X1 U11516 ( .B(n7683), .A(n9213), .S(n10692), .Y(n11389) );
  MUX2X1 U11517 ( .B(n7785), .A(n9315), .S(n10692), .Y(n11388) );
  MUX2X1 U11518 ( .B(n7887), .A(n9417), .S(n10692), .Y(n11392) );
  MUX2X1 U11519 ( .B(n7989), .A(n9519), .S(n10692), .Y(n11391) );
  MUX2X1 U11520 ( .B(n11390), .A(n11387), .S(n10652), .Y(n11401) );
  MUX2X1 U11521 ( .B(n8091), .A(n9621), .S(n10692), .Y(n11395) );
  MUX2X1 U11522 ( .B(n8193), .A(n9723), .S(n10692), .Y(n11394) );
  MUX2X1 U11523 ( .B(n8295), .A(n9825), .S(n10692), .Y(n11398) );
  MUX2X1 U11524 ( .B(n7173), .A(n9927), .S(n10692), .Y(n11397) );
  MUX2X1 U11525 ( .B(n11396), .A(n11393), .S(n10652), .Y(n11400) );
  MUX2X1 U11526 ( .B(n11399), .A(n11384), .S(n10529), .Y(n11783) );
  INVX2 U11527 ( .A(n11783), .Y(n83) );
  MUX2X1 U11528 ( .B(n7278), .A(n8808), .S(n10692), .Y(n11404) );
  MUX2X1 U11529 ( .B(n7380), .A(n8910), .S(n10692), .Y(n11403) );
  MUX2X1 U11530 ( .B(n7482), .A(n9012), .S(n10692), .Y(n11407) );
  MUX2X1 U11531 ( .B(n7584), .A(n9114), .S(n10692), .Y(n11406) );
  MUX2X1 U11532 ( .B(n11405), .A(n11402), .S(n10652), .Y(n11416) );
  MUX2X1 U11533 ( .B(n6972), .A(n8604), .S(n10692), .Y(n11410) );
  MUX2X1 U11534 ( .B(n6768), .A(n8502), .S(n10692), .Y(n11409) );
  MUX2X1 U11535 ( .B(n6870), .A(n8400), .S(n10692), .Y(n11413) );
  MUX2X1 U11536 ( .B(n7074), .A(n8706), .S(n10692), .Y(n11412) );
  MUX2X1 U11537 ( .B(n11411), .A(n11408), .S(n10651), .Y(n11415) );
  MUX2X1 U11538 ( .B(n7686), .A(n9216), .S(n10691), .Y(n11419) );
  MUX2X1 U11539 ( .B(n7788), .A(n9318), .S(n10691), .Y(n11418) );
  MUX2X1 U11540 ( .B(n7890), .A(n9420), .S(n10691), .Y(n11422) );
  MUX2X1 U11541 ( .B(n7992), .A(n9522), .S(n10691), .Y(n11421) );
  MUX2X1 U11542 ( .B(n11420), .A(n11417), .S(n10651), .Y(n11431) );
  MUX2X1 U11543 ( .B(n8094), .A(n9624), .S(n10691), .Y(n11425) );
  MUX2X1 U11544 ( .B(n8196), .A(n9726), .S(n10691), .Y(n11424) );
  MUX2X1 U11545 ( .B(n8298), .A(n9828), .S(n10691), .Y(n11428) );
  MUX2X1 U11546 ( .B(n7176), .A(n9930), .S(n10691), .Y(n11427) );
  MUX2X1 U11547 ( .B(n11426), .A(n11423), .S(n10651), .Y(n11430) );
  MUX2X1 U11548 ( .B(n11429), .A(n11414), .S(n10529), .Y(n11784) );
  INVX2 U11549 ( .A(n11784), .Y(n82) );
  MUX2X1 U11550 ( .B(n7281), .A(n8811), .S(n10691), .Y(n11434) );
  MUX2X1 U11551 ( .B(n7383), .A(n8913), .S(n10691), .Y(n11433) );
  MUX2X1 U11552 ( .B(n7485), .A(n9015), .S(n10691), .Y(n11437) );
  MUX2X1 U11553 ( .B(n7587), .A(n9117), .S(n10691), .Y(n11436) );
  MUX2X1 U11554 ( .B(n11435), .A(n11432), .S(n10651), .Y(n11446) );
  MUX2X1 U11555 ( .B(n6975), .A(n8607), .S(n10691), .Y(n11440) );
  MUX2X1 U11556 ( .B(n6771), .A(n8505), .S(n10691), .Y(n11439) );
  MUX2X1 U11557 ( .B(n6873), .A(n8403), .S(n10691), .Y(n11443) );
  MUX2X1 U11558 ( .B(n7077), .A(n8709), .S(n10691), .Y(n11442) );
  MUX2X1 U11559 ( .B(n11441), .A(n11438), .S(n10651), .Y(n11445) );
  MUX2X1 U11560 ( .B(n7689), .A(n9219), .S(n10691), .Y(n11449) );
  MUX2X1 U11561 ( .B(n7791), .A(n9321), .S(n10690), .Y(n11448) );
  MUX2X1 U11562 ( .B(n7893), .A(n9423), .S(n10690), .Y(n11452) );
  MUX2X1 U11563 ( .B(n7995), .A(n9525), .S(n10690), .Y(n11451) );
  MUX2X1 U11564 ( .B(n11450), .A(n11447), .S(n10651), .Y(n11461) );
  MUX2X1 U11565 ( .B(n8097), .A(n9627), .S(n10690), .Y(n11455) );
  MUX2X1 U11566 ( .B(n8199), .A(n9729), .S(n10690), .Y(n11454) );
  MUX2X1 U11567 ( .B(n8301), .A(n9831), .S(n10690), .Y(n11458) );
  MUX2X1 U11568 ( .B(n7179), .A(n9933), .S(n10690), .Y(n11457) );
  MUX2X1 U11569 ( .B(n11456), .A(n11453), .S(n10651), .Y(n11460) );
  MUX2X1 U11570 ( .B(n11459), .A(n11444), .S(n10529), .Y(n11785) );
  INVX2 U11571 ( .A(n11785), .Y(n81) );
  MUX2X1 U11572 ( .B(n7284), .A(n8814), .S(n10690), .Y(n11464) );
  MUX2X1 U11573 ( .B(n7386), .A(n8916), .S(n10690), .Y(n11463) );
  MUX2X1 U11574 ( .B(n7488), .A(n9018), .S(n10690), .Y(n11467) );
  MUX2X1 U11575 ( .B(n7590), .A(n9120), .S(n10690), .Y(n11466) );
  MUX2X1 U11576 ( .B(n11465), .A(n11462), .S(n10651), .Y(n11476) );
  MUX2X1 U11577 ( .B(n6978), .A(n8610), .S(n10690), .Y(n11470) );
  MUX2X1 U11578 ( .B(n6774), .A(n8508), .S(n10690), .Y(n11469) );
  MUX2X1 U11579 ( .B(n6876), .A(n8406), .S(n10690), .Y(n11473) );
  MUX2X1 U11580 ( .B(n7080), .A(n8712), .S(n10690), .Y(n11472) );
  MUX2X1 U11581 ( .B(n11471), .A(n11468), .S(n10651), .Y(n11475) );
  MUX2X1 U11582 ( .B(n7692), .A(n9222), .S(n10690), .Y(n11479) );
  MUX2X1 U11583 ( .B(n7794), .A(n9324), .S(n10690), .Y(n11478) );
  MUX2X1 U11584 ( .B(n7896), .A(n9426), .S(n10689), .Y(n11482) );
  MUX2X1 U11585 ( .B(n7998), .A(n9528), .S(n10689), .Y(n11481) );
  MUX2X1 U11586 ( .B(n11480), .A(n11477), .S(n10651), .Y(n11491) );
  MUX2X1 U11587 ( .B(n8100), .A(n9630), .S(n10689), .Y(n11485) );
  MUX2X1 U11588 ( .B(n8202), .A(n9732), .S(n10689), .Y(n11484) );
  MUX2X1 U11589 ( .B(n8304), .A(n9834), .S(n10689), .Y(n11488) );
  MUX2X1 U11590 ( .B(n7182), .A(n9936), .S(n10689), .Y(n11487) );
  MUX2X1 U11591 ( .B(n11486), .A(n11483), .S(n10651), .Y(n11490) );
  MUX2X1 U11592 ( .B(n11489), .A(n11474), .S(n10529), .Y(n11786) );
  INVX2 U11593 ( .A(n11786), .Y(n80) );
  MUX2X1 U11594 ( .B(n7287), .A(n8817), .S(n10689), .Y(n11494) );
  MUX2X1 U11595 ( .B(n7389), .A(n8919), .S(n10689), .Y(n11493) );
  MUX2X1 U11596 ( .B(n7491), .A(n9021), .S(n10689), .Y(n11497) );
  MUX2X1 U11597 ( .B(n7593), .A(n9123), .S(n10689), .Y(n11496) );
  MUX2X1 U11598 ( .B(n11495), .A(n11492), .S(n10651), .Y(n11506) );
  MUX2X1 U11599 ( .B(n6981), .A(n8613), .S(n10689), .Y(n11500) );
  MUX2X1 U11600 ( .B(n6777), .A(n8511), .S(n10689), .Y(n11499) );
  MUX2X1 U11601 ( .B(n6879), .A(n8409), .S(n10689), .Y(n11503) );
  MUX2X1 U11602 ( .B(n7083), .A(n8715), .S(n10693), .Y(n11502) );
  MUX2X1 U11603 ( .B(n11501), .A(n11498), .S(n10651), .Y(n11505) );
  MUX2X1 U11604 ( .B(n7695), .A(n9225), .S(n10705), .Y(n11509) );
  MUX2X1 U11605 ( .B(n7797), .A(n9327), .S(n10705), .Y(n11508) );
  MUX2X1 U11606 ( .B(n7899), .A(n9429), .S(n10705), .Y(n11512) );
  MUX2X1 U11607 ( .B(n8001), .A(n9531), .S(n10704), .Y(n11511) );
  MUX2X1 U11608 ( .B(n11510), .A(n11507), .S(n10651), .Y(n11521) );
  MUX2X1 U11609 ( .B(n8103), .A(n9633), .S(n10704), .Y(n11515) );
  MUX2X1 U11610 ( .B(n8205), .A(n9735), .S(n10704), .Y(n11514) );
  MUX2X1 U11611 ( .B(n8307), .A(n9837), .S(n10704), .Y(n11518) );
  MUX2X1 U11612 ( .B(n7185), .A(n9939), .S(n10704), .Y(n11517) );
  MUX2X1 U11613 ( .B(n11516), .A(n11513), .S(n10651), .Y(n11520) );
  MUX2X1 U11614 ( .B(n11519), .A(n11504), .S(n10529), .Y(n11787) );
  INVX2 U11615 ( .A(n11787), .Y(n79) );
  MUX2X1 U11616 ( .B(n7290), .A(n8820), .S(n10704), .Y(n11524) );
  MUX2X1 U11617 ( .B(n7392), .A(n8922), .S(n10704), .Y(n11523) );
  MUX2X1 U11618 ( .B(n7494), .A(n9024), .S(n10704), .Y(n11527) );
  MUX2X1 U11619 ( .B(n7596), .A(n9126), .S(n10704), .Y(n11526) );
  MUX2X1 U11620 ( .B(n11525), .A(n11522), .S(n10651), .Y(n11536) );
  MUX2X1 U11621 ( .B(n6984), .A(n8616), .S(n10704), .Y(n11530) );
  MUX2X1 U11622 ( .B(n6780), .A(n8514), .S(n10704), .Y(n11529) );
  MUX2X1 U11623 ( .B(n6882), .A(n8412), .S(n10704), .Y(n11533) );
  MUX2X1 U11624 ( .B(n7086), .A(n8718), .S(n10704), .Y(n11532) );
  MUX2X1 U11625 ( .B(n11531), .A(n11528), .S(n10653), .Y(n11535) );
  MUX2X1 U11626 ( .B(n7698), .A(n9228), .S(n10704), .Y(n11539) );
  MUX2X1 U11627 ( .B(n7800), .A(n9330), .S(n10704), .Y(n11538) );
  MUX2X1 U11628 ( .B(n7902), .A(n9432), .S(n10704), .Y(n11542) );
  MUX2X1 U11629 ( .B(n8004), .A(n9534), .S(n10704), .Y(n11541) );
  MUX2X1 U11630 ( .B(n11540), .A(n11537), .S(n10651), .Y(n11551) );
  MUX2X1 U11631 ( .B(n8106), .A(n9636), .S(n10703), .Y(n11545) );
  MUX2X1 U11632 ( .B(n8208), .A(n9738), .S(n10703), .Y(n11544) );
  MUX2X1 U11633 ( .B(n8310), .A(n9840), .S(n10703), .Y(n11548) );
  MUX2X1 U11634 ( .B(n7188), .A(n9942), .S(n10703), .Y(n11547) );
  MUX2X1 U11635 ( .B(n11546), .A(n11543), .S(n10650), .Y(n11550) );
  MUX2X1 U11636 ( .B(n11549), .A(n11534), .S(n10529), .Y(n11788) );
  INVX2 U11637 ( .A(n11788), .Y(n78) );
  MUX2X1 U11638 ( .B(n7293), .A(n8823), .S(n10703), .Y(n11554) );
  MUX2X1 U11639 ( .B(n7395), .A(n8925), .S(n10703), .Y(n11553) );
  MUX2X1 U11640 ( .B(n7497), .A(n9027), .S(n10703), .Y(n11557) );
  MUX2X1 U11641 ( .B(n7599), .A(n9129), .S(n10703), .Y(n11556) );
  MUX2X1 U11642 ( .B(n11555), .A(n11552), .S(n10650), .Y(n11566) );
  MUX2X1 U11643 ( .B(n6987), .A(n8619), .S(n10703), .Y(n11560) );
  MUX2X1 U11644 ( .B(n6783), .A(n8517), .S(n10703), .Y(n11559) );
  MUX2X1 U11645 ( .B(n6885), .A(n8415), .S(n10703), .Y(n11563) );
  MUX2X1 U11646 ( .B(n7089), .A(n8721), .S(n10703), .Y(n11562) );
  MUX2X1 U11647 ( .B(n11561), .A(n11558), .S(n10650), .Y(n11565) );
  MUX2X1 U11648 ( .B(n7701), .A(n9231), .S(n10703), .Y(n11569) );
  MUX2X1 U11649 ( .B(n7803), .A(n9333), .S(n10703), .Y(n11568) );
  MUX2X1 U11650 ( .B(n7905), .A(n9435), .S(n10703), .Y(n11572) );
  MUX2X1 U11651 ( .B(n8007), .A(n9537), .S(n10703), .Y(n11571) );
  MUX2X1 U11652 ( .B(n11570), .A(n11567), .S(n10650), .Y(n11581) );
  MUX2X1 U11653 ( .B(n8109), .A(n9639), .S(n10703), .Y(n11575) );
  MUX2X1 U11654 ( .B(n8211), .A(n9741), .S(n10702), .Y(n11574) );
  MUX2X1 U11655 ( .B(n8313), .A(n9843), .S(n10702), .Y(n11578) );
  MUX2X1 U11656 ( .B(n7191), .A(n9945), .S(n10702), .Y(n11577) );
  MUX2X1 U11657 ( .B(n11576), .A(n11573), .S(n10650), .Y(n11580) );
  MUX2X1 U11658 ( .B(n11579), .A(n11564), .S(n10529), .Y(n11789) );
  INVX2 U11659 ( .A(n11789), .Y(n77) );
  MUX2X1 U11660 ( .B(n7296), .A(n8826), .S(n10702), .Y(n11584) );
  MUX2X1 U11661 ( .B(n7398), .A(n8928), .S(n10702), .Y(n11583) );
  MUX2X1 U11662 ( .B(n7500), .A(n9030), .S(n10702), .Y(n11587) );
  MUX2X1 U11663 ( .B(n7602), .A(n9132), .S(n10702), .Y(n11586) );
  MUX2X1 U11664 ( .B(n11585), .A(n11582), .S(n10650), .Y(n11596) );
  MUX2X1 U11665 ( .B(n6990), .A(n8622), .S(n10702), .Y(n11590) );
  MUX2X1 U11666 ( .B(n6786), .A(n8520), .S(n10702), .Y(n11589) );
  MUX2X1 U11667 ( .B(n6888), .A(n8418), .S(n10702), .Y(n11593) );
  MUX2X1 U11668 ( .B(n7092), .A(n8724), .S(n10702), .Y(n11592) );
  MUX2X1 U11669 ( .B(n11591), .A(n11588), .S(n10650), .Y(n11595) );
  MUX2X1 U11670 ( .B(n7704), .A(n9234), .S(n10702), .Y(n11599) );
  MUX2X1 U11671 ( .B(n7806), .A(n9336), .S(n10702), .Y(n11598) );
  MUX2X1 U11672 ( .B(n7908), .A(n9438), .S(n10702), .Y(n11602) );
  MUX2X1 U11673 ( .B(n8010), .A(n9540), .S(n10702), .Y(n11601) );
  MUX2X1 U11674 ( .B(n11600), .A(n11597), .S(n10650), .Y(n11611) );
  MUX2X1 U11675 ( .B(n8112), .A(n9642), .S(n10702), .Y(n11605) );
  MUX2X1 U11676 ( .B(n8214), .A(n9744), .S(n10702), .Y(n11604) );
  MUX2X1 U11677 ( .B(n8316), .A(n9846), .S(n10701), .Y(n11608) );
  MUX2X1 U11678 ( .B(n7194), .A(n9948), .S(n10701), .Y(n11607) );
  MUX2X1 U11679 ( .B(n11606), .A(n11603), .S(n10650), .Y(n11610) );
  MUX2X1 U11680 ( .B(n11609), .A(n11594), .S(n10529), .Y(n11790) );
  INVX2 U11681 ( .A(n11790), .Y(n76) );
  MUX2X1 U11682 ( .B(n7299), .A(n8829), .S(n10701), .Y(n11614) );
  MUX2X1 U11683 ( .B(n7401), .A(n8931), .S(n10701), .Y(n11613) );
  MUX2X1 U11684 ( .B(n7503), .A(n9033), .S(n10701), .Y(n11617) );
  MUX2X1 U11685 ( .B(n7605), .A(n9135), .S(n10701), .Y(n11616) );
  MUX2X1 U11686 ( .B(n11615), .A(n11612), .S(n10650), .Y(n11626) );
  MUX2X1 U11687 ( .B(n6993), .A(n8625), .S(n10701), .Y(n11620) );
  MUX2X1 U11688 ( .B(n6789), .A(n8523), .S(n10701), .Y(n11619) );
  MUX2X1 U11689 ( .B(n6891), .A(n8421), .S(n10701), .Y(n11623) );
  MUX2X1 U11690 ( .B(n7095), .A(n8727), .S(n10701), .Y(n11622) );
  MUX2X1 U11691 ( .B(n11621), .A(n11618), .S(n10650), .Y(n11625) );
  MUX2X1 U11692 ( .B(n7707), .A(n9237), .S(n10701), .Y(n11629) );
  MUX2X1 U11693 ( .B(n7809), .A(n9339), .S(n10701), .Y(n11628) );
  MUX2X1 U11694 ( .B(n7911), .A(n9441), .S(n10701), .Y(n11632) );
  MUX2X1 U11695 ( .B(n8013), .A(n9543), .S(n10701), .Y(n11631) );
  MUX2X1 U11696 ( .B(n11630), .A(n11627), .S(n10650), .Y(n11641) );
  MUX2X1 U11697 ( .B(n8115), .A(n9645), .S(n10701), .Y(n11635) );
  MUX2X1 U11698 ( .B(n8217), .A(n9747), .S(n10701), .Y(n11634) );
  MUX2X1 U11699 ( .B(n8319), .A(n9849), .S(n10700), .Y(n11638) );
  MUX2X1 U11700 ( .B(n7197), .A(n9951), .S(n10700), .Y(n11637) );
  MUX2X1 U11701 ( .B(n11636), .A(n11633), .S(n10650), .Y(n11640) );
  MUX2X1 U11702 ( .B(n11639), .A(n11624), .S(n10529), .Y(n11791) );
  INVX2 U11703 ( .A(n11791), .Y(n75) );
  MUX2X1 U11704 ( .B(n7302), .A(n8832), .S(n10700), .Y(n11644) );
  MUX2X1 U11705 ( .B(n7404), .A(n8934), .S(n10700), .Y(n11643) );
  MUX2X1 U11706 ( .B(n7506), .A(n9036), .S(n10700), .Y(n11647) );
  MUX2X1 U11707 ( .B(n7608), .A(n9138), .S(n10700), .Y(n11646) );
  MUX2X1 U11708 ( .B(n11645), .A(n11642), .S(n10650), .Y(n11656) );
  MUX2X1 U11709 ( .B(n6996), .A(n8628), .S(n10700), .Y(n11650) );
  MUX2X1 U11710 ( .B(n6792), .A(n8526), .S(n10700), .Y(n11649) );
  MUX2X1 U11711 ( .B(n6894), .A(n8424), .S(n10700), .Y(n11653) );
  MUX2X1 U11712 ( .B(n7098), .A(n8730), .S(n10700), .Y(n11652) );
  MUX2X1 U11713 ( .B(n11651), .A(n11648), .S(n10650), .Y(n11655) );
  MUX2X1 U11714 ( .B(n7710), .A(n9240), .S(n10700), .Y(n11659) );
  MUX2X1 U11715 ( .B(n7812), .A(n9342), .S(n10700), .Y(n11658) );
  MUX2X1 U11716 ( .B(n7914), .A(n9444), .S(n10700), .Y(n11662) );
  MUX2X1 U11717 ( .B(n8016), .A(n9546), .S(n10700), .Y(n11661) );
  MUX2X1 U11718 ( .B(n11660), .A(n11657), .S(n10650), .Y(n11671) );
  MUX2X1 U11719 ( .B(n8118), .A(n9648), .S(n10700), .Y(n11665) );
  MUX2X1 U11720 ( .B(n8220), .A(n9750), .S(n10700), .Y(n11664) );
  MUX2X1 U11721 ( .B(n8322), .A(n9852), .S(n10700), .Y(n11668) );
  MUX2X1 U11722 ( .B(n7200), .A(n9954), .S(n10699), .Y(n11667) );
  MUX2X1 U11723 ( .B(n11666), .A(n11663), .S(n10650), .Y(n11670) );
  MUX2X1 U11724 ( .B(n11669), .A(n11654), .S(n10529), .Y(n11792) );
  INVX2 U11725 ( .A(n11792), .Y(n74) );
  MUX2X1 U11726 ( .B(n7305), .A(n8835), .S(n10699), .Y(n11674) );
  MUX2X1 U11727 ( .B(n7407), .A(n8937), .S(n10699), .Y(n11673) );
  MUX2X1 U11728 ( .B(n7509), .A(n9039), .S(n10699), .Y(n11677) );
  MUX2X1 U11729 ( .B(n7611), .A(n9141), .S(n10699), .Y(n11676) );
  MUX2X1 U11730 ( .B(n11675), .A(n11672), .S(n10649), .Y(n11686) );
  MUX2X1 U11731 ( .B(n6999), .A(n8631), .S(n10699), .Y(n11680) );
  MUX2X1 U11732 ( .B(n6795), .A(n8529), .S(n10699), .Y(n11679) );
  MUX2X1 U11733 ( .B(n6897), .A(n8427), .S(n10699), .Y(n11683) );
  MUX2X1 U11734 ( .B(n7101), .A(n8733), .S(n10699), .Y(n11682) );
  MUX2X1 U11735 ( .B(n11681), .A(n11678), .S(n10649), .Y(n11685) );
  MUX2X1 U11736 ( .B(n7713), .A(n9243), .S(n10699), .Y(n11689) );
  MUX2X1 U11737 ( .B(n7815), .A(n9345), .S(n10699), .Y(n11688) );
  MUX2X1 U11738 ( .B(n7917), .A(n9447), .S(n10699), .Y(n11692) );
  MUX2X1 U11739 ( .B(n8019), .A(n9549), .S(n10699), .Y(n11691) );
  MUX2X1 U11740 ( .B(n11690), .A(n11687), .S(n10649), .Y(n11701) );
  MUX2X1 U11741 ( .B(n8121), .A(n9651), .S(n10699), .Y(n11695) );
  MUX2X1 U11742 ( .B(n8223), .A(n9753), .S(n10699), .Y(n11694) );
  MUX2X1 U11743 ( .B(n8325), .A(n9855), .S(n10699), .Y(n11698) );
  MUX2X1 U11744 ( .B(n7203), .A(n9957), .S(n10699), .Y(n11697) );
  MUX2X1 U11745 ( .B(n11696), .A(n11693), .S(n10649), .Y(n11700) );
  MUX2X1 U11746 ( .B(n11699), .A(n11684), .S(n10529), .Y(n11793) );
  INVX2 U11747 ( .A(n11793), .Y(n73) );
  MUX2X1 U11748 ( .B(n7308), .A(n8838), .S(n10698), .Y(n11704) );
  MUX2X1 U11749 ( .B(n7410), .A(n8940), .S(n10698), .Y(n11703) );
  MUX2X1 U11750 ( .B(n7512), .A(n9042), .S(n10698), .Y(n11707) );
  MUX2X1 U11751 ( .B(n7614), .A(n9144), .S(n10698), .Y(n11706) );
  MUX2X1 U11752 ( .B(n11705), .A(n11702), .S(n10649), .Y(n11716) );
  MUX2X1 U11753 ( .B(n7002), .A(n8634), .S(n10698), .Y(n11710) );
  MUX2X1 U11754 ( .B(n6798), .A(n8532), .S(n10698), .Y(n11709) );
  MUX2X1 U11755 ( .B(n6900), .A(n8430), .S(n10698), .Y(n11713) );
  MUX2X1 U11756 ( .B(n7104), .A(n8736), .S(n10698), .Y(n11712) );
  MUX2X1 U11757 ( .B(n11711), .A(n11708), .S(n10649), .Y(n11715) );
  MUX2X1 U11758 ( .B(n7716), .A(n9246), .S(n10698), .Y(n11719) );
  MUX2X1 U11759 ( .B(n7818), .A(n9348), .S(n10698), .Y(n11718) );
  MUX2X1 U11760 ( .B(n7920), .A(n9450), .S(n10698), .Y(n11722) );
  MUX2X1 U11761 ( .B(n8022), .A(n9552), .S(n10698), .Y(n11721) );
  MUX2X1 U11762 ( .B(n11720), .A(n11717), .S(n10649), .Y(n11731) );
  MUX2X1 U11763 ( .B(n8124), .A(n9654), .S(n10698), .Y(n11725) );
  MUX2X1 U11764 ( .B(n8226), .A(n9756), .S(n10698), .Y(n11724) );
  MUX2X1 U11765 ( .B(n8328), .A(n9858), .S(n10698), .Y(n11728) );
  MUX2X1 U11766 ( .B(n7206), .A(n9960), .S(n10698), .Y(n11727) );
  MUX2X1 U11767 ( .B(n11726), .A(n11723), .S(n10649), .Y(n11730) );
  MUX2X1 U11768 ( .B(n11729), .A(n11714), .S(n10529), .Y(n11794) );
  INVX2 U11769 ( .A(n11794), .Y(n72) );
  MUX2X1 U11770 ( .B(n7311), .A(n8841), .S(n10698), .Y(n11734) );
  MUX2X1 U11771 ( .B(n7413), .A(n8943), .S(n10697), .Y(n11733) );
  MUX2X1 U11772 ( .B(n7515), .A(n9045), .S(n10697), .Y(n11737) );
  MUX2X1 U11773 ( .B(n7617), .A(n9147), .S(n10697), .Y(n11736) );
  MUX2X1 U11774 ( .B(n11735), .A(n11732), .S(n10649), .Y(n11746) );
  MUX2X1 U11775 ( .B(n7005), .A(n8637), .S(n10697), .Y(n11740) );
  MUX2X1 U11776 ( .B(n6801), .A(n8535), .S(n10697), .Y(n11739) );
  MUX2X1 U11777 ( .B(n6903), .A(n8433), .S(n10697), .Y(n11743) );
  MUX2X1 U11778 ( .B(n7107), .A(n8739), .S(n10697), .Y(n11742) );
  MUX2X1 U11779 ( .B(n11741), .A(n11738), .S(n10649), .Y(n11745) );
  MUX2X1 U11780 ( .B(n7719), .A(n9249), .S(n10697), .Y(n11749) );
  MUX2X1 U11781 ( .B(n7821), .A(n9351), .S(n10697), .Y(n11748) );
  MUX2X1 U11782 ( .B(n7923), .A(n9453), .S(n10697), .Y(n11752) );
  MUX2X1 U11783 ( .B(n8025), .A(n9555), .S(n10697), .Y(n11751) );
  MUX2X1 U11784 ( .B(n11750), .A(n11747), .S(n10649), .Y(n11761) );
  MUX2X1 U11785 ( .B(n8127), .A(n9657), .S(n10697), .Y(n11755) );
  MUX2X1 U11786 ( .B(n8229), .A(n9759), .S(n10697), .Y(n11754) );
  MUX2X1 U11787 ( .B(n8331), .A(n9861), .S(n10697), .Y(n11758) );
  MUX2X1 U11788 ( .B(n7209), .A(n9963), .S(n10701), .Y(n11757) );
  MUX2X1 U11789 ( .B(n11756), .A(n11753), .S(n10649), .Y(n11760) );
  MUX2X1 U11790 ( .B(n11759), .A(n11744), .S(n10529), .Y(n11795) );
  INVX2 U11791 ( .A(n11795), .Y(n71) );
  INVX1 U11792 ( .A(n3), .Y(r301_B_not_1_) );
  INVX1 U11793 ( .A(rd_ptr_bin_ss[2]), .Y(r301_B_not_2_) );
  INVX1 U11794 ( .A(n5), .Y(r301_B_not_3_) );
  INVX1 U11795 ( .A(n6), .Y(r301_B_not_4_) );
  INVX1 U11796 ( .A(n4), .Y(r301_B_not_5_) );
  XNOR2X1 U11797 ( .A(r301_B_not_0_), .B(n10101), .Y(fillcount[0]) );
  XOR2X1 U11798 ( .A(add_158_carry[5]), .B(n10081), .Y(n38) );
  XOR2X1 U11799 ( .A(add_176_carry[5]), .B(n10047), .Y(n110) );
endmodule


module FIFO_2clk_DATA_WIDTH42_FIFO_DEPTH32_PTR_WIDTH6 ( rclk, wclk, reset, we, 
        re, data_in, empty_bar, full_bar, data_out, fillcount );
  input [41:0] data_in;
  output [41:0] data_out;
  output [5:0] fillcount;
  input rclk, wclk, reset, we, re;
  output empty_bar, full_bar;
  wire   n10, n11, n12, n13, n14, n14681, n14682, n14683, n14684, n14685,
         n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693,
         n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701,
         n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709,
         n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717,
         n14718, n14719, n14720, n14721, n14722, n14723, rd_ptr_bin_5_, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, full_check_4_,
         full_check_3_, n34, n35, n36, n37, n38, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n114, n115,
         n116, n117, n118, n201, n202, n203, n204, n205, n207, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n3072, n3077, n3082, n3087,
         n3089, n3091, n3093, n3095, n3097, n3099, n3101, n3103, n3105, n3107,
         n3109, n3111, n3113, n3115, n3117, n3119, n3121, n3123, n3125, n3127,
         n3129, n3131, n3133, n3135, n3137, n3139, n3141, n3143, n3145, n3147,
         n3149, n3151, n3153, n3155, n3157, n3159, n3161, n3163, n3165, n3167,
         n3169, n3171, n3179, n3184, n3189, n3194, n3196, n3201, n3209, n3210,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, net80703, net80702, net80878,
         net82056, net82055, net82004, net84855, net84771, net80615, net89715,
         net82513, net82512, net82511, net82457, net82147, net82062, net82038,
         net84723, net91760, net91739, net91712, net91816, net92910, net92912,
         net93027, net94407, net94541, net94530, net94529, net94528, net94527,
         net94524, net94521, net94519, net94517, net94515, net94574, net95822,
         net95817, net95818, net95813, net94553, net94546, net84863, net82107,
         net98087, net98077, net84761, net94543, net94487, net91757, net91756,
         net82246, net82074, net82060, net80714, net91711, net82274, net91741,
         net91726, net84864, net84743, net84737, r301_B_not_0_, net94575,
         net92930, net91731, net91715, net91679, net91678, net89699, net84770,
         net84769, net84760, net82261, net82260, net82259, net82166, net82058,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n39, n40, n41, n42, n43, n44, n45, n46, n47, n49, n50, n51,
         n52, n55, n56, n57, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n113, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n206, n208, n268, n796,
         n1228, n1706, n1707, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
         n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
         n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
         n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
         n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
         n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
         n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
         n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433,
         n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443,
         n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
         n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
         n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
         n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
         n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
         n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
         n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
         n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
         n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
         n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
         n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
         n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
         n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
         n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
         n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
         n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
         n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
         n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
         n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
         n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
         n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
         n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
         n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
         n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893,
         n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
         n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
         n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
         n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
         n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
         n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
         n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
         n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
         n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
         n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
         n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
         n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
         n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
         n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
         n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
         n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
         n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
         n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
         n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
         n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
         n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
         n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
         n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
         n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
         n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
         n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
         n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
         n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
         n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
         n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
         n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
         n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,
         n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
         n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
         n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
         n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
         n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
         n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
         n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
         n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
         n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
         n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
         n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
         n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
         n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
         n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,
         n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
         n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,
         n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,
         n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
         n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
         n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
         n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
         n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
         n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
         n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
         n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,
         n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,
         n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
         n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,
         n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
         n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
         n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,
         n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,
         n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
         n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738,
         n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12821, n12822, n12823, n12824, n12825, n12827, n12828,
         n12830, n12831, n12833, n12834, n12836, n12837, n12839, n12840,
         n12842, n12843, n12845, n12846, n12848, n12849, n12851, n12852,
         n12854, n12855, n12857, n12858, n12860, n12861, n12863, n12864,
         n12866, n12867, n12869, n12870, n12872, n12873, n12875, n12876,
         n12878, n12879, n12881, n12882, n12884, n12885, n12887, n12888,
         n12890, n12891, n12893, n12894, n12896, n12897, n12899, n12900,
         n12902, n12903, n12905, n12906, n12908, n12909, n12911, n12912,
         n12914, n12915, n12917, n12918, n12920, n12921, n12923, n12924,
         n12926, n12927, n12929, n12930, n12932, n12933, n12935, n12936,
         n12938, n12939, n12941, n12942, n12944, n12945, n12947, n12948,
         n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956,
         n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964,
         n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972,
         n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980,
         n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988,
         n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996,
         n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004,
         n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012,
         n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020,
         n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028,
         n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036,
         n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044,
         n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052,
         n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060,
         n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068,
         n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076,
         n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084,
         n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092,
         n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100,
         n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108,
         n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116,
         n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124,
         n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132,
         n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140,
         n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148,
         n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156,
         n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164,
         n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172,
         n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180,
         n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188,
         n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196,
         n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204,
         n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212,
         n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220,
         n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228,
         n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236,
         n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244,
         n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252,
         n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260,
         n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268,
         n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276,
         n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284,
         n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292,
         n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300,
         n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308,
         n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316,
         n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324,
         n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332,
         n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340,
         n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348,
         n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356,
         n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364,
         n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372,
         n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380,
         n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388,
         n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396,
         n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404,
         n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412,
         n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420,
         n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428,
         n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436,
         n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444,
         n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452,
         n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460,
         n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468,
         n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476,
         n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484,
         n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492,
         n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500,
         n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508,
         n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516,
         n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524,
         n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532,
         n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540,
         n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548,
         n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556,
         n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564,
         n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572,
         n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580,
         n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588,
         n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596,
         n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604,
         n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612,
         n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620,
         n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628,
         n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636,
         n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644,
         n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652,
         n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660,
         n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668,
         n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676,
         n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684,
         n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692,
         n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700,
         n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708,
         n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716,
         n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724,
         n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732,
         n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740,
         n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748,
         n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756,
         n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764,
         n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772,
         n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780,
         n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788,
         n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796,
         n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804,
         n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812,
         n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820,
         n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828,
         n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836,
         n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844,
         n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852,
         n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860,
         n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868,
         n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876,
         n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884,
         n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892,
         n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900,
         n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908,
         n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916,
         n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924,
         n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932,
         n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940,
         n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948,
         n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956,
         n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964,
         n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972,
         n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980,
         n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988,
         n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996,
         n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004,
         n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012,
         n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020,
         n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028,
         n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036,
         n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044,
         n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052,
         n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060,
         n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068,
         n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076,
         n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084,
         n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092,
         n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100,
         n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108,
         n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116,
         n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124,
         n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132,
         n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140,
         n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148,
         n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156,
         n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164,
         n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172,
         n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180,
         n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188,
         n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196,
         n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204,
         n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212,
         n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220,
         n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228,
         n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236,
         n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244,
         n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252,
         n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260,
         n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268,
         n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276,
         n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284,
         n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292,
         n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300,
         n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308,
         n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316,
         n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324,
         n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332,
         n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340,
         n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348,
         n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356,
         n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364,
         n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372,
         n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380,
         n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388,
         n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396,
         n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404,
         n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412,
         n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420,
         n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428,
         n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436,
         n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444,
         n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452,
         n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460,
         n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468,
         n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476,
         n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484,
         n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492,
         n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500,
         n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508,
         n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516,
         n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524,
         n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532,
         n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540,
         n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548,
         n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556,
         n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564,
         n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572,
         n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580,
         n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588,
         n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596,
         n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604,
         n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612,
         n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620,
         n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628,
         n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636,
         n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644,
         n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652,
         n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660,
         n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668,
         n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676,
         n14677, n14678, n14679, n14680;
  wire   [5:0] wr_ptr_gray;
  wire   [5:0] wr_ptr_gray_ss;
  wire   [5:0] wr_ptr_gray_s;
  wire   [5:0] rd_ptr_gray;
  wire   [5:0] rd_ptr_gray_ss;
  wire   [5:0] rd_ptr_gray_s;
  wire   [5:0] wr_ptr_bin;
  wire   [1343:0] fifo;
  wire   [5:2] add_176_carry;
  wire   [5:2] add_158_carry;

  DFFSR rd_ptr_bin_reg_0_ ( .D(n3212), .CLK(rclk), .R(n13224), .S(1'b1), .Q(
        n10) );
  DFFSR rd_ptr_bin_reg_5_ ( .D(n3209), .CLK(rclk), .R(n13223), .S(1'b1), .Q(
        rd_ptr_bin_5_) );
  DFFSR rd_ptr_gray_reg_5_ ( .D(n12981), .CLK(rclk), .R(n13223), .S(1'b1), .Q(
        rd_ptr_gray[5]) );
  DFFSR rd_ptr_gray_s_reg_5_ ( .D(n187), .CLK(wclk), .R(n13223), .S(1'b1), .Q(
        rd_ptr_gray_s[5]) );
  DFFSR rd_ptr_gray_ss_reg_5_ ( .D(n184), .CLK(wclk), .R(n13223), .S(1'b1), 
        .Q(rd_ptr_gray_ss[5]) );
  DFFSR rd_ptr_gray_reg_4_ ( .D(n15), .CLK(rclk), .R(n13222), .S(1'b1), .Q(
        rd_ptr_gray[4]) );
  DFFSR rd_ptr_gray_s_reg_4_ ( .D(n181), .CLK(wclk), .R(n13222), .S(1'b1), .Q(
        rd_ptr_gray_s[4]) );
  DFFSR rd_ptr_gray_ss_reg_4_ ( .D(n178), .CLK(wclk), .R(n13222), .S(1'b1), 
        .Q(net95822) );
  DFFSR wr_ptr_bin_reg_5_ ( .D(n3201), .CLK(wclk), .R(n13221), .S(1'b1), .Q(
        wr_ptr_bin[5]) );
  DFFSR wr_ptr_gray_reg_5_ ( .D(n12994), .CLK(wclk), .R(n13221), .S(1'b1), .Q(
        wr_ptr_gray[5]) );
  DFFSR wr_ptr_gray_s_reg_5_ ( .D(n175), .CLK(rclk), .R(n13221), .S(1'b1), .Q(
        wr_ptr_gray_s[5]) );
  DFFSR wr_ptr_gray_ss_reg_5_ ( .D(n172), .CLK(rclk), .R(n13221), .S(1'b1), 
        .Q(wr_ptr_gray_ss[5]) );
  DFFSR wr_ptr_bin_reg_0_ ( .D(n3196), .CLK(wclk), .R(n13222), .S(1'b1), .Q(
        wr_ptr_bin[0]) );
  DFFSR wr_ptr_bin_reg_1_ ( .D(n3194), .CLK(wclk), .R(n13222), .S(1'b1), .Q(
        wr_ptr_bin[1]) );
  DFFSR wr_ptr_gray_reg_0_ ( .D(n24), .CLK(wclk), .R(n13222), .S(1'b1), .Q(
        wr_ptr_gray[0]) );
  DFFSR wr_ptr_gray_s_reg_0_ ( .D(n169), .CLK(rclk), .R(n13222), .S(1'b1), .Q(
        wr_ptr_gray_s[0]) );
  DFFSR wr_ptr_gray_ss_reg_0_ ( .D(n166), .CLK(rclk), .R(n13222), .S(1'b1), 
        .Q(wr_ptr_gray_ss[0]) );
  DFFSR wr_ptr_bin_reg_2_ ( .D(n3189), .CLK(wclk), .R(n13222), .S(1'b1), .Q(
        wr_ptr_bin[2]) );
  DFFSR wr_ptr_gray_reg_1_ ( .D(n4557), .CLK(wclk), .R(n13221), .S(1'b1), .Q(
        wr_ptr_gray[1]) );
  DFFSR wr_ptr_gray_s_reg_1_ ( .D(n163), .CLK(rclk), .R(n13221), .S(1'b1), .Q(
        wr_ptr_gray_s[1]) );
  DFFSR wr_ptr_gray_ss_reg_1_ ( .D(n160), .CLK(rclk), .R(n13221), .S(1'b1), 
        .Q(wr_ptr_gray_ss[1]) );
  DFFSR wr_ptr_bin_reg_3_ ( .D(n3184), .CLK(wclk), .R(n13221), .S(1'b1), .Q(
        wr_ptr_bin[3]) );
  DFFSR wr_ptr_gray_reg_2_ ( .D(n22), .CLK(wclk), .R(n13221), .S(1'b1), .Q(
        wr_ptr_gray[2]) );
  DFFSR wr_ptr_gray_s_reg_2_ ( .D(n157), .CLK(rclk), .R(n13221), .S(1'b1), .Q(
        wr_ptr_gray_s[2]) );
  DFFSR wr_ptr_gray_ss_reg_2_ ( .D(n154), .CLK(rclk), .R(n13221), .S(1'b1), 
        .Q(wr_ptr_gray_ss[2]) );
  DFFSR wr_ptr_bin_reg_4_ ( .D(n3179), .CLK(wclk), .R(n13221), .S(1'b1), .Q(
        wr_ptr_bin[4]) );
  DFFSR wr_ptr_gray_reg_3_ ( .D(n21), .CLK(wclk), .R(n13151), .S(1'b1), .Q(
        wr_ptr_gray[3]) );
  DFFSR wr_ptr_gray_s_reg_3_ ( .D(n151), .CLK(rclk), .R(n13151), .S(1'b1), .Q(
        wr_ptr_gray_s[3]) );
  DFFSR wr_ptr_gray_ss_reg_3_ ( .D(n148), .CLK(rclk), .R(n13151), .S(1'b1), 
        .Q(wr_ptr_gray_ss[3]) );
  DFFSR wr_ptr_gray_reg_4_ ( .D(n20), .CLK(wclk), .R(n13151), .S(1'b1), .Q(
        wr_ptr_gray[4]) );
  DFFSR wr_ptr_gray_s_reg_4_ ( .D(n145), .CLK(rclk), .R(n13151), .S(1'b1), .Q(
        wr_ptr_gray_s[4]) );
  DFFSR wr_ptr_gray_ss_reg_4_ ( .D(n142), .CLK(rclk), .R(n13151), .S(1'b1), 
        .Q(wr_ptr_gray_ss[4]) );
  DFFSR data_out_reg_0_ ( .D(n3171), .CLK(rclk), .R(n13146), .S(1'b1), .Q(
        n14723) );
  DFFSR data_out_reg_1_ ( .D(n3169), .CLK(rclk), .R(n13143), .S(1'b1), .Q(
        n14722) );
  DFFSR data_out_reg_2_ ( .D(n3167), .CLK(rclk), .R(n13140), .S(1'b1), .Q(
        n14721) );
  DFFSR data_out_reg_3_ ( .D(n3165), .CLK(rclk), .R(n13138), .S(1'b1), .Q(
        n14720) );
  DFFSR data_out_reg_4_ ( .D(n3163), .CLK(rclk), .R(n13135), .S(1'b1), .Q(
        n14719) );
  DFFSR data_out_reg_5_ ( .D(n3161), .CLK(rclk), .R(n13132), .S(1'b1), .Q(
        n14718) );
  DFFSR data_out_reg_6_ ( .D(n3159), .CLK(rclk), .R(n13129), .S(1'b1), .Q(
        n14717) );
  DFFSR data_out_reg_7_ ( .D(n3157), .CLK(rclk), .R(n13127), .S(1'b1), .Q(
        n14716) );
  DFFSR data_out_reg_8_ ( .D(n3155), .CLK(rclk), .R(n13124), .S(1'b1), .Q(
        n14715) );
  DFFSR data_out_reg_9_ ( .D(n3153), .CLK(rclk), .R(n13121), .S(1'b1), .Q(
        n14714) );
  DFFSR data_out_reg_10_ ( .D(n3151), .CLK(rclk), .R(n13118), .S(1'b1), .Q(
        n14713) );
  DFFSR data_out_reg_11_ ( .D(n3149), .CLK(rclk), .R(n13116), .S(1'b1), .Q(
        n14712) );
  DFFSR data_out_reg_12_ ( .D(n3147), .CLK(rclk), .R(n13113), .S(1'b1), .Q(
        n14711) );
  DFFSR data_out_reg_13_ ( .D(n3145), .CLK(rclk), .R(n13110), .S(1'b1), .Q(
        n14710) );
  DFFSR data_out_reg_14_ ( .D(n3143), .CLK(rclk), .R(n13107), .S(1'b1), .Q(
        n14709) );
  DFFSR data_out_reg_15_ ( .D(n3141), .CLK(rclk), .R(n13105), .S(1'b1), .Q(
        n14708) );
  DFFSR data_out_reg_16_ ( .D(n3139), .CLK(rclk), .R(n13151), .S(1'b1), .Q(
        n14707) );
  DFFSR data_out_reg_17_ ( .D(n3137), .CLK(rclk), .R(n13151), .S(1'b1), .Q(
        n14706) );
  DFFSR data_out_reg_18_ ( .D(n3135), .CLK(rclk), .R(n13150), .S(1'b1), .Q(
        n14705) );
  DFFSR data_out_reg_19_ ( .D(n3133), .CLK(rclk), .R(n13150), .S(1'b1), .Q(
        n14704) );
  DFFSR data_out_reg_20_ ( .D(n3131), .CLK(rclk), .R(n13150), .S(1'b1), .Q(
        n14703) );
  DFFSR data_out_reg_21_ ( .D(n3129), .CLK(rclk), .R(n13150), .S(1'b1), .Q(
        n14702) );
  DFFSR data_out_reg_22_ ( .D(n3127), .CLK(rclk), .R(n13150), .S(1'b1), .Q(
        n14701) );
  DFFSR data_out_reg_23_ ( .D(n3125), .CLK(rclk), .R(n13150), .S(1'b1), .Q(
        n14700) );
  DFFSR data_out_reg_24_ ( .D(n3123), .CLK(rclk), .R(n13150), .S(1'b1), .Q(
        n14699) );
  DFFSR data_out_reg_25_ ( .D(n3121), .CLK(rclk), .R(n13150), .S(1'b1), .Q(
        n14698) );
  DFFSR data_out_reg_26_ ( .D(n3119), .CLK(rclk), .R(n13150), .S(1'b1), .Q(
        n14697) );
  DFFSR data_out_reg_27_ ( .D(n3117), .CLK(rclk), .R(n13150), .S(1'b1), .Q(
        n14696) );
  DFFSR data_out_reg_28_ ( .D(n3115), .CLK(rclk), .R(n13150), .S(1'b1), .Q(
        n14695) );
  DFFSR data_out_reg_29_ ( .D(n3113), .CLK(rclk), .R(n13150), .S(1'b1), .Q(
        n14694) );
  DFFSR data_out_reg_30_ ( .D(n3111), .CLK(rclk), .R(n13149), .S(1'b1), .Q(
        n14693) );
  DFFSR data_out_reg_31_ ( .D(n3109), .CLK(rclk), .R(n13149), .S(1'b1), .Q(
        n14692) );
  DFFSR data_out_reg_32_ ( .D(n3107), .CLK(rclk), .R(n13149), .S(1'b1), .Q(
        n14691) );
  DFFSR data_out_reg_33_ ( .D(n3105), .CLK(rclk), .R(n13149), .S(1'b1), .Q(
        n14690) );
  DFFSR data_out_reg_34_ ( .D(n3103), .CLK(rclk), .R(n13149), .S(1'b1), .Q(
        n14689) );
  DFFSR data_out_reg_35_ ( .D(n3101), .CLK(rclk), .R(n13149), .S(1'b1), .Q(
        n14688) );
  DFFSR data_out_reg_36_ ( .D(n3099), .CLK(rclk), .R(n13149), .S(1'b1), .Q(
        n14687) );
  DFFSR data_out_reg_37_ ( .D(n3097), .CLK(rclk), .R(n13149), .S(1'b1), .Q(
        n14686) );
  DFFSR data_out_reg_38_ ( .D(n3095), .CLK(rclk), .R(n13149), .S(1'b1), .Q(
        n14685) );
  DFFSR data_out_reg_39_ ( .D(n3093), .CLK(rclk), .R(n13149), .S(1'b1), .Q(
        n14684) );
  DFFSR data_out_reg_40_ ( .D(n3091), .CLK(rclk), .R(n13149), .S(1'b1), .Q(
        n14683) );
  DFFSR data_out_reg_41_ ( .D(n3089), .CLK(rclk), .R(n13149), .S(1'b1), .Q(
        n14682) );
  DFFSR rd_ptr_bin_reg_1_ ( .D(n3087), .CLK(rclk), .R(n13224), .S(1'b1), .Q(
        n11) );
  DFFSR rd_ptr_gray_reg_0_ ( .D(n19), .CLK(rclk), .R(n13224), .S(1'b1), .Q(
        rd_ptr_gray[0]) );
  DFFSR rd_ptr_gray_s_reg_0_ ( .D(n139), .CLK(wclk), .R(n13224), .S(1'b1), .Q(
        rd_ptr_gray_s[0]) );
  DFFSR rd_ptr_gray_ss_reg_0_ ( .D(n136), .CLK(wclk), .R(n13224), .S(1'b1), 
        .Q(rd_ptr_gray_ss[0]) );
  DFFSR rd_ptr_bin_reg_2_ ( .D(n3082), .CLK(rclk), .R(n13224), .S(1'b1), .Q(
        n12) );
  DFFSR rd_ptr_gray_reg_1_ ( .D(n18), .CLK(rclk), .R(n13223), .S(1'b1), .Q(
        rd_ptr_gray[1]) );
  DFFSR rd_ptr_gray_s_reg_1_ ( .D(n133), .CLK(wclk), .R(n13223), .S(1'b1), .Q(
        rd_ptr_gray_s[1]) );
  DFFSR rd_ptr_gray_ss_reg_1_ ( .D(n130), .CLK(wclk), .R(n13223), .S(1'b1), 
        .Q(rd_ptr_gray_ss[1]) );
  DFFSR rd_ptr_bin_reg_3_ ( .D(n3077), .CLK(rclk), .R(n13223), .S(1'b1), .Q(
        n13) );
  DFFSR rd_ptr_gray_reg_2_ ( .D(n17), .CLK(rclk), .R(n13223), .S(1'b1), .Q(
        rd_ptr_gray[2]) );
  DFFSR rd_ptr_gray_s_reg_2_ ( .D(n127), .CLK(wclk), .R(n13223), .S(1'b1), .Q(
        rd_ptr_gray_s[2]) );
  DFFSR rd_ptr_gray_ss_reg_2_ ( .D(n124), .CLK(wclk), .R(n13223), .S(1'b1), 
        .Q(rd_ptr_gray_ss[2]) );
  DFFSR rd_ptr_bin_reg_4_ ( .D(n3072), .CLK(rclk), .R(n13223), .S(1'b1), .Q(
        n14) );
  DFFSR rd_ptr_gray_reg_3_ ( .D(n16), .CLK(rclk), .R(n13222), .S(1'b1), .Q(
        rd_ptr_gray[3]) );
  DFFSR rd_ptr_gray_s_reg_3_ ( .D(n121), .CLK(wclk), .R(n13222), .S(1'b1), .Q(
        rd_ptr_gray_s[3]) );
  DFFSR rd_ptr_gray_ss_reg_3_ ( .D(n113), .CLK(wclk), .R(n13222), .S(1'b1), 
        .Q(rd_ptr_gray_ss[3]) );
  DFFSR fifo_reg_0__41_ ( .D(n3213), .CLK(wclk), .R(n13186), .S(1'b1), .Q(
        fifo[1343]) );
  DFFSR fifo_reg_0__40_ ( .D(n3214), .CLK(wclk), .R(n13186), .S(1'b1), .Q(
        fifo[1342]) );
  DFFSR fifo_reg_0__39_ ( .D(n3215), .CLK(wclk), .R(n13186), .S(1'b1), .Q(
        fifo[1341]) );
  DFFSR fifo_reg_0__38_ ( .D(n3216), .CLK(wclk), .R(n13186), .S(1'b1), .Q(
        fifo[1340]) );
  DFFSR fifo_reg_0__37_ ( .D(n3217), .CLK(wclk), .R(n13186), .S(1'b1), .Q(
        fifo[1339]) );
  DFFSR fifo_reg_0__36_ ( .D(n3218), .CLK(wclk), .R(n13186), .S(1'b1), .Q(
        fifo[1338]) );
  DFFSR fifo_reg_0__35_ ( .D(n3219), .CLK(wclk), .R(n13186), .S(1'b1), .Q(
        fifo[1337]) );
  DFFSR fifo_reg_0__34_ ( .D(n3220), .CLK(wclk), .R(n13186), .S(1'b1), .Q(
        fifo[1336]) );
  DFFSR fifo_reg_0__33_ ( .D(n3221), .CLK(wclk), .R(n13187), .S(1'b1), .Q(
        fifo[1335]) );
  DFFSR fifo_reg_0__32_ ( .D(n3222), .CLK(wclk), .R(n13187), .S(1'b1), .Q(
        fifo[1334]) );
  DFFSR fifo_reg_0__31_ ( .D(n3223), .CLK(wclk), .R(n13187), .S(1'b1), .Q(
        fifo[1333]) );
  DFFSR fifo_reg_0__30_ ( .D(n3224), .CLK(wclk), .R(n13187), .S(1'b1), .Q(
        fifo[1332]) );
  DFFSR fifo_reg_0__29_ ( .D(n3225), .CLK(wclk), .R(n13187), .S(1'b1), .Q(
        fifo[1331]) );
  DFFSR fifo_reg_0__28_ ( .D(n3226), .CLK(wclk), .R(n13187), .S(1'b1), .Q(
        fifo[1330]) );
  DFFSR fifo_reg_0__27_ ( .D(n3227), .CLK(wclk), .R(n13187), .S(1'b1), .Q(
        fifo[1329]) );
  DFFSR fifo_reg_0__26_ ( .D(n3228), .CLK(wclk), .R(n13187), .S(1'b1), .Q(
        fifo[1328]) );
  DFFSR fifo_reg_0__25_ ( .D(n3229), .CLK(wclk), .R(n13187), .S(1'b1), .Q(
        fifo[1327]) );
  DFFSR fifo_reg_0__24_ ( .D(n3230), .CLK(wclk), .R(n13187), .S(1'b1), .Q(
        fifo[1326]) );
  DFFSR fifo_reg_0__23_ ( .D(n3231), .CLK(wclk), .R(n13187), .S(1'b1), .Q(
        fifo[1325]) );
  DFFSR fifo_reg_0__22_ ( .D(n3232), .CLK(wclk), .R(n13187), .S(1'b1), .Q(
        fifo[1324]) );
  DFFSR fifo_reg_0__21_ ( .D(n3233), .CLK(wclk), .R(n13188), .S(1'b1), .Q(
        fifo[1323]) );
  DFFSR fifo_reg_0__20_ ( .D(n3234), .CLK(wclk), .R(n13188), .S(1'b1), .Q(
        fifo[1322]) );
  DFFSR fifo_reg_0__19_ ( .D(n3235), .CLK(wclk), .R(n13188), .S(1'b1), .Q(
        fifo[1321]) );
  DFFSR fifo_reg_0__18_ ( .D(n3236), .CLK(wclk), .R(n13188), .S(1'b1), .Q(
        fifo[1320]) );
  DFFSR fifo_reg_0__17_ ( .D(n3237), .CLK(wclk), .R(n13188), .S(1'b1), .Q(
        fifo[1319]) );
  DFFSR fifo_reg_0__16_ ( .D(n3238), .CLK(wclk), .R(n13188), .S(1'b1), .Q(
        fifo[1318]) );
  DFFSR fifo_reg_0__15_ ( .D(n3239), .CLK(wclk), .R(n13105), .S(1'b1), .Q(
        fifo[1317]) );
  DFFSR fifo_reg_0__14_ ( .D(n3240), .CLK(wclk), .R(n13107), .S(1'b1), .Q(
        fifo[1316]) );
  DFFSR fifo_reg_0__13_ ( .D(n3241), .CLK(wclk), .R(n13110), .S(1'b1), .Q(
        fifo[1315]) );
  DFFSR fifo_reg_0__12_ ( .D(n3242), .CLK(wclk), .R(n13113), .S(1'b1), .Q(
        fifo[1314]) );
  DFFSR fifo_reg_0__11_ ( .D(n3243), .CLK(wclk), .R(n13116), .S(1'b1), .Q(
        fifo[1313]) );
  DFFSR fifo_reg_0__10_ ( .D(n3244), .CLK(wclk), .R(n13118), .S(1'b1), .Q(
        fifo[1312]) );
  DFFSR fifo_reg_0__9_ ( .D(n3245), .CLK(wclk), .R(n13121), .S(1'b1), .Q(
        fifo[1311]) );
  DFFSR fifo_reg_0__8_ ( .D(n3246), .CLK(wclk), .R(n13124), .S(1'b1), .Q(
        fifo[1310]) );
  DFFSR fifo_reg_0__7_ ( .D(n3247), .CLK(wclk), .R(n13127), .S(1'b1), .Q(
        fifo[1309]) );
  DFFSR fifo_reg_0__6_ ( .D(n3248), .CLK(wclk), .R(n13129), .S(1'b1), .Q(
        fifo[1308]) );
  DFFSR fifo_reg_0__5_ ( .D(n3249), .CLK(wclk), .R(n13132), .S(1'b1), .Q(
        fifo[1307]) );
  DFFSR fifo_reg_0__4_ ( .D(n3250), .CLK(wclk), .R(n13135), .S(1'b1), .Q(
        fifo[1306]) );
  DFFSR fifo_reg_0__3_ ( .D(n3251), .CLK(wclk), .R(n13138), .S(1'b1), .Q(
        fifo[1305]) );
  DFFSR fifo_reg_0__2_ ( .D(n3252), .CLK(wclk), .R(n13140), .S(1'b1), .Q(
        fifo[1304]) );
  DFFSR fifo_reg_0__1_ ( .D(n3253), .CLK(wclk), .R(n13143), .S(1'b1), .Q(
        fifo[1303]) );
  DFFSR fifo_reg_0__0_ ( .D(n3254), .CLK(wclk), .R(n13146), .S(1'b1), .Q(
        fifo[1302]) );
  DFFSR fifo_reg_1__41_ ( .D(n3255), .CLK(wclk), .R(n13188), .S(1'b1), .Q(
        fifo[1301]) );
  DFFSR fifo_reg_1__40_ ( .D(n3256), .CLK(wclk), .R(n13188), .S(1'b1), .Q(
        fifo[1300]) );
  DFFSR fifo_reg_1__39_ ( .D(n3257), .CLK(wclk), .R(n13188), .S(1'b1), .Q(
        fifo[1299]) );
  DFFSR fifo_reg_1__38_ ( .D(n3258), .CLK(wclk), .R(n13188), .S(1'b1), .Q(
        fifo[1298]) );
  DFFSR fifo_reg_1__37_ ( .D(n3259), .CLK(wclk), .R(n13188), .S(1'b1), .Q(
        fifo[1297]) );
  DFFSR fifo_reg_1__36_ ( .D(n3260), .CLK(wclk), .R(n13188), .S(1'b1), .Q(
        fifo[1296]) );
  DFFSR fifo_reg_1__35_ ( .D(n3261), .CLK(wclk), .R(n13189), .S(1'b1), .Q(
        fifo[1295]) );
  DFFSR fifo_reg_1__34_ ( .D(n3262), .CLK(wclk), .R(n13189), .S(1'b1), .Q(
        fifo[1294]) );
  DFFSR fifo_reg_1__33_ ( .D(n3263), .CLK(wclk), .R(n13189), .S(1'b1), .Q(
        fifo[1293]) );
  DFFSR fifo_reg_1__32_ ( .D(n3264), .CLK(wclk), .R(n13189), .S(1'b1), .Q(
        fifo[1292]) );
  DFFSR fifo_reg_1__31_ ( .D(n3265), .CLK(wclk), .R(n13189), .S(1'b1), .Q(
        fifo[1291]) );
  DFFSR fifo_reg_1__30_ ( .D(n3266), .CLK(wclk), .R(n13189), .S(1'b1), .Q(
        fifo[1290]) );
  DFFSR fifo_reg_1__29_ ( .D(n3267), .CLK(wclk), .R(n13189), .S(1'b1), .Q(
        fifo[1289]) );
  DFFSR fifo_reg_1__28_ ( .D(n3268), .CLK(wclk), .R(n13189), .S(1'b1), .Q(
        fifo[1288]) );
  DFFSR fifo_reg_1__27_ ( .D(n3269), .CLK(wclk), .R(n13189), .S(1'b1), .Q(
        fifo[1287]) );
  DFFSR fifo_reg_1__26_ ( .D(n3270), .CLK(wclk), .R(n13189), .S(1'b1), .Q(
        fifo[1286]) );
  DFFSR fifo_reg_1__25_ ( .D(n3271), .CLK(wclk), .R(n13189), .S(1'b1), .Q(
        fifo[1285]) );
  DFFSR fifo_reg_1__24_ ( .D(n3272), .CLK(wclk), .R(n13189), .S(1'b1), .Q(
        fifo[1284]) );
  DFFSR fifo_reg_1__23_ ( .D(n3273), .CLK(wclk), .R(n13190), .S(1'b1), .Q(
        fifo[1283]) );
  DFFSR fifo_reg_1__22_ ( .D(n3274), .CLK(wclk), .R(n13190), .S(1'b1), .Q(
        fifo[1282]) );
  DFFSR fifo_reg_1__21_ ( .D(n3275), .CLK(wclk), .R(n13190), .S(1'b1), .Q(
        fifo[1281]) );
  DFFSR fifo_reg_1__20_ ( .D(n3276), .CLK(wclk), .R(n13190), .S(1'b1), .Q(
        fifo[1280]) );
  DFFSR fifo_reg_1__19_ ( .D(n3277), .CLK(wclk), .R(n13190), .S(1'b1), .Q(
        fifo[1279]) );
  DFFSR fifo_reg_1__18_ ( .D(n3278), .CLK(wclk), .R(n13190), .S(1'b1), .Q(
        fifo[1278]) );
  DFFSR fifo_reg_1__17_ ( .D(n3279), .CLK(wclk), .R(n13190), .S(1'b1), .Q(
        fifo[1277]) );
  DFFSR fifo_reg_1__16_ ( .D(n3280), .CLK(wclk), .R(n13190), .S(1'b1), .Q(
        fifo[1276]) );
  DFFSR fifo_reg_1__15_ ( .D(n3281), .CLK(wclk), .R(n13105), .S(1'b1), .Q(
        fifo[1275]) );
  DFFSR fifo_reg_1__14_ ( .D(n3282), .CLK(wclk), .R(n13107), .S(1'b1), .Q(
        fifo[1274]) );
  DFFSR fifo_reg_1__13_ ( .D(n3283), .CLK(wclk), .R(n13110), .S(1'b1), .Q(
        fifo[1273]) );
  DFFSR fifo_reg_1__12_ ( .D(n3284), .CLK(wclk), .R(n13113), .S(1'b1), .Q(
        fifo[1272]) );
  DFFSR fifo_reg_1__11_ ( .D(n3285), .CLK(wclk), .R(n13116), .S(1'b1), .Q(
        fifo[1271]) );
  DFFSR fifo_reg_1__10_ ( .D(n3286), .CLK(wclk), .R(n13118), .S(1'b1), .Q(
        fifo[1270]) );
  DFFSR fifo_reg_1__9_ ( .D(n3287), .CLK(wclk), .R(n13121), .S(1'b1), .Q(
        fifo[1269]) );
  DFFSR fifo_reg_1__8_ ( .D(n3288), .CLK(wclk), .R(n13124), .S(1'b1), .Q(
        fifo[1268]) );
  DFFSR fifo_reg_1__7_ ( .D(n3289), .CLK(wclk), .R(n13127), .S(1'b1), .Q(
        fifo[1267]) );
  DFFSR fifo_reg_1__6_ ( .D(n3290), .CLK(wclk), .R(n13129), .S(1'b1), .Q(
        fifo[1266]) );
  DFFSR fifo_reg_1__5_ ( .D(n3291), .CLK(wclk), .R(n13132), .S(1'b1), .Q(
        fifo[1265]) );
  DFFSR fifo_reg_1__4_ ( .D(n3292), .CLK(wclk), .R(n13135), .S(1'b1), .Q(
        fifo[1264]) );
  DFFSR fifo_reg_1__3_ ( .D(n3293), .CLK(wclk), .R(n13138), .S(1'b1), .Q(
        fifo[1263]) );
  DFFSR fifo_reg_1__2_ ( .D(n3294), .CLK(wclk), .R(n13140), .S(1'b1), .Q(
        fifo[1262]) );
  DFFSR fifo_reg_1__1_ ( .D(n3295), .CLK(wclk), .R(n13143), .S(1'b1), .Q(
        fifo[1261]) );
  DFFSR fifo_reg_1__0_ ( .D(n3296), .CLK(wclk), .R(n13146), .S(1'b1), .Q(
        fifo[1260]) );
  DFFSR fifo_reg_2__41_ ( .D(n3297), .CLK(wclk), .R(n13190), .S(1'b1), .Q(
        fifo[1259]) );
  DFFSR fifo_reg_2__40_ ( .D(n3298), .CLK(wclk), .R(n13190), .S(1'b1), .Q(
        fifo[1258]) );
  DFFSR fifo_reg_2__39_ ( .D(n3299), .CLK(wclk), .R(n13190), .S(1'b1), .Q(
        fifo[1257]) );
  DFFSR fifo_reg_2__38_ ( .D(n3300), .CLK(wclk), .R(n13190), .S(1'b1), .Q(
        fifo[1256]) );
  DFFSR fifo_reg_2__37_ ( .D(n3301), .CLK(wclk), .R(n13191), .S(1'b1), .Q(
        fifo[1255]) );
  DFFSR fifo_reg_2__36_ ( .D(n3302), .CLK(wclk), .R(n13191), .S(1'b1), .Q(
        fifo[1254]) );
  DFFSR fifo_reg_2__35_ ( .D(n3303), .CLK(wclk), .R(n13191), .S(1'b1), .Q(
        fifo[1253]) );
  DFFSR fifo_reg_2__34_ ( .D(n3304), .CLK(wclk), .R(n13191), .S(1'b1), .Q(
        fifo[1252]) );
  DFFSR fifo_reg_2__33_ ( .D(n3305), .CLK(wclk), .R(n13191), .S(1'b1), .Q(
        fifo[1251]) );
  DFFSR fifo_reg_2__32_ ( .D(n3306), .CLK(wclk), .R(n13191), .S(1'b1), .Q(
        fifo[1250]) );
  DFFSR fifo_reg_2__31_ ( .D(n3307), .CLK(wclk), .R(n13191), .S(1'b1), .Q(
        fifo[1249]) );
  DFFSR fifo_reg_2__30_ ( .D(n3308), .CLK(wclk), .R(n13191), .S(1'b1), .Q(
        fifo[1248]) );
  DFFSR fifo_reg_2__29_ ( .D(n3309), .CLK(wclk), .R(n13191), .S(1'b1), .Q(
        fifo[1247]) );
  DFFSR fifo_reg_2__28_ ( .D(n3310), .CLK(wclk), .R(n13191), .S(1'b1), .Q(
        fifo[1246]) );
  DFFSR fifo_reg_2__27_ ( .D(n3311), .CLK(wclk), .R(n13191), .S(1'b1), .Q(
        fifo[1245]) );
  DFFSR fifo_reg_2__26_ ( .D(n3312), .CLK(wclk), .R(n13191), .S(1'b1), .Q(
        fifo[1244]) );
  DFFSR fifo_reg_2__25_ ( .D(n3313), .CLK(wclk), .R(n13192), .S(1'b1), .Q(
        fifo[1243]) );
  DFFSR fifo_reg_2__24_ ( .D(n3314), .CLK(wclk), .R(n13192), .S(1'b1), .Q(
        fifo[1242]) );
  DFFSR fifo_reg_2__23_ ( .D(n3315), .CLK(wclk), .R(n13192), .S(1'b1), .Q(
        fifo[1241]) );
  DFFSR fifo_reg_2__22_ ( .D(n3316), .CLK(wclk), .R(n13192), .S(1'b1), .Q(
        fifo[1240]) );
  DFFSR fifo_reg_2__21_ ( .D(n3317), .CLK(wclk), .R(n13192), .S(1'b1), .Q(
        fifo[1239]) );
  DFFSR fifo_reg_2__20_ ( .D(n3318), .CLK(wclk), .R(n13192), .S(1'b1), .Q(
        fifo[1238]) );
  DFFSR fifo_reg_2__19_ ( .D(n3319), .CLK(wclk), .R(n13192), .S(1'b1), .Q(
        fifo[1237]) );
  DFFSR fifo_reg_2__18_ ( .D(n3320), .CLK(wclk), .R(n13192), .S(1'b1), .Q(
        fifo[1236]) );
  DFFSR fifo_reg_2__17_ ( .D(n3321), .CLK(wclk), .R(n13192), .S(1'b1), .Q(
        fifo[1235]) );
  DFFSR fifo_reg_2__16_ ( .D(n3322), .CLK(wclk), .R(n13192), .S(1'b1), .Q(
        fifo[1234]) );
  DFFSR fifo_reg_2__15_ ( .D(n3323), .CLK(wclk), .R(n13105), .S(1'b1), .Q(
        fifo[1233]) );
  DFFSR fifo_reg_2__14_ ( .D(n3324), .CLK(wclk), .R(n13108), .S(1'b1), .Q(
        fifo[1232]) );
  DFFSR fifo_reg_2__13_ ( .D(n3325), .CLK(wclk), .R(n13110), .S(1'b1), .Q(
        fifo[1231]) );
  DFFSR fifo_reg_2__12_ ( .D(n3326), .CLK(wclk), .R(n13113), .S(1'b1), .Q(
        fifo[1230]) );
  DFFSR fifo_reg_2__11_ ( .D(n3327), .CLK(wclk), .R(n13116), .S(1'b1), .Q(
        fifo[1229]) );
  DFFSR fifo_reg_2__10_ ( .D(n3328), .CLK(wclk), .R(n13119), .S(1'b1), .Q(
        fifo[1228]) );
  DFFSR fifo_reg_2__9_ ( .D(n3329), .CLK(wclk), .R(n13121), .S(1'b1), .Q(
        fifo[1227]) );
  DFFSR fifo_reg_2__8_ ( .D(n3330), .CLK(wclk), .R(n13124), .S(1'b1), .Q(
        fifo[1226]) );
  DFFSR fifo_reg_2__7_ ( .D(n3331), .CLK(wclk), .R(n13127), .S(1'b1), .Q(
        fifo[1225]) );
  DFFSR fifo_reg_2__6_ ( .D(n3332), .CLK(wclk), .R(n13130), .S(1'b1), .Q(
        fifo[1224]) );
  DFFSR fifo_reg_2__5_ ( .D(n3333), .CLK(wclk), .R(n13132), .S(1'b1), .Q(
        fifo[1223]) );
  DFFSR fifo_reg_2__4_ ( .D(n3334), .CLK(wclk), .R(n13135), .S(1'b1), .Q(
        fifo[1222]) );
  DFFSR fifo_reg_2__3_ ( .D(n3335), .CLK(wclk), .R(n13138), .S(1'b1), .Q(
        fifo[1221]) );
  DFFSR fifo_reg_2__2_ ( .D(n3336), .CLK(wclk), .R(n13141), .S(1'b1), .Q(
        fifo[1220]) );
  DFFSR fifo_reg_2__1_ ( .D(n3337), .CLK(wclk), .R(n13143), .S(1'b1), .Q(
        fifo[1219]) );
  DFFSR fifo_reg_2__0_ ( .D(n3338), .CLK(wclk), .R(n13146), .S(1'b1), .Q(
        fifo[1218]) );
  DFFSR fifo_reg_3__41_ ( .D(n3339), .CLK(wclk), .R(n13192), .S(1'b1), .Q(
        fifo[1217]) );
  DFFSR fifo_reg_3__40_ ( .D(n3340), .CLK(wclk), .R(n13192), .S(1'b1), .Q(
        fifo[1216]) );
  DFFSR fifo_reg_3__39_ ( .D(n3341), .CLK(wclk), .R(n13193), .S(1'b1), .Q(
        fifo[1215]) );
  DFFSR fifo_reg_3__38_ ( .D(n3342), .CLK(wclk), .R(n13193), .S(1'b1), .Q(
        fifo[1214]) );
  DFFSR fifo_reg_3__37_ ( .D(n3343), .CLK(wclk), .R(n13193), .S(1'b1), .Q(
        fifo[1213]) );
  DFFSR fifo_reg_3__36_ ( .D(n3344), .CLK(wclk), .R(n13193), .S(1'b1), .Q(
        fifo[1212]) );
  DFFSR fifo_reg_3__35_ ( .D(n3345), .CLK(wclk), .R(n13193), .S(1'b1), .Q(
        fifo[1211]) );
  DFFSR fifo_reg_3__34_ ( .D(n3346), .CLK(wclk), .R(n13193), .S(1'b1), .Q(
        fifo[1210]) );
  DFFSR fifo_reg_3__33_ ( .D(n3347), .CLK(wclk), .R(n13193), .S(1'b1), .Q(
        fifo[1209]) );
  DFFSR fifo_reg_3__32_ ( .D(n3348), .CLK(wclk), .R(n13193), .S(1'b1), .Q(
        fifo[1208]) );
  DFFSR fifo_reg_3__31_ ( .D(n3349), .CLK(wclk), .R(n13193), .S(1'b1), .Q(
        fifo[1207]) );
  DFFSR fifo_reg_3__30_ ( .D(n3350), .CLK(wclk), .R(n13193), .S(1'b1), .Q(
        fifo[1206]) );
  DFFSR fifo_reg_3__29_ ( .D(n3351), .CLK(wclk), .R(n13193), .S(1'b1), .Q(
        fifo[1205]) );
  DFFSR fifo_reg_3__28_ ( .D(n3352), .CLK(wclk), .R(n13193), .S(1'b1), .Q(
        fifo[1204]) );
  DFFSR fifo_reg_3__27_ ( .D(n3353), .CLK(wclk), .R(n13194), .S(1'b1), .Q(
        fifo[1203]) );
  DFFSR fifo_reg_3__26_ ( .D(n3354), .CLK(wclk), .R(n13194), .S(1'b1), .Q(
        fifo[1202]) );
  DFFSR fifo_reg_3__25_ ( .D(n3355), .CLK(wclk), .R(n13194), .S(1'b1), .Q(
        fifo[1201]) );
  DFFSR fifo_reg_3__24_ ( .D(n3356), .CLK(wclk), .R(n13194), .S(1'b1), .Q(
        fifo[1200]) );
  DFFSR fifo_reg_3__23_ ( .D(n3357), .CLK(wclk), .R(n13194), .S(1'b1), .Q(
        fifo[1199]) );
  DFFSR fifo_reg_3__22_ ( .D(n3358), .CLK(wclk), .R(n13194), .S(1'b1), .Q(
        fifo[1198]) );
  DFFSR fifo_reg_3__21_ ( .D(n3359), .CLK(wclk), .R(n13194), .S(1'b1), .Q(
        fifo[1197]) );
  DFFSR fifo_reg_3__20_ ( .D(n3360), .CLK(wclk), .R(n13194), .S(1'b1), .Q(
        fifo[1196]) );
  DFFSR fifo_reg_3__19_ ( .D(n3361), .CLK(wclk), .R(n13194), .S(1'b1), .Q(
        fifo[1195]) );
  DFFSR fifo_reg_3__18_ ( .D(n3362), .CLK(wclk), .R(n13194), .S(1'b1), .Q(
        fifo[1194]) );
  DFFSR fifo_reg_3__17_ ( .D(n3363), .CLK(wclk), .R(n13194), .S(1'b1), .Q(
        fifo[1193]) );
  DFFSR fifo_reg_3__16_ ( .D(n3364), .CLK(wclk), .R(n13194), .S(1'b1), .Q(
        fifo[1192]) );
  DFFSR fifo_reg_3__15_ ( .D(n3365), .CLK(wclk), .R(n13105), .S(1'b1), .Q(
        fifo[1191]) );
  DFFSR fifo_reg_3__14_ ( .D(n3366), .CLK(wclk), .R(n13108), .S(1'b1), .Q(
        fifo[1190]) );
  DFFSR fifo_reg_3__13_ ( .D(n3367), .CLK(wclk), .R(n13110), .S(1'b1), .Q(
        fifo[1189]) );
  DFFSR fifo_reg_3__12_ ( .D(n3368), .CLK(wclk), .R(n13113), .S(1'b1), .Q(
        fifo[1188]) );
  DFFSR fifo_reg_3__11_ ( .D(n3369), .CLK(wclk), .R(n13116), .S(1'b1), .Q(
        fifo[1187]) );
  DFFSR fifo_reg_3__10_ ( .D(n3370), .CLK(wclk), .R(n13119), .S(1'b1), .Q(
        fifo[1186]) );
  DFFSR fifo_reg_3__9_ ( .D(n3371), .CLK(wclk), .R(n13121), .S(1'b1), .Q(
        fifo[1185]) );
  DFFSR fifo_reg_3__8_ ( .D(n3372), .CLK(wclk), .R(n13124), .S(1'b1), .Q(
        fifo[1184]) );
  DFFSR fifo_reg_3__7_ ( .D(n3373), .CLK(wclk), .R(n13127), .S(1'b1), .Q(
        fifo[1183]) );
  DFFSR fifo_reg_3__6_ ( .D(n3374), .CLK(wclk), .R(n13130), .S(1'b1), .Q(
        fifo[1182]) );
  DFFSR fifo_reg_3__5_ ( .D(n3375), .CLK(wclk), .R(n13132), .S(1'b1), .Q(
        fifo[1181]) );
  DFFSR fifo_reg_3__4_ ( .D(n3376), .CLK(wclk), .R(n13135), .S(1'b1), .Q(
        fifo[1180]) );
  DFFSR fifo_reg_3__3_ ( .D(n3377), .CLK(wclk), .R(n13138), .S(1'b1), .Q(
        fifo[1179]) );
  DFFSR fifo_reg_3__2_ ( .D(n3378), .CLK(wclk), .R(n13141), .S(1'b1), .Q(
        fifo[1178]) );
  DFFSR fifo_reg_3__1_ ( .D(n3379), .CLK(wclk), .R(n13143), .S(1'b1), .Q(
        fifo[1177]) );
  DFFSR fifo_reg_3__0_ ( .D(n3380), .CLK(wclk), .R(n13146), .S(1'b1), .Q(
        fifo[1176]) );
  DFFSR fifo_reg_4__41_ ( .D(n3381), .CLK(wclk), .R(n13195), .S(1'b1), .Q(
        fifo[1175]) );
  DFFSR fifo_reg_4__40_ ( .D(n3382), .CLK(wclk), .R(n13195), .S(1'b1), .Q(
        fifo[1174]) );
  DFFSR fifo_reg_4__39_ ( .D(n3383), .CLK(wclk), .R(n13195), .S(1'b1), .Q(
        fifo[1173]) );
  DFFSR fifo_reg_4__38_ ( .D(n3384), .CLK(wclk), .R(n13195), .S(1'b1), .Q(
        fifo[1172]) );
  DFFSR fifo_reg_4__37_ ( .D(n3385), .CLK(wclk), .R(n13195), .S(1'b1), .Q(
        fifo[1171]) );
  DFFSR fifo_reg_4__36_ ( .D(n3386), .CLK(wclk), .R(n13195), .S(1'b1), .Q(
        fifo[1170]) );
  DFFSR fifo_reg_4__35_ ( .D(n3387), .CLK(wclk), .R(n13195), .S(1'b1), .Q(
        fifo[1169]) );
  DFFSR fifo_reg_4__34_ ( .D(n3388), .CLK(wclk), .R(n13195), .S(1'b1), .Q(
        fifo[1168]) );
  DFFSR fifo_reg_4__33_ ( .D(n3389), .CLK(wclk), .R(n13195), .S(1'b1), .Q(
        fifo[1167]) );
  DFFSR fifo_reg_4__32_ ( .D(n3390), .CLK(wclk), .R(n13195), .S(1'b1), .Q(
        fifo[1166]) );
  DFFSR fifo_reg_4__31_ ( .D(n3391), .CLK(wclk), .R(n13195), .S(1'b1), .Q(
        fifo[1165]) );
  DFFSR fifo_reg_4__30_ ( .D(n3392), .CLK(wclk), .R(n13195), .S(1'b1), .Q(
        fifo[1164]) );
  DFFSR fifo_reg_4__29_ ( .D(n3393), .CLK(wclk), .R(n13196), .S(1'b1), .Q(
        fifo[1163]) );
  DFFSR fifo_reg_4__28_ ( .D(n3394), .CLK(wclk), .R(n13196), .S(1'b1), .Q(
        fifo[1162]) );
  DFFSR fifo_reg_4__27_ ( .D(n3395), .CLK(wclk), .R(n13196), .S(1'b1), .Q(
        fifo[1161]) );
  DFFSR fifo_reg_4__26_ ( .D(n3396), .CLK(wclk), .R(n13196), .S(1'b1), .Q(
        fifo[1160]) );
  DFFSR fifo_reg_4__25_ ( .D(n3397), .CLK(wclk), .R(n13196), .S(1'b1), .Q(
        fifo[1159]) );
  DFFSR fifo_reg_4__24_ ( .D(n3398), .CLK(wclk), .R(n13196), .S(1'b1), .Q(
        fifo[1158]) );
  DFFSR fifo_reg_4__23_ ( .D(n3399), .CLK(wclk), .R(n13196), .S(1'b1), .Q(
        fifo[1157]) );
  DFFSR fifo_reg_4__22_ ( .D(n3400), .CLK(wclk), .R(n13196), .S(1'b1), .Q(
        fifo[1156]) );
  DFFSR fifo_reg_4__21_ ( .D(n3401), .CLK(wclk), .R(n13196), .S(1'b1), .Q(
        fifo[1155]) );
  DFFSR fifo_reg_4__20_ ( .D(n3402), .CLK(wclk), .R(n13196), .S(1'b1), .Q(
        fifo[1154]) );
  DFFSR fifo_reg_4__19_ ( .D(n3403), .CLK(wclk), .R(n13196), .S(1'b1), .Q(
        fifo[1153]) );
  DFFSR fifo_reg_4__18_ ( .D(n3404), .CLK(wclk), .R(n13196), .S(1'b1), .Q(
        fifo[1152]) );
  DFFSR fifo_reg_4__17_ ( .D(n3405), .CLK(wclk), .R(n13197), .S(1'b1), .Q(
        fifo[1151]) );
  DFFSR fifo_reg_4__16_ ( .D(n3406), .CLK(wclk), .R(n13197), .S(1'b1), .Q(
        fifo[1150]) );
  DFFSR fifo_reg_4__15_ ( .D(n3407), .CLK(wclk), .R(n13105), .S(1'b1), .Q(
        fifo[1149]) );
  DFFSR fifo_reg_4__14_ ( .D(n3408), .CLK(wclk), .R(n13108), .S(1'b1), .Q(
        fifo[1148]) );
  DFFSR fifo_reg_4__13_ ( .D(n3409), .CLK(wclk), .R(n13110), .S(1'b1), .Q(
        fifo[1147]) );
  DFFSR fifo_reg_4__12_ ( .D(n3410), .CLK(wclk), .R(n13113), .S(1'b1), .Q(
        fifo[1146]) );
  DFFSR fifo_reg_4__11_ ( .D(n3411), .CLK(wclk), .R(n13116), .S(1'b1), .Q(
        fifo[1145]) );
  DFFSR fifo_reg_4__10_ ( .D(n3412), .CLK(wclk), .R(n13119), .S(1'b1), .Q(
        fifo[1144]) );
  DFFSR fifo_reg_4__9_ ( .D(n3413), .CLK(wclk), .R(n13121), .S(1'b1), .Q(
        fifo[1143]) );
  DFFSR fifo_reg_4__8_ ( .D(n3414), .CLK(wclk), .R(n13124), .S(1'b1), .Q(
        fifo[1142]) );
  DFFSR fifo_reg_4__7_ ( .D(n3415), .CLK(wclk), .R(n13127), .S(1'b1), .Q(
        fifo[1141]) );
  DFFSR fifo_reg_4__6_ ( .D(n3416), .CLK(wclk), .R(n13130), .S(1'b1), .Q(
        fifo[1140]) );
  DFFSR fifo_reg_4__5_ ( .D(n3417), .CLK(wclk), .R(n13132), .S(1'b1), .Q(
        fifo[1139]) );
  DFFSR fifo_reg_4__4_ ( .D(n3418), .CLK(wclk), .R(n13135), .S(1'b1), .Q(
        fifo[1138]) );
  DFFSR fifo_reg_4__3_ ( .D(n3419), .CLK(wclk), .R(n13138), .S(1'b1), .Q(
        fifo[1137]) );
  DFFSR fifo_reg_4__2_ ( .D(n3420), .CLK(wclk), .R(n13141), .S(1'b1), .Q(
        fifo[1136]) );
  DFFSR fifo_reg_4__1_ ( .D(n3421), .CLK(wclk), .R(n13143), .S(1'b1), .Q(
        fifo[1135]) );
  DFFSR fifo_reg_4__0_ ( .D(n3422), .CLK(wclk), .R(n13146), .S(1'b1), .Q(
        fifo[1134]) );
  DFFSR fifo_reg_5__41_ ( .D(n3423), .CLK(wclk), .R(n13197), .S(1'b1), .Q(
        fifo[1133]) );
  DFFSR fifo_reg_5__40_ ( .D(n3424), .CLK(wclk), .R(n13197), .S(1'b1), .Q(
        fifo[1132]) );
  DFFSR fifo_reg_5__39_ ( .D(n3425), .CLK(wclk), .R(n13197), .S(1'b1), .Q(
        fifo[1131]) );
  DFFSR fifo_reg_5__38_ ( .D(n3426), .CLK(wclk), .R(n13197), .S(1'b1), .Q(
        fifo[1130]) );
  DFFSR fifo_reg_5__37_ ( .D(n3427), .CLK(wclk), .R(n13197), .S(1'b1), .Q(
        fifo[1129]) );
  DFFSR fifo_reg_5__36_ ( .D(n3428), .CLK(wclk), .R(n13197), .S(1'b1), .Q(
        fifo[1128]) );
  DFFSR fifo_reg_5__35_ ( .D(n3429), .CLK(wclk), .R(n13197), .S(1'b1), .Q(
        fifo[1127]) );
  DFFSR fifo_reg_5__34_ ( .D(n3430), .CLK(wclk), .R(n13197), .S(1'b1), .Q(
        fifo[1126]) );
  DFFSR fifo_reg_5__33_ ( .D(n3431), .CLK(wclk), .R(n13197), .S(1'b1), .Q(
        fifo[1125]) );
  DFFSR fifo_reg_5__32_ ( .D(n3432), .CLK(wclk), .R(n13197), .S(1'b1), .Q(
        fifo[1124]) );
  DFFSR fifo_reg_5__31_ ( .D(n3433), .CLK(wclk), .R(n13198), .S(1'b1), .Q(
        fifo[1123]) );
  DFFSR fifo_reg_5__30_ ( .D(n3434), .CLK(wclk), .R(n13198), .S(1'b1), .Q(
        fifo[1122]) );
  DFFSR fifo_reg_5__29_ ( .D(n3435), .CLK(wclk), .R(n13198), .S(1'b1), .Q(
        fifo[1121]) );
  DFFSR fifo_reg_5__28_ ( .D(n3436), .CLK(wclk), .R(n13198), .S(1'b1), .Q(
        fifo[1120]) );
  DFFSR fifo_reg_5__27_ ( .D(n3437), .CLK(wclk), .R(n13198), .S(1'b1), .Q(
        fifo[1119]) );
  DFFSR fifo_reg_5__26_ ( .D(n3438), .CLK(wclk), .R(n13198), .S(1'b1), .Q(
        fifo[1118]) );
  DFFSR fifo_reg_5__25_ ( .D(n3439), .CLK(wclk), .R(n13198), .S(1'b1), .Q(
        fifo[1117]) );
  DFFSR fifo_reg_5__24_ ( .D(n3440), .CLK(wclk), .R(n13198), .S(1'b1), .Q(
        fifo[1116]) );
  DFFSR fifo_reg_5__23_ ( .D(n3441), .CLK(wclk), .R(n13198), .S(1'b1), .Q(
        fifo[1115]) );
  DFFSR fifo_reg_5__22_ ( .D(n3442), .CLK(wclk), .R(n13198), .S(1'b1), .Q(
        fifo[1114]) );
  DFFSR fifo_reg_5__21_ ( .D(n3443), .CLK(wclk), .R(n13198), .S(1'b1), .Q(
        fifo[1113]) );
  DFFSR fifo_reg_5__20_ ( .D(n3444), .CLK(wclk), .R(n13198), .S(1'b1), .Q(
        fifo[1112]) );
  DFFSR fifo_reg_5__19_ ( .D(n3445), .CLK(wclk), .R(n13199), .S(1'b1), .Q(
        fifo[1111]) );
  DFFSR fifo_reg_5__18_ ( .D(n3446), .CLK(wclk), .R(n13199), .S(1'b1), .Q(
        fifo[1110]) );
  DFFSR fifo_reg_5__17_ ( .D(n3447), .CLK(wclk), .R(n13199), .S(1'b1), .Q(
        fifo[1109]) );
  DFFSR fifo_reg_5__16_ ( .D(n3448), .CLK(wclk), .R(n13199), .S(1'b1), .Q(
        fifo[1108]) );
  DFFSR fifo_reg_5__15_ ( .D(n3449), .CLK(wclk), .R(n13105), .S(1'b1), .Q(
        fifo[1107]) );
  DFFSR fifo_reg_5__14_ ( .D(n3450), .CLK(wclk), .R(n13108), .S(1'b1), .Q(
        fifo[1106]) );
  DFFSR fifo_reg_5__13_ ( .D(n3451), .CLK(wclk), .R(n13111), .S(1'b1), .Q(
        fifo[1105]) );
  DFFSR fifo_reg_5__12_ ( .D(n3452), .CLK(wclk), .R(n13113), .S(1'b1), .Q(
        fifo[1104]) );
  DFFSR fifo_reg_5__11_ ( .D(n3453), .CLK(wclk), .R(n13116), .S(1'b1), .Q(
        fifo[1103]) );
  DFFSR fifo_reg_5__10_ ( .D(n3454), .CLK(wclk), .R(n13119), .S(1'b1), .Q(
        fifo[1102]) );
  DFFSR fifo_reg_5__9_ ( .D(n3455), .CLK(wclk), .R(n13122), .S(1'b1), .Q(
        fifo[1101]) );
  DFFSR fifo_reg_5__8_ ( .D(n3456), .CLK(wclk), .R(n13124), .S(1'b1), .Q(
        fifo[1100]) );
  DFFSR fifo_reg_5__7_ ( .D(n3457), .CLK(wclk), .R(n13127), .S(1'b1), .Q(
        fifo[1099]) );
  DFFSR fifo_reg_5__6_ ( .D(n3458), .CLK(wclk), .R(n13130), .S(1'b1), .Q(
        fifo[1098]) );
  DFFSR fifo_reg_5__5_ ( .D(n3459), .CLK(wclk), .R(n13133), .S(1'b1), .Q(
        fifo[1097]) );
  DFFSR fifo_reg_5__4_ ( .D(n3460), .CLK(wclk), .R(n13135), .S(1'b1), .Q(
        fifo[1096]) );
  DFFSR fifo_reg_5__3_ ( .D(n3461), .CLK(wclk), .R(n13138), .S(1'b1), .Q(
        fifo[1095]) );
  DFFSR fifo_reg_5__2_ ( .D(n3462), .CLK(wclk), .R(n13141), .S(1'b1), .Q(
        fifo[1094]) );
  DFFSR fifo_reg_5__1_ ( .D(n3463), .CLK(wclk), .R(n13144), .S(1'b1), .Q(
        fifo[1093]) );
  DFFSR fifo_reg_5__0_ ( .D(n3464), .CLK(wclk), .R(n13146), .S(1'b1), .Q(
        fifo[1092]) );
  DFFSR fifo_reg_6__41_ ( .D(n3465), .CLK(wclk), .R(n13199), .S(1'b1), .Q(
        fifo[1091]) );
  DFFSR fifo_reg_6__40_ ( .D(n3466), .CLK(wclk), .R(n13199), .S(1'b1), .Q(
        fifo[1090]) );
  DFFSR fifo_reg_6__39_ ( .D(n3467), .CLK(wclk), .R(n13199), .S(1'b1), .Q(
        fifo[1089]) );
  DFFSR fifo_reg_6__38_ ( .D(n3468), .CLK(wclk), .R(n13199), .S(1'b1), .Q(
        fifo[1088]) );
  DFFSR fifo_reg_6__37_ ( .D(n3469), .CLK(wclk), .R(n13199), .S(1'b1), .Q(
        fifo[1087]) );
  DFFSR fifo_reg_6__36_ ( .D(n3470), .CLK(wclk), .R(n13199), .S(1'b1), .Q(
        fifo[1086]) );
  DFFSR fifo_reg_6__35_ ( .D(n3471), .CLK(wclk), .R(n13199), .S(1'b1), .Q(
        fifo[1085]) );
  DFFSR fifo_reg_6__34_ ( .D(n3472), .CLK(wclk), .R(n13199), .S(1'b1), .Q(
        fifo[1084]) );
  DFFSR fifo_reg_6__33_ ( .D(n3473), .CLK(wclk), .R(n13200), .S(1'b1), .Q(
        fifo[1083]) );
  DFFSR fifo_reg_6__32_ ( .D(n3474), .CLK(wclk), .R(n13200), .S(1'b1), .Q(
        fifo[1082]) );
  DFFSR fifo_reg_6__31_ ( .D(n3475), .CLK(wclk), .R(n13200), .S(1'b1), .Q(
        fifo[1081]) );
  DFFSR fifo_reg_6__30_ ( .D(n3476), .CLK(wclk), .R(n13200), .S(1'b1), .Q(
        fifo[1080]) );
  DFFSR fifo_reg_6__29_ ( .D(n3477), .CLK(wclk), .R(n13200), .S(1'b1), .Q(
        fifo[1079]) );
  DFFSR fifo_reg_6__28_ ( .D(n3478), .CLK(wclk), .R(n13200), .S(1'b1), .Q(
        fifo[1078]) );
  DFFSR fifo_reg_6__27_ ( .D(n3479), .CLK(wclk), .R(n13200), .S(1'b1), .Q(
        fifo[1077]) );
  DFFSR fifo_reg_6__26_ ( .D(n3480), .CLK(wclk), .R(n13200), .S(1'b1), .Q(
        fifo[1076]) );
  DFFSR fifo_reg_6__25_ ( .D(n3481), .CLK(wclk), .R(n13200), .S(1'b1), .Q(
        fifo[1075]) );
  DFFSR fifo_reg_6__24_ ( .D(n3482), .CLK(wclk), .R(n13200), .S(1'b1), .Q(
        fifo[1074]) );
  DFFSR fifo_reg_6__23_ ( .D(n3483), .CLK(wclk), .R(n13200), .S(1'b1), .Q(
        fifo[1073]) );
  DFFSR fifo_reg_6__22_ ( .D(n3484), .CLK(wclk), .R(n13200), .S(1'b1), .Q(
        fifo[1072]) );
  DFFSR fifo_reg_6__21_ ( .D(n3485), .CLK(wclk), .R(n13201), .S(1'b1), .Q(
        fifo[1071]) );
  DFFSR fifo_reg_6__20_ ( .D(n3486), .CLK(wclk), .R(n13201), .S(1'b1), .Q(
        fifo[1070]) );
  DFFSR fifo_reg_6__19_ ( .D(n3487), .CLK(wclk), .R(n13201), .S(1'b1), .Q(
        fifo[1069]) );
  DFFSR fifo_reg_6__18_ ( .D(n3488), .CLK(wclk), .R(n13201), .S(1'b1), .Q(
        fifo[1068]) );
  DFFSR fifo_reg_6__17_ ( .D(n3489), .CLK(wclk), .R(n13201), .S(1'b1), .Q(
        fifo[1067]) );
  DFFSR fifo_reg_6__16_ ( .D(n3490), .CLK(wclk), .R(n13201), .S(1'b1), .Q(
        fifo[1066]) );
  DFFSR fifo_reg_6__15_ ( .D(n3491), .CLK(wclk), .R(n13105), .S(1'b1), .Q(
        fifo[1065]) );
  DFFSR fifo_reg_6__14_ ( .D(n3492), .CLK(wclk), .R(n13108), .S(1'b1), .Q(
        fifo[1064]) );
  DFFSR fifo_reg_6__13_ ( .D(n3493), .CLK(wclk), .R(n13111), .S(1'b1), .Q(
        fifo[1063]) );
  DFFSR fifo_reg_6__12_ ( .D(n3494), .CLK(wclk), .R(n13113), .S(1'b1), .Q(
        fifo[1062]) );
  DFFSR fifo_reg_6__11_ ( .D(n3495), .CLK(wclk), .R(n13116), .S(1'b1), .Q(
        fifo[1061]) );
  DFFSR fifo_reg_6__10_ ( .D(n3496), .CLK(wclk), .R(n13119), .S(1'b1), .Q(
        fifo[1060]) );
  DFFSR fifo_reg_6__9_ ( .D(n3497), .CLK(wclk), .R(n13122), .S(1'b1), .Q(
        fifo[1059]) );
  DFFSR fifo_reg_6__8_ ( .D(n3498), .CLK(wclk), .R(n13124), .S(1'b1), .Q(
        fifo[1058]) );
  DFFSR fifo_reg_6__7_ ( .D(n3499), .CLK(wclk), .R(n13127), .S(1'b1), .Q(
        fifo[1057]) );
  DFFSR fifo_reg_6__6_ ( .D(n3500), .CLK(wclk), .R(n13130), .S(1'b1), .Q(
        fifo[1056]) );
  DFFSR fifo_reg_6__5_ ( .D(n3501), .CLK(wclk), .R(n13133), .S(1'b1), .Q(
        fifo[1055]) );
  DFFSR fifo_reg_6__4_ ( .D(n3502), .CLK(wclk), .R(n13135), .S(1'b1), .Q(
        fifo[1054]) );
  DFFSR fifo_reg_6__3_ ( .D(n3503), .CLK(wclk), .R(n13138), .S(1'b1), .Q(
        fifo[1053]) );
  DFFSR fifo_reg_6__2_ ( .D(n3504), .CLK(wclk), .R(n13141), .S(1'b1), .Q(
        fifo[1052]) );
  DFFSR fifo_reg_6__1_ ( .D(n3505), .CLK(wclk), .R(n13144), .S(1'b1), .Q(
        fifo[1051]) );
  DFFSR fifo_reg_6__0_ ( .D(n3506), .CLK(wclk), .R(n13146), .S(1'b1), .Q(
        fifo[1050]) );
  DFFSR fifo_reg_7__41_ ( .D(n3507), .CLK(wclk), .R(n13201), .S(1'b1), .Q(
        fifo[1049]) );
  DFFSR fifo_reg_7__40_ ( .D(n3508), .CLK(wclk), .R(n13201), .S(1'b1), .Q(
        fifo[1048]) );
  DFFSR fifo_reg_7__39_ ( .D(n3509), .CLK(wclk), .R(n13201), .S(1'b1), .Q(
        fifo[1047]) );
  DFFSR fifo_reg_7__38_ ( .D(n3510), .CLK(wclk), .R(n13201), .S(1'b1), .Q(
        fifo[1046]) );
  DFFSR fifo_reg_7__37_ ( .D(n3511), .CLK(wclk), .R(n13201), .S(1'b1), .Q(
        fifo[1045]) );
  DFFSR fifo_reg_7__36_ ( .D(n3512), .CLK(wclk), .R(n13201), .S(1'b1), .Q(
        fifo[1044]) );
  DFFSR fifo_reg_7__35_ ( .D(n3513), .CLK(wclk), .R(n13202), .S(1'b1), .Q(
        fifo[1043]) );
  DFFSR fifo_reg_7__34_ ( .D(n3514), .CLK(wclk), .R(n13202), .S(1'b1), .Q(
        fifo[1042]) );
  DFFSR fifo_reg_7__33_ ( .D(n3515), .CLK(wclk), .R(n13202), .S(1'b1), .Q(
        fifo[1041]) );
  DFFSR fifo_reg_7__32_ ( .D(n3516), .CLK(wclk), .R(n13202), .S(1'b1), .Q(
        fifo[1040]) );
  DFFSR fifo_reg_7__31_ ( .D(n3517), .CLK(wclk), .R(n13202), .S(1'b1), .Q(
        fifo[1039]) );
  DFFSR fifo_reg_7__30_ ( .D(n3518), .CLK(wclk), .R(n13202), .S(1'b1), .Q(
        fifo[1038]) );
  DFFSR fifo_reg_7__29_ ( .D(n3519), .CLK(wclk), .R(n13202), .S(1'b1), .Q(
        fifo[1037]) );
  DFFSR fifo_reg_7__28_ ( .D(n3520), .CLK(wclk), .R(n13202), .S(1'b1), .Q(
        fifo[1036]) );
  DFFSR fifo_reg_7__27_ ( .D(n3521), .CLK(wclk), .R(n13202), .S(1'b1), .Q(
        fifo[1035]) );
  DFFSR fifo_reg_7__26_ ( .D(n3522), .CLK(wclk), .R(n13202), .S(1'b1), .Q(
        fifo[1034]) );
  DFFSR fifo_reg_7__25_ ( .D(n3523), .CLK(wclk), .R(n13202), .S(1'b1), .Q(
        fifo[1033]) );
  DFFSR fifo_reg_7__24_ ( .D(n3524), .CLK(wclk), .R(n13202), .S(1'b1), .Q(
        fifo[1032]) );
  DFFSR fifo_reg_7__23_ ( .D(n3525), .CLK(wclk), .R(n13203), .S(1'b1), .Q(
        fifo[1031]) );
  DFFSR fifo_reg_7__22_ ( .D(n3526), .CLK(wclk), .R(n13203), .S(1'b1), .Q(
        fifo[1030]) );
  DFFSR fifo_reg_7__21_ ( .D(n3527), .CLK(wclk), .R(n13203), .S(1'b1), .Q(
        fifo[1029]) );
  DFFSR fifo_reg_7__20_ ( .D(n3528), .CLK(wclk), .R(n13203), .S(1'b1), .Q(
        fifo[1028]) );
  DFFSR fifo_reg_7__19_ ( .D(n3529), .CLK(wclk), .R(n13203), .S(1'b1), .Q(
        fifo[1027]) );
  DFFSR fifo_reg_7__18_ ( .D(n3530), .CLK(wclk), .R(n13203), .S(1'b1), .Q(
        fifo[1026]) );
  DFFSR fifo_reg_7__17_ ( .D(n3531), .CLK(wclk), .R(n13203), .S(1'b1), .Q(
        fifo[1025]) );
  DFFSR fifo_reg_7__16_ ( .D(n3532), .CLK(wclk), .R(n13203), .S(1'b1), .Q(
        fifo[1024]) );
  DFFSR fifo_reg_7__15_ ( .D(n3533), .CLK(wclk), .R(n13105), .S(1'b1), .Q(
        fifo[1023]) );
  DFFSR fifo_reg_7__14_ ( .D(n3534), .CLK(wclk), .R(n13108), .S(1'b1), .Q(
        fifo[1022]) );
  DFFSR fifo_reg_7__13_ ( .D(n3535), .CLK(wclk), .R(n13111), .S(1'b1), .Q(
        fifo[1021]) );
  DFFSR fifo_reg_7__12_ ( .D(n3536), .CLK(wclk), .R(n13113), .S(1'b1), .Q(
        fifo[1020]) );
  DFFSR fifo_reg_7__11_ ( .D(n3537), .CLK(wclk), .R(n13116), .S(1'b1), .Q(
        fifo[1019]) );
  DFFSR fifo_reg_7__10_ ( .D(n3538), .CLK(wclk), .R(n13119), .S(1'b1), .Q(
        fifo[1018]) );
  DFFSR fifo_reg_7__9_ ( .D(n3539), .CLK(wclk), .R(n13122), .S(1'b1), .Q(
        fifo[1017]) );
  DFFSR fifo_reg_7__8_ ( .D(n3540), .CLK(wclk), .R(n13124), .S(1'b1), .Q(
        fifo[1016]) );
  DFFSR fifo_reg_7__7_ ( .D(n3541), .CLK(wclk), .R(n13127), .S(1'b1), .Q(
        fifo[1015]) );
  DFFSR fifo_reg_7__6_ ( .D(n3542), .CLK(wclk), .R(n13130), .S(1'b1), .Q(
        fifo[1014]) );
  DFFSR fifo_reg_7__5_ ( .D(n3543), .CLK(wclk), .R(n13133), .S(1'b1), .Q(
        fifo[1013]) );
  DFFSR fifo_reg_7__4_ ( .D(n3544), .CLK(wclk), .R(n13135), .S(1'b1), .Q(
        fifo[1012]) );
  DFFSR fifo_reg_7__3_ ( .D(n3545), .CLK(wclk), .R(n13138), .S(1'b1), .Q(
        fifo[1011]) );
  DFFSR fifo_reg_7__2_ ( .D(n3546), .CLK(wclk), .R(n13141), .S(1'b1), .Q(
        fifo[1010]) );
  DFFSR fifo_reg_7__1_ ( .D(n3547), .CLK(wclk), .R(n13144), .S(1'b1), .Q(
        fifo[1009]) );
  DFFSR fifo_reg_7__0_ ( .D(n3548), .CLK(wclk), .R(n13146), .S(1'b1), .Q(
        fifo[1008]) );
  DFFSR fifo_reg_8__41_ ( .D(n3549), .CLK(wclk), .R(n13203), .S(1'b1), .Q(
        fifo[1007]) );
  DFFSR fifo_reg_8__40_ ( .D(n3550), .CLK(wclk), .R(n13203), .S(1'b1), .Q(
        fifo[1006]) );
  DFFSR fifo_reg_8__39_ ( .D(n3551), .CLK(wclk), .R(n13203), .S(1'b1), .Q(
        fifo[1005]) );
  DFFSR fifo_reg_8__38_ ( .D(n3552), .CLK(wclk), .R(n13203), .S(1'b1), .Q(
        fifo[1004]) );
  DFFSR fifo_reg_8__37_ ( .D(n3553), .CLK(wclk), .R(n13204), .S(1'b1), .Q(
        fifo[1003]) );
  DFFSR fifo_reg_8__36_ ( .D(n3554), .CLK(wclk), .R(n13204), .S(1'b1), .Q(
        fifo[1002]) );
  DFFSR fifo_reg_8__35_ ( .D(n3555), .CLK(wclk), .R(n13204), .S(1'b1), .Q(
        fifo[1001]) );
  DFFSR fifo_reg_8__34_ ( .D(n3556), .CLK(wclk), .R(n13204), .S(1'b1), .Q(
        fifo[1000]) );
  DFFSR fifo_reg_8__33_ ( .D(n3557), .CLK(wclk), .R(n13204), .S(1'b1), .Q(
        fifo[999]) );
  DFFSR fifo_reg_8__32_ ( .D(n3558), .CLK(wclk), .R(n13204), .S(1'b1), .Q(
        fifo[998]) );
  DFFSR fifo_reg_8__31_ ( .D(n3559), .CLK(wclk), .R(n13204), .S(1'b1), .Q(
        fifo[997]) );
  DFFSR fifo_reg_8__30_ ( .D(n3560), .CLK(wclk), .R(n13204), .S(1'b1), .Q(
        fifo[996]) );
  DFFSR fifo_reg_8__29_ ( .D(n3561), .CLK(wclk), .R(n13204), .S(1'b1), .Q(
        fifo[995]) );
  DFFSR fifo_reg_8__28_ ( .D(n3562), .CLK(wclk), .R(n13204), .S(1'b1), .Q(
        fifo[994]) );
  DFFSR fifo_reg_8__27_ ( .D(n3563), .CLK(wclk), .R(n13204), .S(1'b1), .Q(
        fifo[993]) );
  DFFSR fifo_reg_8__26_ ( .D(n3564), .CLK(wclk), .R(n13204), .S(1'b1), .Q(
        fifo[992]) );
  DFFSR fifo_reg_8__25_ ( .D(n3565), .CLK(wclk), .R(n13205), .S(1'b1), .Q(
        fifo[991]) );
  DFFSR fifo_reg_8__24_ ( .D(n3566), .CLK(wclk), .R(n13205), .S(1'b1), .Q(
        fifo[990]) );
  DFFSR fifo_reg_8__23_ ( .D(n3567), .CLK(wclk), .R(n13205), .S(1'b1), .Q(
        fifo[989]) );
  DFFSR fifo_reg_8__22_ ( .D(n3568), .CLK(wclk), .R(n13205), .S(1'b1), .Q(
        fifo[988]) );
  DFFSR fifo_reg_8__21_ ( .D(n3569), .CLK(wclk), .R(n13205), .S(1'b1), .Q(
        fifo[987]) );
  DFFSR fifo_reg_8__20_ ( .D(n3570), .CLK(wclk), .R(n13205), .S(1'b1), .Q(
        fifo[986]) );
  DFFSR fifo_reg_8__19_ ( .D(n3571), .CLK(wclk), .R(n13205), .S(1'b1), .Q(
        fifo[985]) );
  DFFSR fifo_reg_8__18_ ( .D(n3572), .CLK(wclk), .R(n13205), .S(1'b1), .Q(
        fifo[984]) );
  DFFSR fifo_reg_8__17_ ( .D(n3573), .CLK(wclk), .R(n13205), .S(1'b1), .Q(
        fifo[983]) );
  DFFSR fifo_reg_8__16_ ( .D(n3574), .CLK(wclk), .R(n13205), .S(1'b1), .Q(
        fifo[982]) );
  DFFSR fifo_reg_8__15_ ( .D(n3575), .CLK(wclk), .R(n13105), .S(1'b1), .Q(
        fifo[981]) );
  DFFSR fifo_reg_8__14_ ( .D(n3576), .CLK(wclk), .R(n13108), .S(1'b1), .Q(
        fifo[980]) );
  DFFSR fifo_reg_8__13_ ( .D(n3577), .CLK(wclk), .R(n13111), .S(1'b1), .Q(
        fifo[979]) );
  DFFSR fifo_reg_8__12_ ( .D(n3578), .CLK(wclk), .R(n13114), .S(1'b1), .Q(
        fifo[978]) );
  DFFSR fifo_reg_8__11_ ( .D(n3579), .CLK(wclk), .R(n13116), .S(1'b1), .Q(
        fifo[977]) );
  DFFSR fifo_reg_8__10_ ( .D(n3580), .CLK(wclk), .R(n13119), .S(1'b1), .Q(
        fifo[976]) );
  DFFSR fifo_reg_8__9_ ( .D(n3581), .CLK(wclk), .R(n13122), .S(1'b1), .Q(
        fifo[975]) );
  DFFSR fifo_reg_8__8_ ( .D(n3582), .CLK(wclk), .R(n13125), .S(1'b1), .Q(
        fifo[974]) );
  DFFSR fifo_reg_8__7_ ( .D(n3583), .CLK(wclk), .R(n13127), .S(1'b1), .Q(
        fifo[973]) );
  DFFSR fifo_reg_8__6_ ( .D(n3584), .CLK(wclk), .R(n13130), .S(1'b1), .Q(
        fifo[972]) );
  DFFSR fifo_reg_8__5_ ( .D(n3585), .CLK(wclk), .R(n13133), .S(1'b1), .Q(
        fifo[971]) );
  DFFSR fifo_reg_8__4_ ( .D(n3586), .CLK(wclk), .R(n13136), .S(1'b1), .Q(
        fifo[970]) );
  DFFSR fifo_reg_8__3_ ( .D(n3587), .CLK(wclk), .R(n13138), .S(1'b1), .Q(
        fifo[969]) );
  DFFSR fifo_reg_8__2_ ( .D(n3588), .CLK(wclk), .R(n13141), .S(1'b1), .Q(
        fifo[968]) );
  DFFSR fifo_reg_8__1_ ( .D(n3589), .CLK(wclk), .R(n13144), .S(1'b1), .Q(
        fifo[967]) );
  DFFSR fifo_reg_8__0_ ( .D(n3590), .CLK(wclk), .R(n13147), .S(1'b1), .Q(
        fifo[966]) );
  DFFSR fifo_reg_9__41_ ( .D(n3591), .CLK(wclk), .R(n13205), .S(1'b1), .Q(
        fifo[965]) );
  DFFSR fifo_reg_9__40_ ( .D(n3592), .CLK(wclk), .R(n13205), .S(1'b1), .Q(
        fifo[964]) );
  DFFSR fifo_reg_9__39_ ( .D(n3593), .CLK(wclk), .R(n13206), .S(1'b1), .Q(
        fifo[963]) );
  DFFSR fifo_reg_9__38_ ( .D(n3594), .CLK(wclk), .R(n13206), .S(1'b1), .Q(
        fifo[962]) );
  DFFSR fifo_reg_9__37_ ( .D(n3595), .CLK(wclk), .R(n13206), .S(1'b1), .Q(
        fifo[961]) );
  DFFSR fifo_reg_9__36_ ( .D(n3596), .CLK(wclk), .R(n13206), .S(1'b1), .Q(
        fifo[960]) );
  DFFSR fifo_reg_9__35_ ( .D(n3597), .CLK(wclk), .R(n13206), .S(1'b1), .Q(
        fifo[959]) );
  DFFSR fifo_reg_9__34_ ( .D(n3598), .CLK(wclk), .R(n13206), .S(1'b1), .Q(
        fifo[958]) );
  DFFSR fifo_reg_9__33_ ( .D(n3599), .CLK(wclk), .R(n13206), .S(1'b1), .Q(
        fifo[957]) );
  DFFSR fifo_reg_9__32_ ( .D(n3600), .CLK(wclk), .R(n13206), .S(1'b1), .Q(
        fifo[956]) );
  DFFSR fifo_reg_9__31_ ( .D(n3601), .CLK(wclk), .R(n13206), .S(1'b1), .Q(
        fifo[955]) );
  DFFSR fifo_reg_9__30_ ( .D(n3602), .CLK(wclk), .R(n13206), .S(1'b1), .Q(
        fifo[954]) );
  DFFSR fifo_reg_9__29_ ( .D(n3603), .CLK(wclk), .R(n13206), .S(1'b1), .Q(
        fifo[953]) );
  DFFSR fifo_reg_9__28_ ( .D(n3604), .CLK(wclk), .R(n13206), .S(1'b1), .Q(
        fifo[952]) );
  DFFSR fifo_reg_9__27_ ( .D(n3605), .CLK(wclk), .R(n13207), .S(1'b1), .Q(
        fifo[951]) );
  DFFSR fifo_reg_9__26_ ( .D(n3606), .CLK(wclk), .R(n13207), .S(1'b1), .Q(
        fifo[950]) );
  DFFSR fifo_reg_9__25_ ( .D(n3607), .CLK(wclk), .R(n13207), .S(1'b1), .Q(
        fifo[949]) );
  DFFSR fifo_reg_9__24_ ( .D(n3608), .CLK(wclk), .R(n13207), .S(1'b1), .Q(
        fifo[948]) );
  DFFSR fifo_reg_9__23_ ( .D(n3609), .CLK(wclk), .R(n13207), .S(1'b1), .Q(
        fifo[947]) );
  DFFSR fifo_reg_9__22_ ( .D(n3610), .CLK(wclk), .R(n13207), .S(1'b1), .Q(
        fifo[946]) );
  DFFSR fifo_reg_9__21_ ( .D(n3611), .CLK(wclk), .R(n13207), .S(1'b1), .Q(
        fifo[945]) );
  DFFSR fifo_reg_9__20_ ( .D(n3612), .CLK(wclk), .R(n13207), .S(1'b1), .Q(
        fifo[944]) );
  DFFSR fifo_reg_9__19_ ( .D(n3613), .CLK(wclk), .R(n13207), .S(1'b1), .Q(
        fifo[943]) );
  DFFSR fifo_reg_9__18_ ( .D(n3614), .CLK(wclk), .R(n13207), .S(1'b1), .Q(
        fifo[942]) );
  DFFSR fifo_reg_9__17_ ( .D(n3615), .CLK(wclk), .R(n13207), .S(1'b1), .Q(
        fifo[941]) );
  DFFSR fifo_reg_9__16_ ( .D(n3616), .CLK(wclk), .R(n13207), .S(1'b1), .Q(
        fifo[940]) );
  DFFSR fifo_reg_9__15_ ( .D(n3617), .CLK(wclk), .R(n13105), .S(1'b1), .Q(
        fifo[939]) );
  DFFSR fifo_reg_9__14_ ( .D(n3618), .CLK(wclk), .R(n13108), .S(1'b1), .Q(
        fifo[938]) );
  DFFSR fifo_reg_9__13_ ( .D(n3619), .CLK(wclk), .R(n13111), .S(1'b1), .Q(
        fifo[937]) );
  DFFSR fifo_reg_9__12_ ( .D(n3620), .CLK(wclk), .R(n13114), .S(1'b1), .Q(
        fifo[936]) );
  DFFSR fifo_reg_9__11_ ( .D(n3621), .CLK(wclk), .R(n13116), .S(1'b1), .Q(
        fifo[935]) );
  DFFSR fifo_reg_9__10_ ( .D(n3622), .CLK(wclk), .R(n13119), .S(1'b1), .Q(
        fifo[934]) );
  DFFSR fifo_reg_9__9_ ( .D(n3623), .CLK(wclk), .R(n13122), .S(1'b1), .Q(
        fifo[933]) );
  DFFSR fifo_reg_9__8_ ( .D(n3624), .CLK(wclk), .R(n13125), .S(1'b1), .Q(
        fifo[932]) );
  DFFSR fifo_reg_9__7_ ( .D(n3625), .CLK(wclk), .R(n13127), .S(1'b1), .Q(
        fifo[931]) );
  DFFSR fifo_reg_9__6_ ( .D(n3626), .CLK(wclk), .R(n13130), .S(1'b1), .Q(
        fifo[930]) );
  DFFSR fifo_reg_9__5_ ( .D(n3627), .CLK(wclk), .R(n13133), .S(1'b1), .Q(
        fifo[929]) );
  DFFSR fifo_reg_9__4_ ( .D(n3628), .CLK(wclk), .R(n13136), .S(1'b1), .Q(
        fifo[928]) );
  DFFSR fifo_reg_9__3_ ( .D(n3629), .CLK(wclk), .R(n13138), .S(1'b1), .Q(
        fifo[927]) );
  DFFSR fifo_reg_9__2_ ( .D(n3630), .CLK(wclk), .R(n13141), .S(1'b1), .Q(
        fifo[926]) );
  DFFSR fifo_reg_9__1_ ( .D(n3631), .CLK(wclk), .R(n13144), .S(1'b1), .Q(
        fifo[925]) );
  DFFSR fifo_reg_9__0_ ( .D(n3632), .CLK(wclk), .R(n13147), .S(1'b1), .Q(
        fifo[924]) );
  DFFSR fifo_reg_10__41_ ( .D(n3633), .CLK(wclk), .R(n13208), .S(1'b1), .Q(
        fifo[923]) );
  DFFSR fifo_reg_10__40_ ( .D(n3634), .CLK(wclk), .R(n13208), .S(1'b1), .Q(
        fifo[922]) );
  DFFSR fifo_reg_10__39_ ( .D(n3635), .CLK(wclk), .R(n13208), .S(1'b1), .Q(
        fifo[921]) );
  DFFSR fifo_reg_10__38_ ( .D(n3636), .CLK(wclk), .R(n13208), .S(1'b1), .Q(
        fifo[920]) );
  DFFSR fifo_reg_10__37_ ( .D(n3637), .CLK(wclk), .R(n13208), .S(1'b1), .Q(
        fifo[919]) );
  DFFSR fifo_reg_10__36_ ( .D(n3638), .CLK(wclk), .R(n13208), .S(1'b1), .Q(
        fifo[918]) );
  DFFSR fifo_reg_10__35_ ( .D(n3639), .CLK(wclk), .R(n13208), .S(1'b1), .Q(
        fifo[917]) );
  DFFSR fifo_reg_10__34_ ( .D(n3640), .CLK(wclk), .R(n13208), .S(1'b1), .Q(
        fifo[916]) );
  DFFSR fifo_reg_10__33_ ( .D(n3641), .CLK(wclk), .R(n13208), .S(1'b1), .Q(
        fifo[915]) );
  DFFSR fifo_reg_10__32_ ( .D(n3642), .CLK(wclk), .R(n13208), .S(1'b1), .Q(
        fifo[914]) );
  DFFSR fifo_reg_10__31_ ( .D(n3643), .CLK(wclk), .R(n13208), .S(1'b1), .Q(
        fifo[913]) );
  DFFSR fifo_reg_10__30_ ( .D(n3644), .CLK(wclk), .R(n13208), .S(1'b1), .Q(
        fifo[912]) );
  DFFSR fifo_reg_10__29_ ( .D(n3645), .CLK(wclk), .R(n13209), .S(1'b1), .Q(
        fifo[911]) );
  DFFSR fifo_reg_10__28_ ( .D(n3646), .CLK(wclk), .R(n13209), .S(1'b1), .Q(
        fifo[910]) );
  DFFSR fifo_reg_10__27_ ( .D(n3647), .CLK(wclk), .R(n13209), .S(1'b1), .Q(
        fifo[909]) );
  DFFSR fifo_reg_10__26_ ( .D(n3648), .CLK(wclk), .R(n13209), .S(1'b1), .Q(
        fifo[908]) );
  DFFSR fifo_reg_10__25_ ( .D(n3649), .CLK(wclk), .R(n13209), .S(1'b1), .Q(
        fifo[907]) );
  DFFSR fifo_reg_10__24_ ( .D(n3650), .CLK(wclk), .R(n13209), .S(1'b1), .Q(
        fifo[906]) );
  DFFSR fifo_reg_10__23_ ( .D(n3651), .CLK(wclk), .R(n13209), .S(1'b1), .Q(
        fifo[905]) );
  DFFSR fifo_reg_10__22_ ( .D(n3652), .CLK(wclk), .R(n13209), .S(1'b1), .Q(
        fifo[904]) );
  DFFSR fifo_reg_10__21_ ( .D(n3653), .CLK(wclk), .R(n13209), .S(1'b1), .Q(
        fifo[903]) );
  DFFSR fifo_reg_10__20_ ( .D(n3654), .CLK(wclk), .R(n13209), .S(1'b1), .Q(
        fifo[902]) );
  DFFSR fifo_reg_10__19_ ( .D(n3655), .CLK(wclk), .R(n13209), .S(1'b1), .Q(
        fifo[901]) );
  DFFSR fifo_reg_10__18_ ( .D(n3656), .CLK(wclk), .R(n13209), .S(1'b1), .Q(
        fifo[900]) );
  DFFSR fifo_reg_10__17_ ( .D(n3657), .CLK(wclk), .R(n13210), .S(1'b1), .Q(
        fifo[899]) );
  DFFSR fifo_reg_10__16_ ( .D(n3658), .CLK(wclk), .R(n13210), .S(1'b1), .Q(
        fifo[898]) );
  DFFSR fifo_reg_10__15_ ( .D(n3659), .CLK(wclk), .R(n13105), .S(1'b1), .Q(
        fifo[897]) );
  DFFSR fifo_reg_10__14_ ( .D(n3660), .CLK(wclk), .R(n13108), .S(1'b1), .Q(
        fifo[896]) );
  DFFSR fifo_reg_10__13_ ( .D(n3661), .CLK(wclk), .R(n13111), .S(1'b1), .Q(
        fifo[895]) );
  DFFSR fifo_reg_10__12_ ( .D(n3662), .CLK(wclk), .R(n13114), .S(1'b1), .Q(
        fifo[894]) );
  DFFSR fifo_reg_10__11_ ( .D(n3663), .CLK(wclk), .R(n13116), .S(1'b1), .Q(
        fifo[893]) );
  DFFSR fifo_reg_10__10_ ( .D(n3664), .CLK(wclk), .R(n13119), .S(1'b1), .Q(
        fifo[892]) );
  DFFSR fifo_reg_10__9_ ( .D(n3665), .CLK(wclk), .R(n13122), .S(1'b1), .Q(
        fifo[891]) );
  DFFSR fifo_reg_10__8_ ( .D(n3666), .CLK(wclk), .R(n13125), .S(1'b1), .Q(
        fifo[890]) );
  DFFSR fifo_reg_10__7_ ( .D(n3667), .CLK(wclk), .R(n13127), .S(1'b1), .Q(
        fifo[889]) );
  DFFSR fifo_reg_10__6_ ( .D(n3668), .CLK(wclk), .R(n13130), .S(1'b1), .Q(
        fifo[888]) );
  DFFSR fifo_reg_10__5_ ( .D(n3669), .CLK(wclk), .R(n13133), .S(1'b1), .Q(
        fifo[887]) );
  DFFSR fifo_reg_10__4_ ( .D(n3670), .CLK(wclk), .R(n13136), .S(1'b1), .Q(
        fifo[886]) );
  DFFSR fifo_reg_10__3_ ( .D(n3671), .CLK(wclk), .R(n13138), .S(1'b1), .Q(
        fifo[885]) );
  DFFSR fifo_reg_10__2_ ( .D(n3672), .CLK(wclk), .R(n13141), .S(1'b1), .Q(
        fifo[884]) );
  DFFSR fifo_reg_10__1_ ( .D(n3673), .CLK(wclk), .R(n13144), .S(1'b1), .Q(
        fifo[883]) );
  DFFSR fifo_reg_10__0_ ( .D(n3674), .CLK(wclk), .R(n13147), .S(1'b1), .Q(
        fifo[882]) );
  DFFSR fifo_reg_11__41_ ( .D(n3675), .CLK(wclk), .R(n13210), .S(1'b1), .Q(
        fifo[881]) );
  DFFSR fifo_reg_11__40_ ( .D(n3676), .CLK(wclk), .R(n13210), .S(1'b1), .Q(
        fifo[880]) );
  DFFSR fifo_reg_11__39_ ( .D(n3677), .CLK(wclk), .R(n13210), .S(1'b1), .Q(
        fifo[879]) );
  DFFSR fifo_reg_11__38_ ( .D(n3678), .CLK(wclk), .R(n13210), .S(1'b1), .Q(
        fifo[878]) );
  DFFSR fifo_reg_11__37_ ( .D(n3679), .CLK(wclk), .R(n13210), .S(1'b1), .Q(
        fifo[877]) );
  DFFSR fifo_reg_11__36_ ( .D(n3680), .CLK(wclk), .R(n13210), .S(1'b1), .Q(
        fifo[876]) );
  DFFSR fifo_reg_11__35_ ( .D(n3681), .CLK(wclk), .R(n13210), .S(1'b1), .Q(
        fifo[875]) );
  DFFSR fifo_reg_11__34_ ( .D(n3682), .CLK(wclk), .R(n13210), .S(1'b1), .Q(
        fifo[874]) );
  DFFSR fifo_reg_11__33_ ( .D(n3683), .CLK(wclk), .R(n13210), .S(1'b1), .Q(
        fifo[873]) );
  DFFSR fifo_reg_11__32_ ( .D(n3684), .CLK(wclk), .R(n13210), .S(1'b1), .Q(
        fifo[872]) );
  DFFSR fifo_reg_11__31_ ( .D(n3685), .CLK(wclk), .R(n13211), .S(1'b1), .Q(
        fifo[871]) );
  DFFSR fifo_reg_11__30_ ( .D(n3686), .CLK(wclk), .R(n13211), .S(1'b1), .Q(
        fifo[870]) );
  DFFSR fifo_reg_11__29_ ( .D(n3687), .CLK(wclk), .R(n13211), .S(1'b1), .Q(
        fifo[869]) );
  DFFSR fifo_reg_11__28_ ( .D(n3688), .CLK(wclk), .R(n13211), .S(1'b1), .Q(
        fifo[868]) );
  DFFSR fifo_reg_11__27_ ( .D(n3689), .CLK(wclk), .R(n13211), .S(1'b1), .Q(
        fifo[867]) );
  DFFSR fifo_reg_11__26_ ( .D(n3690), .CLK(wclk), .R(n13211), .S(1'b1), .Q(
        fifo[866]) );
  DFFSR fifo_reg_11__25_ ( .D(n3691), .CLK(wclk), .R(n13211), .S(1'b1), .Q(
        fifo[865]) );
  DFFSR fifo_reg_11__24_ ( .D(n3692), .CLK(wclk), .R(n13211), .S(1'b1), .Q(
        fifo[864]) );
  DFFSR fifo_reg_11__23_ ( .D(n3693), .CLK(wclk), .R(n13211), .S(1'b1), .Q(
        fifo[863]) );
  DFFSR fifo_reg_11__22_ ( .D(n3694), .CLK(wclk), .R(n13211), .S(1'b1), .Q(
        fifo[862]) );
  DFFSR fifo_reg_11__21_ ( .D(n3695), .CLK(wclk), .R(n13211), .S(1'b1), .Q(
        fifo[861]) );
  DFFSR fifo_reg_11__20_ ( .D(n3696), .CLK(wclk), .R(n13211), .S(1'b1), .Q(
        fifo[860]) );
  DFFSR fifo_reg_11__19_ ( .D(n3697), .CLK(wclk), .R(n13212), .S(1'b1), .Q(
        fifo[859]) );
  DFFSR fifo_reg_11__18_ ( .D(n3698), .CLK(wclk), .R(n13212), .S(1'b1), .Q(
        fifo[858]) );
  DFFSR fifo_reg_11__17_ ( .D(n3699), .CLK(wclk), .R(n13212), .S(1'b1), .Q(
        fifo[857]) );
  DFFSR fifo_reg_11__16_ ( .D(n3700), .CLK(wclk), .R(n13212), .S(1'b1), .Q(
        fifo[856]) );
  DFFSR fifo_reg_11__15_ ( .D(n3701), .CLK(wclk), .R(n13106), .S(1'b1), .Q(
        fifo[855]) );
  DFFSR fifo_reg_11__14_ ( .D(n3702), .CLK(wclk), .R(n13108), .S(1'b1), .Q(
        fifo[854]) );
  DFFSR fifo_reg_11__13_ ( .D(n3703), .CLK(wclk), .R(n13111), .S(1'b1), .Q(
        fifo[853]) );
  DFFSR fifo_reg_11__12_ ( .D(n3704), .CLK(wclk), .R(n13114), .S(1'b1), .Q(
        fifo[852]) );
  DFFSR fifo_reg_11__11_ ( .D(n3705), .CLK(wclk), .R(n13117), .S(1'b1), .Q(
        fifo[851]) );
  DFFSR fifo_reg_11__10_ ( .D(n3706), .CLK(wclk), .R(n13119), .S(1'b1), .Q(
        fifo[850]) );
  DFFSR fifo_reg_11__9_ ( .D(n3707), .CLK(wclk), .R(n13122), .S(1'b1), .Q(
        fifo[849]) );
  DFFSR fifo_reg_11__8_ ( .D(n3708), .CLK(wclk), .R(n13125), .S(1'b1), .Q(
        fifo[848]) );
  DFFSR fifo_reg_11__7_ ( .D(n3709), .CLK(wclk), .R(n13128), .S(1'b1), .Q(
        fifo[847]) );
  DFFSR fifo_reg_11__6_ ( .D(n3710), .CLK(wclk), .R(n13130), .S(1'b1), .Q(
        fifo[846]) );
  DFFSR fifo_reg_11__5_ ( .D(n3711), .CLK(wclk), .R(n13133), .S(1'b1), .Q(
        fifo[845]) );
  DFFSR fifo_reg_11__4_ ( .D(n3712), .CLK(wclk), .R(n13136), .S(1'b1), .Q(
        fifo[844]) );
  DFFSR fifo_reg_11__3_ ( .D(n3713), .CLK(wclk), .R(n13139), .S(1'b1), .Q(
        fifo[843]) );
  DFFSR fifo_reg_11__2_ ( .D(n3714), .CLK(wclk), .R(n13141), .S(1'b1), .Q(
        fifo[842]) );
  DFFSR fifo_reg_11__1_ ( .D(n3715), .CLK(wclk), .R(n13144), .S(1'b1), .Q(
        fifo[841]) );
  DFFSR fifo_reg_11__0_ ( .D(n3716), .CLK(wclk), .R(n13147), .S(1'b1), .Q(
        fifo[840]) );
  DFFSR fifo_reg_12__41_ ( .D(n3717), .CLK(wclk), .R(n13212), .S(1'b1), .Q(
        fifo[839]) );
  DFFSR fifo_reg_12__40_ ( .D(n3718), .CLK(wclk), .R(n13212), .S(1'b1), .Q(
        fifo[838]) );
  DFFSR fifo_reg_12__39_ ( .D(n3719), .CLK(wclk), .R(n13212), .S(1'b1), .Q(
        fifo[837]) );
  DFFSR fifo_reg_12__38_ ( .D(n3720), .CLK(wclk), .R(n13212), .S(1'b1), .Q(
        fifo[836]) );
  DFFSR fifo_reg_12__37_ ( .D(n3721), .CLK(wclk), .R(n13212), .S(1'b1), .Q(
        fifo[835]) );
  DFFSR fifo_reg_12__36_ ( .D(n3722), .CLK(wclk), .R(n13212), .S(1'b1), .Q(
        fifo[834]) );
  DFFSR fifo_reg_12__35_ ( .D(n3723), .CLK(wclk), .R(n13212), .S(1'b1), .Q(
        fifo[833]) );
  DFFSR fifo_reg_12__34_ ( .D(n3724), .CLK(wclk), .R(n13212), .S(1'b1), .Q(
        fifo[832]) );
  DFFSR fifo_reg_12__33_ ( .D(n3725), .CLK(wclk), .R(n13213), .S(1'b1), .Q(
        fifo[831]) );
  DFFSR fifo_reg_12__32_ ( .D(n3726), .CLK(wclk), .R(n13213), .S(1'b1), .Q(
        fifo[830]) );
  DFFSR fifo_reg_12__31_ ( .D(n3727), .CLK(wclk), .R(n13213), .S(1'b1), .Q(
        fifo[829]) );
  DFFSR fifo_reg_12__30_ ( .D(n3728), .CLK(wclk), .R(n13213), .S(1'b1), .Q(
        fifo[828]) );
  DFFSR fifo_reg_12__29_ ( .D(n3729), .CLK(wclk), .R(n13213), .S(1'b1), .Q(
        fifo[827]) );
  DFFSR fifo_reg_12__28_ ( .D(n3730), .CLK(wclk), .R(n13213), .S(1'b1), .Q(
        fifo[826]) );
  DFFSR fifo_reg_12__27_ ( .D(n3731), .CLK(wclk), .R(n13213), .S(1'b1), .Q(
        fifo[825]) );
  DFFSR fifo_reg_12__26_ ( .D(n3732), .CLK(wclk), .R(n13213), .S(1'b1), .Q(
        fifo[824]) );
  DFFSR fifo_reg_12__25_ ( .D(n3733), .CLK(wclk), .R(n13213), .S(1'b1), .Q(
        fifo[823]) );
  DFFSR fifo_reg_12__24_ ( .D(n3734), .CLK(wclk), .R(n13213), .S(1'b1), .Q(
        fifo[822]) );
  DFFSR fifo_reg_12__23_ ( .D(n3735), .CLK(wclk), .R(n13213), .S(1'b1), .Q(
        fifo[821]) );
  DFFSR fifo_reg_12__22_ ( .D(n3736), .CLK(wclk), .R(n13213), .S(1'b1), .Q(
        fifo[820]) );
  DFFSR fifo_reg_12__21_ ( .D(n3737), .CLK(wclk), .R(n13214), .S(1'b1), .Q(
        fifo[819]) );
  DFFSR fifo_reg_12__20_ ( .D(n3738), .CLK(wclk), .R(n13214), .S(1'b1), .Q(
        fifo[818]) );
  DFFSR fifo_reg_12__19_ ( .D(n3739), .CLK(wclk), .R(n13214), .S(1'b1), .Q(
        fifo[817]) );
  DFFSR fifo_reg_12__18_ ( .D(n3740), .CLK(wclk), .R(n13214), .S(1'b1), .Q(
        fifo[816]) );
  DFFSR fifo_reg_12__17_ ( .D(n3741), .CLK(wclk), .R(n13214), .S(1'b1), .Q(
        fifo[815]) );
  DFFSR fifo_reg_12__16_ ( .D(n3742), .CLK(wclk), .R(n13214), .S(1'b1), .Q(
        fifo[814]) );
  DFFSR fifo_reg_12__15_ ( .D(n3743), .CLK(wclk), .R(n13106), .S(1'b1), .Q(
        fifo[813]) );
  DFFSR fifo_reg_12__14_ ( .D(n3744), .CLK(wclk), .R(n13108), .S(1'b1), .Q(
        fifo[812]) );
  DFFSR fifo_reg_12__13_ ( .D(n3745), .CLK(wclk), .R(n13111), .S(1'b1), .Q(
        fifo[811]) );
  DFFSR fifo_reg_12__12_ ( .D(n3746), .CLK(wclk), .R(n13114), .S(1'b1), .Q(
        fifo[810]) );
  DFFSR fifo_reg_12__11_ ( .D(n3747), .CLK(wclk), .R(n13117), .S(1'b1), .Q(
        fifo[809]) );
  DFFSR fifo_reg_12__10_ ( .D(n3748), .CLK(wclk), .R(n13119), .S(1'b1), .Q(
        fifo[808]) );
  DFFSR fifo_reg_12__9_ ( .D(n3749), .CLK(wclk), .R(n13122), .S(1'b1), .Q(
        fifo[807]) );
  DFFSR fifo_reg_12__8_ ( .D(n3750), .CLK(wclk), .R(n13125), .S(1'b1), .Q(
        fifo[806]) );
  DFFSR fifo_reg_12__7_ ( .D(n3751), .CLK(wclk), .R(n13128), .S(1'b1), .Q(
        fifo[805]) );
  DFFSR fifo_reg_12__6_ ( .D(n3752), .CLK(wclk), .R(n13130), .S(1'b1), .Q(
        fifo[804]) );
  DFFSR fifo_reg_12__5_ ( .D(n3753), .CLK(wclk), .R(n13133), .S(1'b1), .Q(
        fifo[803]) );
  DFFSR fifo_reg_12__4_ ( .D(n3754), .CLK(wclk), .R(n13136), .S(1'b1), .Q(
        fifo[802]) );
  DFFSR fifo_reg_12__3_ ( .D(n3755), .CLK(wclk), .R(n13139), .S(1'b1), .Q(
        fifo[801]) );
  DFFSR fifo_reg_12__2_ ( .D(n3756), .CLK(wclk), .R(n13141), .S(1'b1), .Q(
        fifo[800]) );
  DFFSR fifo_reg_12__1_ ( .D(n3757), .CLK(wclk), .R(n13144), .S(1'b1), .Q(
        fifo[799]) );
  DFFSR fifo_reg_12__0_ ( .D(n3758), .CLK(wclk), .R(n13147), .S(1'b1), .Q(
        fifo[798]) );
  DFFSR fifo_reg_13__41_ ( .D(n3759), .CLK(wclk), .R(n13214), .S(1'b1), .Q(
        fifo[797]) );
  DFFSR fifo_reg_13__40_ ( .D(n3760), .CLK(wclk), .R(n13214), .S(1'b1), .Q(
        fifo[796]) );
  DFFSR fifo_reg_13__39_ ( .D(n3761), .CLK(wclk), .R(n13214), .S(1'b1), .Q(
        fifo[795]) );
  DFFSR fifo_reg_13__38_ ( .D(n3762), .CLK(wclk), .R(n13214), .S(1'b1), .Q(
        fifo[794]) );
  DFFSR fifo_reg_13__37_ ( .D(n3763), .CLK(wclk), .R(n13214), .S(1'b1), .Q(
        fifo[793]) );
  DFFSR fifo_reg_13__36_ ( .D(n3764), .CLK(wclk), .R(n13214), .S(1'b1), .Q(
        fifo[792]) );
  DFFSR fifo_reg_13__35_ ( .D(n3765), .CLK(wclk), .R(n13215), .S(1'b1), .Q(
        fifo[791]) );
  DFFSR fifo_reg_13__34_ ( .D(n3766), .CLK(wclk), .R(n13215), .S(1'b1), .Q(
        fifo[790]) );
  DFFSR fifo_reg_13__33_ ( .D(n3767), .CLK(wclk), .R(n13215), .S(1'b1), .Q(
        fifo[789]) );
  DFFSR fifo_reg_13__32_ ( .D(n3768), .CLK(wclk), .R(n13215), .S(1'b1), .Q(
        fifo[788]) );
  DFFSR fifo_reg_13__31_ ( .D(n3769), .CLK(wclk), .R(n13215), .S(1'b1), .Q(
        fifo[787]) );
  DFFSR fifo_reg_13__30_ ( .D(n3770), .CLK(wclk), .R(n13215), .S(1'b1), .Q(
        fifo[786]) );
  DFFSR fifo_reg_13__29_ ( .D(n3771), .CLK(wclk), .R(n13215), .S(1'b1), .Q(
        fifo[785]) );
  DFFSR fifo_reg_13__28_ ( .D(n3772), .CLK(wclk), .R(n13215), .S(1'b1), .Q(
        fifo[784]) );
  DFFSR fifo_reg_13__27_ ( .D(n3773), .CLK(wclk), .R(n13215), .S(1'b1), .Q(
        fifo[783]) );
  DFFSR fifo_reg_13__26_ ( .D(n3774), .CLK(wclk), .R(n13215), .S(1'b1), .Q(
        fifo[782]) );
  DFFSR fifo_reg_13__25_ ( .D(n3775), .CLK(wclk), .R(n13215), .S(1'b1), .Q(
        fifo[781]) );
  DFFSR fifo_reg_13__24_ ( .D(n3776), .CLK(wclk), .R(n13215), .S(1'b1), .Q(
        fifo[780]) );
  DFFSR fifo_reg_13__23_ ( .D(n3777), .CLK(wclk), .R(n13216), .S(1'b1), .Q(
        fifo[779]) );
  DFFSR fifo_reg_13__22_ ( .D(n3778), .CLK(wclk), .R(n13216), .S(1'b1), .Q(
        fifo[778]) );
  DFFSR fifo_reg_13__21_ ( .D(n3779), .CLK(wclk), .R(n13216), .S(1'b1), .Q(
        fifo[777]) );
  DFFSR fifo_reg_13__20_ ( .D(n3780), .CLK(wclk), .R(n13216), .S(1'b1), .Q(
        fifo[776]) );
  DFFSR fifo_reg_13__19_ ( .D(n3781), .CLK(wclk), .R(n13216), .S(1'b1), .Q(
        fifo[775]) );
  DFFSR fifo_reg_13__18_ ( .D(n3782), .CLK(wclk), .R(n13216), .S(1'b1), .Q(
        fifo[774]) );
  DFFSR fifo_reg_13__17_ ( .D(n3783), .CLK(wclk), .R(n13216), .S(1'b1), .Q(
        fifo[773]) );
  DFFSR fifo_reg_13__16_ ( .D(n3784), .CLK(wclk), .R(n13216), .S(1'b1), .Q(
        fifo[772]) );
  DFFSR fifo_reg_13__15_ ( .D(n3785), .CLK(wclk), .R(n13106), .S(1'b1), .Q(
        fifo[771]) );
  DFFSR fifo_reg_13__14_ ( .D(n3786), .CLK(wclk), .R(n13108), .S(1'b1), .Q(
        fifo[770]) );
  DFFSR fifo_reg_13__13_ ( .D(n3787), .CLK(wclk), .R(n13111), .S(1'b1), .Q(
        fifo[769]) );
  DFFSR fifo_reg_13__12_ ( .D(n3788), .CLK(wclk), .R(n13114), .S(1'b1), .Q(
        fifo[768]) );
  DFFSR fifo_reg_13__11_ ( .D(n3789), .CLK(wclk), .R(n13117), .S(1'b1), .Q(
        fifo[767]) );
  DFFSR fifo_reg_13__10_ ( .D(n3790), .CLK(wclk), .R(n13119), .S(1'b1), .Q(
        fifo[766]) );
  DFFSR fifo_reg_13__9_ ( .D(n3791), .CLK(wclk), .R(n13122), .S(1'b1), .Q(
        fifo[765]) );
  DFFSR fifo_reg_13__8_ ( .D(n3792), .CLK(wclk), .R(n13125), .S(1'b1), .Q(
        fifo[764]) );
  DFFSR fifo_reg_13__7_ ( .D(n3793), .CLK(wclk), .R(n13128), .S(1'b1), .Q(
        fifo[763]) );
  DFFSR fifo_reg_13__6_ ( .D(n3794), .CLK(wclk), .R(n13130), .S(1'b1), .Q(
        fifo[762]) );
  DFFSR fifo_reg_13__5_ ( .D(n3795), .CLK(wclk), .R(n13133), .S(1'b1), .Q(
        fifo[761]) );
  DFFSR fifo_reg_13__4_ ( .D(n3796), .CLK(wclk), .R(n13136), .S(1'b1), .Q(
        fifo[760]) );
  DFFSR fifo_reg_13__3_ ( .D(n3797), .CLK(wclk), .R(n13139), .S(1'b1), .Q(
        fifo[759]) );
  DFFSR fifo_reg_13__2_ ( .D(n3798), .CLK(wclk), .R(n13141), .S(1'b1), .Q(
        fifo[758]) );
  DFFSR fifo_reg_13__1_ ( .D(n3799), .CLK(wclk), .R(n13144), .S(1'b1), .Q(
        fifo[757]) );
  DFFSR fifo_reg_13__0_ ( .D(n3800), .CLK(wclk), .R(n13147), .S(1'b1), .Q(
        fifo[756]) );
  DFFSR fifo_reg_14__41_ ( .D(n3801), .CLK(wclk), .R(n13216), .S(1'b1), .Q(
        fifo[755]) );
  DFFSR fifo_reg_14__40_ ( .D(n3802), .CLK(wclk), .R(n13216), .S(1'b1), .Q(
        fifo[754]) );
  DFFSR fifo_reg_14__39_ ( .D(n3803), .CLK(wclk), .R(n13216), .S(1'b1), .Q(
        fifo[753]) );
  DFFSR fifo_reg_14__38_ ( .D(n3804), .CLK(wclk), .R(n13216), .S(1'b1), .Q(
        fifo[752]) );
  DFFSR fifo_reg_14__37_ ( .D(n3805), .CLK(wclk), .R(n13217), .S(1'b1), .Q(
        fifo[751]) );
  DFFSR fifo_reg_14__36_ ( .D(n3806), .CLK(wclk), .R(n13217), .S(1'b1), .Q(
        fifo[750]) );
  DFFSR fifo_reg_14__35_ ( .D(n3807), .CLK(wclk), .R(n13217), .S(1'b1), .Q(
        fifo[749]) );
  DFFSR fifo_reg_14__34_ ( .D(n3808), .CLK(wclk), .R(n13217), .S(1'b1), .Q(
        fifo[748]) );
  DFFSR fifo_reg_14__33_ ( .D(n3809), .CLK(wclk), .R(n13217), .S(1'b1), .Q(
        fifo[747]) );
  DFFSR fifo_reg_14__32_ ( .D(n3810), .CLK(wclk), .R(n13217), .S(1'b1), .Q(
        fifo[746]) );
  DFFSR fifo_reg_14__31_ ( .D(n3811), .CLK(wclk), .R(n13217), .S(1'b1), .Q(
        fifo[745]) );
  DFFSR fifo_reg_14__30_ ( .D(n3812), .CLK(wclk), .R(n13217), .S(1'b1), .Q(
        fifo[744]) );
  DFFSR fifo_reg_14__29_ ( .D(n3813), .CLK(wclk), .R(n13217), .S(1'b1), .Q(
        fifo[743]) );
  DFFSR fifo_reg_14__28_ ( .D(n3814), .CLK(wclk), .R(n13217), .S(1'b1), .Q(
        fifo[742]) );
  DFFSR fifo_reg_14__27_ ( .D(n3815), .CLK(wclk), .R(n13217), .S(1'b1), .Q(
        fifo[741]) );
  DFFSR fifo_reg_14__26_ ( .D(n3816), .CLK(wclk), .R(n13217), .S(1'b1), .Q(
        fifo[740]) );
  DFFSR fifo_reg_14__25_ ( .D(n3817), .CLK(wclk), .R(n13218), .S(1'b1), .Q(
        fifo[739]) );
  DFFSR fifo_reg_14__24_ ( .D(n3818), .CLK(wclk), .R(n13218), .S(1'b1), .Q(
        fifo[738]) );
  DFFSR fifo_reg_14__23_ ( .D(n3819), .CLK(wclk), .R(n13218), .S(1'b1), .Q(
        fifo[737]) );
  DFFSR fifo_reg_14__22_ ( .D(n3820), .CLK(wclk), .R(n13218), .S(1'b1), .Q(
        fifo[736]) );
  DFFSR fifo_reg_14__21_ ( .D(n3821), .CLK(wclk), .R(n13218), .S(1'b1), .Q(
        fifo[735]) );
  DFFSR fifo_reg_14__20_ ( .D(n3822), .CLK(wclk), .R(n13218), .S(1'b1), .Q(
        fifo[734]) );
  DFFSR fifo_reg_14__19_ ( .D(n3823), .CLK(wclk), .R(n13218), .S(1'b1), .Q(
        fifo[733]) );
  DFFSR fifo_reg_14__18_ ( .D(n3824), .CLK(wclk), .R(n13218), .S(1'b1), .Q(
        fifo[732]) );
  DFFSR fifo_reg_14__17_ ( .D(n3825), .CLK(wclk), .R(n13218), .S(1'b1), .Q(
        fifo[731]) );
  DFFSR fifo_reg_14__16_ ( .D(n3826), .CLK(wclk), .R(n13218), .S(1'b1), .Q(
        fifo[730]) );
  DFFSR fifo_reg_14__15_ ( .D(n3827), .CLK(wclk), .R(n13106), .S(1'b1), .Q(
        fifo[729]) );
  DFFSR fifo_reg_14__14_ ( .D(n3828), .CLK(wclk), .R(n13109), .S(1'b1), .Q(
        fifo[728]) );
  DFFSR fifo_reg_14__13_ ( .D(n3829), .CLK(wclk), .R(n13111), .S(1'b1), .Q(
        fifo[727]) );
  DFFSR fifo_reg_14__12_ ( .D(n3830), .CLK(wclk), .R(n13114), .S(1'b1), .Q(
        fifo[726]) );
  DFFSR fifo_reg_14__11_ ( .D(n3831), .CLK(wclk), .R(n13117), .S(1'b1), .Q(
        fifo[725]) );
  DFFSR fifo_reg_14__10_ ( .D(n3832), .CLK(wclk), .R(n13120), .S(1'b1), .Q(
        fifo[724]) );
  DFFSR fifo_reg_14__9_ ( .D(n3833), .CLK(wclk), .R(n13122), .S(1'b1), .Q(
        fifo[723]) );
  DFFSR fifo_reg_14__8_ ( .D(n3834), .CLK(wclk), .R(n13125), .S(1'b1), .Q(
        fifo[722]) );
  DFFSR fifo_reg_14__7_ ( .D(n3835), .CLK(wclk), .R(n13128), .S(1'b1), .Q(
        fifo[721]) );
  DFFSR fifo_reg_14__6_ ( .D(n3836), .CLK(wclk), .R(n13131), .S(1'b1), .Q(
        fifo[720]) );
  DFFSR fifo_reg_14__5_ ( .D(n3837), .CLK(wclk), .R(n13133), .S(1'b1), .Q(
        fifo[719]) );
  DFFSR fifo_reg_14__4_ ( .D(n3838), .CLK(wclk), .R(n13136), .S(1'b1), .Q(
        fifo[718]) );
  DFFSR fifo_reg_14__3_ ( .D(n3839), .CLK(wclk), .R(n13139), .S(1'b1), .Q(
        fifo[717]) );
  DFFSR fifo_reg_14__2_ ( .D(n3840), .CLK(wclk), .R(n13142), .S(1'b1), .Q(
        fifo[716]) );
  DFFSR fifo_reg_14__1_ ( .D(n3841), .CLK(wclk), .R(n13144), .S(1'b1), .Q(
        fifo[715]) );
  DFFSR fifo_reg_14__0_ ( .D(n3842), .CLK(wclk), .R(n13147), .S(1'b1), .Q(
        fifo[714]) );
  DFFSR fifo_reg_15__41_ ( .D(n3843), .CLK(wclk), .R(n13218), .S(1'b1), .Q(
        fifo[713]) );
  DFFSR fifo_reg_15__40_ ( .D(n3844), .CLK(wclk), .R(n13218), .S(1'b1), .Q(
        fifo[712]) );
  DFFSR fifo_reg_15__39_ ( .D(n3845), .CLK(wclk), .R(n13219), .S(1'b1), .Q(
        fifo[711]) );
  DFFSR fifo_reg_15__38_ ( .D(n3846), .CLK(wclk), .R(n13219), .S(1'b1), .Q(
        fifo[710]) );
  DFFSR fifo_reg_15__37_ ( .D(n3847), .CLK(wclk), .R(n13219), .S(1'b1), .Q(
        fifo[709]) );
  DFFSR fifo_reg_15__36_ ( .D(n3848), .CLK(wclk), .R(n13219), .S(1'b1), .Q(
        fifo[708]) );
  DFFSR fifo_reg_15__35_ ( .D(n3849), .CLK(wclk), .R(n13219), .S(1'b1), .Q(
        fifo[707]) );
  DFFSR fifo_reg_15__34_ ( .D(n3850), .CLK(wclk), .R(n13219), .S(1'b1), .Q(
        fifo[706]) );
  DFFSR fifo_reg_15__33_ ( .D(n3851), .CLK(wclk), .R(n13219), .S(1'b1), .Q(
        fifo[705]) );
  DFFSR fifo_reg_15__32_ ( .D(n3852), .CLK(wclk), .R(n13219), .S(1'b1), .Q(
        fifo[704]) );
  DFFSR fifo_reg_15__31_ ( .D(n3853), .CLK(wclk), .R(n13219), .S(1'b1), .Q(
        fifo[703]) );
  DFFSR fifo_reg_15__30_ ( .D(n3854), .CLK(wclk), .R(n13219), .S(1'b1), .Q(
        fifo[702]) );
  DFFSR fifo_reg_15__29_ ( .D(n3855), .CLK(wclk), .R(n13219), .S(1'b1), .Q(
        fifo[701]) );
  DFFSR fifo_reg_15__28_ ( .D(n3856), .CLK(wclk), .R(n13219), .S(1'b1), .Q(
        fifo[700]) );
  DFFSR fifo_reg_15__27_ ( .D(n3857), .CLK(wclk), .R(n13220), .S(1'b1), .Q(
        fifo[699]) );
  DFFSR fifo_reg_15__26_ ( .D(n3858), .CLK(wclk), .R(n13220), .S(1'b1), .Q(
        fifo[698]) );
  DFFSR fifo_reg_15__25_ ( .D(n3859), .CLK(wclk), .R(n13220), .S(1'b1), .Q(
        fifo[697]) );
  DFFSR fifo_reg_15__24_ ( .D(n3860), .CLK(wclk), .R(n13220), .S(1'b1), .Q(
        fifo[696]) );
  DFFSR fifo_reg_15__23_ ( .D(n3861), .CLK(wclk), .R(n13220), .S(1'b1), .Q(
        fifo[695]) );
  DFFSR fifo_reg_15__22_ ( .D(n3862), .CLK(wclk), .R(n13220), .S(1'b1), .Q(
        fifo[694]) );
  DFFSR fifo_reg_15__21_ ( .D(n3863), .CLK(wclk), .R(n13220), .S(1'b1), .Q(
        fifo[693]) );
  DFFSR fifo_reg_15__20_ ( .D(n3864), .CLK(wclk), .R(n13220), .S(1'b1), .Q(
        fifo[692]) );
  DFFSR fifo_reg_15__19_ ( .D(n3865), .CLK(wclk), .R(n13220), .S(1'b1), .Q(
        fifo[691]) );
  DFFSR fifo_reg_15__18_ ( .D(n3866), .CLK(wclk), .R(n13220), .S(1'b1), .Q(
        fifo[690]) );
  DFFSR fifo_reg_15__17_ ( .D(n3867), .CLK(wclk), .R(n13220), .S(1'b1), .Q(
        fifo[689]) );
  DFFSR fifo_reg_15__16_ ( .D(n3868), .CLK(wclk), .R(n13220), .S(1'b1), .Q(
        fifo[688]) );
  DFFSR fifo_reg_15__15_ ( .D(n3869), .CLK(wclk), .R(n13106), .S(1'b1), .Q(
        fifo[687]) );
  DFFSR fifo_reg_15__14_ ( .D(n3870), .CLK(wclk), .R(n13109), .S(1'b1), .Q(
        fifo[686]) );
  DFFSR fifo_reg_15__13_ ( .D(n3871), .CLK(wclk), .R(n13111), .S(1'b1), .Q(
        fifo[685]) );
  DFFSR fifo_reg_15__12_ ( .D(n3872), .CLK(wclk), .R(n13114), .S(1'b1), .Q(
        fifo[684]) );
  DFFSR fifo_reg_15__11_ ( .D(n3873), .CLK(wclk), .R(n13117), .S(1'b1), .Q(
        fifo[683]) );
  DFFSR fifo_reg_15__10_ ( .D(n3874), .CLK(wclk), .R(n13120), .S(1'b1), .Q(
        fifo[682]) );
  DFFSR fifo_reg_15__9_ ( .D(n3875), .CLK(wclk), .R(n13122), .S(1'b1), .Q(
        fifo[681]) );
  DFFSR fifo_reg_15__8_ ( .D(n3876), .CLK(wclk), .R(n13125), .S(1'b1), .Q(
        fifo[680]) );
  DFFSR fifo_reg_15__7_ ( .D(n3877), .CLK(wclk), .R(n13128), .S(1'b1), .Q(
        fifo[679]) );
  DFFSR fifo_reg_15__6_ ( .D(n3878), .CLK(wclk), .R(n13131), .S(1'b1), .Q(
        fifo[678]) );
  DFFSR fifo_reg_15__5_ ( .D(n3879), .CLK(wclk), .R(n13133), .S(1'b1), .Q(
        fifo[677]) );
  DFFSR fifo_reg_15__4_ ( .D(n3880), .CLK(wclk), .R(n13136), .S(1'b1), .Q(
        fifo[676]) );
  DFFSR fifo_reg_15__3_ ( .D(n3881), .CLK(wclk), .R(n13139), .S(1'b1), .Q(
        fifo[675]) );
  DFFSR fifo_reg_15__2_ ( .D(n3882), .CLK(wclk), .R(n13142), .S(1'b1), .Q(
        fifo[674]) );
  DFFSR fifo_reg_15__1_ ( .D(n3883), .CLK(wclk), .R(n13144), .S(1'b1), .Q(
        fifo[673]) );
  DFFSR fifo_reg_15__0_ ( .D(n3884), .CLK(wclk), .R(n13147), .S(1'b1), .Q(
        fifo[672]) );
  DFFSR fifo_reg_16__41_ ( .D(n3885), .CLK(wclk), .R(n13169), .S(1'b1), .Q(
        fifo[671]) );
  DFFSR fifo_reg_16__40_ ( .D(n3886), .CLK(wclk), .R(n13169), .S(1'b1), .Q(
        fifo[670]) );
  DFFSR fifo_reg_16__39_ ( .D(n3887), .CLK(wclk), .R(n13169), .S(1'b1), .Q(
        fifo[669]) );
  DFFSR fifo_reg_16__38_ ( .D(n3888), .CLK(wclk), .R(n13169), .S(1'b1), .Q(
        fifo[668]) );
  DFFSR fifo_reg_16__37_ ( .D(n3889), .CLK(wclk), .R(n13169), .S(1'b1), .Q(
        fifo[667]) );
  DFFSR fifo_reg_16__36_ ( .D(n3890), .CLK(wclk), .R(n13169), .S(1'b1), .Q(
        fifo[666]) );
  DFFSR fifo_reg_16__35_ ( .D(n3891), .CLK(wclk), .R(n13169), .S(1'b1), .Q(
        fifo[665]) );
  DFFSR fifo_reg_16__34_ ( .D(n3892), .CLK(wclk), .R(n13169), .S(1'b1), .Q(
        fifo[664]) );
  DFFSR fifo_reg_16__33_ ( .D(n3893), .CLK(wclk), .R(n13169), .S(1'b1), .Q(
        fifo[663]) );
  DFFSR fifo_reg_16__32_ ( .D(n3894), .CLK(wclk), .R(n13169), .S(1'b1), .Q(
        fifo[662]) );
  DFFSR fifo_reg_16__31_ ( .D(n3895), .CLK(wclk), .R(n13169), .S(1'b1), .Q(
        fifo[661]) );
  DFFSR fifo_reg_16__30_ ( .D(n3896), .CLK(wclk), .R(n13169), .S(1'b1), .Q(
        fifo[660]) );
  DFFSR fifo_reg_16__29_ ( .D(n3897), .CLK(wclk), .R(n13170), .S(1'b1), .Q(
        fifo[659]) );
  DFFSR fifo_reg_16__28_ ( .D(n3898), .CLK(wclk), .R(n13170), .S(1'b1), .Q(
        fifo[658]) );
  DFFSR fifo_reg_16__27_ ( .D(n3899), .CLK(wclk), .R(n13170), .S(1'b1), .Q(
        fifo[657]) );
  DFFSR fifo_reg_16__26_ ( .D(n3900), .CLK(wclk), .R(n13170), .S(1'b1), .Q(
        fifo[656]) );
  DFFSR fifo_reg_16__25_ ( .D(n3901), .CLK(wclk), .R(n13170), .S(1'b1), .Q(
        fifo[655]) );
  DFFSR fifo_reg_16__24_ ( .D(n3902), .CLK(wclk), .R(n13170), .S(1'b1), .Q(
        fifo[654]) );
  DFFSR fifo_reg_16__23_ ( .D(n3903), .CLK(wclk), .R(n13170), .S(1'b1), .Q(
        fifo[653]) );
  DFFSR fifo_reg_16__22_ ( .D(n3904), .CLK(wclk), .R(n13170), .S(1'b1), .Q(
        fifo[652]) );
  DFFSR fifo_reg_16__21_ ( .D(n3905), .CLK(wclk), .R(n13170), .S(1'b1), .Q(
        fifo[651]) );
  DFFSR fifo_reg_16__20_ ( .D(n3906), .CLK(wclk), .R(n13170), .S(1'b1), .Q(
        fifo[650]) );
  DFFSR fifo_reg_16__19_ ( .D(n3907), .CLK(wclk), .R(n13170), .S(1'b1), .Q(
        fifo[649]) );
  DFFSR fifo_reg_16__18_ ( .D(n3908), .CLK(wclk), .R(n13170), .S(1'b1), .Q(
        fifo[648]) );
  DFFSR fifo_reg_16__17_ ( .D(n3909), .CLK(wclk), .R(n13171), .S(1'b1), .Q(
        fifo[647]) );
  DFFSR fifo_reg_16__16_ ( .D(n3910), .CLK(wclk), .R(n13171), .S(1'b1), .Q(
        fifo[646]) );
  DFFSR fifo_reg_16__15_ ( .D(n3911), .CLK(wclk), .R(n13106), .S(1'b1), .Q(
        fifo[645]) );
  DFFSR fifo_reg_16__14_ ( .D(n3912), .CLK(wclk), .R(n13109), .S(1'b1), .Q(
        fifo[644]) );
  DFFSR fifo_reg_16__13_ ( .D(n3913), .CLK(wclk), .R(n13111), .S(1'b1), .Q(
        fifo[643]) );
  DFFSR fifo_reg_16__12_ ( .D(n3914), .CLK(wclk), .R(n13114), .S(1'b1), .Q(
        fifo[642]) );
  DFFSR fifo_reg_16__11_ ( .D(n3915), .CLK(wclk), .R(n13117), .S(1'b1), .Q(
        fifo[641]) );
  DFFSR fifo_reg_16__10_ ( .D(n3916), .CLK(wclk), .R(n13120), .S(1'b1), .Q(
        fifo[640]) );
  DFFSR fifo_reg_16__9_ ( .D(n3917), .CLK(wclk), .R(n13122), .S(1'b1), .Q(
        fifo[639]) );
  DFFSR fifo_reg_16__8_ ( .D(n3918), .CLK(wclk), .R(n13125), .S(1'b1), .Q(
        fifo[638]) );
  DFFSR fifo_reg_16__7_ ( .D(n3919), .CLK(wclk), .R(n13128), .S(1'b1), .Q(
        fifo[637]) );
  DFFSR fifo_reg_16__6_ ( .D(n3920), .CLK(wclk), .R(n13131), .S(1'b1), .Q(
        fifo[636]) );
  DFFSR fifo_reg_16__5_ ( .D(n3921), .CLK(wclk), .R(n13133), .S(1'b1), .Q(
        fifo[635]) );
  DFFSR fifo_reg_16__4_ ( .D(n3922), .CLK(wclk), .R(n13136), .S(1'b1), .Q(
        fifo[634]) );
  DFFSR fifo_reg_16__3_ ( .D(n3923), .CLK(wclk), .R(n13139), .S(1'b1), .Q(
        fifo[633]) );
  DFFSR fifo_reg_16__2_ ( .D(n3924), .CLK(wclk), .R(n13142), .S(1'b1), .Q(
        fifo[632]) );
  DFFSR fifo_reg_16__1_ ( .D(n3925), .CLK(wclk), .R(n13144), .S(1'b1), .Q(
        fifo[631]) );
  DFFSR fifo_reg_16__0_ ( .D(n3926), .CLK(wclk), .R(n13147), .S(1'b1), .Q(
        fifo[630]) );
  DFFSR fifo_reg_17__41_ ( .D(n3927), .CLK(wclk), .R(n13171), .S(1'b1), .Q(
        fifo[629]) );
  DFFSR fifo_reg_17__40_ ( .D(n3928), .CLK(wclk), .R(n13171), .S(1'b1), .Q(
        fifo[628]) );
  DFFSR fifo_reg_17__39_ ( .D(n3929), .CLK(wclk), .R(n13171), .S(1'b1), .Q(
        fifo[627]) );
  DFFSR fifo_reg_17__38_ ( .D(n3930), .CLK(wclk), .R(n13171), .S(1'b1), .Q(
        fifo[626]) );
  DFFSR fifo_reg_17__37_ ( .D(n3931), .CLK(wclk), .R(n13171), .S(1'b1), .Q(
        fifo[625]) );
  DFFSR fifo_reg_17__36_ ( .D(n3932), .CLK(wclk), .R(n13171), .S(1'b1), .Q(
        fifo[624]) );
  DFFSR fifo_reg_17__35_ ( .D(n3933), .CLK(wclk), .R(n13171), .S(1'b1), .Q(
        fifo[623]) );
  DFFSR fifo_reg_17__34_ ( .D(n3934), .CLK(wclk), .R(n13171), .S(1'b1), .Q(
        fifo[622]) );
  DFFSR fifo_reg_17__33_ ( .D(n3935), .CLK(wclk), .R(n13171), .S(1'b1), .Q(
        fifo[621]) );
  DFFSR fifo_reg_17__32_ ( .D(n3936), .CLK(wclk), .R(n13171), .S(1'b1), .Q(
        fifo[620]) );
  DFFSR fifo_reg_17__31_ ( .D(n3937), .CLK(wclk), .R(n13172), .S(1'b1), .Q(
        fifo[619]) );
  DFFSR fifo_reg_17__30_ ( .D(n3938), .CLK(wclk), .R(n13172), .S(1'b1), .Q(
        fifo[618]) );
  DFFSR fifo_reg_17__29_ ( .D(n3939), .CLK(wclk), .R(n13172), .S(1'b1), .Q(
        fifo[617]) );
  DFFSR fifo_reg_17__28_ ( .D(n3940), .CLK(wclk), .R(n13172), .S(1'b1), .Q(
        fifo[616]) );
  DFFSR fifo_reg_17__27_ ( .D(n3941), .CLK(wclk), .R(n13172), .S(1'b1), .Q(
        fifo[615]) );
  DFFSR fifo_reg_17__26_ ( .D(n3942), .CLK(wclk), .R(n13172), .S(1'b1), .Q(
        fifo[614]) );
  DFFSR fifo_reg_17__25_ ( .D(n3943), .CLK(wclk), .R(n13172), .S(1'b1), .Q(
        fifo[613]) );
  DFFSR fifo_reg_17__24_ ( .D(n3944), .CLK(wclk), .R(n13172), .S(1'b1), .Q(
        fifo[612]) );
  DFFSR fifo_reg_17__23_ ( .D(n3945), .CLK(wclk), .R(n13172), .S(1'b1), .Q(
        fifo[611]) );
  DFFSR fifo_reg_17__22_ ( .D(n3946), .CLK(wclk), .R(n13172), .S(1'b1), .Q(
        fifo[610]) );
  DFFSR fifo_reg_17__21_ ( .D(n3947), .CLK(wclk), .R(n13172), .S(1'b1), .Q(
        fifo[609]) );
  DFFSR fifo_reg_17__20_ ( .D(n3948), .CLK(wclk), .R(n13172), .S(1'b1), .Q(
        fifo[608]) );
  DFFSR fifo_reg_17__19_ ( .D(n3949), .CLK(wclk), .R(n13173), .S(1'b1), .Q(
        fifo[607]) );
  DFFSR fifo_reg_17__18_ ( .D(n3950), .CLK(wclk), .R(n13173), .S(1'b1), .Q(
        fifo[606]) );
  DFFSR fifo_reg_17__17_ ( .D(n3951), .CLK(wclk), .R(n13173), .S(1'b1), .Q(
        fifo[605]) );
  DFFSR fifo_reg_17__16_ ( .D(n3952), .CLK(wclk), .R(n13173), .S(1'b1), .Q(
        fifo[604]) );
  DFFSR fifo_reg_17__15_ ( .D(n3953), .CLK(wclk), .R(n13106), .S(1'b1), .Q(
        fifo[603]) );
  DFFSR fifo_reg_17__14_ ( .D(n3954), .CLK(wclk), .R(n13109), .S(1'b1), .Q(
        fifo[602]) );
  DFFSR fifo_reg_17__13_ ( .D(n3955), .CLK(wclk), .R(n13112), .S(1'b1), .Q(
        fifo[601]) );
  DFFSR fifo_reg_17__12_ ( .D(n3956), .CLK(wclk), .R(n13114), .S(1'b1), .Q(
        fifo[600]) );
  DFFSR fifo_reg_17__11_ ( .D(n3957), .CLK(wclk), .R(n13117), .S(1'b1), .Q(
        fifo[599]) );
  DFFSR fifo_reg_17__10_ ( .D(n3958), .CLK(wclk), .R(n13120), .S(1'b1), .Q(
        fifo[598]) );
  DFFSR fifo_reg_17__9_ ( .D(n3959), .CLK(wclk), .R(n13123), .S(1'b1), .Q(
        fifo[597]) );
  DFFSR fifo_reg_17__8_ ( .D(n3960), .CLK(wclk), .R(n13125), .S(1'b1), .Q(
        fifo[596]) );
  DFFSR fifo_reg_17__7_ ( .D(n3961), .CLK(wclk), .R(n13128), .S(1'b1), .Q(
        fifo[595]) );
  DFFSR fifo_reg_17__6_ ( .D(n3962), .CLK(wclk), .R(n13131), .S(1'b1), .Q(
        fifo[594]) );
  DFFSR fifo_reg_17__5_ ( .D(n3963), .CLK(wclk), .R(n13134), .S(1'b1), .Q(
        fifo[593]) );
  DFFSR fifo_reg_17__4_ ( .D(n3964), .CLK(wclk), .R(n13136), .S(1'b1), .Q(
        fifo[592]) );
  DFFSR fifo_reg_17__3_ ( .D(n3965), .CLK(wclk), .R(n13139), .S(1'b1), .Q(
        fifo[591]) );
  DFFSR fifo_reg_17__2_ ( .D(n3966), .CLK(wclk), .R(n13142), .S(1'b1), .Q(
        fifo[590]) );
  DFFSR fifo_reg_17__1_ ( .D(n3967), .CLK(wclk), .R(n13145), .S(1'b1), .Q(
        fifo[589]) );
  DFFSR fifo_reg_17__0_ ( .D(n3968), .CLK(wclk), .R(n13147), .S(1'b1), .Q(
        fifo[588]) );
  DFFSR fifo_reg_18__41_ ( .D(n3969), .CLK(wclk), .R(n13173), .S(1'b1), .Q(
        fifo[587]) );
  DFFSR fifo_reg_18__40_ ( .D(n3970), .CLK(wclk), .R(n13173), .S(1'b1), .Q(
        fifo[586]) );
  DFFSR fifo_reg_18__39_ ( .D(n3971), .CLK(wclk), .R(n13173), .S(1'b1), .Q(
        fifo[585]) );
  DFFSR fifo_reg_18__38_ ( .D(n3972), .CLK(wclk), .R(n13173), .S(1'b1), .Q(
        fifo[584]) );
  DFFSR fifo_reg_18__37_ ( .D(n3973), .CLK(wclk), .R(n13173), .S(1'b1), .Q(
        fifo[583]) );
  DFFSR fifo_reg_18__36_ ( .D(n3974), .CLK(wclk), .R(n13173), .S(1'b1), .Q(
        fifo[582]) );
  DFFSR fifo_reg_18__35_ ( .D(n3975), .CLK(wclk), .R(n13173), .S(1'b1), .Q(
        fifo[581]) );
  DFFSR fifo_reg_18__34_ ( .D(n3976), .CLK(wclk), .R(n13173), .S(1'b1), .Q(
        fifo[580]) );
  DFFSR fifo_reg_18__33_ ( .D(n3977), .CLK(wclk), .R(n13174), .S(1'b1), .Q(
        fifo[579]) );
  DFFSR fifo_reg_18__32_ ( .D(n3978), .CLK(wclk), .R(n13174), .S(1'b1), .Q(
        fifo[578]) );
  DFFSR fifo_reg_18__31_ ( .D(n3979), .CLK(wclk), .R(n13174), .S(1'b1), .Q(
        fifo[577]) );
  DFFSR fifo_reg_18__30_ ( .D(n3980), .CLK(wclk), .R(n13174), .S(1'b1), .Q(
        fifo[576]) );
  DFFSR fifo_reg_18__29_ ( .D(n3981), .CLK(wclk), .R(n13174), .S(1'b1), .Q(
        fifo[575]) );
  DFFSR fifo_reg_18__28_ ( .D(n3982), .CLK(wclk), .R(n13174), .S(1'b1), .Q(
        fifo[574]) );
  DFFSR fifo_reg_18__27_ ( .D(n3983), .CLK(wclk), .R(n13174), .S(1'b1), .Q(
        fifo[573]) );
  DFFSR fifo_reg_18__26_ ( .D(n3984), .CLK(wclk), .R(n13174), .S(1'b1), .Q(
        fifo[572]) );
  DFFSR fifo_reg_18__25_ ( .D(n3985), .CLK(wclk), .R(n13174), .S(1'b1), .Q(
        fifo[571]) );
  DFFSR fifo_reg_18__24_ ( .D(n3986), .CLK(wclk), .R(n13174), .S(1'b1), .Q(
        fifo[570]) );
  DFFSR fifo_reg_18__23_ ( .D(n3987), .CLK(wclk), .R(n13174), .S(1'b1), .Q(
        fifo[569]) );
  DFFSR fifo_reg_18__22_ ( .D(n3988), .CLK(wclk), .R(n13174), .S(1'b1), .Q(
        fifo[568]) );
  DFFSR fifo_reg_18__21_ ( .D(n3989), .CLK(wclk), .R(n13175), .S(1'b1), .Q(
        fifo[567]) );
  DFFSR fifo_reg_18__20_ ( .D(n3990), .CLK(wclk), .R(n13175), .S(1'b1), .Q(
        fifo[566]) );
  DFFSR fifo_reg_18__19_ ( .D(n3991), .CLK(wclk), .R(n13175), .S(1'b1), .Q(
        fifo[565]) );
  DFFSR fifo_reg_18__18_ ( .D(n3992), .CLK(wclk), .R(n13175), .S(1'b1), .Q(
        fifo[564]) );
  DFFSR fifo_reg_18__17_ ( .D(n3993), .CLK(wclk), .R(n13175), .S(1'b1), .Q(
        fifo[563]) );
  DFFSR fifo_reg_18__16_ ( .D(n3994), .CLK(wclk), .R(n13175), .S(1'b1), .Q(
        fifo[562]) );
  DFFSR fifo_reg_18__15_ ( .D(n3995), .CLK(wclk), .R(n13106), .S(1'b1), .Q(
        fifo[561]) );
  DFFSR fifo_reg_18__14_ ( .D(n3996), .CLK(wclk), .R(n13109), .S(1'b1), .Q(
        fifo[560]) );
  DFFSR fifo_reg_18__13_ ( .D(n3997), .CLK(wclk), .R(n13112), .S(1'b1), .Q(
        fifo[559]) );
  DFFSR fifo_reg_18__12_ ( .D(n3998), .CLK(wclk), .R(n13114), .S(1'b1), .Q(
        fifo[558]) );
  DFFSR fifo_reg_18__11_ ( .D(n3999), .CLK(wclk), .R(n13117), .S(1'b1), .Q(
        fifo[557]) );
  DFFSR fifo_reg_18__10_ ( .D(n4000), .CLK(wclk), .R(n13120), .S(1'b1), .Q(
        fifo[556]) );
  DFFSR fifo_reg_18__9_ ( .D(n4001), .CLK(wclk), .R(n13123), .S(1'b1), .Q(
        fifo[555]) );
  DFFSR fifo_reg_18__8_ ( .D(n4002), .CLK(wclk), .R(n13125), .S(1'b1), .Q(
        fifo[554]) );
  DFFSR fifo_reg_18__7_ ( .D(n4003), .CLK(wclk), .R(n13128), .S(1'b1), .Q(
        fifo[553]) );
  DFFSR fifo_reg_18__6_ ( .D(n4004), .CLK(wclk), .R(n13131), .S(1'b1), .Q(
        fifo[552]) );
  DFFSR fifo_reg_18__5_ ( .D(n4005), .CLK(wclk), .R(n13134), .S(1'b1), .Q(
        fifo[551]) );
  DFFSR fifo_reg_18__4_ ( .D(n4006), .CLK(wclk), .R(n13136), .S(1'b1), .Q(
        fifo[550]) );
  DFFSR fifo_reg_18__3_ ( .D(n4007), .CLK(wclk), .R(n13139), .S(1'b1), .Q(
        fifo[549]) );
  DFFSR fifo_reg_18__2_ ( .D(n4008), .CLK(wclk), .R(n13142), .S(1'b1), .Q(
        fifo[548]) );
  DFFSR fifo_reg_18__1_ ( .D(n4009), .CLK(wclk), .R(n13145), .S(1'b1), .Q(
        fifo[547]) );
  DFFSR fifo_reg_18__0_ ( .D(n4010), .CLK(wclk), .R(n13147), .S(1'b1), .Q(
        fifo[546]) );
  DFFSR fifo_reg_19__41_ ( .D(n4011), .CLK(wclk), .R(n13175), .S(1'b1), .Q(
        fifo[545]) );
  DFFSR fifo_reg_19__40_ ( .D(n4012), .CLK(wclk), .R(n13175), .S(1'b1), .Q(
        fifo[544]) );
  DFFSR fifo_reg_19__39_ ( .D(n4013), .CLK(wclk), .R(n13175), .S(1'b1), .Q(
        fifo[543]) );
  DFFSR fifo_reg_19__38_ ( .D(n4014), .CLK(wclk), .R(n13175), .S(1'b1), .Q(
        fifo[542]) );
  DFFSR fifo_reg_19__37_ ( .D(n4015), .CLK(wclk), .R(n13175), .S(1'b1), .Q(
        fifo[541]) );
  DFFSR fifo_reg_19__36_ ( .D(n4016), .CLK(wclk), .R(n13175), .S(1'b1), .Q(
        fifo[540]) );
  DFFSR fifo_reg_19__35_ ( .D(n4017), .CLK(wclk), .R(n13176), .S(1'b1), .Q(
        fifo[539]) );
  DFFSR fifo_reg_19__34_ ( .D(n4018), .CLK(wclk), .R(n13176), .S(1'b1), .Q(
        fifo[538]) );
  DFFSR fifo_reg_19__33_ ( .D(n4019), .CLK(wclk), .R(n13176), .S(1'b1), .Q(
        fifo[537]) );
  DFFSR fifo_reg_19__32_ ( .D(n4020), .CLK(wclk), .R(n13176), .S(1'b1), .Q(
        fifo[536]) );
  DFFSR fifo_reg_19__31_ ( .D(n4021), .CLK(wclk), .R(n13176), .S(1'b1), .Q(
        fifo[535]) );
  DFFSR fifo_reg_19__30_ ( .D(n4022), .CLK(wclk), .R(n13176), .S(1'b1), .Q(
        fifo[534]) );
  DFFSR fifo_reg_19__29_ ( .D(n4023), .CLK(wclk), .R(n13176), .S(1'b1), .Q(
        fifo[533]) );
  DFFSR fifo_reg_19__28_ ( .D(n4024), .CLK(wclk), .R(n13176), .S(1'b1), .Q(
        fifo[532]) );
  DFFSR fifo_reg_19__27_ ( .D(n4025), .CLK(wclk), .R(n13176), .S(1'b1), .Q(
        fifo[531]) );
  DFFSR fifo_reg_19__26_ ( .D(n4026), .CLK(wclk), .R(n13176), .S(1'b1), .Q(
        fifo[530]) );
  DFFSR fifo_reg_19__25_ ( .D(n4027), .CLK(wclk), .R(n13176), .S(1'b1), .Q(
        fifo[529]) );
  DFFSR fifo_reg_19__24_ ( .D(n4028), .CLK(wclk), .R(n13176), .S(1'b1), .Q(
        fifo[528]) );
  DFFSR fifo_reg_19__23_ ( .D(n4029), .CLK(wclk), .R(n13177), .S(1'b1), .Q(
        fifo[527]) );
  DFFSR fifo_reg_19__22_ ( .D(n4030), .CLK(wclk), .R(n13177), .S(1'b1), .Q(
        fifo[526]) );
  DFFSR fifo_reg_19__21_ ( .D(n4031), .CLK(wclk), .R(n13177), .S(1'b1), .Q(
        fifo[525]) );
  DFFSR fifo_reg_19__20_ ( .D(n4032), .CLK(wclk), .R(n13177), .S(1'b1), .Q(
        fifo[524]) );
  DFFSR fifo_reg_19__19_ ( .D(n4033), .CLK(wclk), .R(n13177), .S(1'b1), .Q(
        fifo[523]) );
  DFFSR fifo_reg_19__18_ ( .D(n4034), .CLK(wclk), .R(n13177), .S(1'b1), .Q(
        fifo[522]) );
  DFFSR fifo_reg_19__17_ ( .D(n4035), .CLK(wclk), .R(n13177), .S(1'b1), .Q(
        fifo[521]) );
  DFFSR fifo_reg_19__16_ ( .D(n4036), .CLK(wclk), .R(n13177), .S(1'b1), .Q(
        fifo[520]) );
  DFFSR fifo_reg_19__15_ ( .D(n4037), .CLK(wclk), .R(n13106), .S(1'b1), .Q(
        fifo[519]) );
  DFFSR fifo_reg_19__14_ ( .D(n4038), .CLK(wclk), .R(n13109), .S(1'b1), .Q(
        fifo[518]) );
  DFFSR fifo_reg_19__13_ ( .D(n4039), .CLK(wclk), .R(n13112), .S(1'b1), .Q(
        fifo[517]) );
  DFFSR fifo_reg_19__12_ ( .D(n4040), .CLK(wclk), .R(n13114), .S(1'b1), .Q(
        fifo[516]) );
  DFFSR fifo_reg_19__11_ ( .D(n4041), .CLK(wclk), .R(n13117), .S(1'b1), .Q(
        fifo[515]) );
  DFFSR fifo_reg_19__10_ ( .D(n4042), .CLK(wclk), .R(n13120), .S(1'b1), .Q(
        fifo[514]) );
  DFFSR fifo_reg_19__9_ ( .D(n4043), .CLK(wclk), .R(n13123), .S(1'b1), .Q(
        fifo[513]) );
  DFFSR fifo_reg_19__8_ ( .D(n4044), .CLK(wclk), .R(n13125), .S(1'b1), .Q(
        fifo[512]) );
  DFFSR fifo_reg_19__7_ ( .D(n4045), .CLK(wclk), .R(n13128), .S(1'b1), .Q(
        fifo[511]) );
  DFFSR fifo_reg_19__6_ ( .D(n4046), .CLK(wclk), .R(n13131), .S(1'b1), .Q(
        fifo[510]) );
  DFFSR fifo_reg_19__5_ ( .D(n4047), .CLK(wclk), .R(n13134), .S(1'b1), .Q(
        fifo[509]) );
  DFFSR fifo_reg_19__4_ ( .D(n4048), .CLK(wclk), .R(n13136), .S(1'b1), .Q(
        fifo[508]) );
  DFFSR fifo_reg_19__3_ ( .D(n4049), .CLK(wclk), .R(n13139), .S(1'b1), .Q(
        fifo[507]) );
  DFFSR fifo_reg_19__2_ ( .D(n4050), .CLK(wclk), .R(n13142), .S(1'b1), .Q(
        fifo[506]) );
  DFFSR fifo_reg_19__1_ ( .D(n4051), .CLK(wclk), .R(n13145), .S(1'b1), .Q(
        fifo[505]) );
  DFFSR fifo_reg_19__0_ ( .D(n4052), .CLK(wclk), .R(n13147), .S(1'b1), .Q(
        fifo[504]) );
  DFFSR fifo_reg_20__41_ ( .D(n4053), .CLK(wclk), .R(n13177), .S(1'b1), .Q(
        fifo[503]) );
  DFFSR fifo_reg_20__40_ ( .D(n4054), .CLK(wclk), .R(n13177), .S(1'b1), .Q(
        fifo[502]) );
  DFFSR fifo_reg_20__39_ ( .D(n4055), .CLK(wclk), .R(n13177), .S(1'b1), .Q(
        fifo[501]) );
  DFFSR fifo_reg_20__38_ ( .D(n4056), .CLK(wclk), .R(n13177), .S(1'b1), .Q(
        fifo[500]) );
  DFFSR fifo_reg_20__37_ ( .D(n4057), .CLK(wclk), .R(n13178), .S(1'b1), .Q(
        fifo[499]) );
  DFFSR fifo_reg_20__36_ ( .D(n4058), .CLK(wclk), .R(n13178), .S(1'b1), .Q(
        fifo[498]) );
  DFFSR fifo_reg_20__35_ ( .D(n4059), .CLK(wclk), .R(n13178), .S(1'b1), .Q(
        fifo[497]) );
  DFFSR fifo_reg_20__34_ ( .D(n4060), .CLK(wclk), .R(n13178), .S(1'b1), .Q(
        fifo[496]) );
  DFFSR fifo_reg_20__33_ ( .D(n4061), .CLK(wclk), .R(n13178), .S(1'b1), .Q(
        fifo[495]) );
  DFFSR fifo_reg_20__32_ ( .D(n4062), .CLK(wclk), .R(n13178), .S(1'b1), .Q(
        fifo[494]) );
  DFFSR fifo_reg_20__31_ ( .D(n4063), .CLK(wclk), .R(n13178), .S(1'b1), .Q(
        fifo[493]) );
  DFFSR fifo_reg_20__30_ ( .D(n4064), .CLK(wclk), .R(n13178), .S(1'b1), .Q(
        fifo[492]) );
  DFFSR fifo_reg_20__29_ ( .D(n4065), .CLK(wclk), .R(n13178), .S(1'b1), .Q(
        fifo[491]) );
  DFFSR fifo_reg_20__28_ ( .D(n4066), .CLK(wclk), .R(n13178), .S(1'b1), .Q(
        fifo[490]) );
  DFFSR fifo_reg_20__27_ ( .D(n4067), .CLK(wclk), .R(n13178), .S(1'b1), .Q(
        fifo[489]) );
  DFFSR fifo_reg_20__26_ ( .D(n4068), .CLK(wclk), .R(n13178), .S(1'b1), .Q(
        fifo[488]) );
  DFFSR fifo_reg_20__25_ ( .D(n4069), .CLK(wclk), .R(n13179), .S(1'b1), .Q(
        fifo[487]) );
  DFFSR fifo_reg_20__24_ ( .D(n4070), .CLK(wclk), .R(n13179), .S(1'b1), .Q(
        fifo[486]) );
  DFFSR fifo_reg_20__23_ ( .D(n4071), .CLK(wclk), .R(n13179), .S(1'b1), .Q(
        fifo[485]) );
  DFFSR fifo_reg_20__22_ ( .D(n4072), .CLK(wclk), .R(n13179), .S(1'b1), .Q(
        fifo[484]) );
  DFFSR fifo_reg_20__21_ ( .D(n4073), .CLK(wclk), .R(n13179), .S(1'b1), .Q(
        fifo[483]) );
  DFFSR fifo_reg_20__20_ ( .D(n4074), .CLK(wclk), .R(n13179), .S(1'b1), .Q(
        fifo[482]) );
  DFFSR fifo_reg_20__19_ ( .D(n4075), .CLK(wclk), .R(n13179), .S(1'b1), .Q(
        fifo[481]) );
  DFFSR fifo_reg_20__18_ ( .D(n4076), .CLK(wclk), .R(n13179), .S(1'b1), .Q(
        fifo[480]) );
  DFFSR fifo_reg_20__17_ ( .D(n4077), .CLK(wclk), .R(n13179), .S(1'b1), .Q(
        fifo[479]) );
  DFFSR fifo_reg_20__16_ ( .D(n4078), .CLK(wclk), .R(n13179), .S(1'b1), .Q(
        fifo[478]) );
  DFFSR fifo_reg_20__15_ ( .D(n4079), .CLK(wclk), .R(n13106), .S(1'b1), .Q(
        fifo[477]) );
  DFFSR fifo_reg_20__14_ ( .D(n4080), .CLK(wclk), .R(n13109), .S(1'b1), .Q(
        fifo[476]) );
  DFFSR fifo_reg_20__13_ ( .D(n4081), .CLK(wclk), .R(n13112), .S(1'b1), .Q(
        fifo[475]) );
  DFFSR fifo_reg_20__12_ ( .D(n4082), .CLK(wclk), .R(n13115), .S(1'b1), .Q(
        fifo[474]) );
  DFFSR fifo_reg_20__11_ ( .D(n4083), .CLK(wclk), .R(n13117), .S(1'b1), .Q(
        fifo[473]) );
  DFFSR fifo_reg_20__10_ ( .D(n4084), .CLK(wclk), .R(n13120), .S(1'b1), .Q(
        fifo[472]) );
  DFFSR fifo_reg_20__9_ ( .D(n4085), .CLK(wclk), .R(n13123), .S(1'b1), .Q(
        fifo[471]) );
  DFFSR fifo_reg_20__8_ ( .D(n4086), .CLK(wclk), .R(n13126), .S(1'b1), .Q(
        fifo[470]) );
  DFFSR fifo_reg_20__7_ ( .D(n4087), .CLK(wclk), .R(n13128), .S(1'b1), .Q(
        fifo[469]) );
  DFFSR fifo_reg_20__6_ ( .D(n4088), .CLK(wclk), .R(n13131), .S(1'b1), .Q(
        fifo[468]) );
  DFFSR fifo_reg_20__5_ ( .D(n4089), .CLK(wclk), .R(n13134), .S(1'b1), .Q(
        fifo[467]) );
  DFFSR fifo_reg_20__4_ ( .D(n4090), .CLK(wclk), .R(n13137), .S(1'b1), .Q(
        fifo[466]) );
  DFFSR fifo_reg_20__3_ ( .D(n4091), .CLK(wclk), .R(n13139), .S(1'b1), .Q(
        fifo[465]) );
  DFFSR fifo_reg_20__2_ ( .D(n4092), .CLK(wclk), .R(n13142), .S(1'b1), .Q(
        fifo[464]) );
  DFFSR fifo_reg_20__1_ ( .D(n4093), .CLK(wclk), .R(n13145), .S(1'b1), .Q(
        fifo[463]) );
  DFFSR fifo_reg_20__0_ ( .D(n4094), .CLK(wclk), .R(n13148), .S(1'b1), .Q(
        fifo[462]) );
  DFFSR fifo_reg_21__41_ ( .D(n4095), .CLK(wclk), .R(n13179), .S(1'b1), .Q(
        fifo[461]) );
  DFFSR fifo_reg_21__40_ ( .D(n4096), .CLK(wclk), .R(n13179), .S(1'b1), .Q(
        fifo[460]) );
  DFFSR fifo_reg_21__39_ ( .D(n4097), .CLK(wclk), .R(n13180), .S(1'b1), .Q(
        fifo[459]) );
  DFFSR fifo_reg_21__38_ ( .D(n4098), .CLK(wclk), .R(n13180), .S(1'b1), .Q(
        fifo[458]) );
  DFFSR fifo_reg_21__37_ ( .D(n4099), .CLK(wclk), .R(n13180), .S(1'b1), .Q(
        fifo[457]) );
  DFFSR fifo_reg_21__36_ ( .D(n4100), .CLK(wclk), .R(n13180), .S(1'b1), .Q(
        fifo[456]) );
  DFFSR fifo_reg_21__35_ ( .D(n4101), .CLK(wclk), .R(n13180), .S(1'b1), .Q(
        fifo[455]) );
  DFFSR fifo_reg_21__34_ ( .D(n4102), .CLK(wclk), .R(n13180), .S(1'b1), .Q(
        fifo[454]) );
  DFFSR fifo_reg_21__33_ ( .D(n4103), .CLK(wclk), .R(n13180), .S(1'b1), .Q(
        fifo[453]) );
  DFFSR fifo_reg_21__32_ ( .D(n4104), .CLK(wclk), .R(n13180), .S(1'b1), .Q(
        fifo[452]) );
  DFFSR fifo_reg_21__31_ ( .D(n4105), .CLK(wclk), .R(n13180), .S(1'b1), .Q(
        fifo[451]) );
  DFFSR fifo_reg_21__30_ ( .D(n4106), .CLK(wclk), .R(n13180), .S(1'b1), .Q(
        fifo[450]) );
  DFFSR fifo_reg_21__29_ ( .D(n4107), .CLK(wclk), .R(n13180), .S(1'b1), .Q(
        fifo[449]) );
  DFFSR fifo_reg_21__28_ ( .D(n4108), .CLK(wclk), .R(n13180), .S(1'b1), .Q(
        fifo[448]) );
  DFFSR fifo_reg_21__27_ ( .D(n4109), .CLK(wclk), .R(n13181), .S(1'b1), .Q(
        fifo[447]) );
  DFFSR fifo_reg_21__26_ ( .D(n4110), .CLK(wclk), .R(n13181), .S(1'b1), .Q(
        fifo[446]) );
  DFFSR fifo_reg_21__25_ ( .D(n4111), .CLK(wclk), .R(n13181), .S(1'b1), .Q(
        fifo[445]) );
  DFFSR fifo_reg_21__24_ ( .D(n4112), .CLK(wclk), .R(n13181), .S(1'b1), .Q(
        fifo[444]) );
  DFFSR fifo_reg_21__23_ ( .D(n4113), .CLK(wclk), .R(n13181), .S(1'b1), .Q(
        fifo[443]) );
  DFFSR fifo_reg_21__22_ ( .D(n4114), .CLK(wclk), .R(n13181), .S(1'b1), .Q(
        fifo[442]) );
  DFFSR fifo_reg_21__21_ ( .D(n4115), .CLK(wclk), .R(n13181), .S(1'b1), .Q(
        fifo[441]) );
  DFFSR fifo_reg_21__20_ ( .D(n4116), .CLK(wclk), .R(n13181), .S(1'b1), .Q(
        fifo[440]) );
  DFFSR fifo_reg_21__19_ ( .D(n4117), .CLK(wclk), .R(n13181), .S(1'b1), .Q(
        fifo[439]) );
  DFFSR fifo_reg_21__18_ ( .D(n4118), .CLK(wclk), .R(n13181), .S(1'b1), .Q(
        fifo[438]) );
  DFFSR fifo_reg_21__17_ ( .D(n4119), .CLK(wclk), .R(n13181), .S(1'b1), .Q(
        fifo[437]) );
  DFFSR fifo_reg_21__16_ ( .D(n4120), .CLK(wclk), .R(n13181), .S(1'b1), .Q(
        fifo[436]) );
  DFFSR fifo_reg_21__15_ ( .D(n4121), .CLK(wclk), .R(n13106), .S(1'b1), .Q(
        fifo[435]) );
  DFFSR fifo_reg_21__14_ ( .D(n4122), .CLK(wclk), .R(n13109), .S(1'b1), .Q(
        fifo[434]) );
  DFFSR fifo_reg_21__13_ ( .D(n4123), .CLK(wclk), .R(n13112), .S(1'b1), .Q(
        fifo[433]) );
  DFFSR fifo_reg_21__12_ ( .D(n4124), .CLK(wclk), .R(n13115), .S(1'b1), .Q(
        fifo[432]) );
  DFFSR fifo_reg_21__11_ ( .D(n4125), .CLK(wclk), .R(n13117), .S(1'b1), .Q(
        fifo[431]) );
  DFFSR fifo_reg_21__10_ ( .D(n4126), .CLK(wclk), .R(n13120), .S(1'b1), .Q(
        fifo[430]) );
  DFFSR fifo_reg_21__9_ ( .D(n4127), .CLK(wclk), .R(n13123), .S(1'b1), .Q(
        fifo[429]) );
  DFFSR fifo_reg_21__8_ ( .D(n4128), .CLK(wclk), .R(n13126), .S(1'b1), .Q(
        fifo[428]) );
  DFFSR fifo_reg_21__7_ ( .D(n4129), .CLK(wclk), .R(n13128), .S(1'b1), .Q(
        fifo[427]) );
  DFFSR fifo_reg_21__6_ ( .D(n4130), .CLK(wclk), .R(n13131), .S(1'b1), .Q(
        fifo[426]) );
  DFFSR fifo_reg_21__5_ ( .D(n4131), .CLK(wclk), .R(n13134), .S(1'b1), .Q(
        fifo[425]) );
  DFFSR fifo_reg_21__4_ ( .D(n4132), .CLK(wclk), .R(n13137), .S(1'b1), .Q(
        fifo[424]) );
  DFFSR fifo_reg_21__3_ ( .D(n4133), .CLK(wclk), .R(n13139), .S(1'b1), .Q(
        fifo[423]) );
  DFFSR fifo_reg_21__2_ ( .D(n4134), .CLK(wclk), .R(n13142), .S(1'b1), .Q(
        fifo[422]) );
  DFFSR fifo_reg_21__1_ ( .D(n4135), .CLK(wclk), .R(n13145), .S(1'b1), .Q(
        fifo[421]) );
  DFFSR fifo_reg_21__0_ ( .D(n4136), .CLK(wclk), .R(n13148), .S(1'b1), .Q(
        fifo[420]) );
  DFFSR fifo_reg_22__41_ ( .D(n4137), .CLK(wclk), .R(n13182), .S(1'b1), .Q(
        fifo[419]) );
  DFFSR fifo_reg_22__40_ ( .D(n4138), .CLK(wclk), .R(n13182), .S(1'b1), .Q(
        fifo[418]) );
  DFFSR fifo_reg_22__39_ ( .D(n4139), .CLK(wclk), .R(n13182), .S(1'b1), .Q(
        fifo[417]) );
  DFFSR fifo_reg_22__38_ ( .D(n4140), .CLK(wclk), .R(n13182), .S(1'b1), .Q(
        fifo[416]) );
  DFFSR fifo_reg_22__37_ ( .D(n4141), .CLK(wclk), .R(n13182), .S(1'b1), .Q(
        fifo[415]) );
  DFFSR fifo_reg_22__36_ ( .D(n4142), .CLK(wclk), .R(n13182), .S(1'b1), .Q(
        fifo[414]) );
  DFFSR fifo_reg_22__35_ ( .D(n4143), .CLK(wclk), .R(n13182), .S(1'b1), .Q(
        fifo[413]) );
  DFFSR fifo_reg_22__34_ ( .D(n4144), .CLK(wclk), .R(n13182), .S(1'b1), .Q(
        fifo[412]) );
  DFFSR fifo_reg_22__33_ ( .D(n4145), .CLK(wclk), .R(n13182), .S(1'b1), .Q(
        fifo[411]) );
  DFFSR fifo_reg_22__32_ ( .D(n4146), .CLK(wclk), .R(n13182), .S(1'b1), .Q(
        fifo[410]) );
  DFFSR fifo_reg_22__31_ ( .D(n4147), .CLK(wclk), .R(n13182), .S(1'b1), .Q(
        fifo[409]) );
  DFFSR fifo_reg_22__30_ ( .D(n4148), .CLK(wclk), .R(n13182), .S(1'b1), .Q(
        fifo[408]) );
  DFFSR fifo_reg_22__29_ ( .D(n4149), .CLK(wclk), .R(n13183), .S(1'b1), .Q(
        fifo[407]) );
  DFFSR fifo_reg_22__28_ ( .D(n4150), .CLK(wclk), .R(n13183), .S(1'b1), .Q(
        fifo[406]) );
  DFFSR fifo_reg_22__27_ ( .D(n4151), .CLK(wclk), .R(n13183), .S(1'b1), .Q(
        fifo[405]) );
  DFFSR fifo_reg_22__26_ ( .D(n4152), .CLK(wclk), .R(n13183), .S(1'b1), .Q(
        fifo[404]) );
  DFFSR fifo_reg_22__25_ ( .D(n4153), .CLK(wclk), .R(n13183), .S(1'b1), .Q(
        fifo[403]) );
  DFFSR fifo_reg_22__24_ ( .D(n4154), .CLK(wclk), .R(n13183), .S(1'b1), .Q(
        fifo[402]) );
  DFFSR fifo_reg_22__23_ ( .D(n4155), .CLK(wclk), .R(n13183), .S(1'b1), .Q(
        fifo[401]) );
  DFFSR fifo_reg_22__22_ ( .D(n4156), .CLK(wclk), .R(n13183), .S(1'b1), .Q(
        fifo[400]) );
  DFFSR fifo_reg_22__21_ ( .D(n4157), .CLK(wclk), .R(n13183), .S(1'b1), .Q(
        fifo[399]) );
  DFFSR fifo_reg_22__20_ ( .D(n4158), .CLK(wclk), .R(n13183), .S(1'b1), .Q(
        fifo[398]) );
  DFFSR fifo_reg_22__19_ ( .D(n4159), .CLK(wclk), .R(n13183), .S(1'b1), .Q(
        fifo[397]) );
  DFFSR fifo_reg_22__18_ ( .D(n4160), .CLK(wclk), .R(n13183), .S(1'b1), .Q(
        fifo[396]) );
  DFFSR fifo_reg_22__17_ ( .D(n4161), .CLK(wclk), .R(n13184), .S(1'b1), .Q(
        fifo[395]) );
  DFFSR fifo_reg_22__16_ ( .D(n4162), .CLK(wclk), .R(n13184), .S(1'b1), .Q(
        fifo[394]) );
  DFFSR fifo_reg_22__15_ ( .D(n4163), .CLK(wclk), .R(n13106), .S(1'b1), .Q(
        fifo[393]) );
  DFFSR fifo_reg_22__14_ ( .D(n4164), .CLK(wclk), .R(n13109), .S(1'b1), .Q(
        fifo[392]) );
  DFFSR fifo_reg_22__13_ ( .D(n4165), .CLK(wclk), .R(n13112), .S(1'b1), .Q(
        fifo[391]) );
  DFFSR fifo_reg_22__12_ ( .D(n4166), .CLK(wclk), .R(n13115), .S(1'b1), .Q(
        fifo[390]) );
  DFFSR fifo_reg_22__11_ ( .D(n4167), .CLK(wclk), .R(n13117), .S(1'b1), .Q(
        fifo[389]) );
  DFFSR fifo_reg_22__10_ ( .D(n4168), .CLK(wclk), .R(n13120), .S(1'b1), .Q(
        fifo[388]) );
  DFFSR fifo_reg_22__9_ ( .D(n4169), .CLK(wclk), .R(n13123), .S(1'b1), .Q(
        fifo[387]) );
  DFFSR fifo_reg_22__8_ ( .D(n4170), .CLK(wclk), .R(n13126), .S(1'b1), .Q(
        fifo[386]) );
  DFFSR fifo_reg_22__7_ ( .D(n4171), .CLK(wclk), .R(n13128), .S(1'b1), .Q(
        fifo[385]) );
  DFFSR fifo_reg_22__6_ ( .D(n4172), .CLK(wclk), .R(n13131), .S(1'b1), .Q(
        fifo[384]) );
  DFFSR fifo_reg_22__5_ ( .D(n4173), .CLK(wclk), .R(n13134), .S(1'b1), .Q(
        fifo[383]) );
  DFFSR fifo_reg_22__4_ ( .D(n4174), .CLK(wclk), .R(n13137), .S(1'b1), .Q(
        fifo[382]) );
  DFFSR fifo_reg_22__3_ ( .D(n4175), .CLK(wclk), .R(n13139), .S(1'b1), .Q(
        fifo[381]) );
  DFFSR fifo_reg_22__2_ ( .D(n4176), .CLK(wclk), .R(n13142), .S(1'b1), .Q(
        fifo[380]) );
  DFFSR fifo_reg_22__1_ ( .D(n4177), .CLK(wclk), .R(n13145), .S(1'b1), .Q(
        fifo[379]) );
  DFFSR fifo_reg_22__0_ ( .D(n4178), .CLK(wclk), .R(n13148), .S(1'b1), .Q(
        fifo[378]) );
  DFFSR fifo_reg_23__41_ ( .D(n4179), .CLK(wclk), .R(n13184), .S(1'b1), .Q(
        fifo[377]) );
  DFFSR fifo_reg_23__40_ ( .D(n4180), .CLK(wclk), .R(n13184), .S(1'b1), .Q(
        fifo[376]) );
  DFFSR fifo_reg_23__39_ ( .D(n4181), .CLK(wclk), .R(n13184), .S(1'b1), .Q(
        fifo[375]) );
  DFFSR fifo_reg_23__38_ ( .D(n4182), .CLK(wclk), .R(n13184), .S(1'b1), .Q(
        fifo[374]) );
  DFFSR fifo_reg_23__37_ ( .D(n4183), .CLK(wclk), .R(n13184), .S(1'b1), .Q(
        fifo[373]) );
  DFFSR fifo_reg_23__36_ ( .D(n4184), .CLK(wclk), .R(n13184), .S(1'b1), .Q(
        fifo[372]) );
  DFFSR fifo_reg_23__35_ ( .D(n4185), .CLK(wclk), .R(n13184), .S(1'b1), .Q(
        fifo[371]) );
  DFFSR fifo_reg_23__34_ ( .D(n4186), .CLK(wclk), .R(n13184), .S(1'b1), .Q(
        fifo[370]) );
  DFFSR fifo_reg_23__33_ ( .D(n4187), .CLK(wclk), .R(n13184), .S(1'b1), .Q(
        fifo[369]) );
  DFFSR fifo_reg_23__32_ ( .D(n4188), .CLK(wclk), .R(n13184), .S(1'b1), .Q(
        fifo[368]) );
  DFFSR fifo_reg_23__31_ ( .D(n4189), .CLK(wclk), .R(n13185), .S(1'b1), .Q(
        fifo[367]) );
  DFFSR fifo_reg_23__30_ ( .D(n4190), .CLK(wclk), .R(n13185), .S(1'b1), .Q(
        fifo[366]) );
  DFFSR fifo_reg_23__29_ ( .D(n4191), .CLK(wclk), .R(n13185), .S(1'b1), .Q(
        fifo[365]) );
  DFFSR fifo_reg_23__28_ ( .D(n4192), .CLK(wclk), .R(n13185), .S(1'b1), .Q(
        fifo[364]) );
  DFFSR fifo_reg_23__27_ ( .D(n4193), .CLK(wclk), .R(n13185), .S(1'b1), .Q(
        fifo[363]) );
  DFFSR fifo_reg_23__26_ ( .D(n4194), .CLK(wclk), .R(n13185), .S(1'b1), .Q(
        fifo[362]) );
  DFFSR fifo_reg_23__25_ ( .D(n4195), .CLK(wclk), .R(n13185), .S(1'b1), .Q(
        fifo[361]) );
  DFFSR fifo_reg_23__24_ ( .D(n4196), .CLK(wclk), .R(n13185), .S(1'b1), .Q(
        fifo[360]) );
  DFFSR fifo_reg_23__23_ ( .D(n4197), .CLK(wclk), .R(n13185), .S(1'b1), .Q(
        fifo[359]) );
  DFFSR fifo_reg_23__22_ ( .D(n4198), .CLK(wclk), .R(n13185), .S(1'b1), .Q(
        fifo[358]) );
  DFFSR fifo_reg_23__21_ ( .D(n4199), .CLK(wclk), .R(n13185), .S(1'b1), .Q(
        fifo[357]) );
  DFFSR fifo_reg_23__20_ ( .D(n4200), .CLK(wclk), .R(n13185), .S(1'b1), .Q(
        fifo[356]) );
  DFFSR fifo_reg_23__19_ ( .D(n4201), .CLK(wclk), .R(n13186), .S(1'b1), .Q(
        fifo[355]) );
  DFFSR fifo_reg_23__18_ ( .D(n4202), .CLK(wclk), .R(n13186), .S(1'b1), .Q(
        fifo[354]) );
  DFFSR fifo_reg_23__17_ ( .D(n4203), .CLK(wclk), .R(n13186), .S(1'b1), .Q(
        fifo[353]) );
  DFFSR fifo_reg_23__16_ ( .D(n4204), .CLK(wclk), .R(n13186), .S(1'b1), .Q(
        fifo[352]) );
  DFFSR fifo_reg_23__15_ ( .D(n4205), .CLK(wclk), .R(n13107), .S(1'b1), .Q(
        fifo[351]) );
  DFFSR fifo_reg_23__14_ ( .D(n4206), .CLK(wclk), .R(n13109), .S(1'b1), .Q(
        fifo[350]) );
  DFFSR fifo_reg_23__13_ ( .D(n4207), .CLK(wclk), .R(n13112), .S(1'b1), .Q(
        fifo[349]) );
  DFFSR fifo_reg_23__12_ ( .D(n4208), .CLK(wclk), .R(n13115), .S(1'b1), .Q(
        fifo[348]) );
  DFFSR fifo_reg_23__11_ ( .D(n4209), .CLK(wclk), .R(n13118), .S(1'b1), .Q(
        fifo[347]) );
  DFFSR fifo_reg_23__10_ ( .D(n4210), .CLK(wclk), .R(n13120), .S(1'b1), .Q(
        fifo[346]) );
  DFFSR fifo_reg_23__9_ ( .D(n4211), .CLK(wclk), .R(n13123), .S(1'b1), .Q(
        fifo[345]) );
  DFFSR fifo_reg_23__8_ ( .D(n4212), .CLK(wclk), .R(n13126), .S(1'b1), .Q(
        fifo[344]) );
  DFFSR fifo_reg_23__7_ ( .D(n4213), .CLK(wclk), .R(n13129), .S(1'b1), .Q(
        fifo[343]) );
  DFFSR fifo_reg_23__6_ ( .D(n4214), .CLK(wclk), .R(n13131), .S(1'b1), .Q(
        fifo[342]) );
  DFFSR fifo_reg_23__5_ ( .D(n4215), .CLK(wclk), .R(n13134), .S(1'b1), .Q(
        fifo[341]) );
  DFFSR fifo_reg_23__4_ ( .D(n4216), .CLK(wclk), .R(n13137), .S(1'b1), .Q(
        fifo[340]) );
  DFFSR fifo_reg_23__3_ ( .D(n4217), .CLK(wclk), .R(n13140), .S(1'b1), .Q(
        fifo[339]) );
  DFFSR fifo_reg_23__2_ ( .D(n4218), .CLK(wclk), .R(n13142), .S(1'b1), .Q(
        fifo[338]) );
  DFFSR fifo_reg_23__1_ ( .D(n4219), .CLK(wclk), .R(n13145), .S(1'b1), .Q(
        fifo[337]) );
  DFFSR fifo_reg_23__0_ ( .D(n4220), .CLK(wclk), .R(n13148), .S(1'b1), .Q(
        fifo[336]) );
  DFFSR fifo_reg_24__41_ ( .D(n4221), .CLK(wclk), .R(n13151), .S(1'b1), .Q(
        fifo[335]) );
  DFFSR fifo_reg_24__40_ ( .D(n4222), .CLK(wclk), .R(n13151), .S(1'b1), .Q(
        fifo[334]) );
  DFFSR fifo_reg_24__39_ ( .D(n4223), .CLK(wclk), .R(n13151), .S(1'b1), .Q(
        fifo[333]) );
  DFFSR fifo_reg_24__38_ ( .D(n4224), .CLK(wclk), .R(n13151), .S(1'b1), .Q(
        fifo[332]) );
  DFFSR fifo_reg_24__37_ ( .D(n4225), .CLK(wclk), .R(n13152), .S(1'b1), .Q(
        fifo[331]) );
  DFFSR fifo_reg_24__36_ ( .D(n4226), .CLK(wclk), .R(n13152), .S(1'b1), .Q(
        fifo[330]) );
  DFFSR fifo_reg_24__35_ ( .D(n4227), .CLK(wclk), .R(n13152), .S(1'b1), .Q(
        fifo[329]) );
  DFFSR fifo_reg_24__34_ ( .D(n4228), .CLK(wclk), .R(n13152), .S(1'b1), .Q(
        fifo[328]) );
  DFFSR fifo_reg_24__33_ ( .D(n4229), .CLK(wclk), .R(n13152), .S(1'b1), .Q(
        fifo[327]) );
  DFFSR fifo_reg_24__32_ ( .D(n4230), .CLK(wclk), .R(n13152), .S(1'b1), .Q(
        fifo[326]) );
  DFFSR fifo_reg_24__31_ ( .D(n4231), .CLK(wclk), .R(n13152), .S(1'b1), .Q(
        fifo[325]) );
  DFFSR fifo_reg_24__30_ ( .D(n4232), .CLK(wclk), .R(n13152), .S(1'b1), .Q(
        fifo[324]) );
  DFFSR fifo_reg_24__29_ ( .D(n4233), .CLK(wclk), .R(n13152), .S(1'b1), .Q(
        fifo[323]) );
  DFFSR fifo_reg_24__28_ ( .D(n4234), .CLK(wclk), .R(n13152), .S(1'b1), .Q(
        fifo[322]) );
  DFFSR fifo_reg_24__27_ ( .D(n4235), .CLK(wclk), .R(n13152), .S(1'b1), .Q(
        fifo[321]) );
  DFFSR fifo_reg_24__26_ ( .D(n4236), .CLK(wclk), .R(n13152), .S(1'b1), .Q(
        fifo[320]) );
  DFFSR fifo_reg_24__25_ ( .D(n4237), .CLK(wclk), .R(n13153), .S(1'b1), .Q(
        fifo[319]) );
  DFFSR fifo_reg_24__24_ ( .D(n4238), .CLK(wclk), .R(n13153), .S(1'b1), .Q(
        fifo[318]) );
  DFFSR fifo_reg_24__23_ ( .D(n4239), .CLK(wclk), .R(n13153), .S(1'b1), .Q(
        fifo[317]) );
  DFFSR fifo_reg_24__22_ ( .D(n4240), .CLK(wclk), .R(n13153), .S(1'b1), .Q(
        fifo[316]) );
  DFFSR fifo_reg_24__21_ ( .D(n4241), .CLK(wclk), .R(n13153), .S(1'b1), .Q(
        fifo[315]) );
  DFFSR fifo_reg_24__20_ ( .D(n4242), .CLK(wclk), .R(n13153), .S(1'b1), .Q(
        fifo[314]) );
  DFFSR fifo_reg_24__19_ ( .D(n4243), .CLK(wclk), .R(n13153), .S(1'b1), .Q(
        fifo[313]) );
  DFFSR fifo_reg_24__18_ ( .D(n4244), .CLK(wclk), .R(n13153), .S(1'b1), .Q(
        fifo[312]) );
  DFFSR fifo_reg_24__17_ ( .D(n4245), .CLK(wclk), .R(n13153), .S(1'b1), .Q(
        fifo[311]) );
  DFFSR fifo_reg_24__16_ ( .D(n4246), .CLK(wclk), .R(n13153), .S(1'b1), .Q(
        fifo[310]) );
  DFFSR fifo_reg_24__15_ ( .D(n4247), .CLK(wclk), .R(n13107), .S(1'b1), .Q(
        fifo[309]) );
  DFFSR fifo_reg_24__14_ ( .D(n4248), .CLK(wclk), .R(n13109), .S(1'b1), .Q(
        fifo[308]) );
  DFFSR fifo_reg_24__13_ ( .D(n4249), .CLK(wclk), .R(n13112), .S(1'b1), .Q(
        fifo[307]) );
  DFFSR fifo_reg_24__12_ ( .D(n4250), .CLK(wclk), .R(n13115), .S(1'b1), .Q(
        fifo[306]) );
  DFFSR fifo_reg_24__11_ ( .D(n4251), .CLK(wclk), .R(n13118), .S(1'b1), .Q(
        fifo[305]) );
  DFFSR fifo_reg_24__10_ ( .D(n4252), .CLK(wclk), .R(n13120), .S(1'b1), .Q(
        fifo[304]) );
  DFFSR fifo_reg_24__9_ ( .D(n4253), .CLK(wclk), .R(n13123), .S(1'b1), .Q(
        fifo[303]) );
  DFFSR fifo_reg_24__8_ ( .D(n4254), .CLK(wclk), .R(n13126), .S(1'b1), .Q(
        fifo[302]) );
  DFFSR fifo_reg_24__7_ ( .D(n4255), .CLK(wclk), .R(n13129), .S(1'b1), .Q(
        fifo[301]) );
  DFFSR fifo_reg_24__6_ ( .D(n4256), .CLK(wclk), .R(n13131), .S(1'b1), .Q(
        fifo[300]) );
  DFFSR fifo_reg_24__5_ ( .D(n4257), .CLK(wclk), .R(n13134), .S(1'b1), .Q(
        fifo[299]) );
  DFFSR fifo_reg_24__4_ ( .D(n4258), .CLK(wclk), .R(n13137), .S(1'b1), .Q(
        fifo[298]) );
  DFFSR fifo_reg_24__3_ ( .D(n4259), .CLK(wclk), .R(n13140), .S(1'b1), .Q(
        fifo[297]) );
  DFFSR fifo_reg_24__2_ ( .D(n4260), .CLK(wclk), .R(n13142), .S(1'b1), .Q(
        fifo[296]) );
  DFFSR fifo_reg_24__1_ ( .D(n4261), .CLK(wclk), .R(n13145), .S(1'b1), .Q(
        fifo[295]) );
  DFFSR fifo_reg_24__0_ ( .D(n4262), .CLK(wclk), .R(n13148), .S(1'b1), .Q(
        fifo[294]) );
  DFFSR fifo_reg_25__41_ ( .D(n4263), .CLK(wclk), .R(n13153), .S(1'b1), .Q(
        fifo[293]) );
  DFFSR fifo_reg_25__40_ ( .D(n4264), .CLK(wclk), .R(n13153), .S(1'b1), .Q(
        fifo[292]) );
  DFFSR fifo_reg_25__39_ ( .D(n4265), .CLK(wclk), .R(n13154), .S(1'b1), .Q(
        fifo[291]) );
  DFFSR fifo_reg_25__38_ ( .D(n4266), .CLK(wclk), .R(n13154), .S(1'b1), .Q(
        fifo[290]) );
  DFFSR fifo_reg_25__37_ ( .D(n4267), .CLK(wclk), .R(n13154), .S(1'b1), .Q(
        fifo[289]) );
  DFFSR fifo_reg_25__36_ ( .D(n4268), .CLK(wclk), .R(n13154), .S(1'b1), .Q(
        fifo[288]) );
  DFFSR fifo_reg_25__35_ ( .D(n4269), .CLK(wclk), .R(n13154), .S(1'b1), .Q(
        fifo[287]) );
  DFFSR fifo_reg_25__34_ ( .D(n4270), .CLK(wclk), .R(n13154), .S(1'b1), .Q(
        fifo[286]) );
  DFFSR fifo_reg_25__33_ ( .D(n4271), .CLK(wclk), .R(n13154), .S(1'b1), .Q(
        fifo[285]) );
  DFFSR fifo_reg_25__32_ ( .D(n4272), .CLK(wclk), .R(n13154), .S(1'b1), .Q(
        fifo[284]) );
  DFFSR fifo_reg_25__31_ ( .D(n4273), .CLK(wclk), .R(n13154), .S(1'b1), .Q(
        fifo[283]) );
  DFFSR fifo_reg_25__30_ ( .D(n4274), .CLK(wclk), .R(n13154), .S(1'b1), .Q(
        fifo[282]) );
  DFFSR fifo_reg_25__29_ ( .D(n4275), .CLK(wclk), .R(n13154), .S(1'b1), .Q(
        fifo[281]) );
  DFFSR fifo_reg_25__28_ ( .D(n4276), .CLK(wclk), .R(n13154), .S(1'b1), .Q(
        fifo[280]) );
  DFFSR fifo_reg_25__27_ ( .D(n4277), .CLK(wclk), .R(n13155), .S(1'b1), .Q(
        fifo[279]) );
  DFFSR fifo_reg_25__26_ ( .D(n4278), .CLK(wclk), .R(n13155), .S(1'b1), .Q(
        fifo[278]) );
  DFFSR fifo_reg_25__25_ ( .D(n4279), .CLK(wclk), .R(n13155), .S(1'b1), .Q(
        fifo[277]) );
  DFFSR fifo_reg_25__24_ ( .D(n4280), .CLK(wclk), .R(n13155), .S(1'b1), .Q(
        fifo[276]) );
  DFFSR fifo_reg_25__23_ ( .D(n4281), .CLK(wclk), .R(n13155), .S(1'b1), .Q(
        fifo[275]) );
  DFFSR fifo_reg_25__22_ ( .D(n4282), .CLK(wclk), .R(n13155), .S(1'b1), .Q(
        fifo[274]) );
  DFFSR fifo_reg_25__21_ ( .D(n4283), .CLK(wclk), .R(n13155), .S(1'b1), .Q(
        fifo[273]) );
  DFFSR fifo_reg_25__20_ ( .D(n4284), .CLK(wclk), .R(n13155), .S(1'b1), .Q(
        fifo[272]) );
  DFFSR fifo_reg_25__19_ ( .D(n4285), .CLK(wclk), .R(n13155), .S(1'b1), .Q(
        fifo[271]) );
  DFFSR fifo_reg_25__18_ ( .D(n4286), .CLK(wclk), .R(n13155), .S(1'b1), .Q(
        fifo[270]) );
  DFFSR fifo_reg_25__17_ ( .D(n4287), .CLK(wclk), .R(n13155), .S(1'b1), .Q(
        fifo[269]) );
  DFFSR fifo_reg_25__16_ ( .D(n4288), .CLK(wclk), .R(n13155), .S(1'b1), .Q(
        fifo[268]) );
  DFFSR fifo_reg_25__15_ ( .D(n4289), .CLK(wclk), .R(n13107), .S(1'b1), .Q(
        fifo[267]) );
  DFFSR fifo_reg_25__14_ ( .D(n4290), .CLK(wclk), .R(n13109), .S(1'b1), .Q(
        fifo[266]) );
  DFFSR fifo_reg_25__13_ ( .D(n4291), .CLK(wclk), .R(n13112), .S(1'b1), .Q(
        fifo[265]) );
  DFFSR fifo_reg_25__12_ ( .D(n4292), .CLK(wclk), .R(n13115), .S(1'b1), .Q(
        fifo[264]) );
  DFFSR fifo_reg_25__11_ ( .D(n4293), .CLK(wclk), .R(n13118), .S(1'b1), .Q(
        fifo[263]) );
  DFFSR fifo_reg_25__10_ ( .D(n4294), .CLK(wclk), .R(n13120), .S(1'b1), .Q(
        fifo[262]) );
  DFFSR fifo_reg_25__9_ ( .D(n4295), .CLK(wclk), .R(n13123), .S(1'b1), .Q(
        fifo[261]) );
  DFFSR fifo_reg_25__8_ ( .D(n4296), .CLK(wclk), .R(n13126), .S(1'b1), .Q(
        fifo[260]) );
  DFFSR fifo_reg_25__7_ ( .D(n4297), .CLK(wclk), .R(n13129), .S(1'b1), .Q(
        fifo[259]) );
  DFFSR fifo_reg_25__6_ ( .D(n4298), .CLK(wclk), .R(n13131), .S(1'b1), .Q(
        fifo[258]) );
  DFFSR fifo_reg_25__5_ ( .D(n4299), .CLK(wclk), .R(n13134), .S(1'b1), .Q(
        fifo[257]) );
  DFFSR fifo_reg_25__4_ ( .D(n4300), .CLK(wclk), .R(n13137), .S(1'b1), .Q(
        fifo[256]) );
  DFFSR fifo_reg_25__3_ ( .D(n4301), .CLK(wclk), .R(n13140), .S(1'b1), .Q(
        fifo[255]) );
  DFFSR fifo_reg_25__2_ ( .D(n4302), .CLK(wclk), .R(n13142), .S(1'b1), .Q(
        fifo[254]) );
  DFFSR fifo_reg_25__1_ ( .D(n4303), .CLK(wclk), .R(n13145), .S(1'b1), .Q(
        fifo[253]) );
  DFFSR fifo_reg_25__0_ ( .D(n4304), .CLK(wclk), .R(n13148), .S(1'b1), .Q(
        fifo[252]) );
  DFFSR fifo_reg_26__41_ ( .D(n4305), .CLK(wclk), .R(n13156), .S(1'b1), .Q(
        fifo[251]) );
  DFFSR fifo_reg_26__40_ ( .D(n4306), .CLK(wclk), .R(n13156), .S(1'b1), .Q(
        fifo[250]) );
  DFFSR fifo_reg_26__39_ ( .D(n4307), .CLK(wclk), .R(n13156), .S(1'b1), .Q(
        fifo[249]) );
  DFFSR fifo_reg_26__38_ ( .D(n4308), .CLK(wclk), .R(n13156), .S(1'b1), .Q(
        fifo[248]) );
  DFFSR fifo_reg_26__37_ ( .D(n4309), .CLK(wclk), .R(n13156), .S(1'b1), .Q(
        fifo[247]) );
  DFFSR fifo_reg_26__36_ ( .D(n4310), .CLK(wclk), .R(n13156), .S(1'b1), .Q(
        fifo[246]) );
  DFFSR fifo_reg_26__35_ ( .D(n4311), .CLK(wclk), .R(n13156), .S(1'b1), .Q(
        fifo[245]) );
  DFFSR fifo_reg_26__34_ ( .D(n4312), .CLK(wclk), .R(n13156), .S(1'b1), .Q(
        fifo[244]) );
  DFFSR fifo_reg_26__33_ ( .D(n4313), .CLK(wclk), .R(n13156), .S(1'b1), .Q(
        fifo[243]) );
  DFFSR fifo_reg_26__32_ ( .D(n4314), .CLK(wclk), .R(n13156), .S(1'b1), .Q(
        fifo[242]) );
  DFFSR fifo_reg_26__31_ ( .D(n4315), .CLK(wclk), .R(n13156), .S(1'b1), .Q(
        fifo[241]) );
  DFFSR fifo_reg_26__30_ ( .D(n4316), .CLK(wclk), .R(n13156), .S(1'b1), .Q(
        fifo[240]) );
  DFFSR fifo_reg_26__29_ ( .D(n4317), .CLK(wclk), .R(n13157), .S(1'b1), .Q(
        fifo[239]) );
  DFFSR fifo_reg_26__28_ ( .D(n4318), .CLK(wclk), .R(n13157), .S(1'b1), .Q(
        fifo[238]) );
  DFFSR fifo_reg_26__27_ ( .D(n4319), .CLK(wclk), .R(n13157), .S(1'b1), .Q(
        fifo[237]) );
  DFFSR fifo_reg_26__26_ ( .D(n4320), .CLK(wclk), .R(n13157), .S(1'b1), .Q(
        fifo[236]) );
  DFFSR fifo_reg_26__25_ ( .D(n4321), .CLK(wclk), .R(n13157), .S(1'b1), .Q(
        fifo[235]) );
  DFFSR fifo_reg_26__24_ ( .D(n4322), .CLK(wclk), .R(n13157), .S(1'b1), .Q(
        fifo[234]) );
  DFFSR fifo_reg_26__23_ ( .D(n4323), .CLK(wclk), .R(n13157), .S(1'b1), .Q(
        fifo[233]) );
  DFFSR fifo_reg_26__22_ ( .D(n4324), .CLK(wclk), .R(n13157), .S(1'b1), .Q(
        fifo[232]) );
  DFFSR fifo_reg_26__21_ ( .D(n4325), .CLK(wclk), .R(n13157), .S(1'b1), .Q(
        fifo[231]) );
  DFFSR fifo_reg_26__20_ ( .D(n4326), .CLK(wclk), .R(n13157), .S(1'b1), .Q(
        fifo[230]) );
  DFFSR fifo_reg_26__19_ ( .D(n4327), .CLK(wclk), .R(n13157), .S(1'b1), .Q(
        fifo[229]) );
  DFFSR fifo_reg_26__18_ ( .D(n4328), .CLK(wclk), .R(n13157), .S(1'b1), .Q(
        fifo[228]) );
  DFFSR fifo_reg_26__17_ ( .D(n4329), .CLK(wclk), .R(n13158), .S(1'b1), .Q(
        fifo[227]) );
  DFFSR fifo_reg_26__16_ ( .D(n4330), .CLK(wclk), .R(n13158), .S(1'b1), .Q(
        fifo[226]) );
  DFFSR fifo_reg_26__15_ ( .D(n4331), .CLK(wclk), .R(n13107), .S(1'b1), .Q(
        fifo[225]) );
  DFFSR fifo_reg_26__14_ ( .D(n4332), .CLK(wclk), .R(n13110), .S(1'b1), .Q(
        fifo[224]) );
  DFFSR fifo_reg_26__13_ ( .D(n4333), .CLK(wclk), .R(n13112), .S(1'b1), .Q(
        fifo[223]) );
  DFFSR fifo_reg_26__12_ ( .D(n4334), .CLK(wclk), .R(n13115), .S(1'b1), .Q(
        fifo[222]) );
  DFFSR fifo_reg_26__11_ ( .D(n4335), .CLK(wclk), .R(n13118), .S(1'b1), .Q(
        fifo[221]) );
  DFFSR fifo_reg_26__10_ ( .D(n4336), .CLK(wclk), .R(n13121), .S(1'b1), .Q(
        fifo[220]) );
  DFFSR fifo_reg_26__9_ ( .D(n4337), .CLK(wclk), .R(n13123), .S(1'b1), .Q(
        fifo[219]) );
  DFFSR fifo_reg_26__8_ ( .D(n4338), .CLK(wclk), .R(n13126), .S(1'b1), .Q(
        fifo[218]) );
  DFFSR fifo_reg_26__7_ ( .D(n4339), .CLK(wclk), .R(n13129), .S(1'b1), .Q(
        fifo[217]) );
  DFFSR fifo_reg_26__6_ ( .D(n4340), .CLK(wclk), .R(n13132), .S(1'b1), .Q(
        fifo[216]) );
  DFFSR fifo_reg_26__5_ ( .D(n4341), .CLK(wclk), .R(n13134), .S(1'b1), .Q(
        fifo[215]) );
  DFFSR fifo_reg_26__4_ ( .D(n4342), .CLK(wclk), .R(n13137), .S(1'b1), .Q(
        fifo[214]) );
  DFFSR fifo_reg_26__3_ ( .D(n4343), .CLK(wclk), .R(n13140), .S(1'b1), .Q(
        fifo[213]) );
  DFFSR fifo_reg_26__2_ ( .D(n4344), .CLK(wclk), .R(n13143), .S(1'b1), .Q(
        fifo[212]) );
  DFFSR fifo_reg_26__1_ ( .D(n4345), .CLK(wclk), .R(n13145), .S(1'b1), .Q(
        fifo[211]) );
  DFFSR fifo_reg_26__0_ ( .D(n4346), .CLK(wclk), .R(n13148), .S(1'b1), .Q(
        fifo[210]) );
  DFFSR fifo_reg_27__41_ ( .D(n4347), .CLK(wclk), .R(n13158), .S(1'b1), .Q(
        fifo[209]) );
  DFFSR fifo_reg_27__40_ ( .D(n4348), .CLK(wclk), .R(n13158), .S(1'b1), .Q(
        fifo[208]) );
  DFFSR fifo_reg_27__39_ ( .D(n4349), .CLK(wclk), .R(n13158), .S(1'b1), .Q(
        fifo[207]) );
  DFFSR fifo_reg_27__38_ ( .D(n4350), .CLK(wclk), .R(n13158), .S(1'b1), .Q(
        fifo[206]) );
  DFFSR fifo_reg_27__37_ ( .D(n4351), .CLK(wclk), .R(n13158), .S(1'b1), .Q(
        fifo[205]) );
  DFFSR fifo_reg_27__36_ ( .D(n4352), .CLK(wclk), .R(n13158), .S(1'b1), .Q(
        fifo[204]) );
  DFFSR fifo_reg_27__35_ ( .D(n4353), .CLK(wclk), .R(n13158), .S(1'b1), .Q(
        fifo[203]) );
  DFFSR fifo_reg_27__34_ ( .D(n4354), .CLK(wclk), .R(n13158), .S(1'b1), .Q(
        fifo[202]) );
  DFFSR fifo_reg_27__33_ ( .D(n4355), .CLK(wclk), .R(n13158), .S(1'b1), .Q(
        fifo[201]) );
  DFFSR fifo_reg_27__32_ ( .D(n4356), .CLK(wclk), .R(n13158), .S(1'b1), .Q(
        fifo[200]) );
  DFFSR fifo_reg_27__31_ ( .D(n4357), .CLK(wclk), .R(n13159), .S(1'b1), .Q(
        fifo[199]) );
  DFFSR fifo_reg_27__30_ ( .D(n4358), .CLK(wclk), .R(n13159), .S(1'b1), .Q(
        fifo[198]) );
  DFFSR fifo_reg_27__29_ ( .D(n4359), .CLK(wclk), .R(n13159), .S(1'b1), .Q(
        fifo[197]) );
  DFFSR fifo_reg_27__28_ ( .D(n4360), .CLK(wclk), .R(n13159), .S(1'b1), .Q(
        fifo[196]) );
  DFFSR fifo_reg_27__27_ ( .D(n4361), .CLK(wclk), .R(n13159), .S(1'b1), .Q(
        fifo[195]) );
  DFFSR fifo_reg_27__26_ ( .D(n4362), .CLK(wclk), .R(n13159), .S(1'b1), .Q(
        fifo[194]) );
  DFFSR fifo_reg_27__25_ ( .D(n4363), .CLK(wclk), .R(n13159), .S(1'b1), .Q(
        fifo[193]) );
  DFFSR fifo_reg_27__24_ ( .D(n4364), .CLK(wclk), .R(n13159), .S(1'b1), .Q(
        fifo[192]) );
  DFFSR fifo_reg_27__23_ ( .D(n4365), .CLK(wclk), .R(n13159), .S(1'b1), .Q(
        fifo[191]) );
  DFFSR fifo_reg_27__22_ ( .D(n4366), .CLK(wclk), .R(n13159), .S(1'b1), .Q(
        fifo[190]) );
  DFFSR fifo_reg_27__21_ ( .D(n4367), .CLK(wclk), .R(n13159), .S(1'b1), .Q(
        fifo[189]) );
  DFFSR fifo_reg_27__20_ ( .D(n4368), .CLK(wclk), .R(n13159), .S(1'b1), .Q(
        fifo[188]) );
  DFFSR fifo_reg_27__19_ ( .D(n4369), .CLK(wclk), .R(n13160), .S(1'b1), .Q(
        fifo[187]) );
  DFFSR fifo_reg_27__18_ ( .D(n4370), .CLK(wclk), .R(n13160), .S(1'b1), .Q(
        fifo[186]) );
  DFFSR fifo_reg_27__17_ ( .D(n4371), .CLK(wclk), .R(n13160), .S(1'b1), .Q(
        fifo[185]) );
  DFFSR fifo_reg_27__16_ ( .D(n4372), .CLK(wclk), .R(n13160), .S(1'b1), .Q(
        fifo[184]) );
  DFFSR fifo_reg_27__15_ ( .D(n4373), .CLK(wclk), .R(n13107), .S(1'b1), .Q(
        fifo[183]) );
  DFFSR fifo_reg_27__14_ ( .D(n4374), .CLK(wclk), .R(n13110), .S(1'b1), .Q(
        fifo[182]) );
  DFFSR fifo_reg_27__13_ ( .D(n4375), .CLK(wclk), .R(n13112), .S(1'b1), .Q(
        fifo[181]) );
  DFFSR fifo_reg_27__12_ ( .D(n4376), .CLK(wclk), .R(n13115), .S(1'b1), .Q(
        fifo[180]) );
  DFFSR fifo_reg_27__11_ ( .D(n4377), .CLK(wclk), .R(n13118), .S(1'b1), .Q(
        fifo[179]) );
  DFFSR fifo_reg_27__10_ ( .D(n4378), .CLK(wclk), .R(n13121), .S(1'b1), .Q(
        fifo[178]) );
  DFFSR fifo_reg_27__9_ ( .D(n4379), .CLK(wclk), .R(n13123), .S(1'b1), .Q(
        fifo[177]) );
  DFFSR fifo_reg_27__8_ ( .D(n4380), .CLK(wclk), .R(n13126), .S(1'b1), .Q(
        fifo[176]) );
  DFFSR fifo_reg_27__7_ ( .D(n4381), .CLK(wclk), .R(n13129), .S(1'b1), .Q(
        fifo[175]) );
  DFFSR fifo_reg_27__6_ ( .D(n4382), .CLK(wclk), .R(n13132), .S(1'b1), .Q(
        fifo[174]) );
  DFFSR fifo_reg_27__5_ ( .D(n4383), .CLK(wclk), .R(n13134), .S(1'b1), .Q(
        fifo[173]) );
  DFFSR fifo_reg_27__4_ ( .D(n4384), .CLK(wclk), .R(n13137), .S(1'b1), .Q(
        fifo[172]) );
  DFFSR fifo_reg_27__3_ ( .D(n4385), .CLK(wclk), .R(n13140), .S(1'b1), .Q(
        fifo[171]) );
  DFFSR fifo_reg_27__2_ ( .D(n4386), .CLK(wclk), .R(n13143), .S(1'b1), .Q(
        fifo[170]) );
  DFFSR fifo_reg_27__1_ ( .D(n4387), .CLK(wclk), .R(n13145), .S(1'b1), .Q(
        fifo[169]) );
  DFFSR fifo_reg_27__0_ ( .D(n4388), .CLK(wclk), .R(n13148), .S(1'b1), .Q(
        fifo[168]) );
  DFFSR fifo_reg_28__41_ ( .D(n4389), .CLK(wclk), .R(n13160), .S(1'b1), .Q(
        fifo[167]) );
  DFFSR fifo_reg_28__40_ ( .D(n4390), .CLK(wclk), .R(n13160), .S(1'b1), .Q(
        fifo[166]) );
  DFFSR fifo_reg_28__39_ ( .D(n4391), .CLK(wclk), .R(n13160), .S(1'b1), .Q(
        fifo[165]) );
  DFFSR fifo_reg_28__38_ ( .D(n4392), .CLK(wclk), .R(n13160), .S(1'b1), .Q(
        fifo[164]) );
  DFFSR fifo_reg_28__37_ ( .D(n4393), .CLK(wclk), .R(n13160), .S(1'b1), .Q(
        fifo[163]) );
  DFFSR fifo_reg_28__36_ ( .D(n4394), .CLK(wclk), .R(n13160), .S(1'b1), .Q(
        fifo[162]) );
  DFFSR fifo_reg_28__35_ ( .D(n4395), .CLK(wclk), .R(n13160), .S(1'b1), .Q(
        fifo[161]) );
  DFFSR fifo_reg_28__34_ ( .D(n4396), .CLK(wclk), .R(n13160), .S(1'b1), .Q(
        fifo[160]) );
  DFFSR fifo_reg_28__33_ ( .D(n4397), .CLK(wclk), .R(n13161), .S(1'b1), .Q(
        fifo[159]) );
  DFFSR fifo_reg_28__32_ ( .D(n4398), .CLK(wclk), .R(n13161), .S(1'b1), .Q(
        fifo[158]) );
  DFFSR fifo_reg_28__31_ ( .D(n4399), .CLK(wclk), .R(n13161), .S(1'b1), .Q(
        fifo[157]) );
  DFFSR fifo_reg_28__30_ ( .D(n4400), .CLK(wclk), .R(n13161), .S(1'b1), .Q(
        fifo[156]) );
  DFFSR fifo_reg_28__29_ ( .D(n4401), .CLK(wclk), .R(n13161), .S(1'b1), .Q(
        fifo[155]) );
  DFFSR fifo_reg_28__28_ ( .D(n4402), .CLK(wclk), .R(n13161), .S(1'b1), .Q(
        fifo[154]) );
  DFFSR fifo_reg_28__27_ ( .D(n4403), .CLK(wclk), .R(n13161), .S(1'b1), .Q(
        fifo[153]) );
  DFFSR fifo_reg_28__26_ ( .D(n4404), .CLK(wclk), .R(n13161), .S(1'b1), .Q(
        fifo[152]) );
  DFFSR fifo_reg_28__25_ ( .D(n4405), .CLK(wclk), .R(n13161), .S(1'b1), .Q(
        fifo[151]) );
  DFFSR fifo_reg_28__24_ ( .D(n4406), .CLK(wclk), .R(n13161), .S(1'b1), .Q(
        fifo[150]) );
  DFFSR fifo_reg_28__23_ ( .D(n4407), .CLK(wclk), .R(n13161), .S(1'b1), .Q(
        fifo[149]) );
  DFFSR fifo_reg_28__22_ ( .D(n4408), .CLK(wclk), .R(n13161), .S(1'b1), .Q(
        fifo[148]) );
  DFFSR fifo_reg_28__21_ ( .D(n4409), .CLK(wclk), .R(n13162), .S(1'b1), .Q(
        fifo[147]) );
  DFFSR fifo_reg_28__20_ ( .D(n4410), .CLK(wclk), .R(n13162), .S(1'b1), .Q(
        fifo[146]) );
  DFFSR fifo_reg_28__19_ ( .D(n4411), .CLK(wclk), .R(n13162), .S(1'b1), .Q(
        fifo[145]) );
  DFFSR fifo_reg_28__18_ ( .D(n4412), .CLK(wclk), .R(n13162), .S(1'b1), .Q(
        fifo[144]) );
  DFFSR fifo_reg_28__17_ ( .D(n4413), .CLK(wclk), .R(n13162), .S(1'b1), .Q(
        fifo[143]) );
  DFFSR fifo_reg_28__16_ ( .D(n4414), .CLK(wclk), .R(n13162), .S(1'b1), .Q(
        fifo[142]) );
  DFFSR fifo_reg_28__15_ ( .D(n4415), .CLK(wclk), .R(n13107), .S(1'b1), .Q(
        fifo[141]) );
  DFFSR fifo_reg_28__14_ ( .D(n4416), .CLK(wclk), .R(n13110), .S(1'b1), .Q(
        fifo[140]) );
  DFFSR fifo_reg_28__13_ ( .D(n4417), .CLK(wclk), .R(n13112), .S(1'b1), .Q(
        fifo[139]) );
  DFFSR fifo_reg_28__12_ ( .D(n4418), .CLK(wclk), .R(n13115), .S(1'b1), .Q(
        fifo[138]) );
  DFFSR fifo_reg_28__11_ ( .D(n4419), .CLK(wclk), .R(n13118), .S(1'b1), .Q(
        fifo[137]) );
  DFFSR fifo_reg_28__10_ ( .D(n4420), .CLK(wclk), .R(n13121), .S(1'b1), .Q(
        fifo[136]) );
  DFFSR fifo_reg_28__9_ ( .D(n4421), .CLK(wclk), .R(n13123), .S(1'b1), .Q(
        fifo[135]) );
  DFFSR fifo_reg_28__8_ ( .D(n4422), .CLK(wclk), .R(n13126), .S(1'b1), .Q(
        fifo[134]) );
  DFFSR fifo_reg_28__7_ ( .D(n4423), .CLK(wclk), .R(n13129), .S(1'b1), .Q(
        fifo[133]) );
  DFFSR fifo_reg_28__6_ ( .D(n4424), .CLK(wclk), .R(n13132), .S(1'b1), .Q(
        fifo[132]) );
  DFFSR fifo_reg_28__5_ ( .D(n4425), .CLK(wclk), .R(n13134), .S(1'b1), .Q(
        fifo[131]) );
  DFFSR fifo_reg_28__4_ ( .D(n4426), .CLK(wclk), .R(n13137), .S(1'b1), .Q(
        fifo[130]) );
  DFFSR fifo_reg_28__3_ ( .D(n4427), .CLK(wclk), .R(n13140), .S(1'b1), .Q(
        fifo[129]) );
  DFFSR fifo_reg_28__2_ ( .D(n4428), .CLK(wclk), .R(n13143), .S(1'b1), .Q(
        fifo[128]) );
  DFFSR fifo_reg_28__1_ ( .D(n4429), .CLK(wclk), .R(n13145), .S(1'b1), .Q(
        fifo[127]) );
  DFFSR fifo_reg_28__0_ ( .D(n4430), .CLK(wclk), .R(n13148), .S(1'b1), .Q(
        fifo[126]) );
  DFFSR fifo_reg_29__41_ ( .D(n4431), .CLK(wclk), .R(n13162), .S(1'b1), .Q(
        fifo[125]) );
  DFFSR fifo_reg_29__40_ ( .D(n4432), .CLK(wclk), .R(n13162), .S(1'b1), .Q(
        fifo[124]) );
  DFFSR fifo_reg_29__39_ ( .D(n4433), .CLK(wclk), .R(n13162), .S(1'b1), .Q(
        fifo[123]) );
  DFFSR fifo_reg_29__38_ ( .D(n4434), .CLK(wclk), .R(n13162), .S(1'b1), .Q(
        fifo[122]) );
  DFFSR fifo_reg_29__37_ ( .D(n4435), .CLK(wclk), .R(n13162), .S(1'b1), .Q(
        fifo[121]) );
  DFFSR fifo_reg_29__36_ ( .D(n4436), .CLK(wclk), .R(n13162), .S(1'b1), .Q(
        fifo[120]) );
  DFFSR fifo_reg_29__35_ ( .D(n4437), .CLK(wclk), .R(n13163), .S(1'b1), .Q(
        fifo[119]) );
  DFFSR fifo_reg_29__34_ ( .D(n4438), .CLK(wclk), .R(n13163), .S(1'b1), .Q(
        fifo[118]) );
  DFFSR fifo_reg_29__33_ ( .D(n4439), .CLK(wclk), .R(n13163), .S(1'b1), .Q(
        fifo[117]) );
  DFFSR fifo_reg_29__32_ ( .D(n4440), .CLK(wclk), .R(n13163), .S(1'b1), .Q(
        fifo[116]) );
  DFFSR fifo_reg_29__31_ ( .D(n4441), .CLK(wclk), .R(n13163), .S(1'b1), .Q(
        fifo[115]) );
  DFFSR fifo_reg_29__30_ ( .D(n4442), .CLK(wclk), .R(n13163), .S(1'b1), .Q(
        fifo[114]) );
  DFFSR fifo_reg_29__29_ ( .D(n4443), .CLK(wclk), .R(n13163), .S(1'b1), .Q(
        fifo[113]) );
  DFFSR fifo_reg_29__28_ ( .D(n4444), .CLK(wclk), .R(n13163), .S(1'b1), .Q(
        fifo[112]) );
  DFFSR fifo_reg_29__27_ ( .D(n4445), .CLK(wclk), .R(n13163), .S(1'b1), .Q(
        fifo[111]) );
  DFFSR fifo_reg_29__26_ ( .D(n4446), .CLK(wclk), .R(n13163), .S(1'b1), .Q(
        fifo[110]) );
  DFFSR fifo_reg_29__25_ ( .D(n4447), .CLK(wclk), .R(n13163), .S(1'b1), .Q(
        fifo[109]) );
  DFFSR fifo_reg_29__24_ ( .D(n4448), .CLK(wclk), .R(n13163), .S(1'b1), .Q(
        fifo[108]) );
  DFFSR fifo_reg_29__23_ ( .D(n4449), .CLK(wclk), .R(n13164), .S(1'b1), .Q(
        fifo[107]) );
  DFFSR fifo_reg_29__22_ ( .D(n4450), .CLK(wclk), .R(n13164), .S(1'b1), .Q(
        fifo[106]) );
  DFFSR fifo_reg_29__21_ ( .D(n4451), .CLK(wclk), .R(n13164), .S(1'b1), .Q(
        fifo[105]) );
  DFFSR fifo_reg_29__20_ ( .D(n4452), .CLK(wclk), .R(n13164), .S(1'b1), .Q(
        fifo[104]) );
  DFFSR fifo_reg_29__19_ ( .D(n4453), .CLK(wclk), .R(n13164), .S(1'b1), .Q(
        fifo[103]) );
  DFFSR fifo_reg_29__18_ ( .D(n4454), .CLK(wclk), .R(n13164), .S(1'b1), .Q(
        fifo[102]) );
  DFFSR fifo_reg_29__17_ ( .D(n4455), .CLK(wclk), .R(n13164), .S(1'b1), .Q(
        fifo[101]) );
  DFFSR fifo_reg_29__16_ ( .D(n4456), .CLK(wclk), .R(n13164), .S(1'b1), .Q(
        fifo[100]) );
  DFFSR fifo_reg_29__15_ ( .D(n4457), .CLK(wclk), .R(n13107), .S(1'b1), .Q(
        fifo[99]) );
  DFFSR fifo_reg_29__14_ ( .D(n4458), .CLK(wclk), .R(n13110), .S(1'b1), .Q(
        fifo[98]) );
  DFFSR fifo_reg_29__13_ ( .D(n4459), .CLK(wclk), .R(n13113), .S(1'b1), .Q(
        fifo[97]) );
  DFFSR fifo_reg_29__12_ ( .D(n4460), .CLK(wclk), .R(n13115), .S(1'b1), .Q(
        fifo[96]) );
  DFFSR fifo_reg_29__11_ ( .D(n4461), .CLK(wclk), .R(n13118), .S(1'b1), .Q(
        fifo[95]) );
  DFFSR fifo_reg_29__10_ ( .D(n4462), .CLK(wclk), .R(n13121), .S(1'b1), .Q(
        fifo[94]) );
  DFFSR fifo_reg_29__9_ ( .D(n4463), .CLK(wclk), .R(n13124), .S(1'b1), .Q(
        fifo[93]) );
  DFFSR fifo_reg_29__8_ ( .D(n4464), .CLK(wclk), .R(n13126), .S(1'b1), .Q(
        fifo[92]) );
  DFFSR fifo_reg_29__7_ ( .D(n4465), .CLK(wclk), .R(n13129), .S(1'b1), .Q(
        fifo[91]) );
  DFFSR fifo_reg_29__6_ ( .D(n4466), .CLK(wclk), .R(n13132), .S(1'b1), .Q(
        fifo[90]) );
  DFFSR fifo_reg_29__5_ ( .D(n4467), .CLK(wclk), .R(n13135), .S(1'b1), .Q(
        fifo[89]) );
  DFFSR fifo_reg_29__4_ ( .D(n4468), .CLK(wclk), .R(n13137), .S(1'b1), .Q(
        fifo[88]) );
  DFFSR fifo_reg_29__3_ ( .D(n4469), .CLK(wclk), .R(n13140), .S(1'b1), .Q(
        fifo[87]) );
  DFFSR fifo_reg_29__2_ ( .D(n4470), .CLK(wclk), .R(n13143), .S(1'b1), .Q(
        fifo[86]) );
  DFFSR fifo_reg_29__1_ ( .D(n4471), .CLK(wclk), .R(n13146), .S(1'b1), .Q(
        fifo[85]) );
  DFFSR fifo_reg_29__0_ ( .D(n4472), .CLK(wclk), .R(n13148), .S(1'b1), .Q(
        fifo[84]) );
  DFFSR fifo_reg_30__41_ ( .D(n4473), .CLK(wclk), .R(n13164), .S(1'b1), .Q(
        fifo[83]) );
  DFFSR fifo_reg_30__40_ ( .D(n4474), .CLK(wclk), .R(n13164), .S(1'b1), .Q(
        fifo[82]) );
  DFFSR fifo_reg_30__39_ ( .D(n4475), .CLK(wclk), .R(n13164), .S(1'b1), .Q(
        fifo[81]) );
  DFFSR fifo_reg_30__38_ ( .D(n4476), .CLK(wclk), .R(n13164), .S(1'b1), .Q(
        fifo[80]) );
  DFFSR fifo_reg_30__37_ ( .D(n4477), .CLK(wclk), .R(n13165), .S(1'b1), .Q(
        fifo[79]) );
  DFFSR fifo_reg_30__36_ ( .D(n4478), .CLK(wclk), .R(n13165), .S(1'b1), .Q(
        fifo[78]) );
  DFFSR fifo_reg_30__35_ ( .D(n4479), .CLK(wclk), .R(n13165), .S(1'b1), .Q(
        fifo[77]) );
  DFFSR fifo_reg_30__34_ ( .D(n4480), .CLK(wclk), .R(n13165), .S(1'b1), .Q(
        fifo[76]) );
  DFFSR fifo_reg_30__33_ ( .D(n4481), .CLK(wclk), .R(n13165), .S(1'b1), .Q(
        fifo[75]) );
  DFFSR fifo_reg_30__32_ ( .D(n4482), .CLK(wclk), .R(n13165), .S(1'b1), .Q(
        fifo[74]) );
  DFFSR fifo_reg_30__31_ ( .D(n4483), .CLK(wclk), .R(n13165), .S(1'b1), .Q(
        fifo[73]) );
  DFFSR fifo_reg_30__30_ ( .D(n4484), .CLK(wclk), .R(n13165), .S(1'b1), .Q(
        fifo[72]) );
  DFFSR fifo_reg_30__29_ ( .D(n4485), .CLK(wclk), .R(n13165), .S(1'b1), .Q(
        fifo[71]) );
  DFFSR fifo_reg_30__28_ ( .D(n4486), .CLK(wclk), .R(n13165), .S(1'b1), .Q(
        fifo[70]) );
  DFFSR fifo_reg_30__27_ ( .D(n4487), .CLK(wclk), .R(n13165), .S(1'b1), .Q(
        fifo[69]) );
  DFFSR fifo_reg_30__26_ ( .D(n4488), .CLK(wclk), .R(n13165), .S(1'b1), .Q(
        fifo[68]) );
  DFFSR fifo_reg_30__25_ ( .D(n4489), .CLK(wclk), .R(n13166), .S(1'b1), .Q(
        fifo[67]) );
  DFFSR fifo_reg_30__24_ ( .D(n4490), .CLK(wclk), .R(n13166), .S(1'b1), .Q(
        fifo[66]) );
  DFFSR fifo_reg_30__23_ ( .D(n4491), .CLK(wclk), .R(n13166), .S(1'b1), .Q(
        fifo[65]) );
  DFFSR fifo_reg_30__22_ ( .D(n4492), .CLK(wclk), .R(n13166), .S(1'b1), .Q(
        fifo[64]) );
  DFFSR fifo_reg_30__21_ ( .D(n4493), .CLK(wclk), .R(n13166), .S(1'b1), .Q(
        fifo[63]) );
  DFFSR fifo_reg_30__20_ ( .D(n4494), .CLK(wclk), .R(n13166), .S(1'b1), .Q(
        fifo[62]) );
  DFFSR fifo_reg_30__19_ ( .D(n4495), .CLK(wclk), .R(n13166), .S(1'b1), .Q(
        fifo[61]) );
  DFFSR fifo_reg_30__18_ ( .D(n4496), .CLK(wclk), .R(n13166), .S(1'b1), .Q(
        fifo[60]) );
  DFFSR fifo_reg_30__17_ ( .D(n4497), .CLK(wclk), .R(n13166), .S(1'b1), .Q(
        fifo[59]) );
  DFFSR fifo_reg_30__16_ ( .D(n4498), .CLK(wclk), .R(n13166), .S(1'b1), .Q(
        fifo[58]) );
  DFFSR fifo_reg_30__15_ ( .D(n4499), .CLK(wclk), .R(n13107), .S(1'b1), .Q(
        fifo[57]) );
  DFFSR fifo_reg_30__14_ ( .D(n4500), .CLK(wclk), .R(n13110), .S(1'b1), .Q(
        fifo[56]) );
  DFFSR fifo_reg_30__13_ ( .D(n4501), .CLK(wclk), .R(n13113), .S(1'b1), .Q(
        fifo[55]) );
  DFFSR fifo_reg_30__12_ ( .D(n4502), .CLK(wclk), .R(n13115), .S(1'b1), .Q(
        fifo[54]) );
  DFFSR fifo_reg_30__11_ ( .D(n4503), .CLK(wclk), .R(n13118), .S(1'b1), .Q(
        fifo[53]) );
  DFFSR fifo_reg_30__10_ ( .D(n4504), .CLK(wclk), .R(n13121), .S(1'b1), .Q(
        fifo[52]) );
  DFFSR fifo_reg_30__9_ ( .D(n4505), .CLK(wclk), .R(n13124), .S(1'b1), .Q(
        fifo[51]) );
  DFFSR fifo_reg_30__8_ ( .D(n4506), .CLK(wclk), .R(n13126), .S(1'b1), .Q(
        fifo[50]) );
  DFFSR fifo_reg_30__7_ ( .D(n4507), .CLK(wclk), .R(n13129), .S(1'b1), .Q(
        fifo[49]) );
  DFFSR fifo_reg_30__6_ ( .D(n4508), .CLK(wclk), .R(n13132), .S(1'b1), .Q(
        fifo[48]) );
  DFFSR fifo_reg_30__5_ ( .D(n4509), .CLK(wclk), .R(n13135), .S(1'b1), .Q(
        fifo[47]) );
  DFFSR fifo_reg_30__4_ ( .D(n4510), .CLK(wclk), .R(n13137), .S(1'b1), .Q(
        fifo[46]) );
  DFFSR fifo_reg_30__3_ ( .D(n4511), .CLK(wclk), .R(n13140), .S(1'b1), .Q(
        fifo[45]) );
  DFFSR fifo_reg_30__2_ ( .D(n4512), .CLK(wclk), .R(n13143), .S(1'b1), .Q(
        fifo[44]) );
  DFFSR fifo_reg_30__1_ ( .D(n4513), .CLK(wclk), .R(n13146), .S(1'b1), .Q(
        fifo[43]) );
  DFFSR fifo_reg_30__0_ ( .D(n4514), .CLK(wclk), .R(n13148), .S(1'b1), .Q(
        fifo[42]) );
  DFFSR fifo_reg_31__41_ ( .D(n4515), .CLK(wclk), .R(n13166), .S(1'b1), .Q(
        fifo[41]) );
  DFFSR fifo_reg_31__40_ ( .D(n4516), .CLK(wclk), .R(n13166), .S(1'b1), .Q(
        fifo[40]) );
  DFFSR fifo_reg_31__39_ ( .D(n4517), .CLK(wclk), .R(n13167), .S(1'b1), .Q(
        fifo[39]) );
  DFFSR fifo_reg_31__38_ ( .D(n4518), .CLK(wclk), .R(n13167), .S(1'b1), .Q(
        fifo[38]) );
  DFFSR fifo_reg_31__37_ ( .D(n4519), .CLK(wclk), .R(n13167), .S(1'b1), .Q(
        fifo[37]) );
  DFFSR fifo_reg_31__36_ ( .D(n4520), .CLK(wclk), .R(n13167), .S(1'b1), .Q(
        fifo[36]) );
  DFFSR fifo_reg_31__35_ ( .D(n4521), .CLK(wclk), .R(n13167), .S(1'b1), .Q(
        fifo[35]) );
  DFFSR fifo_reg_31__34_ ( .D(n4522), .CLK(wclk), .R(n13167), .S(1'b1), .Q(
        fifo[34]) );
  DFFSR fifo_reg_31__33_ ( .D(n4523), .CLK(wclk), .R(n13167), .S(1'b1), .Q(
        fifo[33]) );
  DFFSR fifo_reg_31__32_ ( .D(n4524), .CLK(wclk), .R(n13167), .S(1'b1), .Q(
        fifo[32]) );
  DFFSR fifo_reg_31__31_ ( .D(n4525), .CLK(wclk), .R(n13167), .S(1'b1), .Q(
        fifo[31]) );
  DFFSR fifo_reg_31__30_ ( .D(n4526), .CLK(wclk), .R(n13167), .S(1'b1), .Q(
        fifo[30]) );
  DFFSR fifo_reg_31__29_ ( .D(n4527), .CLK(wclk), .R(n13167), .S(1'b1), .Q(
        fifo[29]) );
  DFFSR fifo_reg_31__28_ ( .D(n4528), .CLK(wclk), .R(n13167), .S(1'b1), .Q(
        fifo[28]) );
  DFFSR fifo_reg_31__27_ ( .D(n4529), .CLK(wclk), .R(n13168), .S(1'b1), .Q(
        fifo[27]) );
  DFFSR fifo_reg_31__26_ ( .D(n4530), .CLK(wclk), .R(n13168), .S(1'b1), .Q(
        fifo[26]) );
  DFFSR fifo_reg_31__25_ ( .D(n4531), .CLK(wclk), .R(n13168), .S(1'b1), .Q(
        fifo[25]) );
  DFFSR fifo_reg_31__24_ ( .D(n4532), .CLK(wclk), .R(n13168), .S(1'b1), .Q(
        fifo[24]) );
  DFFSR fifo_reg_31__23_ ( .D(n4533), .CLK(wclk), .R(n13168), .S(1'b1), .Q(
        fifo[23]) );
  DFFSR fifo_reg_31__22_ ( .D(n4534), .CLK(wclk), .R(n13168), .S(1'b1), .Q(
        fifo[22]) );
  DFFSR fifo_reg_31__21_ ( .D(n4535), .CLK(wclk), .R(n13168), .S(1'b1), .Q(
        fifo[21]) );
  DFFSR fifo_reg_31__20_ ( .D(n4536), .CLK(wclk), .R(n13168), .S(1'b1), .Q(
        fifo[20]) );
  DFFSR fifo_reg_31__19_ ( .D(n4537), .CLK(wclk), .R(n13168), .S(1'b1), .Q(
        fifo[19]) );
  DFFSR fifo_reg_31__18_ ( .D(n4538), .CLK(wclk), .R(n13168), .S(1'b1), .Q(
        fifo[18]) );
  DFFSR fifo_reg_31__17_ ( .D(n4539), .CLK(wclk), .R(n13168), .S(1'b1), .Q(
        fifo[17]) );
  DFFSR fifo_reg_31__16_ ( .D(n4540), .CLK(wclk), .R(n13168), .S(1'b1), .Q(
        fifo[16]) );
  DFFSR fifo_reg_31__15_ ( .D(n4541), .CLK(wclk), .R(n13107), .S(1'b1), .Q(
        fifo[15]) );
  DFFSR fifo_reg_31__14_ ( .D(n4542), .CLK(wclk), .R(n13110), .S(1'b1), .Q(
        fifo[14]) );
  DFFSR fifo_reg_31__13_ ( .D(n4543), .CLK(wclk), .R(n13113), .S(1'b1), .Q(
        fifo[13]) );
  DFFSR fifo_reg_31__12_ ( .D(n4544), .CLK(wclk), .R(n13115), .S(1'b1), .Q(
        fifo[12]) );
  DFFSR fifo_reg_31__11_ ( .D(n4545), .CLK(wclk), .R(n13118), .S(1'b1), .Q(
        fifo[11]) );
  DFFSR fifo_reg_31__10_ ( .D(n4546), .CLK(wclk), .R(n13121), .S(1'b1), .Q(
        fifo[10]) );
  DFFSR fifo_reg_31__9_ ( .D(n4547), .CLK(wclk), .R(n13124), .S(1'b1), .Q(
        fifo[9]) );
  DFFSR fifo_reg_31__8_ ( .D(n4548), .CLK(wclk), .R(n13126), .S(1'b1), .Q(
        fifo[8]) );
  DFFSR fifo_reg_31__7_ ( .D(n4549), .CLK(wclk), .R(n13129), .S(1'b1), .Q(
        fifo[7]) );
  DFFSR fifo_reg_31__6_ ( .D(n4550), .CLK(wclk), .R(n13132), .S(1'b1), .Q(
        fifo[6]) );
  DFFSR fifo_reg_31__5_ ( .D(n4551), .CLK(wclk), .R(n13135), .S(1'b1), .Q(
        fifo[5]) );
  DFFSR fifo_reg_31__4_ ( .D(n4552), .CLK(wclk), .R(n13137), .S(1'b1), .Q(
        fifo[4]) );
  DFFSR fifo_reg_31__3_ ( .D(n4553), .CLK(wclk), .R(n13140), .S(1'b1), .Q(
        fifo[3]) );
  DFFSR fifo_reg_31__2_ ( .D(n4554), .CLK(wclk), .R(n13143), .S(1'b1), .Q(
        fifo[2]) );
  DFFSR fifo_reg_31__1_ ( .D(n4555), .CLK(wclk), .R(n13146), .S(1'b1), .Q(
        fifo[1]) );
  DFFSR fifo_reg_31__0_ ( .D(n4556), .CLK(wclk), .R(n13148), .S(1'b1), .Q(
        fifo[0]) );
  OAI21X1 U9 ( .A(n201), .B(n202), .C(n8625), .Y(n3072) );
  INVX1 U11 ( .A(n13101), .Y(n202) );
  OAI21X1 U12 ( .A(n201), .B(n204), .C(n8622), .Y(n3077) );
  INVX1 U14 ( .A(n13104), .Y(n204) );
  OAI21X1 U15 ( .A(n201), .B(n13276), .C(n8619), .Y(n3082) );
  OAI21X1 U17 ( .A(n201), .B(n13304), .C(n8616), .Y(n3087) );
  INVX1 U19 ( .A(n210), .Y(n3089) );
  AOI22X1 U20 ( .A(data_out[41]), .B(n13047), .C(n71), .D(n201), .Y(n210) );
  INVX1 U21 ( .A(n212), .Y(n3091) );
  AOI22X1 U22 ( .A(data_out[40]), .B(n13047), .C(n72), .D(n201), .Y(n212) );
  INVX1 U23 ( .A(n213), .Y(n3093) );
  AOI22X1 U24 ( .A(data_out[39]), .B(n13047), .C(n73), .D(n201), .Y(n213) );
  INVX1 U25 ( .A(n214), .Y(n3095) );
  AOI22X1 U26 ( .A(data_out[38]), .B(n13047), .C(n74), .D(n201), .Y(n214) );
  INVX1 U27 ( .A(n215), .Y(n3097) );
  AOI22X1 U28 ( .A(data_out[37]), .B(n13047), .C(n75), .D(n201), .Y(n215) );
  INVX1 U29 ( .A(n216), .Y(n3099) );
  AOI22X1 U30 ( .A(data_out[36]), .B(n13047), .C(n76), .D(n201), .Y(n216) );
  INVX1 U31 ( .A(n217), .Y(n3101) );
  AOI22X1 U32 ( .A(data_out[35]), .B(n13047), .C(n77), .D(n201), .Y(n217) );
  INVX1 U33 ( .A(n218), .Y(n3103) );
  AOI22X1 U34 ( .A(data_out[34]), .B(n13047), .C(n78), .D(n201), .Y(n218) );
  INVX1 U35 ( .A(n219), .Y(n3105) );
  AOI22X1 U36 ( .A(data_out[33]), .B(n13047), .C(n79), .D(n201), .Y(n219) );
  INVX1 U37 ( .A(n220), .Y(n3107) );
  AOI22X1 U38 ( .A(data_out[32]), .B(n13047), .C(n80), .D(n201), .Y(n220) );
  INVX1 U39 ( .A(n221), .Y(n3109) );
  AOI22X1 U40 ( .A(data_out[31]), .B(n13047), .C(n81), .D(n201), .Y(n221) );
  INVX1 U41 ( .A(n222), .Y(n3111) );
  AOI22X1 U42 ( .A(data_out[30]), .B(n13047), .C(n82), .D(n201), .Y(n222) );
  INVX1 U43 ( .A(n223), .Y(n3113) );
  AOI22X1 U44 ( .A(data_out[29]), .B(n13047), .C(n83), .D(n201), .Y(n223) );
  INVX1 U45 ( .A(n224), .Y(n3115) );
  AOI22X1 U46 ( .A(data_out[28]), .B(n13047), .C(n84), .D(n201), .Y(n224) );
  INVX1 U47 ( .A(n225), .Y(n3117) );
  AOI22X1 U48 ( .A(data_out[27]), .B(n13047), .C(n85), .D(n201), .Y(n225) );
  INVX1 U49 ( .A(n226), .Y(n3119) );
  AOI22X1 U50 ( .A(data_out[26]), .B(n13047), .C(n86), .D(n201), .Y(n226) );
  INVX1 U51 ( .A(n227), .Y(n3121) );
  AOI22X1 U52 ( .A(data_out[25]), .B(n13047), .C(n87), .D(n201), .Y(n227) );
  INVX1 U53 ( .A(n228), .Y(n3123) );
  AOI22X1 U54 ( .A(data_out[24]), .B(n13047), .C(n88), .D(n201), .Y(n228) );
  INVX1 U55 ( .A(n229), .Y(n3125) );
  AOI22X1 U56 ( .A(data_out[23]), .B(n13047), .C(n89), .D(n201), .Y(n229) );
  INVX1 U57 ( .A(n230), .Y(n3127) );
  AOI22X1 U58 ( .A(data_out[22]), .B(n13047), .C(n90), .D(n201), .Y(n230) );
  INVX1 U59 ( .A(n231), .Y(n3129) );
  AOI22X1 U60 ( .A(data_out[21]), .B(n13047), .C(n91), .D(n201), .Y(n231) );
  INVX1 U61 ( .A(n232), .Y(n3131) );
  AOI22X1 U62 ( .A(data_out[20]), .B(n13047), .C(n92), .D(n201), .Y(n232) );
  INVX1 U63 ( .A(n233), .Y(n3133) );
  AOI22X1 U64 ( .A(data_out[19]), .B(n13047), .C(n93), .D(n201), .Y(n233) );
  INVX1 U65 ( .A(n234), .Y(n3135) );
  AOI22X1 U66 ( .A(data_out[18]), .B(n13047), .C(n94), .D(n201), .Y(n234) );
  INVX1 U67 ( .A(n235), .Y(n3137) );
  AOI22X1 U68 ( .A(data_out[17]), .B(n13047), .C(n95), .D(n201), .Y(n235) );
  INVX1 U69 ( .A(n236), .Y(n3139) );
  AOI22X1 U70 ( .A(data_out[16]), .B(n13047), .C(n96), .D(n201), .Y(n236) );
  INVX1 U71 ( .A(n237), .Y(n3141) );
  AOI22X1 U72 ( .A(data_out[15]), .B(n13047), .C(n97), .D(n201), .Y(n237) );
  INVX1 U73 ( .A(n238), .Y(n3143) );
  AOI22X1 U74 ( .A(data_out[14]), .B(n13047), .C(n98), .D(n201), .Y(n238) );
  INVX1 U75 ( .A(n239), .Y(n3145) );
  AOI22X1 U76 ( .A(data_out[13]), .B(n13047), .C(n99), .D(n201), .Y(n239) );
  INVX1 U77 ( .A(n240), .Y(n3147) );
  AOI22X1 U78 ( .A(data_out[12]), .B(n13047), .C(n100), .D(n201), .Y(n240) );
  INVX1 U79 ( .A(n241), .Y(n3149) );
  AOI22X1 U80 ( .A(data_out[11]), .B(n13047), .C(n101), .D(n201), .Y(n241) );
  INVX1 U81 ( .A(n242), .Y(n3151) );
  AOI22X1 U82 ( .A(data_out[10]), .B(n13047), .C(n102), .D(n201), .Y(n242) );
  INVX1 U83 ( .A(n243), .Y(n3153) );
  AOI22X1 U84 ( .A(data_out[9]), .B(n13047), .C(n103), .D(n201), .Y(n243) );
  INVX1 U85 ( .A(n244), .Y(n3155) );
  AOI22X1 U86 ( .A(data_out[8]), .B(n13047), .C(n104), .D(n201), .Y(n244) );
  INVX1 U87 ( .A(n245), .Y(n3157) );
  AOI22X1 U88 ( .A(data_out[7]), .B(n13047), .C(n105), .D(n201), .Y(n245) );
  INVX1 U89 ( .A(n246), .Y(n3159) );
  AOI22X1 U90 ( .A(data_out[6]), .B(n13047), .C(n106), .D(n201), .Y(n246) );
  INVX1 U91 ( .A(n247), .Y(n3161) );
  AOI22X1 U92 ( .A(data_out[5]), .B(n13047), .C(n107), .D(n201), .Y(n247) );
  INVX1 U93 ( .A(n248), .Y(n3163) );
  AOI22X1 U94 ( .A(data_out[4]), .B(n13047), .C(n108), .D(n201), .Y(n248) );
  INVX1 U95 ( .A(n249), .Y(n3165) );
  AOI22X1 U96 ( .A(data_out[3]), .B(n13047), .C(n109), .D(n201), .Y(n249) );
  INVX1 U97 ( .A(n250), .Y(n3167) );
  AOI22X1 U98 ( .A(data_out[2]), .B(n13047), .C(n110), .D(n201), .Y(n250) );
  INVX1 U99 ( .A(n251), .Y(n3169) );
  AOI22X1 U100 ( .A(data_out[1]), .B(n13047), .C(n111), .D(n201), .Y(n251) );
  INVX1 U101 ( .A(n252), .Y(n3171) );
  AOI22X1 U102 ( .A(data_out[0]), .B(n13047), .C(n112), .D(n201), .Y(n252) );
  OAI21X1 U103 ( .A(n253), .B(n254), .C(n8613), .Y(n3179) );
  OAI21X1 U105 ( .A(n253), .B(n256), .C(n8610), .Y(n3184) );
  OAI21X1 U107 ( .A(n253), .B(n258), .C(n8607), .Y(n3189) );
  OAI21X1 U109 ( .A(n253), .B(n260), .C(n8604), .Y(n3194) );
  OAI21X1 U111 ( .A(n253), .B(n262), .C(n4560), .Y(n3196) );
  OAI21X1 U113 ( .A(n253), .B(n264), .C(n8601), .Y(n3201) );
  INVX1 U115 ( .A(n12994), .Y(n264) );
  OAI21X1 U116 ( .A(n201), .B(n266), .C(n8598), .Y(n3209) );
  INVX1 U118 ( .A(reset), .Y(n3210) );
  OAI21X1 U119 ( .A(n201), .B(n13356), .C(n8595), .Y(n3212) );
  INVX1 U121 ( .A(n13047), .Y(n201) );
  OAI21X1 U123 ( .A(n270), .B(n271), .C(n8592), .Y(n3213) );
  OAI21X1 U125 ( .A(n270), .B(n273), .C(n8589), .Y(n3214) );
  OAI21X1 U127 ( .A(n270), .B(n275), .C(n8586), .Y(n3215) );
  OAI21X1 U129 ( .A(n270), .B(n277), .C(n8583), .Y(n3216) );
  OAI21X1 U131 ( .A(n270), .B(n279), .C(n8580), .Y(n3217) );
  OAI21X1 U133 ( .A(n270), .B(n281), .C(n8577), .Y(n3218) );
  OAI21X1 U135 ( .A(n270), .B(n283), .C(n8574), .Y(n3219) );
  OAI21X1 U137 ( .A(n270), .B(n285), .C(n8571), .Y(n3220) );
  OAI21X1 U139 ( .A(n270), .B(n287), .C(n8568), .Y(n3221) );
  OAI21X1 U141 ( .A(n270), .B(n289), .C(n8565), .Y(n3222) );
  OAI21X1 U143 ( .A(n270), .B(n291), .C(n8562), .Y(n3223) );
  OAI21X1 U145 ( .A(n270), .B(n293), .C(n8559), .Y(n3224) );
  OAI21X1 U147 ( .A(n270), .B(n295), .C(n8556), .Y(n3225) );
  OAI21X1 U149 ( .A(n270), .B(n297), .C(n8553), .Y(n3226) );
  OAI21X1 U151 ( .A(n270), .B(n299), .C(n8550), .Y(n3227) );
  OAI21X1 U153 ( .A(n270), .B(n301), .C(n8547), .Y(n3228) );
  OAI21X1 U155 ( .A(n270), .B(n303), .C(n8544), .Y(n3229) );
  OAI21X1 U157 ( .A(n270), .B(n305), .C(n8541), .Y(n3230) );
  OAI21X1 U159 ( .A(n270), .B(n307), .C(n8538), .Y(n3231) );
  OAI21X1 U161 ( .A(n270), .B(n309), .C(n8535), .Y(n3232) );
  OAI21X1 U163 ( .A(n270), .B(n311), .C(n8532), .Y(n3233) );
  OAI21X1 U165 ( .A(n270), .B(n313), .C(n8529), .Y(n3234) );
  OAI21X1 U167 ( .A(n270), .B(n315), .C(n8526), .Y(n3235) );
  OAI21X1 U169 ( .A(n270), .B(n317), .C(n8523), .Y(n3236) );
  OAI21X1 U171 ( .A(n270), .B(n319), .C(n8520), .Y(n3237) );
  OAI21X1 U173 ( .A(n270), .B(n321), .C(n8517), .Y(n3238) );
  OAI21X1 U175 ( .A(n270), .B(n323), .C(n8514), .Y(n3239) );
  OAI21X1 U177 ( .A(n270), .B(n325), .C(n8511), .Y(n3240) );
  OAI21X1 U179 ( .A(n270), .B(n327), .C(n8508), .Y(n3241) );
  OAI21X1 U181 ( .A(n270), .B(n329), .C(n8505), .Y(n3242) );
  OAI21X1 U183 ( .A(n270), .B(n331), .C(n8502), .Y(n3243) );
  OAI21X1 U185 ( .A(n270), .B(n333), .C(n8499), .Y(n3244) );
  OAI21X1 U187 ( .A(n270), .B(n335), .C(n8496), .Y(n3245) );
  OAI21X1 U189 ( .A(n270), .B(n337), .C(n8493), .Y(n3246) );
  OAI21X1 U191 ( .A(n270), .B(n339), .C(n8490), .Y(n3247) );
  OAI21X1 U193 ( .A(n270), .B(n341), .C(n8487), .Y(n3248) );
  OAI21X1 U195 ( .A(n270), .B(n343), .C(n8484), .Y(n3249) );
  OAI21X1 U197 ( .A(n270), .B(n345), .C(n8481), .Y(n3250) );
  OAI21X1 U199 ( .A(n270), .B(n347), .C(n8478), .Y(n3251) );
  OAI21X1 U201 ( .A(n270), .B(n349), .C(n8475), .Y(n3252) );
  OAI21X1 U203 ( .A(n270), .B(n351), .C(n8472), .Y(n3253) );
  OAI21X1 U205 ( .A(n270), .B(n353), .C(n8469), .Y(n3254) );
  OAI21X1 U208 ( .A(n271), .B(n357), .C(n8466), .Y(n3255) );
  OAI21X1 U210 ( .A(n273), .B(n357), .C(n8463), .Y(n3256) );
  OAI21X1 U212 ( .A(n275), .B(n357), .C(n8460), .Y(n3257) );
  OAI21X1 U214 ( .A(n277), .B(n357), .C(n8457), .Y(n3258) );
  OAI21X1 U216 ( .A(n279), .B(n357), .C(n8454), .Y(n3259) );
  OAI21X1 U218 ( .A(n281), .B(n357), .C(n8451), .Y(n3260) );
  OAI21X1 U220 ( .A(n283), .B(n357), .C(n8448), .Y(n3261) );
  OAI21X1 U222 ( .A(n285), .B(n357), .C(n8445), .Y(n3262) );
  OAI21X1 U224 ( .A(n287), .B(n357), .C(n8442), .Y(n3263) );
  OAI21X1 U226 ( .A(n289), .B(n357), .C(n8439), .Y(n3264) );
  OAI21X1 U228 ( .A(n291), .B(n357), .C(n8436), .Y(n3265) );
  OAI21X1 U230 ( .A(n293), .B(n357), .C(n8433), .Y(n3266) );
  OAI21X1 U232 ( .A(n295), .B(n357), .C(n8430), .Y(n3267) );
  OAI21X1 U234 ( .A(n297), .B(n357), .C(n8427), .Y(n3268) );
  OAI21X1 U236 ( .A(n299), .B(n357), .C(n8424), .Y(n3269) );
  OAI21X1 U238 ( .A(n301), .B(n357), .C(n8421), .Y(n3270) );
  OAI21X1 U240 ( .A(n303), .B(n357), .C(n8418), .Y(n3271) );
  OAI21X1 U242 ( .A(n305), .B(n357), .C(n8415), .Y(n3272) );
  OAI21X1 U244 ( .A(n307), .B(n357), .C(n8412), .Y(n3273) );
  OAI21X1 U246 ( .A(n309), .B(n357), .C(n8409), .Y(n3274) );
  OAI21X1 U248 ( .A(n311), .B(n357), .C(n8406), .Y(n3275) );
  OAI21X1 U250 ( .A(n313), .B(n357), .C(n8403), .Y(n3276) );
  OAI21X1 U252 ( .A(n315), .B(n357), .C(n8400), .Y(n3277) );
  OAI21X1 U254 ( .A(n317), .B(n357), .C(n8397), .Y(n3278) );
  OAI21X1 U256 ( .A(n319), .B(n357), .C(n8394), .Y(n3279) );
  OAI21X1 U258 ( .A(n321), .B(n357), .C(n8391), .Y(n3280) );
  OAI21X1 U260 ( .A(n323), .B(n357), .C(n8388), .Y(n3281) );
  OAI21X1 U262 ( .A(n325), .B(n357), .C(n8385), .Y(n3282) );
  OAI21X1 U264 ( .A(n327), .B(n357), .C(n8382), .Y(n3283) );
  OAI21X1 U266 ( .A(n329), .B(n357), .C(n8379), .Y(n3284) );
  OAI21X1 U268 ( .A(n331), .B(n357), .C(n8376), .Y(n3285) );
  OAI21X1 U270 ( .A(n333), .B(n357), .C(n8373), .Y(n3286) );
  OAI21X1 U272 ( .A(n335), .B(n357), .C(n8370), .Y(n3287) );
  OAI21X1 U274 ( .A(n337), .B(n357), .C(n8367), .Y(n3288) );
  OAI21X1 U276 ( .A(n339), .B(n357), .C(n8364), .Y(n3289) );
  OAI21X1 U278 ( .A(n341), .B(n357), .C(n8361), .Y(n3290) );
  OAI21X1 U280 ( .A(n343), .B(n357), .C(n8358), .Y(n3291) );
  OAI21X1 U282 ( .A(n345), .B(n357), .C(n8355), .Y(n3292) );
  OAI21X1 U284 ( .A(n347), .B(n357), .C(n8352), .Y(n3293) );
  OAI21X1 U286 ( .A(n349), .B(n357), .C(n8349), .Y(n3294) );
  OAI21X1 U288 ( .A(n351), .B(n357), .C(n8346), .Y(n3295) );
  OAI21X1 U290 ( .A(n353), .B(n357), .C(n8343), .Y(n3296) );
  OAI21X1 U293 ( .A(n271), .B(n8676), .C(n8340), .Y(n3297) );
  OAI21X1 U295 ( .A(n273), .B(n8696), .C(n8337), .Y(n3298) );
  OAI21X1 U297 ( .A(n275), .B(n13042), .C(n8334), .Y(n3299) );
  OAI21X1 U299 ( .A(n277), .B(n8688), .C(n8331), .Y(n3300) );
  OAI21X1 U301 ( .A(n279), .B(n8678), .C(n8328), .Y(n3301) );
  OAI21X1 U303 ( .A(n281), .B(n13042), .C(n8325), .Y(n3302) );
  OAI21X1 U305 ( .A(n283), .B(n8708), .C(n8322), .Y(n3303) );
  OAI21X1 U307 ( .A(n285), .B(n13043), .C(n8319), .Y(n3304) );
  OAI21X1 U309 ( .A(n287), .B(n13042), .C(n8316), .Y(n3305) );
  OAI21X1 U311 ( .A(n289), .B(n12971), .C(n8313), .Y(n3306) );
  OAI21X1 U313 ( .A(n291), .B(n13024), .C(n8310), .Y(n3307) );
  OAI21X1 U315 ( .A(n293), .B(n13042), .C(n8307), .Y(n3308) );
  OAI21X1 U317 ( .A(n295), .B(n13043), .C(n8304), .Y(n3309) );
  OAI21X1 U319 ( .A(n297), .B(n13024), .C(n8301), .Y(n3310) );
  OAI21X1 U321 ( .A(n299), .B(n13042), .C(n8298), .Y(n3311) );
  OAI21X1 U323 ( .A(n301), .B(n12960), .C(n8295), .Y(n3312) );
  OAI21X1 U325 ( .A(n303), .B(n13043), .C(n8292), .Y(n3313) );
  OAI21X1 U327 ( .A(n305), .B(n13042), .C(n8289), .Y(n3314) );
  OAI21X1 U329 ( .A(n307), .B(n8720), .C(n8286), .Y(n3315) );
  OAI21X1 U331 ( .A(n309), .B(n13024), .C(n8283), .Y(n3316) );
  OAI21X1 U333 ( .A(n311), .B(n13042), .C(n8280), .Y(n3317) );
  OAI21X1 U335 ( .A(n313), .B(n13043), .C(n8277), .Y(n3318) );
  OAI21X1 U337 ( .A(n315), .B(n12988), .C(n8274), .Y(n3319) );
  OAI21X1 U339 ( .A(n317), .B(n13042), .C(n8271), .Y(n3320) );
  OAI21X1 U341 ( .A(n319), .B(n13024), .C(n8268), .Y(n3321) );
  OAI21X1 U343 ( .A(n321), .B(n8770), .C(n8265), .Y(n3322) );
  OAI21X1 U345 ( .A(n323), .B(n13042), .C(n8262), .Y(n3323) );
  OAI21X1 U347 ( .A(n325), .B(n12988), .C(n8259), .Y(n3324) );
  OAI21X1 U349 ( .A(n327), .B(n10798), .C(n8256), .Y(n3325) );
  OAI21X1 U351 ( .A(n329), .B(n13042), .C(n8253), .Y(n3326) );
  OAI21X1 U353 ( .A(n331), .B(n13043), .C(n8250), .Y(n3327) );
  OAI21X1 U355 ( .A(n333), .B(n12971), .C(n8247), .Y(n3328) );
  OAI21X1 U357 ( .A(n335), .B(n13042), .C(n8244), .Y(n3329) );
  OAI21X1 U359 ( .A(n337), .B(n13024), .C(n8241), .Y(n3330) );
  OAI21X1 U361 ( .A(n339), .B(n13024), .C(n8238), .Y(n3331) );
  OAI21X1 U363 ( .A(n341), .B(n13042), .C(n8235), .Y(n3332) );
  OAI21X1 U365 ( .A(n343), .B(n12971), .C(n8232), .Y(n3333) );
  OAI21X1 U367 ( .A(n345), .B(n12988), .C(n8229), .Y(n3334) );
  OAI21X1 U369 ( .A(n347), .B(n13042), .C(n8226), .Y(n3335) );
  OAI21X1 U371 ( .A(n349), .B(n8690), .C(n8223), .Y(n3336) );
  OAI21X1 U373 ( .A(n351), .B(n8684), .C(n8220), .Y(n3337) );
  OAI21X1 U375 ( .A(n353), .B(n13042), .C(n8217), .Y(n3338) );
  OAI21X1 U378 ( .A(n271), .B(n445), .C(n8214), .Y(n3339) );
  OAI21X1 U380 ( .A(n273), .B(n445), .C(n8211), .Y(n3340) );
  OAI21X1 U382 ( .A(n275), .B(n445), .C(n8208), .Y(n3341) );
  OAI21X1 U384 ( .A(n277), .B(n445), .C(n8205), .Y(n3342) );
  OAI21X1 U386 ( .A(n279), .B(n445), .C(n8202), .Y(n3343) );
  OAI21X1 U388 ( .A(n281), .B(n445), .C(n8199), .Y(n3344) );
  OAI21X1 U390 ( .A(n283), .B(n445), .C(n8196), .Y(n3345) );
  OAI21X1 U392 ( .A(n285), .B(n445), .C(n8193), .Y(n3346) );
  OAI21X1 U394 ( .A(n287), .B(n445), .C(n8190), .Y(n3347) );
  OAI21X1 U396 ( .A(n289), .B(n445), .C(n8187), .Y(n3348) );
  OAI21X1 U398 ( .A(n291), .B(n445), .C(n8184), .Y(n3349) );
  OAI21X1 U400 ( .A(n293), .B(n445), .C(n8181), .Y(n3350) );
  OAI21X1 U402 ( .A(n295), .B(n445), .C(n8178), .Y(n3351) );
  OAI21X1 U404 ( .A(n297), .B(n445), .C(n8175), .Y(n3352) );
  OAI21X1 U406 ( .A(n299), .B(n445), .C(n8172), .Y(n3353) );
  OAI21X1 U408 ( .A(n301), .B(n445), .C(n8169), .Y(n3354) );
  OAI21X1 U410 ( .A(n303), .B(n445), .C(n8166), .Y(n3355) );
  OAI21X1 U412 ( .A(n305), .B(n445), .C(n8163), .Y(n3356) );
  OAI21X1 U414 ( .A(n307), .B(n445), .C(n8160), .Y(n3357) );
  OAI21X1 U416 ( .A(n309), .B(n445), .C(n8157), .Y(n3358) );
  OAI21X1 U418 ( .A(n311), .B(n445), .C(n8154), .Y(n3359) );
  OAI21X1 U420 ( .A(n313), .B(n445), .C(n8151), .Y(n3360) );
  OAI21X1 U422 ( .A(n315), .B(n445), .C(n8148), .Y(n3361) );
  OAI21X1 U424 ( .A(n317), .B(n445), .C(n8145), .Y(n3362) );
  OAI21X1 U426 ( .A(n319), .B(n445), .C(n8142), .Y(n3363) );
  OAI21X1 U428 ( .A(n321), .B(n445), .C(n8139), .Y(n3364) );
  OAI21X1 U430 ( .A(n323), .B(n445), .C(n8136), .Y(n3365) );
  OAI21X1 U432 ( .A(n325), .B(n445), .C(n8133), .Y(n3366) );
  OAI21X1 U434 ( .A(n327), .B(n445), .C(n8130), .Y(n3367) );
  OAI21X1 U436 ( .A(n329), .B(n445), .C(n8127), .Y(n3368) );
  OAI21X1 U438 ( .A(n331), .B(n445), .C(n8124), .Y(n3369) );
  OAI21X1 U440 ( .A(n333), .B(n445), .C(n8121), .Y(n3370) );
  OAI21X1 U442 ( .A(n335), .B(n445), .C(n8118), .Y(n3371) );
  OAI21X1 U444 ( .A(n337), .B(n445), .C(n8115), .Y(n3372) );
  OAI21X1 U446 ( .A(n339), .B(n445), .C(n8112), .Y(n3373) );
  OAI21X1 U448 ( .A(n341), .B(n445), .C(n8109), .Y(n3374) );
  OAI21X1 U450 ( .A(n343), .B(n445), .C(n8106), .Y(n3375) );
  OAI21X1 U452 ( .A(n345), .B(n445), .C(n8103), .Y(n3376) );
  OAI21X1 U454 ( .A(n347), .B(n445), .C(n8100), .Y(n3377) );
  OAI21X1 U456 ( .A(n349), .B(n445), .C(n8097), .Y(n3378) );
  OAI21X1 U458 ( .A(n351), .B(n445), .C(n8094), .Y(n3379) );
  OAI21X1 U460 ( .A(n353), .B(n445), .C(n8091), .Y(n3380) );
  OAI21X1 U463 ( .A(n271), .B(n489), .C(n8088), .Y(n3381) );
  OAI21X1 U465 ( .A(n273), .B(n489), .C(n8085), .Y(n3382) );
  OAI21X1 U467 ( .A(n275), .B(n489), .C(n8082), .Y(n3383) );
  OAI21X1 U469 ( .A(n277), .B(n489), .C(n8079), .Y(n3384) );
  OAI21X1 U471 ( .A(n279), .B(n489), .C(n8076), .Y(n3385) );
  OAI21X1 U473 ( .A(n281), .B(n489), .C(n8073), .Y(n3386) );
  OAI21X1 U475 ( .A(n283), .B(n489), .C(n8070), .Y(n3387) );
  OAI21X1 U477 ( .A(n285), .B(n489), .C(n8067), .Y(n3388) );
  OAI21X1 U479 ( .A(n287), .B(n489), .C(n8064), .Y(n3389) );
  OAI21X1 U481 ( .A(n289), .B(n489), .C(n8061), .Y(n3390) );
  OAI21X1 U483 ( .A(n291), .B(n489), .C(n8058), .Y(n3391) );
  OAI21X1 U485 ( .A(n293), .B(n489), .C(n8055), .Y(n3392) );
  OAI21X1 U487 ( .A(n295), .B(n489), .C(n8052), .Y(n3393) );
  OAI21X1 U489 ( .A(n297), .B(n489), .C(n8049), .Y(n3394) );
  OAI21X1 U491 ( .A(n299), .B(n489), .C(n8046), .Y(n3395) );
  OAI21X1 U493 ( .A(n301), .B(n489), .C(n8043), .Y(n3396) );
  OAI21X1 U495 ( .A(n303), .B(n489), .C(n8040), .Y(n3397) );
  OAI21X1 U497 ( .A(n305), .B(n489), .C(n8037), .Y(n3398) );
  OAI21X1 U499 ( .A(n307), .B(n489), .C(n8034), .Y(n3399) );
  OAI21X1 U501 ( .A(n309), .B(n489), .C(n8031), .Y(n3400) );
  OAI21X1 U503 ( .A(n311), .B(n489), .C(n8028), .Y(n3401) );
  OAI21X1 U505 ( .A(n313), .B(n489), .C(n8025), .Y(n3402) );
  OAI21X1 U507 ( .A(n315), .B(n489), .C(n8022), .Y(n3403) );
  OAI21X1 U509 ( .A(n317), .B(n489), .C(n8019), .Y(n3404) );
  OAI21X1 U511 ( .A(n319), .B(n489), .C(n8016), .Y(n3405) );
  OAI21X1 U513 ( .A(n321), .B(n489), .C(n8013), .Y(n3406) );
  OAI21X1 U515 ( .A(n323), .B(n489), .C(n8010), .Y(n3407) );
  OAI21X1 U517 ( .A(n325), .B(n489), .C(n8007), .Y(n3408) );
  OAI21X1 U519 ( .A(n327), .B(n489), .C(n8004), .Y(n3409) );
  OAI21X1 U521 ( .A(n329), .B(n489), .C(n8001), .Y(n3410) );
  OAI21X1 U523 ( .A(n331), .B(n489), .C(n7998), .Y(n3411) );
  OAI21X1 U525 ( .A(n333), .B(n489), .C(n7995), .Y(n3412) );
  OAI21X1 U527 ( .A(n335), .B(n489), .C(n7992), .Y(n3413) );
  OAI21X1 U529 ( .A(n337), .B(n489), .C(n7989), .Y(n3414) );
  OAI21X1 U531 ( .A(n339), .B(n489), .C(n7986), .Y(n3415) );
  OAI21X1 U533 ( .A(n341), .B(n489), .C(n7983), .Y(n3416) );
  OAI21X1 U535 ( .A(n343), .B(n489), .C(n7980), .Y(n3417) );
  OAI21X1 U537 ( .A(n345), .B(n489), .C(n7977), .Y(n3418) );
  OAI21X1 U539 ( .A(n347), .B(n489), .C(n7974), .Y(n3419) );
  OAI21X1 U541 ( .A(n349), .B(n489), .C(n7971), .Y(n3420) );
  OAI21X1 U543 ( .A(n351), .B(n489), .C(n7968), .Y(n3421) );
  OAI21X1 U545 ( .A(n353), .B(n489), .C(n7965), .Y(n3422) );
  OAI21X1 U548 ( .A(n271), .B(n533), .C(n7962), .Y(n3423) );
  OAI21X1 U550 ( .A(n273), .B(n533), .C(n7959), .Y(n3424) );
  OAI21X1 U552 ( .A(n275), .B(n533), .C(n7956), .Y(n3425) );
  OAI21X1 U554 ( .A(n277), .B(n533), .C(n7953), .Y(n3426) );
  OAI21X1 U556 ( .A(n279), .B(n533), .C(n7950), .Y(n3427) );
  OAI21X1 U558 ( .A(n281), .B(n533), .C(n7947), .Y(n3428) );
  OAI21X1 U560 ( .A(n283), .B(n533), .C(n7944), .Y(n3429) );
  OAI21X1 U562 ( .A(n285), .B(n533), .C(n7941), .Y(n3430) );
  OAI21X1 U564 ( .A(n287), .B(n533), .C(n7938), .Y(n3431) );
  OAI21X1 U566 ( .A(n289), .B(n533), .C(n7935), .Y(n3432) );
  OAI21X1 U568 ( .A(n291), .B(n533), .C(n7932), .Y(n3433) );
  OAI21X1 U570 ( .A(n293), .B(n533), .C(n7929), .Y(n3434) );
  OAI21X1 U572 ( .A(n295), .B(n533), .C(n7926), .Y(n3435) );
  OAI21X1 U574 ( .A(n297), .B(n533), .C(n7923), .Y(n3436) );
  OAI21X1 U576 ( .A(n299), .B(n533), .C(n7920), .Y(n3437) );
  OAI21X1 U578 ( .A(n301), .B(n533), .C(n7917), .Y(n3438) );
  OAI21X1 U580 ( .A(n303), .B(n533), .C(n7914), .Y(n3439) );
  OAI21X1 U582 ( .A(n305), .B(n533), .C(n7911), .Y(n3440) );
  OAI21X1 U584 ( .A(n307), .B(n533), .C(n7908), .Y(n3441) );
  OAI21X1 U586 ( .A(n309), .B(n533), .C(n7905), .Y(n3442) );
  OAI21X1 U588 ( .A(n311), .B(n533), .C(n7902), .Y(n3443) );
  OAI21X1 U590 ( .A(n313), .B(n533), .C(n7899), .Y(n3444) );
  OAI21X1 U592 ( .A(n315), .B(n533), .C(n7896), .Y(n3445) );
  OAI21X1 U594 ( .A(n317), .B(n533), .C(n7893), .Y(n3446) );
  OAI21X1 U596 ( .A(n319), .B(n533), .C(n7890), .Y(n3447) );
  OAI21X1 U598 ( .A(n321), .B(n533), .C(n7887), .Y(n3448) );
  OAI21X1 U600 ( .A(n323), .B(n533), .C(n7884), .Y(n3449) );
  OAI21X1 U602 ( .A(n325), .B(n533), .C(n7881), .Y(n3450) );
  OAI21X1 U604 ( .A(n327), .B(n533), .C(n7878), .Y(n3451) );
  OAI21X1 U606 ( .A(n329), .B(n533), .C(n7875), .Y(n3452) );
  OAI21X1 U608 ( .A(n331), .B(n533), .C(n7872), .Y(n3453) );
  OAI21X1 U610 ( .A(n333), .B(n533), .C(n7869), .Y(n3454) );
  OAI21X1 U612 ( .A(n335), .B(n533), .C(n7866), .Y(n3455) );
  OAI21X1 U614 ( .A(n337), .B(n533), .C(n7863), .Y(n3456) );
  OAI21X1 U616 ( .A(n339), .B(n533), .C(n7860), .Y(n3457) );
  OAI21X1 U618 ( .A(n341), .B(n533), .C(n7857), .Y(n3458) );
  OAI21X1 U620 ( .A(n343), .B(n533), .C(n7854), .Y(n3459) );
  OAI21X1 U622 ( .A(n345), .B(n533), .C(n7851), .Y(n3460) );
  OAI21X1 U624 ( .A(n347), .B(n533), .C(n7848), .Y(n3461) );
  OAI21X1 U626 ( .A(n349), .B(n533), .C(n7845), .Y(n3462) );
  OAI21X1 U628 ( .A(n351), .B(n533), .C(n7842), .Y(n3463) );
  OAI21X1 U630 ( .A(n353), .B(n533), .C(n7839), .Y(n3464) );
  OAI21X1 U633 ( .A(n271), .B(n577), .C(n7836), .Y(n3465) );
  OAI21X1 U635 ( .A(n273), .B(n577), .C(n7833), .Y(n3466) );
  OAI21X1 U637 ( .A(n275), .B(n577), .C(n7830), .Y(n3467) );
  OAI21X1 U639 ( .A(n277), .B(n577), .C(n7827), .Y(n3468) );
  OAI21X1 U641 ( .A(n279), .B(n577), .C(n7824), .Y(n3469) );
  OAI21X1 U643 ( .A(n281), .B(n577), .C(n7821), .Y(n3470) );
  OAI21X1 U645 ( .A(n283), .B(n577), .C(n7818), .Y(n3471) );
  OAI21X1 U647 ( .A(n285), .B(n577), .C(n7815), .Y(n3472) );
  OAI21X1 U649 ( .A(n287), .B(n577), .C(n7812), .Y(n3473) );
  OAI21X1 U651 ( .A(n289), .B(n577), .C(n7809), .Y(n3474) );
  OAI21X1 U653 ( .A(n291), .B(n577), .C(n7806), .Y(n3475) );
  OAI21X1 U655 ( .A(n293), .B(n577), .C(n7803), .Y(n3476) );
  OAI21X1 U657 ( .A(n295), .B(n577), .C(n7800), .Y(n3477) );
  OAI21X1 U659 ( .A(n297), .B(n577), .C(n7797), .Y(n3478) );
  OAI21X1 U661 ( .A(n299), .B(n577), .C(n7794), .Y(n3479) );
  OAI21X1 U663 ( .A(n301), .B(n577), .C(n7791), .Y(n3480) );
  OAI21X1 U665 ( .A(n303), .B(n577), .C(n7788), .Y(n3481) );
  OAI21X1 U667 ( .A(n305), .B(n577), .C(n7785), .Y(n3482) );
  OAI21X1 U669 ( .A(n307), .B(n577), .C(n7782), .Y(n3483) );
  OAI21X1 U671 ( .A(n309), .B(n577), .C(n7779), .Y(n3484) );
  OAI21X1 U673 ( .A(n311), .B(n577), .C(n7776), .Y(n3485) );
  OAI21X1 U675 ( .A(n313), .B(n577), .C(n7773), .Y(n3486) );
  OAI21X1 U677 ( .A(n315), .B(n577), .C(n7770), .Y(n3487) );
  OAI21X1 U679 ( .A(n317), .B(n577), .C(n7767), .Y(n3488) );
  OAI21X1 U681 ( .A(n319), .B(n577), .C(n7764), .Y(n3489) );
  OAI21X1 U683 ( .A(n321), .B(n577), .C(n7761), .Y(n3490) );
  OAI21X1 U685 ( .A(n323), .B(n577), .C(n7758), .Y(n3491) );
  OAI21X1 U687 ( .A(n325), .B(n577), .C(n7755), .Y(n3492) );
  OAI21X1 U689 ( .A(n327), .B(n577), .C(n7752), .Y(n3493) );
  OAI21X1 U691 ( .A(n329), .B(n577), .C(n7749), .Y(n3494) );
  OAI21X1 U693 ( .A(n331), .B(n577), .C(n7746), .Y(n3495) );
  OAI21X1 U695 ( .A(n333), .B(n577), .C(n7743), .Y(n3496) );
  OAI21X1 U697 ( .A(n335), .B(n577), .C(n7740), .Y(n3497) );
  OAI21X1 U699 ( .A(n337), .B(n577), .C(n7737), .Y(n3498) );
  OAI21X1 U701 ( .A(n339), .B(n577), .C(n7734), .Y(n3499) );
  OAI21X1 U703 ( .A(n341), .B(n577), .C(n7731), .Y(n3500) );
  OAI21X1 U705 ( .A(n343), .B(n577), .C(n7728), .Y(n3501) );
  OAI21X1 U707 ( .A(n345), .B(n577), .C(n7725), .Y(n3502) );
  OAI21X1 U709 ( .A(n347), .B(n577), .C(n7722), .Y(n3503) );
  OAI21X1 U711 ( .A(n349), .B(n577), .C(n7719), .Y(n3504) );
  OAI21X1 U713 ( .A(n351), .B(n577), .C(n7716), .Y(n3505) );
  OAI21X1 U715 ( .A(n353), .B(n577), .C(n7713), .Y(n3506) );
  OAI21X1 U718 ( .A(n271), .B(n621), .C(n7710), .Y(n3507) );
  OAI21X1 U720 ( .A(n273), .B(n621), .C(n7707), .Y(n3508) );
  OAI21X1 U722 ( .A(n275), .B(n621), .C(n7704), .Y(n3509) );
  OAI21X1 U724 ( .A(n277), .B(n621), .C(n7701), .Y(n3510) );
  OAI21X1 U726 ( .A(n279), .B(n621), .C(n7698), .Y(n3511) );
  OAI21X1 U728 ( .A(n281), .B(n621), .C(n7695), .Y(n3512) );
  OAI21X1 U730 ( .A(n283), .B(n621), .C(n7692), .Y(n3513) );
  OAI21X1 U732 ( .A(n285), .B(n621), .C(n7689), .Y(n3514) );
  OAI21X1 U734 ( .A(n287), .B(n621), .C(n7686), .Y(n3515) );
  OAI21X1 U736 ( .A(n289), .B(n621), .C(n7683), .Y(n3516) );
  OAI21X1 U738 ( .A(n291), .B(n621), .C(n7680), .Y(n3517) );
  OAI21X1 U740 ( .A(n293), .B(n621), .C(n7677), .Y(n3518) );
  OAI21X1 U742 ( .A(n295), .B(n621), .C(n7674), .Y(n3519) );
  OAI21X1 U744 ( .A(n297), .B(n621), .C(n7671), .Y(n3520) );
  OAI21X1 U746 ( .A(n299), .B(n621), .C(n7668), .Y(n3521) );
  OAI21X1 U748 ( .A(n301), .B(n621), .C(n7665), .Y(n3522) );
  OAI21X1 U750 ( .A(n303), .B(n621), .C(n7662), .Y(n3523) );
  OAI21X1 U752 ( .A(n305), .B(n621), .C(n7659), .Y(n3524) );
  OAI21X1 U754 ( .A(n307), .B(n621), .C(n7656), .Y(n3525) );
  OAI21X1 U756 ( .A(n309), .B(n621), .C(n7653), .Y(n3526) );
  OAI21X1 U758 ( .A(n311), .B(n621), .C(n7650), .Y(n3527) );
  OAI21X1 U760 ( .A(n313), .B(n621), .C(n7647), .Y(n3528) );
  OAI21X1 U762 ( .A(n315), .B(n621), .C(n7644), .Y(n3529) );
  OAI21X1 U764 ( .A(n317), .B(n621), .C(n7641), .Y(n3530) );
  OAI21X1 U766 ( .A(n319), .B(n621), .C(n7638), .Y(n3531) );
  OAI21X1 U768 ( .A(n321), .B(n621), .C(n7635), .Y(n3532) );
  OAI21X1 U770 ( .A(n323), .B(n621), .C(n7632), .Y(n3533) );
  OAI21X1 U772 ( .A(n325), .B(n621), .C(n7629), .Y(n3534) );
  OAI21X1 U774 ( .A(n327), .B(n621), .C(n7626), .Y(n3535) );
  OAI21X1 U776 ( .A(n329), .B(n621), .C(n7623), .Y(n3536) );
  OAI21X1 U778 ( .A(n331), .B(n621), .C(n7620), .Y(n3537) );
  OAI21X1 U780 ( .A(n333), .B(n621), .C(n7617), .Y(n3538) );
  OAI21X1 U782 ( .A(n335), .B(n621), .C(n7614), .Y(n3539) );
  OAI21X1 U784 ( .A(n337), .B(n621), .C(n7611), .Y(n3540) );
  OAI21X1 U786 ( .A(n339), .B(n621), .C(n7608), .Y(n3541) );
  OAI21X1 U788 ( .A(n341), .B(n621), .C(n7605), .Y(n3542) );
  OAI21X1 U790 ( .A(n343), .B(n621), .C(n7602), .Y(n3543) );
  OAI21X1 U792 ( .A(n345), .B(n621), .C(n7599), .Y(n3544) );
  OAI21X1 U794 ( .A(n347), .B(n621), .C(n7596), .Y(n3545) );
  OAI21X1 U796 ( .A(n349), .B(n621), .C(n7593), .Y(n3546) );
  OAI21X1 U798 ( .A(n351), .B(n621), .C(n7590), .Y(n3547) );
  OAI21X1 U800 ( .A(n353), .B(n621), .C(n7587), .Y(n3548) );
  NAND3X1 U804 ( .A(n256), .B(n254), .C(n253), .Y(n665) );
  OAI21X1 U805 ( .A(n271), .B(n666), .C(n7584), .Y(n3549) );
  OAI21X1 U807 ( .A(n273), .B(n666), .C(n7581), .Y(n3550) );
  OAI21X1 U809 ( .A(n275), .B(n666), .C(n7578), .Y(n3551) );
  OAI21X1 U811 ( .A(n277), .B(n666), .C(n7575), .Y(n3552) );
  OAI21X1 U813 ( .A(n279), .B(n666), .C(n7572), .Y(n3553) );
  OAI21X1 U815 ( .A(n281), .B(n666), .C(n7569), .Y(n3554) );
  OAI21X1 U817 ( .A(n283), .B(n666), .C(n7566), .Y(n3555) );
  OAI21X1 U819 ( .A(n285), .B(n666), .C(n7563), .Y(n3556) );
  OAI21X1 U821 ( .A(n287), .B(n666), .C(n7560), .Y(n3557) );
  OAI21X1 U823 ( .A(n289), .B(n666), .C(n7557), .Y(n3558) );
  OAI21X1 U825 ( .A(n291), .B(n666), .C(n7554), .Y(n3559) );
  OAI21X1 U827 ( .A(n293), .B(n666), .C(n7551), .Y(n3560) );
  OAI21X1 U829 ( .A(n295), .B(n666), .C(n7548), .Y(n3561) );
  OAI21X1 U831 ( .A(n297), .B(n666), .C(n7545), .Y(n3562) );
  OAI21X1 U833 ( .A(n299), .B(n666), .C(n7542), .Y(n3563) );
  OAI21X1 U835 ( .A(n301), .B(n666), .C(n7539), .Y(n3564) );
  OAI21X1 U837 ( .A(n303), .B(n666), .C(n7536), .Y(n3565) );
  OAI21X1 U839 ( .A(n305), .B(n666), .C(n7533), .Y(n3566) );
  OAI21X1 U841 ( .A(n307), .B(n666), .C(n7530), .Y(n3567) );
  OAI21X1 U843 ( .A(n309), .B(n666), .C(n7527), .Y(n3568) );
  OAI21X1 U845 ( .A(n311), .B(n666), .C(n7524), .Y(n3569) );
  OAI21X1 U847 ( .A(n313), .B(n666), .C(n7521), .Y(n3570) );
  OAI21X1 U849 ( .A(n315), .B(n666), .C(n7518), .Y(n3571) );
  OAI21X1 U851 ( .A(n317), .B(n666), .C(n7515), .Y(n3572) );
  OAI21X1 U853 ( .A(n319), .B(n666), .C(n7512), .Y(n3573) );
  OAI21X1 U855 ( .A(n321), .B(n666), .C(n7509), .Y(n3574) );
  OAI21X1 U857 ( .A(n323), .B(n666), .C(n7506), .Y(n3575) );
  OAI21X1 U859 ( .A(n325), .B(n666), .C(n7503), .Y(n3576) );
  OAI21X1 U861 ( .A(n327), .B(n666), .C(n7500), .Y(n3577) );
  OAI21X1 U863 ( .A(n329), .B(n666), .C(n7497), .Y(n3578) );
  OAI21X1 U865 ( .A(n331), .B(n666), .C(n7494), .Y(n3579) );
  OAI21X1 U867 ( .A(n333), .B(n666), .C(n7491), .Y(n3580) );
  OAI21X1 U869 ( .A(n335), .B(n666), .C(n7488), .Y(n3581) );
  OAI21X1 U871 ( .A(n337), .B(n666), .C(n7485), .Y(n3582) );
  OAI21X1 U873 ( .A(n339), .B(n666), .C(n7482), .Y(n3583) );
  OAI21X1 U875 ( .A(n341), .B(n666), .C(n7479), .Y(n3584) );
  OAI21X1 U877 ( .A(n343), .B(n666), .C(n7476), .Y(n3585) );
  OAI21X1 U879 ( .A(n345), .B(n666), .C(n7473), .Y(n3586) );
  OAI21X1 U881 ( .A(n347), .B(n666), .C(n7470), .Y(n3587) );
  OAI21X1 U883 ( .A(n349), .B(n666), .C(n7467), .Y(n3588) );
  OAI21X1 U885 ( .A(n351), .B(n666), .C(n7464), .Y(n3589) );
  OAI21X1 U887 ( .A(n353), .B(n666), .C(n7461), .Y(n3590) );
  OAI21X1 U890 ( .A(n271), .B(n710), .C(n7458), .Y(n3591) );
  OAI21X1 U892 ( .A(n273), .B(n710), .C(n7455), .Y(n3592) );
  OAI21X1 U894 ( .A(n275), .B(n710), .C(n7452), .Y(n3593) );
  OAI21X1 U896 ( .A(n277), .B(n710), .C(n7449), .Y(n3594) );
  OAI21X1 U898 ( .A(n279), .B(n710), .C(n7446), .Y(n3595) );
  OAI21X1 U900 ( .A(n281), .B(n710), .C(n7443), .Y(n3596) );
  OAI21X1 U902 ( .A(n283), .B(n710), .C(n7440), .Y(n3597) );
  OAI21X1 U904 ( .A(n285), .B(n710), .C(n7437), .Y(n3598) );
  OAI21X1 U906 ( .A(n287), .B(n710), .C(n7434), .Y(n3599) );
  OAI21X1 U908 ( .A(n289), .B(n710), .C(n7431), .Y(n3600) );
  OAI21X1 U910 ( .A(n291), .B(n710), .C(n7428), .Y(n3601) );
  OAI21X1 U912 ( .A(n293), .B(n710), .C(n7425), .Y(n3602) );
  OAI21X1 U914 ( .A(n295), .B(n710), .C(n7422), .Y(n3603) );
  OAI21X1 U916 ( .A(n297), .B(n710), .C(n7419), .Y(n3604) );
  OAI21X1 U918 ( .A(n299), .B(n710), .C(n7416), .Y(n3605) );
  OAI21X1 U920 ( .A(n301), .B(n710), .C(n7413), .Y(n3606) );
  OAI21X1 U922 ( .A(n303), .B(n710), .C(n7410), .Y(n3607) );
  OAI21X1 U924 ( .A(n305), .B(n710), .C(n7407), .Y(n3608) );
  OAI21X1 U926 ( .A(n307), .B(n710), .C(n7404), .Y(n3609) );
  OAI21X1 U928 ( .A(n309), .B(n710), .C(n7401), .Y(n3610) );
  OAI21X1 U930 ( .A(n311), .B(n710), .C(n7398), .Y(n3611) );
  OAI21X1 U932 ( .A(n313), .B(n710), .C(n7395), .Y(n3612) );
  OAI21X1 U934 ( .A(n315), .B(n710), .C(n7392), .Y(n3613) );
  OAI21X1 U936 ( .A(n317), .B(n710), .C(n7389), .Y(n3614) );
  OAI21X1 U938 ( .A(n319), .B(n710), .C(n7386), .Y(n3615) );
  OAI21X1 U940 ( .A(n321), .B(n710), .C(n7383), .Y(n3616) );
  OAI21X1 U942 ( .A(n323), .B(n710), .C(n7380), .Y(n3617) );
  OAI21X1 U944 ( .A(n325), .B(n710), .C(n7377), .Y(n3618) );
  OAI21X1 U946 ( .A(n327), .B(n710), .C(n7374), .Y(n3619) );
  OAI21X1 U948 ( .A(n329), .B(n710), .C(n7371), .Y(n3620) );
  OAI21X1 U950 ( .A(n331), .B(n710), .C(n7368), .Y(n3621) );
  OAI21X1 U952 ( .A(n333), .B(n710), .C(n7365), .Y(n3622) );
  OAI21X1 U954 ( .A(n335), .B(n710), .C(n7362), .Y(n3623) );
  OAI21X1 U956 ( .A(n337), .B(n710), .C(n7359), .Y(n3624) );
  OAI21X1 U958 ( .A(n339), .B(n710), .C(n7356), .Y(n3625) );
  OAI21X1 U960 ( .A(n341), .B(n710), .C(n7353), .Y(n3626) );
  OAI21X1 U962 ( .A(n343), .B(n710), .C(n7350), .Y(n3627) );
  OAI21X1 U964 ( .A(n345), .B(n710), .C(n7347), .Y(n3628) );
  OAI21X1 U966 ( .A(n347), .B(n710), .C(n7344), .Y(n3629) );
  OAI21X1 U968 ( .A(n349), .B(n710), .C(n7341), .Y(n3630) );
  OAI21X1 U970 ( .A(n351), .B(n710), .C(n7338), .Y(n3631) );
  OAI21X1 U972 ( .A(n353), .B(n710), .C(n7335), .Y(n3632) );
  OAI21X1 U975 ( .A(n271), .B(n753), .C(n7332), .Y(n3633) );
  OAI21X1 U977 ( .A(n273), .B(n753), .C(n7329), .Y(n3634) );
  OAI21X1 U979 ( .A(n275), .B(n753), .C(n7326), .Y(n3635) );
  OAI21X1 U981 ( .A(n277), .B(n753), .C(n7323), .Y(n3636) );
  OAI21X1 U983 ( .A(n279), .B(n753), .C(n7320), .Y(n3637) );
  OAI21X1 U985 ( .A(n281), .B(n753), .C(n7317), .Y(n3638) );
  OAI21X1 U987 ( .A(n283), .B(n753), .C(n7314), .Y(n3639) );
  OAI21X1 U989 ( .A(n285), .B(n753), .C(n7311), .Y(n3640) );
  OAI21X1 U991 ( .A(n287), .B(n753), .C(n7308), .Y(n3641) );
  OAI21X1 U993 ( .A(n289), .B(n753), .C(n7305), .Y(n3642) );
  OAI21X1 U995 ( .A(n291), .B(n753), .C(n7302), .Y(n3643) );
  OAI21X1 U997 ( .A(n293), .B(n753), .C(n7299), .Y(n3644) );
  OAI21X1 U999 ( .A(n295), .B(n753), .C(n7296), .Y(n3645) );
  OAI21X1 U1001 ( .A(n297), .B(n753), .C(n7293), .Y(n3646) );
  OAI21X1 U1003 ( .A(n299), .B(n753), .C(n7290), .Y(n3647) );
  OAI21X1 U1005 ( .A(n301), .B(n753), .C(n7287), .Y(n3648) );
  OAI21X1 U1007 ( .A(n303), .B(n753), .C(n7284), .Y(n3649) );
  OAI21X1 U1009 ( .A(n305), .B(n753), .C(n7281), .Y(n3650) );
  OAI21X1 U1011 ( .A(n307), .B(n753), .C(n7278), .Y(n3651) );
  OAI21X1 U1013 ( .A(n309), .B(n753), .C(n7275), .Y(n3652) );
  OAI21X1 U1015 ( .A(n311), .B(n753), .C(n7272), .Y(n3653) );
  OAI21X1 U1017 ( .A(n313), .B(n753), .C(n7269), .Y(n3654) );
  OAI21X1 U1019 ( .A(n315), .B(n753), .C(n7266), .Y(n3655) );
  OAI21X1 U1021 ( .A(n317), .B(n753), .C(n7263), .Y(n3656) );
  OAI21X1 U1023 ( .A(n319), .B(n753), .C(n7260), .Y(n3657) );
  OAI21X1 U1025 ( .A(n321), .B(n753), .C(n7257), .Y(n3658) );
  OAI21X1 U1027 ( .A(n323), .B(n753), .C(n7254), .Y(n3659) );
  OAI21X1 U1029 ( .A(n325), .B(n753), .C(n7251), .Y(n3660) );
  OAI21X1 U1031 ( .A(n327), .B(n753), .C(n7248), .Y(n3661) );
  OAI21X1 U1033 ( .A(n329), .B(n753), .C(n7245), .Y(n3662) );
  OAI21X1 U1035 ( .A(n331), .B(n753), .C(n7242), .Y(n3663) );
  OAI21X1 U1037 ( .A(n333), .B(n753), .C(n7239), .Y(n3664) );
  OAI21X1 U1039 ( .A(n335), .B(n753), .C(n7236), .Y(n3665) );
  OAI21X1 U1041 ( .A(n337), .B(n753), .C(n7233), .Y(n3666) );
  OAI21X1 U1043 ( .A(n339), .B(n753), .C(n7230), .Y(n3667) );
  OAI21X1 U1045 ( .A(n341), .B(n753), .C(n7227), .Y(n3668) );
  OAI21X1 U1047 ( .A(n343), .B(n753), .C(n7224), .Y(n3669) );
  OAI21X1 U1049 ( .A(n345), .B(n753), .C(n7221), .Y(n3670) );
  OAI21X1 U1051 ( .A(n347), .B(n753), .C(n7218), .Y(n3671) );
  OAI21X1 U1053 ( .A(n349), .B(n753), .C(n7215), .Y(n3672) );
  OAI21X1 U1055 ( .A(n351), .B(n753), .C(n7212), .Y(n3673) );
  OAI21X1 U1057 ( .A(n353), .B(n753), .C(n7209), .Y(n3674) );
  OAI21X1 U1060 ( .A(n271), .B(n12961), .C(n7206), .Y(n3675) );
  OAI21X1 U1062 ( .A(n273), .B(n8700), .C(n7203), .Y(n3676) );
  OAI21X1 U1064 ( .A(n275), .B(n13038), .C(n7200), .Y(n3677) );
  OAI21X1 U1066 ( .A(n277), .B(n8674), .C(n7197), .Y(n3678) );
  OAI21X1 U1068 ( .A(n279), .B(n8718), .C(n7194), .Y(n3679) );
  OAI21X1 U1070 ( .A(n281), .B(n13038), .C(n7191), .Y(n3680) );
  OAI21X1 U1072 ( .A(n283), .B(n8680), .C(n7188), .Y(n3681) );
  OAI21X1 U1074 ( .A(n285), .B(n13039), .C(n7185), .Y(n3682) );
  OAI21X1 U1076 ( .A(n287), .B(n13038), .C(n7182), .Y(n3683) );
  OAI21X1 U1078 ( .A(n289), .B(n12973), .C(n7179), .Y(n3684) );
  OAI21X1 U1080 ( .A(n291), .B(n13025), .C(n7176), .Y(n3685) );
  OAI21X1 U1082 ( .A(n293), .B(n13038), .C(n7173), .Y(n3686) );
  OAI21X1 U1084 ( .A(n295), .B(n13040), .C(n7170), .Y(n3687) );
  OAI21X1 U1086 ( .A(n297), .B(n13025), .C(n7167), .Y(n3688) );
  OAI21X1 U1088 ( .A(n299), .B(n13038), .C(n7164), .Y(n3689) );
  OAI21X1 U1090 ( .A(n301), .B(n8692), .C(n7161), .Y(n3690) );
  OAI21X1 U1092 ( .A(n303), .B(n13039), .C(n7158), .Y(n3691) );
  OAI21X1 U1094 ( .A(n305), .B(n13038), .C(n7155), .Y(n3692) );
  OAI21X1 U1096 ( .A(n307), .B(n8775), .C(n7152), .Y(n3693) );
  OAI21X1 U1098 ( .A(n309), .B(n13025), .C(n7149), .Y(n3694) );
  OAI21X1 U1100 ( .A(n311), .B(n13038), .C(n7146), .Y(n3695) );
  OAI21X1 U1102 ( .A(n313), .B(n13040), .C(n7143), .Y(n3696) );
  OAI21X1 U1104 ( .A(n315), .B(n12986), .C(n7140), .Y(n3697) );
  OAI21X1 U1106 ( .A(n317), .B(n13038), .C(n7137), .Y(n3698) );
  OAI21X1 U1108 ( .A(n319), .B(n13025), .C(n7134), .Y(n3699) );
  OAI21X1 U1110 ( .A(n321), .B(n8712), .C(n7131), .Y(n3700) );
  OAI21X1 U1112 ( .A(n323), .B(n13038), .C(n7128), .Y(n3701) );
  OAI21X1 U1114 ( .A(n325), .B(n12986), .C(n7125), .Y(n3702) );
  OAI21X1 U1116 ( .A(n327), .B(n8698), .C(n7122), .Y(n3703) );
  OAI21X1 U1118 ( .A(n329), .B(n13038), .C(n7119), .Y(n3704) );
  OAI21X1 U1120 ( .A(n331), .B(n13039), .C(n7116), .Y(n3705) );
  OAI21X1 U1122 ( .A(n333), .B(n13040), .C(n7113), .Y(n3706) );
  OAI21X1 U1124 ( .A(n335), .B(n13038), .C(n7110), .Y(n3707) );
  OAI21X1 U1126 ( .A(n337), .B(n13025), .C(n7107), .Y(n3708) );
  OAI21X1 U1128 ( .A(n339), .B(n13025), .C(n7104), .Y(n3709) );
  OAI21X1 U1130 ( .A(n341), .B(n13038), .C(n7101), .Y(n3710) );
  OAI21X1 U1132 ( .A(n343), .B(n12973), .C(n7098), .Y(n3711) );
  OAI21X1 U1134 ( .A(n345), .B(n12986), .C(n7095), .Y(n3712) );
  OAI21X1 U1136 ( .A(n347), .B(n13038), .C(n7092), .Y(n3713) );
  OAI21X1 U1138 ( .A(n349), .B(n8722), .C(n7089), .Y(n3714) );
  OAI21X1 U1140 ( .A(n351), .B(n10800), .C(n7086), .Y(n3715) );
  OAI21X1 U1142 ( .A(n353), .B(n13038), .C(n7083), .Y(n3716) );
  OAI21X1 U1145 ( .A(n271), .B(n839), .C(n7080), .Y(n3717) );
  OAI21X1 U1147 ( .A(n273), .B(n839), .C(n7077), .Y(n3718) );
  OAI21X1 U1149 ( .A(n275), .B(n839), .C(n7074), .Y(n3719) );
  OAI21X1 U1151 ( .A(n277), .B(n839), .C(n7071), .Y(n3720) );
  OAI21X1 U1153 ( .A(n279), .B(n839), .C(n7068), .Y(n3721) );
  OAI21X1 U1155 ( .A(n281), .B(n839), .C(n7065), .Y(n3722) );
  OAI21X1 U1157 ( .A(n283), .B(n839), .C(n7062), .Y(n3723) );
  OAI21X1 U1159 ( .A(n285), .B(n839), .C(n7059), .Y(n3724) );
  OAI21X1 U1161 ( .A(n287), .B(n839), .C(n7056), .Y(n3725) );
  OAI21X1 U1163 ( .A(n289), .B(n839), .C(n7053), .Y(n3726) );
  OAI21X1 U1165 ( .A(n291), .B(n839), .C(n7050), .Y(n3727) );
  OAI21X1 U1167 ( .A(n293), .B(n839), .C(n7047), .Y(n3728) );
  OAI21X1 U1169 ( .A(n295), .B(n839), .C(n7044), .Y(n3729) );
  OAI21X1 U1171 ( .A(n297), .B(n839), .C(n7041), .Y(n3730) );
  OAI21X1 U1173 ( .A(n299), .B(n839), .C(n7038), .Y(n3731) );
  OAI21X1 U1175 ( .A(n301), .B(n839), .C(n7035), .Y(n3732) );
  OAI21X1 U1177 ( .A(n303), .B(n839), .C(n7032), .Y(n3733) );
  OAI21X1 U1179 ( .A(n305), .B(n839), .C(n7029), .Y(n3734) );
  OAI21X1 U1181 ( .A(n307), .B(n839), .C(n7026), .Y(n3735) );
  OAI21X1 U1183 ( .A(n309), .B(n839), .C(n7023), .Y(n3736) );
  OAI21X1 U1185 ( .A(n311), .B(n839), .C(n7020), .Y(n3737) );
  OAI21X1 U1187 ( .A(n313), .B(n839), .C(n7017), .Y(n3738) );
  OAI21X1 U1189 ( .A(n315), .B(n839), .C(n7014), .Y(n3739) );
  OAI21X1 U1191 ( .A(n317), .B(n839), .C(n7011), .Y(n3740) );
  OAI21X1 U1193 ( .A(n319), .B(n839), .C(n7008), .Y(n3741) );
  OAI21X1 U1195 ( .A(n321), .B(n839), .C(n7005), .Y(n3742) );
  OAI21X1 U1197 ( .A(n323), .B(n839), .C(n7002), .Y(n3743) );
  OAI21X1 U1199 ( .A(n325), .B(n839), .C(n6999), .Y(n3744) );
  OAI21X1 U1201 ( .A(n327), .B(n839), .C(n6996), .Y(n3745) );
  OAI21X1 U1203 ( .A(n329), .B(n839), .C(n6993), .Y(n3746) );
  OAI21X1 U1205 ( .A(n331), .B(n839), .C(n6990), .Y(n3747) );
  OAI21X1 U1207 ( .A(n333), .B(n839), .C(n6987), .Y(n3748) );
  OAI21X1 U1209 ( .A(n335), .B(n839), .C(n6984), .Y(n3749) );
  OAI21X1 U1211 ( .A(n337), .B(n839), .C(n6981), .Y(n3750) );
  OAI21X1 U1213 ( .A(n339), .B(n839), .C(n6978), .Y(n3751) );
  OAI21X1 U1215 ( .A(n341), .B(n839), .C(n6975), .Y(n3752) );
  OAI21X1 U1217 ( .A(n343), .B(n839), .C(n6972), .Y(n3753) );
  OAI21X1 U1219 ( .A(n345), .B(n839), .C(n6969), .Y(n3754) );
  OAI21X1 U1221 ( .A(n347), .B(n839), .C(n6966), .Y(n3755) );
  OAI21X1 U1223 ( .A(n349), .B(n839), .C(n6963), .Y(n3756) );
  OAI21X1 U1225 ( .A(n351), .B(n839), .C(n6960), .Y(n3757) );
  OAI21X1 U1227 ( .A(n353), .B(n839), .C(n6957), .Y(n3758) );
  OAI21X1 U1230 ( .A(n271), .B(n882), .C(n6954), .Y(n3759) );
  OAI21X1 U1232 ( .A(n273), .B(n882), .C(n6951), .Y(n3760) );
  OAI21X1 U1234 ( .A(n275), .B(n882), .C(n6948), .Y(n3761) );
  OAI21X1 U1236 ( .A(n277), .B(n882), .C(n6945), .Y(n3762) );
  OAI21X1 U1238 ( .A(n279), .B(n882), .C(n6942), .Y(n3763) );
  OAI21X1 U1240 ( .A(n281), .B(n882), .C(n6939), .Y(n3764) );
  OAI21X1 U1242 ( .A(n283), .B(n882), .C(n6936), .Y(n3765) );
  OAI21X1 U1244 ( .A(n285), .B(n882), .C(n6933), .Y(n3766) );
  OAI21X1 U1246 ( .A(n287), .B(n882), .C(n6930), .Y(n3767) );
  OAI21X1 U1248 ( .A(n289), .B(n882), .C(n6927), .Y(n3768) );
  OAI21X1 U1250 ( .A(n291), .B(n882), .C(n6924), .Y(n3769) );
  OAI21X1 U1252 ( .A(n293), .B(n882), .C(n6921), .Y(n3770) );
  OAI21X1 U1254 ( .A(n295), .B(n882), .C(n6918), .Y(n3771) );
  OAI21X1 U1256 ( .A(n297), .B(n882), .C(n6915), .Y(n3772) );
  OAI21X1 U1258 ( .A(n299), .B(n882), .C(n6912), .Y(n3773) );
  OAI21X1 U1260 ( .A(n301), .B(n882), .C(n6909), .Y(n3774) );
  OAI21X1 U1262 ( .A(n303), .B(n882), .C(n6906), .Y(n3775) );
  OAI21X1 U1264 ( .A(n305), .B(n882), .C(n6903), .Y(n3776) );
  OAI21X1 U1266 ( .A(n307), .B(n882), .C(n6900), .Y(n3777) );
  OAI21X1 U1268 ( .A(n309), .B(n882), .C(n6897), .Y(n3778) );
  OAI21X1 U1270 ( .A(n311), .B(n882), .C(n6894), .Y(n3779) );
  OAI21X1 U1272 ( .A(n313), .B(n882), .C(n6891), .Y(n3780) );
  OAI21X1 U1274 ( .A(n315), .B(n882), .C(n6888), .Y(n3781) );
  OAI21X1 U1276 ( .A(n317), .B(n882), .C(n6885), .Y(n3782) );
  OAI21X1 U1278 ( .A(n319), .B(n882), .C(n6882), .Y(n3783) );
  OAI21X1 U1280 ( .A(n321), .B(n882), .C(n6879), .Y(n3784) );
  OAI21X1 U1282 ( .A(n323), .B(n882), .C(n6876), .Y(n3785) );
  OAI21X1 U1284 ( .A(n325), .B(n882), .C(n6873), .Y(n3786) );
  OAI21X1 U1286 ( .A(n327), .B(n882), .C(n6870), .Y(n3787) );
  OAI21X1 U1288 ( .A(n329), .B(n882), .C(n6867), .Y(n3788) );
  OAI21X1 U1290 ( .A(n331), .B(n882), .C(n6864), .Y(n3789) );
  OAI21X1 U1292 ( .A(n333), .B(n882), .C(n6861), .Y(n3790) );
  OAI21X1 U1294 ( .A(n335), .B(n882), .C(n6858), .Y(n3791) );
  OAI21X1 U1296 ( .A(n337), .B(n882), .C(n6855), .Y(n3792) );
  OAI21X1 U1298 ( .A(n339), .B(n882), .C(n6852), .Y(n3793) );
  OAI21X1 U1300 ( .A(n341), .B(n882), .C(n6849), .Y(n3794) );
  OAI21X1 U1302 ( .A(n343), .B(n882), .C(n6846), .Y(n3795) );
  OAI21X1 U1304 ( .A(n345), .B(n882), .C(n6843), .Y(n3796) );
  OAI21X1 U1306 ( .A(n347), .B(n882), .C(n6840), .Y(n3797) );
  OAI21X1 U1308 ( .A(n349), .B(n882), .C(n6837), .Y(n3798) );
  OAI21X1 U1310 ( .A(n351), .B(n882), .C(n6834), .Y(n3799) );
  OAI21X1 U1312 ( .A(n353), .B(n882), .C(n6831), .Y(n3800) );
  OAI21X1 U1315 ( .A(n271), .B(n925), .C(n6828), .Y(n3801) );
  OAI21X1 U1317 ( .A(n273), .B(n925), .C(n6825), .Y(n3802) );
  OAI21X1 U1319 ( .A(n275), .B(n925), .C(n6822), .Y(n3803) );
  OAI21X1 U1321 ( .A(n277), .B(n925), .C(n6819), .Y(n3804) );
  OAI21X1 U1323 ( .A(n279), .B(n925), .C(n6816), .Y(n3805) );
  OAI21X1 U1325 ( .A(n281), .B(n925), .C(n6813), .Y(n3806) );
  OAI21X1 U1327 ( .A(n283), .B(n925), .C(n6810), .Y(n3807) );
  OAI21X1 U1329 ( .A(n285), .B(n925), .C(n6807), .Y(n3808) );
  OAI21X1 U1331 ( .A(n287), .B(n925), .C(n6804), .Y(n3809) );
  OAI21X1 U1333 ( .A(n289), .B(n925), .C(n6801), .Y(n3810) );
  OAI21X1 U1335 ( .A(n291), .B(n925), .C(n6798), .Y(n3811) );
  OAI21X1 U1337 ( .A(n293), .B(n925), .C(n6795), .Y(n3812) );
  OAI21X1 U1339 ( .A(n295), .B(n925), .C(n6792), .Y(n3813) );
  OAI21X1 U1341 ( .A(n297), .B(n925), .C(n6789), .Y(n3814) );
  OAI21X1 U1343 ( .A(n299), .B(n925), .C(n6786), .Y(n3815) );
  OAI21X1 U1345 ( .A(n301), .B(n925), .C(n6783), .Y(n3816) );
  OAI21X1 U1347 ( .A(n303), .B(n925), .C(n6780), .Y(n3817) );
  OAI21X1 U1349 ( .A(n305), .B(n925), .C(n6777), .Y(n3818) );
  OAI21X1 U1351 ( .A(n307), .B(n925), .C(n6774), .Y(n3819) );
  OAI21X1 U1353 ( .A(n309), .B(n925), .C(n6771), .Y(n3820) );
  OAI21X1 U1355 ( .A(n311), .B(n925), .C(n6768), .Y(n3821) );
  OAI21X1 U1357 ( .A(n313), .B(n925), .C(n6765), .Y(n3822) );
  OAI21X1 U1359 ( .A(n315), .B(n925), .C(n6762), .Y(n3823) );
  OAI21X1 U1361 ( .A(n317), .B(n925), .C(n6759), .Y(n3824) );
  OAI21X1 U1363 ( .A(n319), .B(n925), .C(n6756), .Y(n3825) );
  OAI21X1 U1365 ( .A(n321), .B(n925), .C(n6753), .Y(n3826) );
  OAI21X1 U1367 ( .A(n323), .B(n925), .C(n6750), .Y(n3827) );
  OAI21X1 U1369 ( .A(n325), .B(n925), .C(n6747), .Y(n3828) );
  OAI21X1 U1371 ( .A(n327), .B(n925), .C(n6744), .Y(n3829) );
  OAI21X1 U1373 ( .A(n329), .B(n925), .C(n6741), .Y(n3830) );
  OAI21X1 U1375 ( .A(n331), .B(n925), .C(n6738), .Y(n3831) );
  OAI21X1 U1377 ( .A(n333), .B(n925), .C(n6735), .Y(n3832) );
  OAI21X1 U1379 ( .A(n335), .B(n925), .C(n6732), .Y(n3833) );
  OAI21X1 U1381 ( .A(n337), .B(n925), .C(n6729), .Y(n3834) );
  OAI21X1 U1383 ( .A(n339), .B(n925), .C(n6726), .Y(n3835) );
  OAI21X1 U1385 ( .A(n341), .B(n925), .C(n6723), .Y(n3836) );
  OAI21X1 U1387 ( .A(n343), .B(n925), .C(n6720), .Y(n3837) );
  OAI21X1 U1389 ( .A(n345), .B(n925), .C(n6717), .Y(n3838) );
  OAI21X1 U1391 ( .A(n347), .B(n925), .C(n6714), .Y(n3839) );
  OAI21X1 U1393 ( .A(n349), .B(n925), .C(n6711), .Y(n3840) );
  OAI21X1 U1395 ( .A(n351), .B(n925), .C(n6708), .Y(n3841) );
  OAI21X1 U1397 ( .A(n353), .B(n925), .C(n6705), .Y(n3842) );
  OAI21X1 U1400 ( .A(n271), .B(n968), .C(n6702), .Y(n3843) );
  OAI21X1 U1402 ( .A(n273), .B(n968), .C(n6699), .Y(n3844) );
  OAI21X1 U1404 ( .A(n275), .B(n968), .C(n6696), .Y(n3845) );
  OAI21X1 U1406 ( .A(n277), .B(n968), .C(n6693), .Y(n3846) );
  OAI21X1 U1408 ( .A(n279), .B(n968), .C(n6690), .Y(n3847) );
  OAI21X1 U1410 ( .A(n281), .B(n968), .C(n6687), .Y(n3848) );
  OAI21X1 U1412 ( .A(n283), .B(n968), .C(n6684), .Y(n3849) );
  OAI21X1 U1414 ( .A(n285), .B(n968), .C(n6681), .Y(n3850) );
  OAI21X1 U1416 ( .A(n287), .B(n968), .C(n6678), .Y(n3851) );
  OAI21X1 U1418 ( .A(n289), .B(n968), .C(n6675), .Y(n3852) );
  OAI21X1 U1420 ( .A(n291), .B(n968), .C(n6672), .Y(n3853) );
  OAI21X1 U1422 ( .A(n293), .B(n968), .C(n6669), .Y(n3854) );
  OAI21X1 U1424 ( .A(n295), .B(n968), .C(n6666), .Y(n3855) );
  OAI21X1 U1426 ( .A(n297), .B(n968), .C(n6663), .Y(n3856) );
  OAI21X1 U1428 ( .A(n299), .B(n968), .C(n6660), .Y(n3857) );
  OAI21X1 U1430 ( .A(n301), .B(n968), .C(n6657), .Y(n3858) );
  OAI21X1 U1432 ( .A(n303), .B(n968), .C(n6654), .Y(n3859) );
  OAI21X1 U1434 ( .A(n305), .B(n968), .C(n6651), .Y(n3860) );
  OAI21X1 U1436 ( .A(n307), .B(n968), .C(n6648), .Y(n3861) );
  OAI21X1 U1438 ( .A(n309), .B(n968), .C(n6645), .Y(n3862) );
  OAI21X1 U1440 ( .A(n311), .B(n968), .C(n6642), .Y(n3863) );
  OAI21X1 U1442 ( .A(n313), .B(n968), .C(n6639), .Y(n3864) );
  OAI21X1 U1444 ( .A(n315), .B(n968), .C(n6636), .Y(n3865) );
  OAI21X1 U1446 ( .A(n317), .B(n968), .C(n6633), .Y(n3866) );
  OAI21X1 U1448 ( .A(n319), .B(n968), .C(n6630), .Y(n3867) );
  OAI21X1 U1450 ( .A(n321), .B(n968), .C(n6627), .Y(n3868) );
  OAI21X1 U1452 ( .A(n323), .B(n968), .C(n6624), .Y(n3869) );
  OAI21X1 U1454 ( .A(n325), .B(n968), .C(n6621), .Y(n3870) );
  OAI21X1 U1456 ( .A(n327), .B(n968), .C(n6618), .Y(n3871) );
  OAI21X1 U1458 ( .A(n329), .B(n968), .C(n6615), .Y(n3872) );
  OAI21X1 U1460 ( .A(n331), .B(n968), .C(n6612), .Y(n3873) );
  OAI21X1 U1462 ( .A(n333), .B(n968), .C(n6609), .Y(n3874) );
  OAI21X1 U1464 ( .A(n335), .B(n968), .C(n6606), .Y(n3875) );
  OAI21X1 U1466 ( .A(n337), .B(n968), .C(n6603), .Y(n3876) );
  OAI21X1 U1468 ( .A(n339), .B(n968), .C(n6600), .Y(n3877) );
  OAI21X1 U1470 ( .A(n341), .B(n968), .C(n6597), .Y(n3878) );
  OAI21X1 U1472 ( .A(n343), .B(n968), .C(n6594), .Y(n3879) );
  OAI21X1 U1474 ( .A(n345), .B(n968), .C(n6591), .Y(n3880) );
  OAI21X1 U1476 ( .A(n347), .B(n968), .C(n6588), .Y(n3881) );
  OAI21X1 U1478 ( .A(n349), .B(n968), .C(n6585), .Y(n3882) );
  OAI21X1 U1480 ( .A(n351), .B(n968), .C(n6582), .Y(n3883) );
  OAI21X1 U1482 ( .A(n353), .B(n968), .C(n6579), .Y(n3884) );
  NAND3X1 U1486 ( .A(n253), .B(n254), .C(n13011), .Y(n1011) );
  INVX1 U1487 ( .A(n13019), .Y(n254) );
  OAI21X1 U1488 ( .A(n271), .B(n1012), .C(n6576), .Y(n3885) );
  OAI21X1 U1490 ( .A(n273), .B(n1012), .C(n6573), .Y(n3886) );
  OAI21X1 U1492 ( .A(n275), .B(n1012), .C(n6570), .Y(n3887) );
  OAI21X1 U1494 ( .A(n277), .B(n1012), .C(n6567), .Y(n3888) );
  OAI21X1 U1496 ( .A(n279), .B(n1012), .C(n6564), .Y(n3889) );
  OAI21X1 U1498 ( .A(n281), .B(n1012), .C(n6561), .Y(n3890) );
  OAI21X1 U1500 ( .A(n283), .B(n1012), .C(n6558), .Y(n3891) );
  OAI21X1 U1502 ( .A(n285), .B(n1012), .C(n6555), .Y(n3892) );
  OAI21X1 U1504 ( .A(n287), .B(n1012), .C(n6552), .Y(n3893) );
  OAI21X1 U1506 ( .A(n289), .B(n1012), .C(n6549), .Y(n3894) );
  OAI21X1 U1508 ( .A(n291), .B(n1012), .C(n6546), .Y(n3895) );
  OAI21X1 U1510 ( .A(n293), .B(n1012), .C(n6543), .Y(n3896) );
  OAI21X1 U1512 ( .A(n295), .B(n1012), .C(n6540), .Y(n3897) );
  OAI21X1 U1514 ( .A(n297), .B(n1012), .C(n6537), .Y(n3898) );
  OAI21X1 U1516 ( .A(n299), .B(n1012), .C(n6534), .Y(n3899) );
  OAI21X1 U1518 ( .A(n301), .B(n1012), .C(n6531), .Y(n3900) );
  OAI21X1 U1520 ( .A(n303), .B(n1012), .C(n6528), .Y(n3901) );
  OAI21X1 U1522 ( .A(n305), .B(n1012), .C(n6525), .Y(n3902) );
  OAI21X1 U1524 ( .A(n307), .B(n1012), .C(n6522), .Y(n3903) );
  OAI21X1 U1526 ( .A(n309), .B(n1012), .C(n6519), .Y(n3904) );
  OAI21X1 U1528 ( .A(n311), .B(n1012), .C(n6516), .Y(n3905) );
  OAI21X1 U1530 ( .A(n313), .B(n1012), .C(n6513), .Y(n3906) );
  OAI21X1 U1532 ( .A(n315), .B(n1012), .C(n6510), .Y(n3907) );
  OAI21X1 U1534 ( .A(n317), .B(n1012), .C(n6507), .Y(n3908) );
  OAI21X1 U1536 ( .A(n319), .B(n1012), .C(n6504), .Y(n3909) );
  OAI21X1 U1538 ( .A(n321), .B(n1012), .C(n6501), .Y(n3910) );
  OAI21X1 U1540 ( .A(n323), .B(n1012), .C(n6498), .Y(n3911) );
  OAI21X1 U1542 ( .A(n325), .B(n1012), .C(n6495), .Y(n3912) );
  OAI21X1 U1544 ( .A(n327), .B(n1012), .C(n6492), .Y(n3913) );
  OAI21X1 U1546 ( .A(n329), .B(n1012), .C(n6489), .Y(n3914) );
  OAI21X1 U1548 ( .A(n331), .B(n1012), .C(n6486), .Y(n3915) );
  OAI21X1 U1550 ( .A(n333), .B(n1012), .C(n6483), .Y(n3916) );
  OAI21X1 U1552 ( .A(n335), .B(n1012), .C(n6480), .Y(n3917) );
  OAI21X1 U1554 ( .A(n337), .B(n1012), .C(n6477), .Y(n3918) );
  OAI21X1 U1556 ( .A(n339), .B(n1012), .C(n6474), .Y(n3919) );
  OAI21X1 U1558 ( .A(n341), .B(n1012), .C(n6471), .Y(n3920) );
  OAI21X1 U1560 ( .A(n343), .B(n1012), .C(n6468), .Y(n3921) );
  OAI21X1 U1562 ( .A(n345), .B(n1012), .C(n6465), .Y(n3922) );
  OAI21X1 U1564 ( .A(n347), .B(n1012), .C(n6462), .Y(n3923) );
  OAI21X1 U1566 ( .A(n349), .B(n1012), .C(n6459), .Y(n3924) );
  OAI21X1 U1568 ( .A(n351), .B(n1012), .C(n6456), .Y(n3925) );
  OAI21X1 U1570 ( .A(n353), .B(n1012), .C(n6453), .Y(n3926) );
  OAI21X1 U1573 ( .A(n271), .B(n1056), .C(n6450), .Y(n3927) );
  OAI21X1 U1575 ( .A(n273), .B(n1056), .C(n6447), .Y(n3928) );
  OAI21X1 U1577 ( .A(n275), .B(n1056), .C(n6444), .Y(n3929) );
  OAI21X1 U1579 ( .A(n277), .B(n1056), .C(n6441), .Y(n3930) );
  OAI21X1 U1581 ( .A(n279), .B(n1056), .C(n6438), .Y(n3931) );
  OAI21X1 U1583 ( .A(n281), .B(n1056), .C(n6435), .Y(n3932) );
  OAI21X1 U1585 ( .A(n283), .B(n1056), .C(n6432), .Y(n3933) );
  OAI21X1 U1587 ( .A(n285), .B(n1056), .C(n6429), .Y(n3934) );
  OAI21X1 U1589 ( .A(n287), .B(n1056), .C(n6426), .Y(n3935) );
  OAI21X1 U1591 ( .A(n289), .B(n1056), .C(n6423), .Y(n3936) );
  OAI21X1 U1593 ( .A(n291), .B(n1056), .C(n6420), .Y(n3937) );
  OAI21X1 U1595 ( .A(n293), .B(n1056), .C(n6417), .Y(n3938) );
  OAI21X1 U1597 ( .A(n295), .B(n1056), .C(n6414), .Y(n3939) );
  OAI21X1 U1599 ( .A(n297), .B(n1056), .C(n6411), .Y(n3940) );
  OAI21X1 U1601 ( .A(n299), .B(n1056), .C(n6408), .Y(n3941) );
  OAI21X1 U1603 ( .A(n301), .B(n1056), .C(n6405), .Y(n3942) );
  OAI21X1 U1605 ( .A(n303), .B(n1056), .C(n6402), .Y(n3943) );
  OAI21X1 U1607 ( .A(n305), .B(n1056), .C(n6399), .Y(n3944) );
  OAI21X1 U1609 ( .A(n307), .B(n1056), .C(n6396), .Y(n3945) );
  OAI21X1 U1611 ( .A(n309), .B(n1056), .C(n6393), .Y(n3946) );
  OAI21X1 U1613 ( .A(n311), .B(n1056), .C(n6390), .Y(n3947) );
  OAI21X1 U1615 ( .A(n313), .B(n1056), .C(n6387), .Y(n3948) );
  OAI21X1 U1617 ( .A(n315), .B(n1056), .C(n6384), .Y(n3949) );
  OAI21X1 U1619 ( .A(n317), .B(n1056), .C(n6381), .Y(n3950) );
  OAI21X1 U1621 ( .A(n319), .B(n1056), .C(n6378), .Y(n3951) );
  OAI21X1 U1623 ( .A(n321), .B(n1056), .C(n6375), .Y(n3952) );
  OAI21X1 U1625 ( .A(n323), .B(n1056), .C(n6372), .Y(n3953) );
  OAI21X1 U1627 ( .A(n325), .B(n1056), .C(n6369), .Y(n3954) );
  OAI21X1 U1629 ( .A(n327), .B(n1056), .C(n6366), .Y(n3955) );
  OAI21X1 U1631 ( .A(n329), .B(n1056), .C(n6363), .Y(n3956) );
  OAI21X1 U1633 ( .A(n331), .B(n1056), .C(n6360), .Y(n3957) );
  OAI21X1 U1635 ( .A(n333), .B(n1056), .C(n6357), .Y(n3958) );
  OAI21X1 U1637 ( .A(n335), .B(n1056), .C(n6354), .Y(n3959) );
  OAI21X1 U1639 ( .A(n337), .B(n1056), .C(n6351), .Y(n3960) );
  OAI21X1 U1641 ( .A(n339), .B(n1056), .C(n6348), .Y(n3961) );
  OAI21X1 U1643 ( .A(n341), .B(n1056), .C(n6345), .Y(n3962) );
  OAI21X1 U1645 ( .A(n343), .B(n1056), .C(n6342), .Y(n3963) );
  OAI21X1 U1647 ( .A(n345), .B(n1056), .C(n6339), .Y(n3964) );
  OAI21X1 U1649 ( .A(n347), .B(n1056), .C(n6336), .Y(n3965) );
  OAI21X1 U1651 ( .A(n349), .B(n1056), .C(n6333), .Y(n3966) );
  OAI21X1 U1653 ( .A(n351), .B(n1056), .C(n6330), .Y(n3967) );
  OAI21X1 U1655 ( .A(n353), .B(n1056), .C(n6327), .Y(n3968) );
  OAI21X1 U1658 ( .A(n271), .B(n1099), .C(n6324), .Y(n3969) );
  OAI21X1 U1660 ( .A(n273), .B(n1099), .C(n6321), .Y(n3970) );
  OAI21X1 U1662 ( .A(n275), .B(n1099), .C(n6318), .Y(n3971) );
  OAI21X1 U1664 ( .A(n277), .B(n1099), .C(n6315), .Y(n3972) );
  OAI21X1 U1666 ( .A(n279), .B(n1099), .C(n6312), .Y(n3973) );
  OAI21X1 U1668 ( .A(n281), .B(n1099), .C(n6309), .Y(n3974) );
  OAI21X1 U1670 ( .A(n283), .B(n1099), .C(n6306), .Y(n3975) );
  OAI21X1 U1672 ( .A(n285), .B(n1099), .C(n6303), .Y(n3976) );
  OAI21X1 U1674 ( .A(n287), .B(n1099), .C(n6300), .Y(n3977) );
  OAI21X1 U1676 ( .A(n289), .B(n1099), .C(n6297), .Y(n3978) );
  OAI21X1 U1678 ( .A(n291), .B(n1099), .C(n6294), .Y(n3979) );
  OAI21X1 U1680 ( .A(n293), .B(n1099), .C(n6291), .Y(n3980) );
  OAI21X1 U1682 ( .A(n295), .B(n1099), .C(n6288), .Y(n3981) );
  OAI21X1 U1684 ( .A(n297), .B(n1099), .C(n6285), .Y(n3982) );
  OAI21X1 U1686 ( .A(n299), .B(n1099), .C(n6282), .Y(n3983) );
  OAI21X1 U1688 ( .A(n301), .B(n1099), .C(n6279), .Y(n3984) );
  OAI21X1 U1690 ( .A(n303), .B(n1099), .C(n6276), .Y(n3985) );
  OAI21X1 U1692 ( .A(n305), .B(n1099), .C(n6273), .Y(n3986) );
  OAI21X1 U1694 ( .A(n307), .B(n1099), .C(n6270), .Y(n3987) );
  OAI21X1 U1696 ( .A(n309), .B(n1099), .C(n6267), .Y(n3988) );
  OAI21X1 U1698 ( .A(n311), .B(n1099), .C(n6264), .Y(n3989) );
  OAI21X1 U1700 ( .A(n313), .B(n1099), .C(n6261), .Y(n3990) );
  OAI21X1 U1702 ( .A(n315), .B(n1099), .C(n6258), .Y(n3991) );
  OAI21X1 U1704 ( .A(n317), .B(n1099), .C(n6255), .Y(n3992) );
  OAI21X1 U1706 ( .A(n319), .B(n1099), .C(n6252), .Y(n3993) );
  OAI21X1 U1708 ( .A(n321), .B(n1099), .C(n6249), .Y(n3994) );
  OAI21X1 U1710 ( .A(n323), .B(n1099), .C(n6246), .Y(n3995) );
  OAI21X1 U1712 ( .A(n325), .B(n1099), .C(n6243), .Y(n3996) );
  OAI21X1 U1714 ( .A(n327), .B(n1099), .C(n6240), .Y(n3997) );
  OAI21X1 U1716 ( .A(n329), .B(n1099), .C(n6237), .Y(n3998) );
  OAI21X1 U1718 ( .A(n331), .B(n1099), .C(n6234), .Y(n3999) );
  OAI21X1 U1720 ( .A(n333), .B(n1099), .C(n6231), .Y(n4000) );
  OAI21X1 U1722 ( .A(n335), .B(n1099), .C(n6228), .Y(n4001) );
  OAI21X1 U1724 ( .A(n337), .B(n1099), .C(n6225), .Y(n4002) );
  OAI21X1 U1726 ( .A(n339), .B(n1099), .C(n6222), .Y(n4003) );
  OAI21X1 U1728 ( .A(n341), .B(n1099), .C(n6219), .Y(n4004) );
  OAI21X1 U1730 ( .A(n343), .B(n1099), .C(n6216), .Y(n4005) );
  OAI21X1 U1732 ( .A(n345), .B(n1099), .C(n6213), .Y(n4006) );
  OAI21X1 U1734 ( .A(n347), .B(n1099), .C(n6210), .Y(n4007) );
  OAI21X1 U1736 ( .A(n349), .B(n1099), .C(n6207), .Y(n4008) );
  OAI21X1 U1738 ( .A(n351), .B(n1099), .C(n6204), .Y(n4009) );
  OAI21X1 U1740 ( .A(n353), .B(n1099), .C(n6201), .Y(n4010) );
  OAI21X1 U1743 ( .A(n271), .B(n1142), .C(n6198), .Y(n4011) );
  OAI21X1 U1745 ( .A(n273), .B(n1142), .C(n6195), .Y(n4012) );
  OAI21X1 U1747 ( .A(n275), .B(n1142), .C(n6192), .Y(n4013) );
  OAI21X1 U1749 ( .A(n277), .B(n1142), .C(n6189), .Y(n4014) );
  OAI21X1 U1751 ( .A(n279), .B(n1142), .C(n6186), .Y(n4015) );
  OAI21X1 U1753 ( .A(n281), .B(n1142), .C(n6183), .Y(n4016) );
  OAI21X1 U1755 ( .A(n283), .B(n1142), .C(n6180), .Y(n4017) );
  OAI21X1 U1757 ( .A(n285), .B(n1142), .C(n6177), .Y(n4018) );
  OAI21X1 U1759 ( .A(n287), .B(n1142), .C(n6174), .Y(n4019) );
  OAI21X1 U1761 ( .A(n289), .B(n1142), .C(n6171), .Y(n4020) );
  OAI21X1 U1763 ( .A(n291), .B(n1142), .C(n6168), .Y(n4021) );
  OAI21X1 U1765 ( .A(n293), .B(n1142), .C(n6165), .Y(n4022) );
  OAI21X1 U1767 ( .A(n295), .B(n1142), .C(n6162), .Y(n4023) );
  OAI21X1 U1769 ( .A(n297), .B(n1142), .C(n6159), .Y(n4024) );
  OAI21X1 U1771 ( .A(n299), .B(n1142), .C(n6156), .Y(n4025) );
  OAI21X1 U1773 ( .A(n301), .B(n1142), .C(n6153), .Y(n4026) );
  OAI21X1 U1775 ( .A(n303), .B(n1142), .C(n6150), .Y(n4027) );
  OAI21X1 U1777 ( .A(n305), .B(n1142), .C(n6147), .Y(n4028) );
  OAI21X1 U1779 ( .A(n307), .B(n1142), .C(n6144), .Y(n4029) );
  OAI21X1 U1781 ( .A(n309), .B(n1142), .C(n6141), .Y(n4030) );
  OAI21X1 U1783 ( .A(n311), .B(n1142), .C(n6138), .Y(n4031) );
  OAI21X1 U1785 ( .A(n313), .B(n1142), .C(n6135), .Y(n4032) );
  OAI21X1 U1787 ( .A(n315), .B(n1142), .C(n6132), .Y(n4033) );
  OAI21X1 U1789 ( .A(n317), .B(n1142), .C(n6129), .Y(n4034) );
  OAI21X1 U1791 ( .A(n319), .B(n1142), .C(n6126), .Y(n4035) );
  OAI21X1 U1793 ( .A(n321), .B(n1142), .C(n6123), .Y(n4036) );
  OAI21X1 U1795 ( .A(n323), .B(n1142), .C(n6120), .Y(n4037) );
  OAI21X1 U1797 ( .A(n325), .B(n1142), .C(n6117), .Y(n4038) );
  OAI21X1 U1799 ( .A(n327), .B(n1142), .C(n6114), .Y(n4039) );
  OAI21X1 U1801 ( .A(n329), .B(n1142), .C(n6111), .Y(n4040) );
  OAI21X1 U1803 ( .A(n331), .B(n1142), .C(n6108), .Y(n4041) );
  OAI21X1 U1805 ( .A(n333), .B(n1142), .C(n6105), .Y(n4042) );
  OAI21X1 U1807 ( .A(n335), .B(n1142), .C(n6102), .Y(n4043) );
  OAI21X1 U1809 ( .A(n337), .B(n1142), .C(n6099), .Y(n4044) );
  OAI21X1 U1811 ( .A(n339), .B(n1142), .C(n6096), .Y(n4045) );
  OAI21X1 U1813 ( .A(n341), .B(n1142), .C(n6093), .Y(n4046) );
  OAI21X1 U1815 ( .A(n343), .B(n1142), .C(n6090), .Y(n4047) );
  OAI21X1 U1817 ( .A(n345), .B(n1142), .C(n6087), .Y(n4048) );
  OAI21X1 U1819 ( .A(n347), .B(n1142), .C(n6084), .Y(n4049) );
  OAI21X1 U1821 ( .A(n349), .B(n1142), .C(n6081), .Y(n4050) );
  OAI21X1 U1823 ( .A(n351), .B(n1142), .C(n6078), .Y(n4051) );
  OAI21X1 U1825 ( .A(n353), .B(n1142), .C(n6075), .Y(n4052) );
  OAI21X1 U1828 ( .A(n271), .B(n1185), .C(n6072), .Y(n4053) );
  OAI21X1 U1830 ( .A(n273), .B(n1185), .C(n6069), .Y(n4054) );
  OAI21X1 U1832 ( .A(n275), .B(n1185), .C(n6066), .Y(n4055) );
  OAI21X1 U1834 ( .A(n277), .B(n1185), .C(n6063), .Y(n4056) );
  OAI21X1 U1836 ( .A(n279), .B(n1185), .C(n6060), .Y(n4057) );
  OAI21X1 U1838 ( .A(n281), .B(n1185), .C(n6057), .Y(n4058) );
  OAI21X1 U1840 ( .A(n283), .B(n1185), .C(n6054), .Y(n4059) );
  OAI21X1 U1842 ( .A(n285), .B(n1185), .C(n6051), .Y(n4060) );
  OAI21X1 U1844 ( .A(n287), .B(n1185), .C(n6048), .Y(n4061) );
  OAI21X1 U1846 ( .A(n289), .B(n1185), .C(n6045), .Y(n4062) );
  OAI21X1 U1848 ( .A(n291), .B(n1185), .C(n6042), .Y(n4063) );
  OAI21X1 U1850 ( .A(n293), .B(n1185), .C(n6039), .Y(n4064) );
  OAI21X1 U1852 ( .A(n295), .B(n1185), .C(n6036), .Y(n4065) );
  OAI21X1 U1854 ( .A(n297), .B(n1185), .C(n6033), .Y(n4066) );
  OAI21X1 U1856 ( .A(n299), .B(n1185), .C(n6030), .Y(n4067) );
  OAI21X1 U1858 ( .A(n301), .B(n1185), .C(n6027), .Y(n4068) );
  OAI21X1 U1860 ( .A(n303), .B(n1185), .C(n6024), .Y(n4069) );
  OAI21X1 U1862 ( .A(n305), .B(n1185), .C(n6021), .Y(n4070) );
  OAI21X1 U1864 ( .A(n307), .B(n1185), .C(n6018), .Y(n4071) );
  OAI21X1 U1866 ( .A(n309), .B(n1185), .C(n6015), .Y(n4072) );
  OAI21X1 U1868 ( .A(n311), .B(n1185), .C(n6012), .Y(n4073) );
  OAI21X1 U1870 ( .A(n313), .B(n1185), .C(n6009), .Y(n4074) );
  OAI21X1 U1872 ( .A(n315), .B(n1185), .C(n6006), .Y(n4075) );
  OAI21X1 U1874 ( .A(n317), .B(n1185), .C(n6003), .Y(n4076) );
  OAI21X1 U1876 ( .A(n319), .B(n1185), .C(n6000), .Y(n4077) );
  OAI21X1 U1878 ( .A(n321), .B(n1185), .C(n5997), .Y(n4078) );
  OAI21X1 U1880 ( .A(n323), .B(n1185), .C(n5994), .Y(n4079) );
  OAI21X1 U1882 ( .A(n325), .B(n1185), .C(n5991), .Y(n4080) );
  OAI21X1 U1884 ( .A(n327), .B(n1185), .C(n5988), .Y(n4081) );
  OAI21X1 U1886 ( .A(n329), .B(n1185), .C(n5985), .Y(n4082) );
  OAI21X1 U1888 ( .A(n331), .B(n1185), .C(n5982), .Y(n4083) );
  OAI21X1 U1890 ( .A(n333), .B(n1185), .C(n5979), .Y(n4084) );
  OAI21X1 U1892 ( .A(n335), .B(n1185), .C(n5976), .Y(n4085) );
  OAI21X1 U1894 ( .A(n337), .B(n1185), .C(n5973), .Y(n4086) );
  OAI21X1 U1896 ( .A(n339), .B(n1185), .C(n5970), .Y(n4087) );
  OAI21X1 U1898 ( .A(n341), .B(n1185), .C(n5967), .Y(n4088) );
  OAI21X1 U1900 ( .A(n343), .B(n1185), .C(n5964), .Y(n4089) );
  OAI21X1 U1902 ( .A(n345), .B(n1185), .C(n5961), .Y(n4090) );
  OAI21X1 U1904 ( .A(n347), .B(n1185), .C(n5958), .Y(n4091) );
  OAI21X1 U1906 ( .A(n349), .B(n1185), .C(n5955), .Y(n4092) );
  OAI21X1 U1908 ( .A(n351), .B(n1185), .C(n5952), .Y(n4093) );
  OAI21X1 U1910 ( .A(n353), .B(n1185), .C(n5949), .Y(n4094) );
  OAI21X1 U1913 ( .A(n271), .B(n12962), .C(n5946), .Y(n4095) );
  OAI21X1 U1915 ( .A(n273), .B(n8704), .C(n5943), .Y(n4096) );
  OAI21X1 U1917 ( .A(n275), .B(n13034), .C(n5940), .Y(n4097) );
  OAI21X1 U1919 ( .A(n277), .B(n8672), .C(n5937), .Y(n4098) );
  OAI21X1 U1921 ( .A(n279), .B(n8716), .C(n5934), .Y(n4099) );
  OAI21X1 U1923 ( .A(n281), .B(n13034), .C(n5931), .Y(n4100) );
  OAI21X1 U1925 ( .A(n283), .B(n8682), .C(n5928), .Y(n4101) );
  OAI21X1 U1927 ( .A(n285), .B(n13035), .C(n5925), .Y(n4102) );
  OAI21X1 U1929 ( .A(n287), .B(n13034), .C(n5922), .Y(n4103) );
  OAI21X1 U1931 ( .A(n289), .B(n12975), .C(n5919), .Y(n4104) );
  OAI21X1 U1933 ( .A(n291), .B(n13026), .C(n5916), .Y(n4105) );
  OAI21X1 U1935 ( .A(n293), .B(n13034), .C(n5913), .Y(n4106) );
  OAI21X1 U1937 ( .A(n295), .B(n13036), .C(n5910), .Y(n4107) );
  OAI21X1 U1939 ( .A(n297), .B(n13026), .C(n5907), .Y(n4108) );
  OAI21X1 U1941 ( .A(n299), .B(n13034), .C(n5904), .Y(n4109) );
  OAI21X1 U1943 ( .A(n301), .B(n8694), .C(n5901), .Y(n4110) );
  OAI21X1 U1945 ( .A(n303), .B(n13035), .C(n5898), .Y(n4111) );
  OAI21X1 U1947 ( .A(n305), .B(n13034), .C(n5895), .Y(n4112) );
  OAI21X1 U1949 ( .A(n307), .B(n8772), .C(n5892), .Y(n4113) );
  OAI21X1 U1951 ( .A(n309), .B(n13026), .C(n5889), .Y(n4114) );
  OAI21X1 U1953 ( .A(n311), .B(n13034), .C(n5886), .Y(n4115) );
  OAI21X1 U1955 ( .A(n313), .B(n13036), .C(n5883), .Y(n4116) );
  OAI21X1 U1957 ( .A(n315), .B(n12984), .C(n5880), .Y(n4117) );
  OAI21X1 U1959 ( .A(n317), .B(n13034), .C(n5877), .Y(n4118) );
  OAI21X1 U1961 ( .A(n319), .B(n13026), .C(n5874), .Y(n4119) );
  OAI21X1 U1963 ( .A(n321), .B(n8710), .C(n5871), .Y(n4120) );
  OAI21X1 U1965 ( .A(n323), .B(n13034), .C(n5868), .Y(n4121) );
  OAI21X1 U1967 ( .A(n325), .B(n12984), .C(n5865), .Y(n4122) );
  OAI21X1 U1969 ( .A(n327), .B(n8702), .C(n5862), .Y(n4123) );
  OAI21X1 U1971 ( .A(n329), .B(n13034), .C(n5859), .Y(n4124) );
  OAI21X1 U1973 ( .A(n331), .B(n13035), .C(n5856), .Y(n4125) );
  OAI21X1 U1975 ( .A(n333), .B(n13036), .C(n5853), .Y(n4126) );
  OAI21X1 U1977 ( .A(n335), .B(n13034), .C(n5850), .Y(n4127) );
  OAI21X1 U1979 ( .A(n337), .B(n13026), .C(n5847), .Y(n4128) );
  OAI21X1 U1981 ( .A(n339), .B(n13026), .C(n5844), .Y(n4129) );
  OAI21X1 U1983 ( .A(n341), .B(n13034), .C(n5841), .Y(n4130) );
  OAI21X1 U1985 ( .A(n343), .B(n12975), .C(n5838), .Y(n4131) );
  OAI21X1 U1987 ( .A(n345), .B(n12984), .C(n5835), .Y(n4132) );
  OAI21X1 U1989 ( .A(n347), .B(n13034), .C(n5832), .Y(n4133) );
  OAI21X1 U1991 ( .A(n349), .B(n8724), .C(n5829), .Y(n4134) );
  OAI21X1 U1993 ( .A(n351), .B(n10802), .C(n5826), .Y(n4135) );
  OAI21X1 U1995 ( .A(n353), .B(n13034), .C(n5823), .Y(n4136) );
  OAI21X1 U1998 ( .A(n271), .B(n1271), .C(n5820), .Y(n4137) );
  OAI21X1 U2000 ( .A(n273), .B(n1271), .C(n5817), .Y(n4138) );
  OAI21X1 U2002 ( .A(n275), .B(n1271), .C(n5814), .Y(n4139) );
  OAI21X1 U2004 ( .A(n277), .B(n1271), .C(n5811), .Y(n4140) );
  OAI21X1 U2006 ( .A(n279), .B(n1271), .C(n5808), .Y(n4141) );
  OAI21X1 U2008 ( .A(n281), .B(n1271), .C(n5805), .Y(n4142) );
  OAI21X1 U2010 ( .A(n283), .B(n1271), .C(n5802), .Y(n4143) );
  OAI21X1 U2012 ( .A(n285), .B(n1271), .C(n5799), .Y(n4144) );
  OAI21X1 U2014 ( .A(n287), .B(n1271), .C(n5796), .Y(n4145) );
  OAI21X1 U2016 ( .A(n289), .B(n1271), .C(n5793), .Y(n4146) );
  OAI21X1 U2018 ( .A(n291), .B(n1271), .C(n5790), .Y(n4147) );
  OAI21X1 U2020 ( .A(n293), .B(n1271), .C(n5787), .Y(n4148) );
  OAI21X1 U2022 ( .A(n295), .B(n1271), .C(n5784), .Y(n4149) );
  OAI21X1 U2024 ( .A(n297), .B(n1271), .C(n5781), .Y(n4150) );
  OAI21X1 U2026 ( .A(n299), .B(n1271), .C(n5778), .Y(n4151) );
  OAI21X1 U2028 ( .A(n301), .B(n1271), .C(n5775), .Y(n4152) );
  OAI21X1 U2030 ( .A(n303), .B(n1271), .C(n5772), .Y(n4153) );
  OAI21X1 U2032 ( .A(n305), .B(n1271), .C(n5769), .Y(n4154) );
  OAI21X1 U2034 ( .A(n307), .B(n1271), .C(n5766), .Y(n4155) );
  OAI21X1 U2036 ( .A(n309), .B(n1271), .C(n5763), .Y(n4156) );
  OAI21X1 U2038 ( .A(n311), .B(n1271), .C(n5760), .Y(n4157) );
  OAI21X1 U2040 ( .A(n313), .B(n1271), .C(n5757), .Y(n4158) );
  OAI21X1 U2042 ( .A(n315), .B(n1271), .C(n5754), .Y(n4159) );
  OAI21X1 U2044 ( .A(n317), .B(n1271), .C(n5751), .Y(n4160) );
  OAI21X1 U2046 ( .A(n319), .B(n1271), .C(n5748), .Y(n4161) );
  OAI21X1 U2048 ( .A(n321), .B(n1271), .C(n5745), .Y(n4162) );
  OAI21X1 U2050 ( .A(n323), .B(n1271), .C(n5742), .Y(n4163) );
  OAI21X1 U2052 ( .A(n325), .B(n1271), .C(n5739), .Y(n4164) );
  OAI21X1 U2054 ( .A(n327), .B(n1271), .C(n5736), .Y(n4165) );
  OAI21X1 U2056 ( .A(n329), .B(n1271), .C(n5733), .Y(n4166) );
  OAI21X1 U2058 ( .A(n331), .B(n1271), .C(n5730), .Y(n4167) );
  OAI21X1 U2060 ( .A(n333), .B(n1271), .C(n5727), .Y(n4168) );
  OAI21X1 U2062 ( .A(n335), .B(n1271), .C(n5724), .Y(n4169) );
  OAI21X1 U2064 ( .A(n337), .B(n1271), .C(n5721), .Y(n4170) );
  OAI21X1 U2066 ( .A(n339), .B(n1271), .C(n5718), .Y(n4171) );
  OAI21X1 U2068 ( .A(n341), .B(n1271), .C(n5715), .Y(n4172) );
  OAI21X1 U2070 ( .A(n343), .B(n1271), .C(n5712), .Y(n4173) );
  OAI21X1 U2072 ( .A(n345), .B(n1271), .C(n5709), .Y(n4174) );
  OAI21X1 U2074 ( .A(n347), .B(n1271), .C(n5706), .Y(n4175) );
  OAI21X1 U2076 ( .A(n349), .B(n1271), .C(n5703), .Y(n4176) );
  OAI21X1 U2078 ( .A(n351), .B(n1271), .C(n5700), .Y(n4177) );
  OAI21X1 U2080 ( .A(n353), .B(n1271), .C(n5697), .Y(n4178) );
  OAI21X1 U2083 ( .A(n271), .B(n1314), .C(n5694), .Y(n4179) );
  OAI21X1 U2085 ( .A(n273), .B(n1314), .C(n5691), .Y(n4180) );
  OAI21X1 U2087 ( .A(n275), .B(n1314), .C(n5688), .Y(n4181) );
  OAI21X1 U2089 ( .A(n277), .B(n1314), .C(n5685), .Y(n4182) );
  OAI21X1 U2091 ( .A(n279), .B(n1314), .C(n5682), .Y(n4183) );
  OAI21X1 U2093 ( .A(n281), .B(n1314), .C(n5679), .Y(n4184) );
  OAI21X1 U2095 ( .A(n283), .B(n1314), .C(n5676), .Y(n4185) );
  OAI21X1 U2097 ( .A(n285), .B(n1314), .C(n5673), .Y(n4186) );
  OAI21X1 U2099 ( .A(n287), .B(n1314), .C(n5670), .Y(n4187) );
  OAI21X1 U2101 ( .A(n289), .B(n1314), .C(n5667), .Y(n4188) );
  OAI21X1 U2103 ( .A(n291), .B(n1314), .C(n5664), .Y(n4189) );
  OAI21X1 U2105 ( .A(n293), .B(n1314), .C(n5661), .Y(n4190) );
  OAI21X1 U2107 ( .A(n295), .B(n1314), .C(n5658), .Y(n4191) );
  OAI21X1 U2109 ( .A(n297), .B(n1314), .C(n5655), .Y(n4192) );
  OAI21X1 U2111 ( .A(n299), .B(n1314), .C(n5652), .Y(n4193) );
  OAI21X1 U2113 ( .A(n301), .B(n1314), .C(n5649), .Y(n4194) );
  OAI21X1 U2115 ( .A(n303), .B(n1314), .C(n5646), .Y(n4195) );
  OAI21X1 U2117 ( .A(n305), .B(n1314), .C(n5643), .Y(n4196) );
  OAI21X1 U2119 ( .A(n307), .B(n1314), .C(n5640), .Y(n4197) );
  OAI21X1 U2121 ( .A(n309), .B(n1314), .C(n5637), .Y(n4198) );
  OAI21X1 U2123 ( .A(n311), .B(n1314), .C(n5634), .Y(n4199) );
  OAI21X1 U2125 ( .A(n313), .B(n1314), .C(n5631), .Y(n4200) );
  OAI21X1 U2127 ( .A(n315), .B(n1314), .C(n5628), .Y(n4201) );
  OAI21X1 U2129 ( .A(n317), .B(n1314), .C(n5625), .Y(n4202) );
  OAI21X1 U2131 ( .A(n319), .B(n1314), .C(n5622), .Y(n4203) );
  OAI21X1 U2133 ( .A(n321), .B(n1314), .C(n5619), .Y(n4204) );
  OAI21X1 U2135 ( .A(n323), .B(n1314), .C(n5616), .Y(n4205) );
  OAI21X1 U2137 ( .A(n325), .B(n1314), .C(n5613), .Y(n4206) );
  OAI21X1 U2139 ( .A(n327), .B(n1314), .C(n5610), .Y(n4207) );
  OAI21X1 U2141 ( .A(n329), .B(n1314), .C(n5607), .Y(n4208) );
  OAI21X1 U2143 ( .A(n331), .B(n1314), .C(n5604), .Y(n4209) );
  OAI21X1 U2145 ( .A(n333), .B(n1314), .C(n5601), .Y(n4210) );
  OAI21X1 U2147 ( .A(n335), .B(n1314), .C(n5598), .Y(n4211) );
  OAI21X1 U2149 ( .A(n337), .B(n1314), .C(n5595), .Y(n4212) );
  OAI21X1 U2151 ( .A(n339), .B(n1314), .C(n5592), .Y(n4213) );
  OAI21X1 U2153 ( .A(n341), .B(n1314), .C(n5589), .Y(n4214) );
  OAI21X1 U2155 ( .A(n343), .B(n1314), .C(n5586), .Y(n4215) );
  OAI21X1 U2157 ( .A(n345), .B(n1314), .C(n5583), .Y(n4216) );
  OAI21X1 U2159 ( .A(n347), .B(n1314), .C(n5580), .Y(n4217) );
  OAI21X1 U2161 ( .A(n349), .B(n1314), .C(n5577), .Y(n4218) );
  OAI21X1 U2163 ( .A(n351), .B(n1314), .C(n5574), .Y(n4219) );
  OAI21X1 U2165 ( .A(n353), .B(n1314), .C(n5571), .Y(n4220) );
  NAND3X1 U2169 ( .A(n253), .B(n256), .C(n13020), .Y(n1357) );
  INVX1 U2170 ( .A(n13011), .Y(n256) );
  OAI21X1 U2171 ( .A(n271), .B(n1358), .C(n5568), .Y(n4221) );
  OAI21X1 U2173 ( .A(n273), .B(n1358), .C(n5565), .Y(n4222) );
  OAI21X1 U2175 ( .A(n275), .B(n1358), .C(n5562), .Y(n4223) );
  OAI21X1 U2177 ( .A(n277), .B(n1358), .C(n5559), .Y(n4224) );
  OAI21X1 U2179 ( .A(n279), .B(n1358), .C(n5556), .Y(n4225) );
  OAI21X1 U2181 ( .A(n281), .B(n1358), .C(n5553), .Y(n4226) );
  OAI21X1 U2183 ( .A(n283), .B(n1358), .C(n5550), .Y(n4227) );
  OAI21X1 U2185 ( .A(n285), .B(n1358), .C(n5547), .Y(n4228) );
  OAI21X1 U2187 ( .A(n287), .B(n1358), .C(n5544), .Y(n4229) );
  OAI21X1 U2189 ( .A(n289), .B(n1358), .C(n5541), .Y(n4230) );
  OAI21X1 U2191 ( .A(n291), .B(n1358), .C(n5538), .Y(n4231) );
  OAI21X1 U2193 ( .A(n293), .B(n1358), .C(n5535), .Y(n4232) );
  OAI21X1 U2195 ( .A(n295), .B(n1358), .C(n5532), .Y(n4233) );
  OAI21X1 U2197 ( .A(n297), .B(n1358), .C(n5529), .Y(n4234) );
  OAI21X1 U2199 ( .A(n299), .B(n1358), .C(n5526), .Y(n4235) );
  OAI21X1 U2201 ( .A(n301), .B(n1358), .C(n5523), .Y(n4236) );
  OAI21X1 U2203 ( .A(n303), .B(n1358), .C(n5520), .Y(n4237) );
  OAI21X1 U2205 ( .A(n305), .B(n1358), .C(n5517), .Y(n4238) );
  OAI21X1 U2207 ( .A(n307), .B(n1358), .C(n5514), .Y(n4239) );
  OAI21X1 U2209 ( .A(n309), .B(n1358), .C(n5511), .Y(n4240) );
  OAI21X1 U2211 ( .A(n311), .B(n1358), .C(n5508), .Y(n4241) );
  OAI21X1 U2213 ( .A(n313), .B(n1358), .C(n5505), .Y(n4242) );
  OAI21X1 U2215 ( .A(n315), .B(n1358), .C(n5502), .Y(n4243) );
  OAI21X1 U2217 ( .A(n317), .B(n1358), .C(n5499), .Y(n4244) );
  OAI21X1 U2219 ( .A(n319), .B(n1358), .C(n5496), .Y(n4245) );
  OAI21X1 U2221 ( .A(n321), .B(n1358), .C(n5493), .Y(n4246) );
  OAI21X1 U2223 ( .A(n323), .B(n1358), .C(n5490), .Y(n4247) );
  OAI21X1 U2225 ( .A(n325), .B(n1358), .C(n5487), .Y(n4248) );
  OAI21X1 U2227 ( .A(n327), .B(n1358), .C(n5484), .Y(n4249) );
  OAI21X1 U2229 ( .A(n329), .B(n1358), .C(n5481), .Y(n4250) );
  OAI21X1 U2231 ( .A(n331), .B(n1358), .C(n5478), .Y(n4251) );
  OAI21X1 U2233 ( .A(n333), .B(n1358), .C(n5475), .Y(n4252) );
  OAI21X1 U2235 ( .A(n335), .B(n1358), .C(n5472), .Y(n4253) );
  OAI21X1 U2237 ( .A(n337), .B(n1358), .C(n5469), .Y(n4254) );
  OAI21X1 U2239 ( .A(n339), .B(n1358), .C(n5466), .Y(n4255) );
  OAI21X1 U2241 ( .A(n341), .B(n1358), .C(n5463), .Y(n4256) );
  OAI21X1 U2243 ( .A(n343), .B(n1358), .C(n5460), .Y(n4257) );
  OAI21X1 U2245 ( .A(n345), .B(n1358), .C(n5457), .Y(n4258) );
  OAI21X1 U2247 ( .A(n347), .B(n1358), .C(n5454), .Y(n4259) );
  OAI21X1 U2249 ( .A(n349), .B(n1358), .C(n5451), .Y(n4260) );
  OAI21X1 U2251 ( .A(n351), .B(n1358), .C(n5448), .Y(n4261) );
  OAI21X1 U2253 ( .A(n353), .B(n1358), .C(n5445), .Y(n4262) );
  NOR3X1 U2256 ( .A(n13015), .B(n68), .C(n13030), .Y(n355) );
  OAI21X1 U2257 ( .A(n271), .B(n1402), .C(n5442), .Y(n4263) );
  OAI21X1 U2259 ( .A(n273), .B(n1402), .C(n5439), .Y(n4264) );
  OAI21X1 U2261 ( .A(n275), .B(n1402), .C(n5436), .Y(n4265) );
  OAI21X1 U2263 ( .A(n277), .B(n1402), .C(n5433), .Y(n4266) );
  OAI21X1 U2265 ( .A(n279), .B(n1402), .C(n5430), .Y(n4267) );
  OAI21X1 U2267 ( .A(n281), .B(n1402), .C(n5427), .Y(n4268) );
  OAI21X1 U2269 ( .A(n283), .B(n1402), .C(n5424), .Y(n4269) );
  OAI21X1 U2271 ( .A(n285), .B(n1402), .C(n5421), .Y(n4270) );
  OAI21X1 U2273 ( .A(n287), .B(n1402), .C(n5418), .Y(n4271) );
  OAI21X1 U2275 ( .A(n289), .B(n1402), .C(n5415), .Y(n4272) );
  OAI21X1 U2277 ( .A(n291), .B(n1402), .C(n5412), .Y(n4273) );
  OAI21X1 U2279 ( .A(n293), .B(n1402), .C(n5409), .Y(n4274) );
  OAI21X1 U2281 ( .A(n295), .B(n1402), .C(n5406), .Y(n4275) );
  OAI21X1 U2283 ( .A(n297), .B(n1402), .C(n5403), .Y(n4276) );
  OAI21X1 U2285 ( .A(n299), .B(n1402), .C(n5400), .Y(n4277) );
  OAI21X1 U2287 ( .A(n301), .B(n1402), .C(n5397), .Y(n4278) );
  OAI21X1 U2289 ( .A(n303), .B(n1402), .C(n5394), .Y(n4279) );
  OAI21X1 U2291 ( .A(n305), .B(n1402), .C(n5391), .Y(n4280) );
  OAI21X1 U2293 ( .A(n307), .B(n1402), .C(n5388), .Y(n4281) );
  OAI21X1 U2295 ( .A(n309), .B(n1402), .C(n5385), .Y(n4282) );
  OAI21X1 U2297 ( .A(n311), .B(n1402), .C(n5382), .Y(n4283) );
  OAI21X1 U2299 ( .A(n313), .B(n1402), .C(n5379), .Y(n4284) );
  OAI21X1 U2301 ( .A(n315), .B(n1402), .C(n5376), .Y(n4285) );
  OAI21X1 U2303 ( .A(n317), .B(n1402), .C(n5373), .Y(n4286) );
  OAI21X1 U2305 ( .A(n319), .B(n1402), .C(n5370), .Y(n4287) );
  OAI21X1 U2307 ( .A(n321), .B(n1402), .C(n5367), .Y(n4288) );
  OAI21X1 U2309 ( .A(n323), .B(n1402), .C(n5364), .Y(n4289) );
  OAI21X1 U2311 ( .A(n325), .B(n1402), .C(n5361), .Y(n4290) );
  OAI21X1 U2313 ( .A(n327), .B(n1402), .C(n5358), .Y(n4291) );
  OAI21X1 U2315 ( .A(n329), .B(n1402), .C(n5355), .Y(n4292) );
  OAI21X1 U2317 ( .A(n331), .B(n1402), .C(n5352), .Y(n4293) );
  OAI21X1 U2319 ( .A(n333), .B(n1402), .C(n5349), .Y(n4294) );
  OAI21X1 U2321 ( .A(n335), .B(n1402), .C(n5346), .Y(n4295) );
  OAI21X1 U2323 ( .A(n337), .B(n1402), .C(n5343), .Y(n4296) );
  OAI21X1 U2325 ( .A(n339), .B(n1402), .C(n5340), .Y(n4297) );
  OAI21X1 U2327 ( .A(n341), .B(n1402), .C(n5337), .Y(n4298) );
  OAI21X1 U2329 ( .A(n343), .B(n1402), .C(n5334), .Y(n4299) );
  OAI21X1 U2331 ( .A(n345), .B(n1402), .C(n5331), .Y(n4300) );
  OAI21X1 U2333 ( .A(n347), .B(n1402), .C(n5328), .Y(n4301) );
  OAI21X1 U2335 ( .A(n349), .B(n1402), .C(n5325), .Y(n4302) );
  OAI21X1 U2337 ( .A(n351), .B(n1402), .C(n5322), .Y(n4303) );
  OAI21X1 U2339 ( .A(n353), .B(n1402), .C(n5319), .Y(n4304) );
  NOR3X1 U2342 ( .A(n13015), .B(n68), .C(n262), .Y(n400) );
  OAI21X1 U2343 ( .A(n271), .B(n1445), .C(n5316), .Y(n4305) );
  OAI21X1 U2345 ( .A(n273), .B(n1445), .C(n5313), .Y(n4306) );
  OAI21X1 U2347 ( .A(n275), .B(n1445), .C(n5310), .Y(n4307) );
  OAI21X1 U2349 ( .A(n277), .B(n1445), .C(n5307), .Y(n4308) );
  OAI21X1 U2351 ( .A(n279), .B(n1445), .C(n5304), .Y(n4309) );
  OAI21X1 U2353 ( .A(n281), .B(n1445), .C(n5301), .Y(n4310) );
  OAI21X1 U2355 ( .A(n283), .B(n1445), .C(n5298), .Y(n4311) );
  OAI21X1 U2357 ( .A(n285), .B(n1445), .C(n5295), .Y(n4312) );
  OAI21X1 U2359 ( .A(n287), .B(n1445), .C(n5292), .Y(n4313) );
  OAI21X1 U2361 ( .A(n289), .B(n1445), .C(n5289), .Y(n4314) );
  OAI21X1 U2363 ( .A(n291), .B(n1445), .C(n5286), .Y(n4315) );
  OAI21X1 U2365 ( .A(n293), .B(n1445), .C(n5283), .Y(n4316) );
  OAI21X1 U2367 ( .A(n295), .B(n1445), .C(n5280), .Y(n4317) );
  OAI21X1 U2369 ( .A(n297), .B(n1445), .C(n5277), .Y(n4318) );
  OAI21X1 U2371 ( .A(n299), .B(n1445), .C(n5274), .Y(n4319) );
  OAI21X1 U2373 ( .A(n301), .B(n1445), .C(n5271), .Y(n4320) );
  OAI21X1 U2375 ( .A(n303), .B(n1445), .C(n5268), .Y(n4321) );
  OAI21X1 U2377 ( .A(n305), .B(n1445), .C(n5265), .Y(n4322) );
  OAI21X1 U2379 ( .A(n307), .B(n1445), .C(n5262), .Y(n4323) );
  OAI21X1 U2381 ( .A(n309), .B(n1445), .C(n5259), .Y(n4324) );
  OAI21X1 U2383 ( .A(n311), .B(n1445), .C(n5256), .Y(n4325) );
  OAI21X1 U2385 ( .A(n313), .B(n1445), .C(n5253), .Y(n4326) );
  OAI21X1 U2387 ( .A(n315), .B(n1445), .C(n5250), .Y(n4327) );
  OAI21X1 U2389 ( .A(n317), .B(n1445), .C(n5247), .Y(n4328) );
  OAI21X1 U2391 ( .A(n319), .B(n1445), .C(n5244), .Y(n4329) );
  OAI21X1 U2393 ( .A(n321), .B(n1445), .C(n5241), .Y(n4330) );
  OAI21X1 U2395 ( .A(n323), .B(n1445), .C(n5238), .Y(n4331) );
  OAI21X1 U2397 ( .A(n325), .B(n1445), .C(n5235), .Y(n4332) );
  OAI21X1 U2399 ( .A(n327), .B(n1445), .C(n5232), .Y(n4333) );
  OAI21X1 U2401 ( .A(n329), .B(n1445), .C(n5229), .Y(n4334) );
  OAI21X1 U2403 ( .A(n331), .B(n1445), .C(n5226), .Y(n4335) );
  OAI21X1 U2405 ( .A(n333), .B(n1445), .C(n5223), .Y(n4336) );
  OAI21X1 U2407 ( .A(n335), .B(n1445), .C(n5220), .Y(n4337) );
  OAI21X1 U2409 ( .A(n337), .B(n1445), .C(n5217), .Y(n4338) );
  OAI21X1 U2411 ( .A(n339), .B(n1445), .C(n5214), .Y(n4339) );
  OAI21X1 U2413 ( .A(n341), .B(n1445), .C(n5211), .Y(n4340) );
  OAI21X1 U2415 ( .A(n343), .B(n1445), .C(n5208), .Y(n4341) );
  OAI21X1 U2417 ( .A(n345), .B(n1445), .C(n5205), .Y(n4342) );
  OAI21X1 U2419 ( .A(n347), .B(n1445), .C(n5202), .Y(n4343) );
  OAI21X1 U2421 ( .A(n349), .B(n1445), .C(n5199), .Y(n4344) );
  OAI21X1 U2423 ( .A(n351), .B(n1445), .C(n5196), .Y(n4345) );
  OAI21X1 U2425 ( .A(n353), .B(n1445), .C(n5193), .Y(n4346) );
  OAI21X1 U2429 ( .A(n271), .B(n1489), .C(n5190), .Y(n4347) );
  OAI21X1 U2431 ( .A(n273), .B(n1489), .C(n5187), .Y(n4348) );
  OAI21X1 U2433 ( .A(n275), .B(n1489), .C(n5184), .Y(n4349) );
  OAI21X1 U2435 ( .A(n277), .B(n1489), .C(n5181), .Y(n4350) );
  OAI21X1 U2437 ( .A(n279), .B(n1489), .C(n5178), .Y(n4351) );
  OAI21X1 U2439 ( .A(n281), .B(n1489), .C(n5175), .Y(n4352) );
  OAI21X1 U2441 ( .A(n283), .B(n1489), .C(n5172), .Y(n4353) );
  OAI21X1 U2443 ( .A(n285), .B(n1489), .C(n5169), .Y(n4354) );
  OAI21X1 U2445 ( .A(n287), .B(n1489), .C(n5166), .Y(n4355) );
  OAI21X1 U2447 ( .A(n289), .B(n1489), .C(n5163), .Y(n4356) );
  OAI21X1 U2449 ( .A(n291), .B(n1489), .C(n5160), .Y(n4357) );
  OAI21X1 U2451 ( .A(n293), .B(n1489), .C(n5157), .Y(n4358) );
  OAI21X1 U2453 ( .A(n295), .B(n1489), .C(n5154), .Y(n4359) );
  OAI21X1 U2455 ( .A(n297), .B(n1489), .C(n5151), .Y(n4360) );
  OAI21X1 U2457 ( .A(n299), .B(n1489), .C(n5148), .Y(n4361) );
  OAI21X1 U2459 ( .A(n301), .B(n1489), .C(n5145), .Y(n4362) );
  OAI21X1 U2461 ( .A(n303), .B(n1489), .C(n5142), .Y(n4363) );
  OAI21X1 U2463 ( .A(n305), .B(n1489), .C(n5139), .Y(n4364) );
  OAI21X1 U2465 ( .A(n307), .B(n1489), .C(n5136), .Y(n4365) );
  OAI21X1 U2467 ( .A(n309), .B(n1489), .C(n5133), .Y(n4366) );
  OAI21X1 U2469 ( .A(n311), .B(n1489), .C(n5130), .Y(n4367) );
  OAI21X1 U2471 ( .A(n313), .B(n1489), .C(n5127), .Y(n4368) );
  OAI21X1 U2473 ( .A(n315), .B(n1489), .C(n5124), .Y(n4369) );
  OAI21X1 U2475 ( .A(n317), .B(n1489), .C(n5121), .Y(n4370) );
  OAI21X1 U2477 ( .A(n319), .B(n1489), .C(n5118), .Y(n4371) );
  OAI21X1 U2479 ( .A(n321), .B(n1489), .C(n5115), .Y(n4372) );
  OAI21X1 U2481 ( .A(n323), .B(n1489), .C(n5112), .Y(n4373) );
  OAI21X1 U2483 ( .A(n325), .B(n1489), .C(n5109), .Y(n4374) );
  OAI21X1 U2485 ( .A(n327), .B(n1489), .C(n5106), .Y(n4375) );
  OAI21X1 U2487 ( .A(n329), .B(n1489), .C(n5103), .Y(n4376) );
  OAI21X1 U2489 ( .A(n331), .B(n1489), .C(n5100), .Y(n4377) );
  OAI21X1 U2491 ( .A(n333), .B(n1489), .C(n5097), .Y(n4378) );
  OAI21X1 U2493 ( .A(n335), .B(n1489), .C(n5094), .Y(n4379) );
  OAI21X1 U2495 ( .A(n337), .B(n1489), .C(n5091), .Y(n4380) );
  OAI21X1 U2497 ( .A(n339), .B(n1489), .C(n5088), .Y(n4381) );
  OAI21X1 U2499 ( .A(n341), .B(n1489), .C(n5085), .Y(n4382) );
  OAI21X1 U2501 ( .A(n343), .B(n1489), .C(n5082), .Y(n4383) );
  OAI21X1 U2503 ( .A(n345), .B(n1489), .C(n5079), .Y(n4384) );
  OAI21X1 U2505 ( .A(n347), .B(n1489), .C(n5076), .Y(n4385) );
  OAI21X1 U2507 ( .A(n349), .B(n1489), .C(n5073), .Y(n4386) );
  OAI21X1 U2509 ( .A(n351), .B(n1489), .C(n5070), .Y(n4387) );
  OAI21X1 U2511 ( .A(n353), .B(n1489), .C(n5067), .Y(n4388) );
  OAI21X1 U2515 ( .A(n271), .B(n13032), .C(n5064), .Y(n4389) );
  OAI21X1 U2517 ( .A(n273), .B(n13045), .C(n5061), .Y(n4390) );
  OAI21X1 U2519 ( .A(n275), .B(n12949), .C(n5058), .Y(n4391) );
  OAI21X1 U2521 ( .A(n277), .B(n13045), .C(n5055), .Y(n4392) );
  OAI21X1 U2523 ( .A(n279), .B(n12992), .C(n5052), .Y(n4393) );
  OAI21X1 U2525 ( .A(n281), .B(n13045), .C(n5049), .Y(n4394) );
  OAI21X1 U2527 ( .A(n283), .B(n13032), .C(n5046), .Y(n4395) );
  OAI21X1 U2529 ( .A(n285), .B(n13045), .C(n5043), .Y(n4396) );
  OAI21X1 U2531 ( .A(n287), .B(n12990), .C(n5040), .Y(n4397) );
  OAI21X1 U2533 ( .A(n289), .B(n13045), .C(n5037), .Y(n4398) );
  OAI21X1 U2535 ( .A(n291), .B(n8686), .C(n5034), .Y(n4399) );
  OAI21X1 U2537 ( .A(n293), .B(n13045), .C(n5031), .Y(n4400) );
  OAI21X1 U2539 ( .A(n295), .B(n13032), .C(n5028), .Y(n4401) );
  OAI21X1 U2541 ( .A(n297), .B(n13045), .C(n5025), .Y(n4402) );
  OAI21X1 U2543 ( .A(n299), .B(n12969), .C(n5022), .Y(n4403) );
  OAI21X1 U2545 ( .A(n301), .B(n13045), .C(n5019), .Y(n4404) );
  OAI21X1 U2547 ( .A(n303), .B(n12949), .C(n5016), .Y(n4405) );
  OAI21X1 U2549 ( .A(n305), .B(n13045), .C(n5013), .Y(n4406) );
  OAI21X1 U2551 ( .A(n307), .B(n13032), .C(n5010), .Y(n4407) );
  OAI21X1 U2553 ( .A(n309), .B(n13045), .C(n5007), .Y(n4408) );
  OAI21X1 U2555 ( .A(n311), .B(n12992), .C(n5004), .Y(n4409) );
  OAI21X1 U2557 ( .A(n313), .B(n13045), .C(n5001), .Y(n4410) );
  OAI21X1 U2559 ( .A(n315), .B(n12990), .C(n4998), .Y(n4411) );
  OAI21X1 U2561 ( .A(n317), .B(n13045), .C(n4995), .Y(n4412) );
  OAI21X1 U2563 ( .A(n319), .B(n13032), .C(n4992), .Y(n4413) );
  OAI21X1 U2565 ( .A(n321), .B(n13045), .C(n4989), .Y(n4414) );
  OAI21X1 U2567 ( .A(n323), .B(n12992), .C(n4986), .Y(n4415) );
  OAI21X1 U2569 ( .A(n325), .B(n13045), .C(n4983), .Y(n4416) );
  OAI21X1 U2571 ( .A(n327), .B(n10796), .C(n4980), .Y(n4417) );
  OAI21X1 U2573 ( .A(n329), .B(n13045), .C(n4977), .Y(n4418) );
  OAI21X1 U2575 ( .A(n331), .B(n13032), .C(n4974), .Y(n4419) );
  OAI21X1 U2577 ( .A(n333), .B(n13045), .C(n4971), .Y(n4420) );
  OAI21X1 U2579 ( .A(n335), .B(n8714), .C(n4968), .Y(n4421) );
  OAI21X1 U2581 ( .A(n337), .B(n13045), .C(n4965), .Y(n4422) );
  OAI21X1 U2583 ( .A(n339), .B(n12967), .C(n4962), .Y(n4423) );
  OAI21X1 U2585 ( .A(n341), .B(n13045), .C(n4959), .Y(n4424) );
  OAI21X1 U2587 ( .A(n343), .B(n13032), .C(n4956), .Y(n4425) );
  OAI21X1 U2589 ( .A(n345), .B(n13045), .C(n4953), .Y(n4426) );
  OAI21X1 U2591 ( .A(n347), .B(n8706), .C(n4950), .Y(n4427) );
  OAI21X1 U2593 ( .A(n349), .B(n13045), .C(n4947), .Y(n4428) );
  OAI21X1 U2595 ( .A(n351), .B(n12990), .C(n4944), .Y(n4429) );
  OAI21X1 U2597 ( .A(n353), .B(n13045), .C(n4941), .Y(n4430) );
  OAI21X1 U2601 ( .A(n271), .B(n1576), .C(n4938), .Y(n4431) );
  OAI21X1 U2603 ( .A(n273), .B(n1576), .C(n4935), .Y(n4432) );
  OAI21X1 U2605 ( .A(n275), .B(n1576), .C(n4932), .Y(n4433) );
  OAI21X1 U2607 ( .A(n277), .B(n1576), .C(n4929), .Y(n4434) );
  OAI21X1 U2609 ( .A(n279), .B(n1576), .C(n4926), .Y(n4435) );
  OAI21X1 U2611 ( .A(n281), .B(n1576), .C(n4923), .Y(n4436) );
  OAI21X1 U2613 ( .A(n283), .B(n1576), .C(n4920), .Y(n4437) );
  OAI21X1 U2615 ( .A(n285), .B(n1576), .C(n4917), .Y(n4438) );
  OAI21X1 U2617 ( .A(n287), .B(n1576), .C(n4914), .Y(n4439) );
  OAI21X1 U2619 ( .A(n289), .B(n1576), .C(n4911), .Y(n4440) );
  OAI21X1 U2621 ( .A(n291), .B(n1576), .C(n4908), .Y(n4441) );
  OAI21X1 U2623 ( .A(n293), .B(n1576), .C(n4905), .Y(n4442) );
  OAI21X1 U2625 ( .A(n295), .B(n1576), .C(n4902), .Y(n4443) );
  OAI21X1 U2627 ( .A(n297), .B(n1576), .C(n4899), .Y(n4444) );
  OAI21X1 U2629 ( .A(n299), .B(n1576), .C(n4896), .Y(n4445) );
  OAI21X1 U2631 ( .A(n301), .B(n1576), .C(n4893), .Y(n4446) );
  OAI21X1 U2633 ( .A(n303), .B(n1576), .C(n4890), .Y(n4447) );
  OAI21X1 U2635 ( .A(n305), .B(n1576), .C(n4887), .Y(n4448) );
  OAI21X1 U2637 ( .A(n307), .B(n1576), .C(n4884), .Y(n4449) );
  OAI21X1 U2639 ( .A(n309), .B(n1576), .C(n4881), .Y(n4450) );
  OAI21X1 U2641 ( .A(n311), .B(n1576), .C(n4878), .Y(n4451) );
  OAI21X1 U2643 ( .A(n313), .B(n1576), .C(n4875), .Y(n4452) );
  OAI21X1 U2645 ( .A(n315), .B(n1576), .C(n4872), .Y(n4453) );
  OAI21X1 U2647 ( .A(n317), .B(n1576), .C(n4869), .Y(n4454) );
  OAI21X1 U2649 ( .A(n319), .B(n1576), .C(n4866), .Y(n4455) );
  OAI21X1 U2651 ( .A(n321), .B(n1576), .C(n4863), .Y(n4456) );
  OAI21X1 U2653 ( .A(n323), .B(n1576), .C(n4860), .Y(n4457) );
  OAI21X1 U2655 ( .A(n325), .B(n1576), .C(n4857), .Y(n4458) );
  OAI21X1 U2657 ( .A(n327), .B(n1576), .C(n4854), .Y(n4459) );
  OAI21X1 U2659 ( .A(n329), .B(n1576), .C(n4851), .Y(n4460) );
  OAI21X1 U2661 ( .A(n331), .B(n1576), .C(n4848), .Y(n4461) );
  OAI21X1 U2663 ( .A(n333), .B(n1576), .C(n4845), .Y(n4462) );
  OAI21X1 U2665 ( .A(n335), .B(n1576), .C(n4842), .Y(n4463) );
  OAI21X1 U2667 ( .A(n337), .B(n1576), .C(n4839), .Y(n4464) );
  OAI21X1 U2669 ( .A(n339), .B(n1576), .C(n4836), .Y(n4465) );
  OAI21X1 U2671 ( .A(n341), .B(n1576), .C(n4833), .Y(n4466) );
  OAI21X1 U2673 ( .A(n343), .B(n1576), .C(n4830), .Y(n4467) );
  OAI21X1 U2675 ( .A(n345), .B(n1576), .C(n4827), .Y(n4468) );
  OAI21X1 U2677 ( .A(n347), .B(n1576), .C(n4824), .Y(n4469) );
  OAI21X1 U2679 ( .A(n349), .B(n1576), .C(n4821), .Y(n4470) );
  OAI21X1 U2681 ( .A(n351), .B(n1576), .C(n4818), .Y(n4471) );
  OAI21X1 U2683 ( .A(n353), .B(n1576), .C(n4815), .Y(n4472) );
  OAI21X1 U2687 ( .A(n271), .B(n1619), .C(n4812), .Y(n4473) );
  OAI21X1 U2689 ( .A(n273), .B(n1619), .C(n4809), .Y(n4474) );
  OAI21X1 U2691 ( .A(n275), .B(n1619), .C(n4806), .Y(n4475) );
  OAI21X1 U2693 ( .A(n277), .B(n1619), .C(n4803), .Y(n4476) );
  OAI21X1 U2695 ( .A(n279), .B(n1619), .C(n4800), .Y(n4477) );
  OAI21X1 U2697 ( .A(n281), .B(n1619), .C(n4797), .Y(n4478) );
  OAI21X1 U2699 ( .A(n283), .B(n1619), .C(n4794), .Y(n4479) );
  OAI21X1 U2701 ( .A(n285), .B(n1619), .C(n4791), .Y(n4480) );
  OAI21X1 U2703 ( .A(n287), .B(n1619), .C(n4788), .Y(n4481) );
  OAI21X1 U2705 ( .A(n289), .B(n1619), .C(n4785), .Y(n4482) );
  OAI21X1 U2707 ( .A(n291), .B(n1619), .C(n4782), .Y(n4483) );
  OAI21X1 U2709 ( .A(n293), .B(n1619), .C(n4779), .Y(n4484) );
  OAI21X1 U2711 ( .A(n295), .B(n1619), .C(n4776), .Y(n4485) );
  OAI21X1 U2713 ( .A(n297), .B(n1619), .C(n4773), .Y(n4486) );
  OAI21X1 U2715 ( .A(n299), .B(n1619), .C(n4770), .Y(n4487) );
  OAI21X1 U2717 ( .A(n301), .B(n1619), .C(n4767), .Y(n4488) );
  OAI21X1 U2719 ( .A(n303), .B(n1619), .C(n4764), .Y(n4489) );
  OAI21X1 U2721 ( .A(n305), .B(n1619), .C(n4761), .Y(n4490) );
  OAI21X1 U2723 ( .A(n307), .B(n1619), .C(n4758), .Y(n4491) );
  OAI21X1 U2725 ( .A(n309), .B(n1619), .C(n4755), .Y(n4492) );
  OAI21X1 U2727 ( .A(n311), .B(n1619), .C(n4752), .Y(n4493) );
  OAI21X1 U2729 ( .A(n313), .B(n1619), .C(n4749), .Y(n4494) );
  OAI21X1 U2731 ( .A(n315), .B(n1619), .C(n4746), .Y(n4495) );
  OAI21X1 U2733 ( .A(n317), .B(n1619), .C(n4743), .Y(n4496) );
  OAI21X1 U2735 ( .A(n319), .B(n1619), .C(n4740), .Y(n4497) );
  OAI21X1 U2737 ( .A(n321), .B(n1619), .C(n4737), .Y(n4498) );
  OAI21X1 U2739 ( .A(n323), .B(n1619), .C(n4734), .Y(n4499) );
  OAI21X1 U2741 ( .A(n325), .B(n1619), .C(n4731), .Y(n4500) );
  OAI21X1 U2743 ( .A(n327), .B(n1619), .C(n4728), .Y(n4501) );
  OAI21X1 U2745 ( .A(n329), .B(n1619), .C(n4725), .Y(n4502) );
  OAI21X1 U2747 ( .A(n331), .B(n1619), .C(n4722), .Y(n4503) );
  OAI21X1 U2749 ( .A(n333), .B(n1619), .C(n4719), .Y(n4504) );
  OAI21X1 U2751 ( .A(n335), .B(n1619), .C(n4716), .Y(n4505) );
  OAI21X1 U2753 ( .A(n337), .B(n1619), .C(n4713), .Y(n4506) );
  OAI21X1 U2755 ( .A(n339), .B(n1619), .C(n4710), .Y(n4507) );
  OAI21X1 U2757 ( .A(n341), .B(n1619), .C(n4707), .Y(n4508) );
  OAI21X1 U2759 ( .A(n343), .B(n1619), .C(n4704), .Y(n4509) );
  OAI21X1 U2761 ( .A(n345), .B(n1619), .C(n4701), .Y(n4510) );
  OAI21X1 U2763 ( .A(n347), .B(n1619), .C(n4698), .Y(n4511) );
  OAI21X1 U2765 ( .A(n349), .B(n1619), .C(n4695), .Y(n4512) );
  OAI21X1 U2767 ( .A(n351), .B(n1619), .C(n4692), .Y(n4513) );
  OAI21X1 U2769 ( .A(n353), .B(n1619), .C(n4689), .Y(n4514) );
  NOR3X1 U2772 ( .A(n258), .B(n13030), .C(n260), .Y(n620) );
  OAI21X1 U2773 ( .A(n271), .B(n1662), .C(n4686), .Y(n4515) );
  INVX1 U2775 ( .A(data_in[41]), .Y(n271) );
  OAI21X1 U2776 ( .A(n273), .B(n1662), .C(n4683), .Y(n4516) );
  INVX1 U2778 ( .A(data_in[40]), .Y(n273) );
  OAI21X1 U2779 ( .A(n275), .B(n1662), .C(n4680), .Y(n4517) );
  INVX1 U2781 ( .A(data_in[39]), .Y(n275) );
  OAI21X1 U2782 ( .A(n277), .B(n1662), .C(n4677), .Y(n4518) );
  INVX1 U2784 ( .A(data_in[38]), .Y(n277) );
  OAI21X1 U2785 ( .A(n279), .B(n1662), .C(n4674), .Y(n4519) );
  INVX1 U2787 ( .A(data_in[37]), .Y(n279) );
  OAI21X1 U2788 ( .A(n281), .B(n1662), .C(n4671), .Y(n4520) );
  INVX1 U2790 ( .A(data_in[36]), .Y(n281) );
  OAI21X1 U2791 ( .A(n283), .B(n1662), .C(n4668), .Y(n4521) );
  INVX1 U2793 ( .A(data_in[35]), .Y(n283) );
  OAI21X1 U2794 ( .A(n285), .B(n1662), .C(n4665), .Y(n4522) );
  INVX1 U2796 ( .A(data_in[34]), .Y(n285) );
  OAI21X1 U2797 ( .A(n287), .B(n1662), .C(n4662), .Y(n4523) );
  INVX1 U2799 ( .A(data_in[33]), .Y(n287) );
  OAI21X1 U2800 ( .A(n289), .B(n1662), .C(n4659), .Y(n4524) );
  INVX1 U2802 ( .A(data_in[32]), .Y(n289) );
  OAI21X1 U2803 ( .A(n291), .B(n1662), .C(n4656), .Y(n4525) );
  INVX1 U2805 ( .A(data_in[31]), .Y(n291) );
  OAI21X1 U2806 ( .A(n293), .B(n1662), .C(n4653), .Y(n4526) );
  INVX1 U2808 ( .A(data_in[30]), .Y(n293) );
  OAI21X1 U2809 ( .A(n295), .B(n1662), .C(n4650), .Y(n4527) );
  INVX1 U2811 ( .A(data_in[29]), .Y(n295) );
  OAI21X1 U2812 ( .A(n297), .B(n1662), .C(n4647), .Y(n4528) );
  INVX1 U2814 ( .A(data_in[28]), .Y(n297) );
  OAI21X1 U2815 ( .A(n299), .B(n1662), .C(n4644), .Y(n4529) );
  INVX1 U2817 ( .A(data_in[27]), .Y(n299) );
  OAI21X1 U2818 ( .A(n301), .B(n1662), .C(n4641), .Y(n4530) );
  INVX1 U2820 ( .A(data_in[26]), .Y(n301) );
  OAI21X1 U2821 ( .A(n303), .B(n1662), .C(n4638), .Y(n4531) );
  INVX1 U2823 ( .A(data_in[25]), .Y(n303) );
  OAI21X1 U2824 ( .A(n305), .B(n1662), .C(n4635), .Y(n4532) );
  INVX1 U2826 ( .A(data_in[24]), .Y(n305) );
  OAI21X1 U2827 ( .A(n307), .B(n1662), .C(n4632), .Y(n4533) );
  INVX1 U2829 ( .A(data_in[23]), .Y(n307) );
  OAI21X1 U2830 ( .A(n309), .B(n1662), .C(n4629), .Y(n4534) );
  INVX1 U2832 ( .A(data_in[22]), .Y(n309) );
  OAI21X1 U2833 ( .A(n311), .B(n1662), .C(n4626), .Y(n4535) );
  INVX1 U2835 ( .A(data_in[21]), .Y(n311) );
  OAI21X1 U2836 ( .A(n313), .B(n1662), .C(n4623), .Y(n4536) );
  INVX1 U2838 ( .A(data_in[20]), .Y(n313) );
  OAI21X1 U2839 ( .A(n315), .B(n1662), .C(n4620), .Y(n4537) );
  INVX1 U2841 ( .A(data_in[19]), .Y(n315) );
  OAI21X1 U2842 ( .A(n317), .B(n1662), .C(n4617), .Y(n4538) );
  INVX1 U2844 ( .A(data_in[18]), .Y(n317) );
  OAI21X1 U2845 ( .A(n319), .B(n1662), .C(n4614), .Y(n4539) );
  INVX1 U2847 ( .A(data_in[17]), .Y(n319) );
  OAI21X1 U2848 ( .A(n321), .B(n1662), .C(n4611), .Y(n4540) );
  INVX1 U2850 ( .A(data_in[16]), .Y(n321) );
  OAI21X1 U2851 ( .A(n323), .B(n1662), .C(n4608), .Y(n4541) );
  INVX1 U2853 ( .A(data_in[15]), .Y(n323) );
  OAI21X1 U2854 ( .A(n325), .B(n1662), .C(n4605), .Y(n4542) );
  INVX1 U2856 ( .A(data_in[14]), .Y(n325) );
  OAI21X1 U2857 ( .A(n327), .B(n1662), .C(n4602), .Y(n4543) );
  INVX1 U2859 ( .A(data_in[13]), .Y(n327) );
  OAI21X1 U2860 ( .A(n329), .B(n1662), .C(n4599), .Y(n4544) );
  INVX1 U2862 ( .A(data_in[12]), .Y(n329) );
  OAI21X1 U2863 ( .A(n331), .B(n1662), .C(n4596), .Y(n4545) );
  INVX1 U2865 ( .A(data_in[11]), .Y(n331) );
  OAI21X1 U2866 ( .A(n333), .B(n1662), .C(n4593), .Y(n4546) );
  INVX1 U2868 ( .A(data_in[10]), .Y(n333) );
  OAI21X1 U2869 ( .A(n335), .B(n1662), .C(n4590), .Y(n4547) );
  INVX1 U2871 ( .A(data_in[9]), .Y(n335) );
  OAI21X1 U2872 ( .A(n337), .B(n1662), .C(n4587), .Y(n4548) );
  INVX1 U2874 ( .A(data_in[8]), .Y(n337) );
  OAI21X1 U2875 ( .A(n339), .B(n1662), .C(n4584), .Y(n4549) );
  INVX1 U2877 ( .A(data_in[7]), .Y(n339) );
  OAI21X1 U2878 ( .A(n341), .B(n1662), .C(n4581), .Y(n4550) );
  INVX1 U2880 ( .A(data_in[6]), .Y(n341) );
  OAI21X1 U2881 ( .A(n343), .B(n1662), .C(n4578), .Y(n4551) );
  INVX1 U2883 ( .A(data_in[5]), .Y(n343) );
  OAI21X1 U2884 ( .A(n345), .B(n1662), .C(n4575), .Y(n4552) );
  INVX1 U2886 ( .A(data_in[4]), .Y(n345) );
  OAI21X1 U2887 ( .A(n347), .B(n1662), .C(n4572), .Y(n4553) );
  INVX1 U2889 ( .A(data_in[3]), .Y(n347) );
  OAI21X1 U2890 ( .A(n349), .B(n1662), .C(n4569), .Y(n4554) );
  INVX1 U2892 ( .A(data_in[2]), .Y(n349) );
  OAI21X1 U2893 ( .A(n351), .B(n1662), .C(n4566), .Y(n4555) );
  INVX1 U2895 ( .A(data_in[1]), .Y(n351) );
  OAI21X1 U2896 ( .A(n353), .B(n1662), .C(n4563), .Y(n4556) );
  NOR3X1 U2899 ( .A(n260), .B(n258), .C(n262), .Y(n664) );
  INVX1 U2900 ( .A(n13029), .Y(n262) );
  NAND3X1 U2902 ( .A(n13022), .B(n253), .C(n13011), .Y(n1705) );
  INVX1 U2904 ( .A(data_in[0]), .Y(n353) );
  XOR2X1 U2905 ( .A(n13016), .B(n13029), .Y(n24) );
  INVX1 U2908 ( .A(n68), .Y(n258) );
  INVX1 U2910 ( .A(n13015), .Y(n260) );
  XOR2X1 U2911 ( .A(n13011), .B(n68), .Y(n22) );
  XOR2X1 U2912 ( .A(n13019), .B(n13011), .Y(n21) );
  XOR2X1 U2913 ( .A(n12995), .B(n13022), .Y(n20) );
  XOR2X1 U2914 ( .A(n13283), .B(n13316), .Y(n19) );
  XOR2X1 U2915 ( .A(n13265), .B(n13283), .Y(n18) );
  XOR2X1 U2916 ( .A(n13104), .B(n13265), .Y(n17) );
  XOR2X1 U2917 ( .A(n13101), .B(n13104), .Y(n16) );
  XOR2X1 U2918 ( .A(n12981), .B(n13101), .Y(n15) );
  NAND3X1 U2922 ( .A(n193), .B(n1709), .C(n8731), .Y(n14681) );
  XOR2X1 U2924 ( .A(n13100), .B(n1713), .Y(n1712) );
  XOR2X1 U2925 ( .A(n13103), .B(n1714), .Y(n1711) );
  XOR2X1 U2926 ( .A(n266), .B(n12964), .Y(n1709) );
  INVX1 U2927 ( .A(n12981), .Y(n266) );
  AOI22X1 U2928 ( .A(n1715), .B(n199), .C(n1717), .D(n8726), .Y(n1708) );
  NAND3X1 U2929 ( .A(n1719), .B(n13277), .C(n1720), .Y(n1718) );
  XOR2X1 U2930 ( .A(n13369), .B(n1721), .Y(n1720) );
  XOR2X1 U2933 ( .A(n12978), .B(n13311), .Y(n1719) );
  NAND3X1 U2935 ( .A(n1722), .B(n1723), .C(n13275), .Y(n1716) );
  XOR2X1 U2936 ( .A(n12978), .B(n13283), .Y(n1723) );
  XOR2X1 U2937 ( .A(n13316), .B(n1721), .Y(n1722) );
  XOR2X1 U2938 ( .A(n12978), .B(n8743), .Y(n1721) );
  INVX1 U2939 ( .A(n1717), .Y(n1715) );
  XNOR2X1 U2940 ( .A(n1714), .B(n8734), .Y(n1717) );
  XOR2X1 U2941 ( .A(n1713), .B(n8740), .Y(n1714) );
  XOR2X1 U2942 ( .A(n12964), .B(n8737), .Y(n1713) );
  HAX1 add_176_U1_1_1 ( .A(n13283), .B(n13355), .YC(add_176_carry[2]), .YS(
        n114) );
  HAX1 add_176_U1_1_2 ( .A(n13265), .B(add_176_carry[2]), .YC(add_176_carry[3]), .YS(n115) );
  HAX1 add_176_U1_1_3 ( .A(n13104), .B(add_176_carry[3]), .YC(add_176_carry[4]), .YS(n116) );
  HAX1 add_176_U1_1_4 ( .A(n13101), .B(add_176_carry[4]), .YC(add_176_carry[5]), .YS(n117) );
  HAX1 add_158_U1_1_1 ( .A(n13016), .B(n13029), .YC(add_158_carry[2]), .YS(n34) );
  HAX1 add_158_U1_1_2 ( .A(n68), .B(add_158_carry[2]), .YC(add_158_carry[3]), 
        .YS(n35) );
  HAX1 add_158_U1_1_3 ( .A(n13011), .B(add_158_carry[3]), .YC(add_158_carry[4]), .YS(n36) );
  HAX1 add_158_U1_1_4 ( .A(n13021), .B(add_158_carry[4]), .YC(add_158_carry[5]), .YS(n37) );
  INVX1 U3 ( .A(n3), .Y(n1) );
  XOR2X1 U4 ( .A(n13065), .B(net84863), .Y(fillcount[5]) );
  INVX1 U5 ( .A(r301_B_not_0_), .Y(n2) );
  AND2X2 U6 ( .A(net94574), .B(net91739), .Y(n3) );
  XNOR2X1 U7 ( .A(n32), .B(n206), .Y(net82274) );
  BUFX2 U8 ( .A(net92912), .Y(n4) );
  INVX1 U10 ( .A(net98087), .Y(net94543) );
  AND2X2 U13 ( .A(n2), .B(n30), .Y(n5) );
  INVX1 U16 ( .A(n5), .Y(net91678) );
  OAI21X1 U18 ( .A(n7), .B(net91760), .C(net94407), .Y(n6) );
  INVX1 U104 ( .A(n6), .Y(n13067) );
  INVX8 U106 ( .A(net91739), .Y(n7) );
  OAI21X1 U108 ( .A(net91678), .B(n9), .C(n13056), .Y(n8) );
  INVX1 U110 ( .A(n8), .Y(n13059) );
  INVX1 U112 ( .A(n60), .Y(n9) );
  INVX1 U114 ( .A(n13053), .Y(n25) );
  AND2X2 U117 ( .A(n51), .B(fillcount[5]), .Y(n26) );
  BUFX2 U120 ( .A(n13058), .Y(n27) );
  BUFX2 U122 ( .A(n12952), .Y(n28) );
  INVX1 U124 ( .A(n64), .Y(n29) );
  INVX4 U126 ( .A(net82457), .Y(net82062) );
  NOR3X1 U128 ( .A(net91712), .B(n8670), .C(n13028), .Y(n30) );
  XOR2X1 U130 ( .A(n67), .B(n12952), .Y(n31) );
  XNOR2X1 U132 ( .A(n31), .B(n13052), .Y(net98077) );
  XOR2X1 U134 ( .A(net98087), .B(n66), .Y(n32) );
  INVX1 U136 ( .A(n64), .Y(n13052) );
  OR2X2 U138 ( .A(n12976), .B(net94515), .Y(net94524) );
  INVX1 U140 ( .A(net94524), .Y(n33) );
  AND2X2 U142 ( .A(net94553), .B(n25), .Y(n8669) );
  AND2X2 U144 ( .A(net82147), .B(net82062), .Y(n12976) );
  INVX1 U146 ( .A(n12976), .Y(n39) );
  OR2X2 U148 ( .A(n52), .B(n13057), .Y(n13056) );
  AND2X2 U150 ( .A(net94541), .B(n13020), .Y(net94529) );
  INVX1 U152 ( .A(net94529), .Y(n40) );
  AND2X2 U154 ( .A(net82511), .B(net82512), .Y(net82513) );
  INVX1 U156 ( .A(net82513), .Y(n41) );
  AND2X2 U158 ( .A(n13059), .B(net84769), .Y(net82260) );
  INVX1 U160 ( .A(net82260), .Y(n42) );
  AND2X2 U162 ( .A(n32), .B(net84737), .Y(net84743) );
  INVX1 U164 ( .A(net84743), .Y(n43) );
  AND2X2 U166 ( .A(net82055), .B(net82056), .Y(n13097) );
  INVX1 U168 ( .A(n13097), .Y(n44) );
  BUFX2 U170 ( .A(n13064), .Y(n45) );
  AND2X2 U172 ( .A(net84770), .B(net82259), .Y(net82261) );
  INVX1 U174 ( .A(net82261), .Y(n46) );
  AND2X2 U176 ( .A(n13068), .B(net84855), .Y(n13098) );
  INVX1 U178 ( .A(n13098), .Y(n47) );
  BUFX2 U180 ( .A(n14681), .Y(empty_bar) );
  BUFX2 U182 ( .A(net84760), .Y(n49) );
  OR2X2 U184 ( .A(fillcount[4]), .B(net92930), .Y(net82166) );
  INVX1 U186 ( .A(net82166), .Y(n50) );
  OR2X2 U188 ( .A(fillcount[3]), .B(fillcount[2]), .Y(net80714) );
  INVX1 U190 ( .A(net80714), .Y(n51) );
  AND2X2 U192 ( .A(n62), .B(n13055), .Y(n13054) );
  INVX1 U194 ( .A(n13054), .Y(n52) );
  AND2X2 U196 ( .A(n46), .B(n42), .Y(full_check_4_) );
  INVX1 U198 ( .A(full_check_4_), .Y(fillcount[4]) );
  AND2X2 U200 ( .A(n47), .B(n44), .Y(full_check_3_) );
  INVX1 U202 ( .A(full_check_3_), .Y(fillcount[3]) );
  AND2X2 U204 ( .A(net91739), .B(n57), .Y(n13066) );
  INVX1 U206 ( .A(n13066), .Y(n55) );
  AND2X2 U207 ( .A(net94521), .B(n8669), .Y(n13063) );
  INVX1 U209 ( .A(n13063), .Y(n56) );
  AND2X2 U211 ( .A(net92912), .B(net84737), .Y(n13053) );
  INVX1 U213 ( .A(net84743), .Y(n57) );
  AND2X2 U215 ( .A(n26), .B(n50), .Y(n13058) );
  INVX1 U217 ( .A(n13058), .Y(full_bar) );
  INVX1 U219 ( .A(n27), .Y(n59) );
  AND2X2 U221 ( .A(net84771), .B(net91739), .Y(net91741) );
  INVX1 U223 ( .A(n3), .Y(n60) );
  INVX1 U225 ( .A(net91741), .Y(n61) );
  AND2X2 U227 ( .A(n43), .B(net91739), .Y(net91726) );
  INVX1 U229 ( .A(net91726), .Y(n62) );
  INVX1 U231 ( .A(net91726), .Y(n63) );
  AND2X2 U233 ( .A(n190), .B(n45), .Y(n13065) );
  BUFX2 U235 ( .A(rd_ptr_gray_ss[3]), .Y(n64) );
  BUFX2 U237 ( .A(rd_ptr_gray_ss[2]), .Y(n65) );
  BUFX2 U239 ( .A(rd_ptr_gray_ss[1]), .Y(n66) );
  BUFX2 U241 ( .A(rd_ptr_gray_ss[5]), .Y(n67) );
  BUFX2 U243 ( .A(wr_ptr_bin[2]), .Y(n68) );
  INVX1 U245 ( .A(n67), .Y(net95813) );
  INVX1 U247 ( .A(n12976), .Y(n69) );
  INVX1 U249 ( .A(n119), .Y(n70) );
  INVX1 U251 ( .A(n70), .Y(n113) );
  BUFX2 U253 ( .A(rd_ptr_gray_s[3]), .Y(n119) );
  INVX1 U255 ( .A(n122), .Y(n120) );
  INVX1 U257 ( .A(n120), .Y(n121) );
  BUFX2 U259 ( .A(rd_ptr_gray[3]), .Y(n122) );
  INVX1 U261 ( .A(n125), .Y(n123) );
  INVX1 U263 ( .A(n123), .Y(n124) );
  BUFX2 U265 ( .A(rd_ptr_gray_s[2]), .Y(n125) );
  INVX1 U267 ( .A(n128), .Y(n126) );
  INVX1 U269 ( .A(n126), .Y(n127) );
  BUFX2 U271 ( .A(rd_ptr_gray[2]), .Y(n128) );
  INVX1 U273 ( .A(n131), .Y(n129) );
  INVX1 U275 ( .A(n129), .Y(n130) );
  BUFX2 U277 ( .A(rd_ptr_gray_s[1]), .Y(n131) );
  INVX1 U279 ( .A(n134), .Y(n132) );
  INVX1 U281 ( .A(n132), .Y(n133) );
  BUFX2 U283 ( .A(rd_ptr_gray[1]), .Y(n134) );
  INVX1 U285 ( .A(n137), .Y(n135) );
  INVX1 U287 ( .A(n135), .Y(n136) );
  BUFX2 U289 ( .A(rd_ptr_gray_s[0]), .Y(n137) );
  INVX1 U291 ( .A(n140), .Y(n138) );
  INVX1 U292 ( .A(n138), .Y(n139) );
  BUFX2 U294 ( .A(rd_ptr_gray[0]), .Y(n140) );
  INVX1 U296 ( .A(n143), .Y(n141) );
  INVX1 U298 ( .A(n141), .Y(n142) );
  BUFX2 U300 ( .A(wr_ptr_gray_s[4]), .Y(n143) );
  INVX1 U302 ( .A(n146), .Y(n144) );
  INVX1 U304 ( .A(n144), .Y(n145) );
  BUFX2 U306 ( .A(wr_ptr_gray[4]), .Y(n146) );
  INVX1 U308 ( .A(n149), .Y(n147) );
  INVX1 U310 ( .A(n147), .Y(n148) );
  BUFX2 U312 ( .A(wr_ptr_gray_s[3]), .Y(n149) );
  INVX1 U314 ( .A(n152), .Y(n150) );
  INVX1 U316 ( .A(n150), .Y(n151) );
  BUFX2 U318 ( .A(wr_ptr_gray[3]), .Y(n152) );
  INVX1 U320 ( .A(n155), .Y(n153) );
  INVX1 U322 ( .A(n153), .Y(n154) );
  BUFX2 U324 ( .A(wr_ptr_gray_s[2]), .Y(n155) );
  INVX1 U326 ( .A(n158), .Y(n156) );
  INVX1 U328 ( .A(n156), .Y(n157) );
  BUFX2 U330 ( .A(wr_ptr_gray[2]), .Y(n158) );
  INVX1 U332 ( .A(n161), .Y(n159) );
  INVX1 U334 ( .A(n159), .Y(n160) );
  BUFX2 U336 ( .A(wr_ptr_gray_s[1]), .Y(n161) );
  INVX1 U338 ( .A(n164), .Y(n162) );
  INVX1 U340 ( .A(n162), .Y(n163) );
  BUFX2 U342 ( .A(wr_ptr_gray[1]), .Y(n164) );
  INVX1 U344 ( .A(n167), .Y(n165) );
  INVX1 U346 ( .A(n165), .Y(n166) );
  BUFX2 U348 ( .A(wr_ptr_gray_s[0]), .Y(n167) );
  INVX1 U350 ( .A(n170), .Y(n168) );
  INVX1 U352 ( .A(n168), .Y(n169) );
  BUFX2 U354 ( .A(wr_ptr_gray[0]), .Y(n170) );
  INVX1 U356 ( .A(n173), .Y(n171) );
  INVX1 U358 ( .A(n171), .Y(n172) );
  BUFX2 U360 ( .A(wr_ptr_gray_s[5]), .Y(n173) );
  INVX1 U362 ( .A(n176), .Y(n174) );
  INVX1 U364 ( .A(n174), .Y(n175) );
  BUFX2 U366 ( .A(wr_ptr_gray[5]), .Y(n176) );
  INVX1 U368 ( .A(n179), .Y(n177) );
  INVX1 U370 ( .A(n177), .Y(n178) );
  BUFX2 U372 ( .A(rd_ptr_gray_s[4]), .Y(n179) );
  INVX1 U374 ( .A(n182), .Y(n180) );
  INVX1 U376 ( .A(n180), .Y(n181) );
  BUFX2 U377 ( .A(rd_ptr_gray[4]), .Y(n182) );
  INVX1 U379 ( .A(n185), .Y(n183) );
  INVX1 U381 ( .A(n183), .Y(n184) );
  BUFX2 U383 ( .A(rd_ptr_gray_s[5]), .Y(n185) );
  INVX1 U385 ( .A(n188), .Y(n186) );
  INVX1 U387 ( .A(n186), .Y(n187) );
  BUFX2 U389 ( .A(rd_ptr_gray[5]), .Y(n188) );
  INVX1 U391 ( .A(n191), .Y(n189) );
  INVX1 U393 ( .A(n189), .Y(n190) );
  BUFX2 U395 ( .A(net94530), .Y(n191) );
  INVX1 U397 ( .A(n194), .Y(n192) );
  INVX1 U399 ( .A(n192), .Y(n193) );
  BUFX2 U401 ( .A(n1708), .Y(n194) );
  INVX1 U403 ( .A(n197), .Y(n195) );
  INVX1 U405 ( .A(n195), .Y(n196) );
  BUFX2 U407 ( .A(n33), .Y(n197) );
  INVX1 U409 ( .A(n200), .Y(n198) );
  INVX1 U411 ( .A(n198), .Y(n199) );
  BUFX2 U413 ( .A(n1716), .Y(n200) );
  INVX1 U415 ( .A(n208), .Y(n206) );
  BUFX2 U417 ( .A(rd_ptr_gray_ss[0]), .Y(n208) );
  INVX1 U419 ( .A(n57), .Y(net92910) );
  AND2X1 U421 ( .A(n1055), .B(n664), .Y(n13090) );
  AND2X1 U423 ( .A(n1055), .B(n620), .Y(n13088) );
  AND2X1 U425 ( .A(n1055), .B(n400), .Y(n13086) );
  AND2X1 U427 ( .A(n1055), .B(n12998), .Y(n13096) );
  AND2X1 U429 ( .A(n1055), .B(n13004), .Y(n13094) );
  AND2X1 U431 ( .A(n1055), .B(n13007), .Y(n13092) );
  AND2X1 U433 ( .A(n709), .B(n12998), .Y(n13095) );
  AND2X1 U435 ( .A(n709), .B(n13001), .Y(n13093) );
  AND2X1 U437 ( .A(n709), .B(n13007), .Y(n13091) );
  AND2X1 U439 ( .A(n709), .B(n664), .Y(n13089) );
  AND2X1 U441 ( .A(n709), .B(n620), .Y(n13087) );
  AND2X1 U443 ( .A(n709), .B(n400), .Y(n13085) );
  AND2X1 U445 ( .A(n12998), .B(n356), .Y(n13075) );
  AND2X1 U447 ( .A(n13001), .B(n356), .Y(n13074) );
  AND2X1 U449 ( .A(n13004), .B(n356), .Y(n13073) );
  AND2X1 U451 ( .A(n400), .B(n356), .Y(n13072) );
  AND2X1 U453 ( .A(n664), .B(n356), .Y(n13071) );
  AND2X1 U455 ( .A(n620), .B(n356), .Y(n13070) );
  AND2X1 U457 ( .A(n1055), .B(n13001), .Y(n8773) );
  INVX1 U459 ( .A(n8773), .Y(n268) );
  AND2X1 U461 ( .A(n709), .B(n13004), .Y(n8776) );
  INVX1 U462 ( .A(n8776), .Y(n796) );
  AND2X1 U464 ( .A(n1401), .B(n12998), .Y(n1532) );
  INVX1 U466 ( .A(n1532), .Y(n1228) );
  AND2X1 U468 ( .A(n13007), .B(n356), .Y(n401) );
  INVX1 U470 ( .A(n401), .Y(n1706) );
  INVX1 U472 ( .A(n4558), .Y(n1707) );
  INVX1 U474 ( .A(n1707), .Y(n4557) );
  AND2X1 U476 ( .A(n12958), .B(n12955), .Y(n23) );
  INVX1 U478 ( .A(n23), .Y(n4558) );
  INVX1 U480 ( .A(n4561), .Y(n4559) );
  INVX1 U482 ( .A(n4559), .Y(n4560) );
  AND2X1 U484 ( .A(n253), .B(net82004), .Y(n263) );
  INVX1 U486 ( .A(n263), .Y(n4561) );
  INVX1 U488 ( .A(n4564), .Y(n4562) );
  INVX1 U490 ( .A(n4562), .Y(n4563) );
  AND2X1 U492 ( .A(n10804), .B(n1662), .Y(n1704) );
  INVX1 U494 ( .A(n1704), .Y(n4564) );
  INVX1 U496 ( .A(n4567), .Y(n4565) );
  INVX1 U498 ( .A(n4565), .Y(n4566) );
  AND2X1 U500 ( .A(n10807), .B(n1662), .Y(n1703) );
  INVX1 U502 ( .A(n1703), .Y(n4567) );
  INVX1 U504 ( .A(n4570), .Y(n4568) );
  INVX1 U506 ( .A(n4568), .Y(n4569) );
  AND2X1 U508 ( .A(n10810), .B(n1662), .Y(n1702) );
  INVX1 U510 ( .A(n1702), .Y(n4570) );
  INVX1 U512 ( .A(n4573), .Y(n4571) );
  INVX1 U514 ( .A(n4571), .Y(n4572) );
  AND2X1 U516 ( .A(n10813), .B(n1662), .Y(n1701) );
  INVX1 U518 ( .A(n1701), .Y(n4573) );
  INVX1 U520 ( .A(n4576), .Y(n4574) );
  INVX1 U522 ( .A(n4574), .Y(n4575) );
  AND2X1 U524 ( .A(n10816), .B(n1662), .Y(n1700) );
  INVX1 U526 ( .A(n1700), .Y(n4576) );
  INVX1 U528 ( .A(n4579), .Y(n4577) );
  INVX1 U530 ( .A(n4577), .Y(n4578) );
  AND2X1 U532 ( .A(n10819), .B(n1662), .Y(n1699) );
  INVX1 U534 ( .A(n1699), .Y(n4579) );
  INVX1 U536 ( .A(n4582), .Y(n4580) );
  INVX1 U538 ( .A(n4580), .Y(n4581) );
  AND2X1 U540 ( .A(n10822), .B(n1662), .Y(n1698) );
  INVX1 U542 ( .A(n1698), .Y(n4582) );
  INVX1 U544 ( .A(n4585), .Y(n4583) );
  INVX1 U546 ( .A(n4583), .Y(n4584) );
  AND2X1 U547 ( .A(n10825), .B(n1662), .Y(n1697) );
  INVX1 U549 ( .A(n1697), .Y(n4585) );
  INVX1 U551 ( .A(n4588), .Y(n4586) );
  INVX1 U553 ( .A(n4586), .Y(n4587) );
  AND2X1 U555 ( .A(n10828), .B(n1662), .Y(n1696) );
  INVX1 U557 ( .A(n1696), .Y(n4588) );
  INVX1 U559 ( .A(n4591), .Y(n4589) );
  INVX1 U561 ( .A(n4589), .Y(n4590) );
  AND2X1 U563 ( .A(n10831), .B(n1662), .Y(n1695) );
  INVX1 U565 ( .A(n1695), .Y(n4591) );
  INVX1 U567 ( .A(n4594), .Y(n4592) );
  INVX1 U569 ( .A(n4592), .Y(n4593) );
  AND2X1 U571 ( .A(n10834), .B(n1662), .Y(n1694) );
  INVX1 U573 ( .A(n1694), .Y(n4594) );
  INVX1 U575 ( .A(n4597), .Y(n4595) );
  INVX1 U577 ( .A(n4595), .Y(n4596) );
  AND2X1 U579 ( .A(n10837), .B(n1662), .Y(n1693) );
  INVX1 U581 ( .A(n1693), .Y(n4597) );
  INVX1 U583 ( .A(n4600), .Y(n4598) );
  INVX1 U585 ( .A(n4598), .Y(n4599) );
  AND2X1 U587 ( .A(n10840), .B(n1662), .Y(n1692) );
  INVX1 U589 ( .A(n1692), .Y(n4600) );
  INVX1 U591 ( .A(n4603), .Y(n4601) );
  INVX1 U593 ( .A(n4601), .Y(n4602) );
  AND2X1 U595 ( .A(n10843), .B(n1662), .Y(n1691) );
  INVX1 U597 ( .A(n1691), .Y(n4603) );
  INVX1 U599 ( .A(n4606), .Y(n4604) );
  INVX1 U601 ( .A(n4604), .Y(n4605) );
  AND2X1 U603 ( .A(n10846), .B(n1662), .Y(n1690) );
  INVX1 U605 ( .A(n1690), .Y(n4606) );
  INVX1 U607 ( .A(n4609), .Y(n4607) );
  INVX1 U609 ( .A(n4607), .Y(n4608) );
  AND2X1 U611 ( .A(n10849), .B(n1662), .Y(n1689) );
  INVX1 U613 ( .A(n1689), .Y(n4609) );
  INVX1 U615 ( .A(n4612), .Y(n4610) );
  INVX1 U617 ( .A(n4610), .Y(n4611) );
  AND2X1 U619 ( .A(n10852), .B(n1662), .Y(n1688) );
  INVX1 U621 ( .A(n1688), .Y(n4612) );
  INVX1 U623 ( .A(n4615), .Y(n4613) );
  INVX1 U625 ( .A(n4613), .Y(n4614) );
  AND2X1 U627 ( .A(n10855), .B(n1662), .Y(n1687) );
  INVX1 U629 ( .A(n1687), .Y(n4615) );
  INVX1 U631 ( .A(n4618), .Y(n4616) );
  INVX1 U632 ( .A(n4616), .Y(n4617) );
  AND2X1 U634 ( .A(n10858), .B(n1662), .Y(n1686) );
  INVX1 U636 ( .A(n1686), .Y(n4618) );
  INVX1 U638 ( .A(n4621), .Y(n4619) );
  INVX1 U640 ( .A(n4619), .Y(n4620) );
  AND2X1 U642 ( .A(n10861), .B(n1662), .Y(n1685) );
  INVX1 U644 ( .A(n1685), .Y(n4621) );
  INVX1 U646 ( .A(n4624), .Y(n4622) );
  INVX1 U648 ( .A(n4622), .Y(n4623) );
  AND2X1 U650 ( .A(n10864), .B(n1662), .Y(n1684) );
  INVX1 U652 ( .A(n1684), .Y(n4624) );
  INVX1 U654 ( .A(n4627), .Y(n4625) );
  INVX1 U656 ( .A(n4625), .Y(n4626) );
  AND2X1 U658 ( .A(n10867), .B(n1662), .Y(n1683) );
  INVX1 U660 ( .A(n1683), .Y(n4627) );
  INVX1 U662 ( .A(n4630), .Y(n4628) );
  INVX1 U664 ( .A(n4628), .Y(n4629) );
  AND2X1 U666 ( .A(n10870), .B(n1662), .Y(n1682) );
  INVX1 U668 ( .A(n1682), .Y(n4630) );
  INVX1 U670 ( .A(n4633), .Y(n4631) );
  INVX1 U672 ( .A(n4631), .Y(n4632) );
  AND2X1 U674 ( .A(n10873), .B(n1662), .Y(n1681) );
  INVX1 U676 ( .A(n1681), .Y(n4633) );
  INVX1 U678 ( .A(n4636), .Y(n4634) );
  INVX1 U680 ( .A(n4634), .Y(n4635) );
  AND2X1 U682 ( .A(n10876), .B(n1662), .Y(n1680) );
  INVX1 U684 ( .A(n1680), .Y(n4636) );
  INVX1 U686 ( .A(n4639), .Y(n4637) );
  INVX1 U688 ( .A(n4637), .Y(n4638) );
  AND2X1 U690 ( .A(n10879), .B(n1662), .Y(n1679) );
  INVX1 U692 ( .A(n1679), .Y(n4639) );
  INVX1 U694 ( .A(n4642), .Y(n4640) );
  INVX1 U696 ( .A(n4640), .Y(n4641) );
  AND2X1 U698 ( .A(n10882), .B(n1662), .Y(n1678) );
  INVX1 U700 ( .A(n1678), .Y(n4642) );
  INVX1 U702 ( .A(n4645), .Y(n4643) );
  INVX1 U704 ( .A(n4643), .Y(n4644) );
  AND2X1 U706 ( .A(n10885), .B(n1662), .Y(n1677) );
  INVX1 U708 ( .A(n1677), .Y(n4645) );
  INVX1 U710 ( .A(n4648), .Y(n4646) );
  INVX1 U712 ( .A(n4646), .Y(n4647) );
  AND2X1 U714 ( .A(n10888), .B(n1662), .Y(n1676) );
  INVX1 U716 ( .A(n1676), .Y(n4648) );
  INVX1 U717 ( .A(n4651), .Y(n4649) );
  INVX1 U719 ( .A(n4649), .Y(n4650) );
  AND2X1 U721 ( .A(n10891), .B(n1662), .Y(n1675) );
  INVX1 U723 ( .A(n1675), .Y(n4651) );
  INVX1 U725 ( .A(n4654), .Y(n4652) );
  INVX1 U727 ( .A(n4652), .Y(n4653) );
  AND2X1 U729 ( .A(n10894), .B(n1662), .Y(n1674) );
  INVX1 U731 ( .A(n1674), .Y(n4654) );
  INVX1 U733 ( .A(n4657), .Y(n4655) );
  INVX1 U735 ( .A(n4655), .Y(n4656) );
  AND2X1 U737 ( .A(n10897), .B(n1662), .Y(n1673) );
  INVX1 U739 ( .A(n1673), .Y(n4657) );
  INVX1 U741 ( .A(n4660), .Y(n4658) );
  INVX1 U743 ( .A(n4658), .Y(n4659) );
  AND2X1 U745 ( .A(n10900), .B(n1662), .Y(n1672) );
  INVX1 U747 ( .A(n1672), .Y(n4660) );
  INVX1 U749 ( .A(n4663), .Y(n4661) );
  INVX1 U751 ( .A(n4661), .Y(n4662) );
  AND2X1 U753 ( .A(n10903), .B(n1662), .Y(n1671) );
  INVX1 U755 ( .A(n1671), .Y(n4663) );
  INVX1 U757 ( .A(n4666), .Y(n4664) );
  INVX1 U759 ( .A(n4664), .Y(n4665) );
  AND2X1 U761 ( .A(n10906), .B(n1662), .Y(n1670) );
  INVX1 U763 ( .A(n1670), .Y(n4666) );
  INVX1 U765 ( .A(n4669), .Y(n4667) );
  INVX1 U767 ( .A(n4667), .Y(n4668) );
  AND2X1 U769 ( .A(n10909), .B(n1662), .Y(n1669) );
  INVX1 U771 ( .A(n1669), .Y(n4669) );
  INVX1 U773 ( .A(n4672), .Y(n4670) );
  INVX1 U775 ( .A(n4670), .Y(n4671) );
  AND2X1 U777 ( .A(n10912), .B(n1662), .Y(n1668) );
  INVX1 U779 ( .A(n1668), .Y(n4672) );
  INVX1 U781 ( .A(n4675), .Y(n4673) );
  INVX1 U783 ( .A(n4673), .Y(n4674) );
  AND2X1 U785 ( .A(n10915), .B(n1662), .Y(n1667) );
  INVX1 U787 ( .A(n1667), .Y(n4675) );
  INVX1 U789 ( .A(n4678), .Y(n4676) );
  INVX1 U791 ( .A(n4676), .Y(n4677) );
  AND2X1 U793 ( .A(n10918), .B(n1662), .Y(n1666) );
  INVX1 U795 ( .A(n1666), .Y(n4678) );
  INVX1 U797 ( .A(n4681), .Y(n4679) );
  INVX1 U799 ( .A(n4679), .Y(n4680) );
  AND2X1 U801 ( .A(n10921), .B(n1662), .Y(n1665) );
  INVX1 U802 ( .A(n1665), .Y(n4681) );
  INVX1 U803 ( .A(n4684), .Y(n4682) );
  INVX1 U806 ( .A(n4682), .Y(n4683) );
  AND2X1 U808 ( .A(n10924), .B(n1662), .Y(n1664) );
  INVX1 U810 ( .A(n1664), .Y(n4684) );
  INVX1 U812 ( .A(n4687), .Y(n4685) );
  INVX1 U814 ( .A(n4685), .Y(n4686) );
  AND2X1 U816 ( .A(n10927), .B(n1662), .Y(n1663) );
  INVX1 U818 ( .A(n1663), .Y(n4687) );
  INVX1 U820 ( .A(n4690), .Y(n4688) );
  INVX1 U822 ( .A(n4688), .Y(n4689) );
  AND2X1 U824 ( .A(n8780), .B(n1619), .Y(n1661) );
  INVX1 U826 ( .A(n1661), .Y(n4690) );
  INVX1 U828 ( .A(n4693), .Y(n4691) );
  INVX1 U830 ( .A(n4691), .Y(n4692) );
  AND2X1 U832 ( .A(n8783), .B(n1619), .Y(n1660) );
  INVX1 U834 ( .A(n1660), .Y(n4693) );
  INVX1 U836 ( .A(n4696), .Y(n4694) );
  INVX1 U838 ( .A(n4694), .Y(n4695) );
  AND2X1 U840 ( .A(n8786), .B(n1619), .Y(n1659) );
  INVX1 U842 ( .A(n1659), .Y(n4696) );
  INVX1 U844 ( .A(n4699), .Y(n4697) );
  INVX1 U846 ( .A(n4697), .Y(n4698) );
  AND2X1 U848 ( .A(n8789), .B(n1619), .Y(n1658) );
  INVX1 U850 ( .A(n1658), .Y(n4699) );
  INVX1 U852 ( .A(n4702), .Y(n4700) );
  INVX1 U854 ( .A(n4700), .Y(n4701) );
  AND2X1 U856 ( .A(n8792), .B(n1619), .Y(n1657) );
  INVX1 U858 ( .A(n1657), .Y(n4702) );
  INVX1 U860 ( .A(n4705), .Y(n4703) );
  INVX1 U862 ( .A(n4703), .Y(n4704) );
  AND2X1 U864 ( .A(n8795), .B(n1619), .Y(n1656) );
  INVX1 U866 ( .A(n1656), .Y(n4705) );
  INVX1 U868 ( .A(n4708), .Y(n4706) );
  INVX1 U870 ( .A(n4706), .Y(n4707) );
  AND2X1 U872 ( .A(n8798), .B(n1619), .Y(n1655) );
  INVX1 U874 ( .A(n1655), .Y(n4708) );
  INVX1 U876 ( .A(n4711), .Y(n4709) );
  INVX1 U878 ( .A(n4709), .Y(n4710) );
  AND2X1 U880 ( .A(n8801), .B(n1619), .Y(n1654) );
  INVX1 U882 ( .A(n1654), .Y(n4711) );
  INVX1 U884 ( .A(n4714), .Y(n4712) );
  INVX1 U886 ( .A(n4712), .Y(n4713) );
  AND2X1 U888 ( .A(n8804), .B(n1619), .Y(n1653) );
  INVX1 U889 ( .A(n1653), .Y(n4714) );
  INVX1 U891 ( .A(n4717), .Y(n4715) );
  INVX1 U893 ( .A(n4715), .Y(n4716) );
  AND2X1 U895 ( .A(n8807), .B(n1619), .Y(n1652) );
  INVX1 U897 ( .A(n1652), .Y(n4717) );
  INVX1 U899 ( .A(n4720), .Y(n4718) );
  INVX1 U901 ( .A(n4718), .Y(n4719) );
  AND2X1 U903 ( .A(n8810), .B(n1619), .Y(n1651) );
  INVX1 U905 ( .A(n1651), .Y(n4720) );
  INVX1 U907 ( .A(n4723), .Y(n4721) );
  INVX1 U909 ( .A(n4721), .Y(n4722) );
  AND2X1 U911 ( .A(n8813), .B(n1619), .Y(n1650) );
  INVX1 U913 ( .A(n1650), .Y(n4723) );
  INVX1 U915 ( .A(n4726), .Y(n4724) );
  INVX1 U917 ( .A(n4724), .Y(n4725) );
  AND2X1 U919 ( .A(n8816), .B(n1619), .Y(n1649) );
  INVX1 U921 ( .A(n1649), .Y(n4726) );
  INVX1 U923 ( .A(n4729), .Y(n4727) );
  INVX1 U925 ( .A(n4727), .Y(n4728) );
  AND2X1 U927 ( .A(n8819), .B(n1619), .Y(n1648) );
  INVX1 U929 ( .A(n1648), .Y(n4729) );
  INVX1 U931 ( .A(n4732), .Y(n4730) );
  INVX1 U933 ( .A(n4730), .Y(n4731) );
  AND2X1 U935 ( .A(n8822), .B(n1619), .Y(n1647) );
  INVX1 U937 ( .A(n1647), .Y(n4732) );
  INVX1 U939 ( .A(n4735), .Y(n4733) );
  INVX1 U941 ( .A(n4733), .Y(n4734) );
  AND2X1 U943 ( .A(n8825), .B(n1619), .Y(n1646) );
  INVX1 U945 ( .A(n1646), .Y(n4735) );
  INVX1 U947 ( .A(n4738), .Y(n4736) );
  INVX1 U949 ( .A(n4736), .Y(n4737) );
  AND2X1 U951 ( .A(n8828), .B(n1619), .Y(n1645) );
  INVX1 U953 ( .A(n1645), .Y(n4738) );
  INVX1 U955 ( .A(n4741), .Y(n4739) );
  INVX1 U957 ( .A(n4739), .Y(n4740) );
  AND2X1 U959 ( .A(n8831), .B(n1619), .Y(n1644) );
  INVX1 U961 ( .A(n1644), .Y(n4741) );
  INVX1 U963 ( .A(n4744), .Y(n4742) );
  INVX1 U965 ( .A(n4742), .Y(n4743) );
  AND2X1 U967 ( .A(n8834), .B(n1619), .Y(n1643) );
  INVX1 U969 ( .A(n1643), .Y(n4744) );
  INVX1 U971 ( .A(n4747), .Y(n4745) );
  INVX1 U973 ( .A(n4745), .Y(n4746) );
  AND2X1 U974 ( .A(n8837), .B(n1619), .Y(n1642) );
  INVX1 U976 ( .A(n1642), .Y(n4747) );
  INVX1 U978 ( .A(n4750), .Y(n4748) );
  INVX1 U980 ( .A(n4748), .Y(n4749) );
  AND2X1 U982 ( .A(n8840), .B(n1619), .Y(n1641) );
  INVX1 U984 ( .A(n1641), .Y(n4750) );
  INVX1 U986 ( .A(n4753), .Y(n4751) );
  INVX1 U988 ( .A(n4751), .Y(n4752) );
  AND2X1 U990 ( .A(n8843), .B(n1619), .Y(n1640) );
  INVX1 U992 ( .A(n1640), .Y(n4753) );
  INVX1 U994 ( .A(n4756), .Y(n4754) );
  INVX1 U996 ( .A(n4754), .Y(n4755) );
  AND2X1 U998 ( .A(n8846), .B(n1619), .Y(n1639) );
  INVX1 U1000 ( .A(n1639), .Y(n4756) );
  INVX1 U1002 ( .A(n4759), .Y(n4757) );
  INVX1 U1004 ( .A(n4757), .Y(n4758) );
  AND2X1 U1006 ( .A(n8849), .B(n1619), .Y(n1638) );
  INVX1 U1008 ( .A(n1638), .Y(n4759) );
  INVX1 U1010 ( .A(n4762), .Y(n4760) );
  INVX1 U1012 ( .A(n4760), .Y(n4761) );
  AND2X1 U1014 ( .A(n8852), .B(n1619), .Y(n1637) );
  INVX1 U1016 ( .A(n1637), .Y(n4762) );
  INVX1 U1018 ( .A(n4765), .Y(n4763) );
  INVX1 U1020 ( .A(n4763), .Y(n4764) );
  AND2X1 U1022 ( .A(n8855), .B(n1619), .Y(n1636) );
  INVX1 U1024 ( .A(n1636), .Y(n4765) );
  INVX1 U1026 ( .A(n4768), .Y(n4766) );
  INVX1 U1028 ( .A(n4766), .Y(n4767) );
  AND2X1 U1030 ( .A(n8858), .B(n1619), .Y(n1635) );
  INVX1 U1032 ( .A(n1635), .Y(n4768) );
  INVX1 U1034 ( .A(n4771), .Y(n4769) );
  INVX1 U1036 ( .A(n4769), .Y(n4770) );
  AND2X1 U1038 ( .A(n8861), .B(n1619), .Y(n1634) );
  INVX1 U1040 ( .A(n1634), .Y(n4771) );
  INVX1 U1042 ( .A(n4774), .Y(n4772) );
  INVX1 U1044 ( .A(n4772), .Y(n4773) );
  AND2X1 U1046 ( .A(n8864), .B(n1619), .Y(n1633) );
  INVX1 U1048 ( .A(n1633), .Y(n4774) );
  INVX1 U1050 ( .A(n4777), .Y(n4775) );
  INVX1 U1052 ( .A(n4775), .Y(n4776) );
  AND2X1 U1054 ( .A(n8867), .B(n1619), .Y(n1632) );
  INVX1 U1056 ( .A(n1632), .Y(n4777) );
  INVX1 U1058 ( .A(n4780), .Y(n4778) );
  INVX1 U1059 ( .A(n4778), .Y(n4779) );
  AND2X1 U1061 ( .A(n8870), .B(n1619), .Y(n1631) );
  INVX1 U1063 ( .A(n1631), .Y(n4780) );
  INVX1 U1065 ( .A(n4783), .Y(n4781) );
  INVX1 U1067 ( .A(n4781), .Y(n4782) );
  AND2X1 U1069 ( .A(n8873), .B(n1619), .Y(n1630) );
  INVX1 U1071 ( .A(n1630), .Y(n4783) );
  INVX1 U1073 ( .A(n4786), .Y(n4784) );
  INVX1 U1075 ( .A(n4784), .Y(n4785) );
  AND2X1 U1077 ( .A(n8876), .B(n1619), .Y(n1629) );
  INVX1 U1079 ( .A(n1629), .Y(n4786) );
  INVX1 U1081 ( .A(n4789), .Y(n4787) );
  INVX1 U1083 ( .A(n4787), .Y(n4788) );
  AND2X1 U1085 ( .A(n8879), .B(n1619), .Y(n1628) );
  INVX1 U1087 ( .A(n1628), .Y(n4789) );
  INVX1 U1089 ( .A(n4792), .Y(n4790) );
  INVX1 U1091 ( .A(n4790), .Y(n4791) );
  AND2X1 U1093 ( .A(n8882), .B(n1619), .Y(n1627) );
  INVX1 U1095 ( .A(n1627), .Y(n4792) );
  INVX1 U1097 ( .A(n4795), .Y(n4793) );
  INVX1 U1099 ( .A(n4793), .Y(n4794) );
  AND2X1 U1101 ( .A(n8885), .B(n1619), .Y(n1626) );
  INVX1 U1103 ( .A(n1626), .Y(n4795) );
  INVX1 U1105 ( .A(n4798), .Y(n4796) );
  INVX1 U1107 ( .A(n4796), .Y(n4797) );
  AND2X1 U1109 ( .A(n8888), .B(n1619), .Y(n1625) );
  INVX1 U1111 ( .A(n1625), .Y(n4798) );
  INVX1 U1113 ( .A(n4801), .Y(n4799) );
  INVX1 U1115 ( .A(n4799), .Y(n4800) );
  AND2X1 U1117 ( .A(n8891), .B(n1619), .Y(n1624) );
  INVX1 U1119 ( .A(n1624), .Y(n4801) );
  INVX1 U1121 ( .A(n4804), .Y(n4802) );
  INVX1 U1123 ( .A(n4802), .Y(n4803) );
  AND2X1 U1125 ( .A(n8894), .B(n1619), .Y(n1623) );
  INVX1 U1127 ( .A(n1623), .Y(n4804) );
  INVX1 U1129 ( .A(n4807), .Y(n4805) );
  INVX1 U1131 ( .A(n4805), .Y(n4806) );
  AND2X1 U1133 ( .A(n8897), .B(n1619), .Y(n1622) );
  INVX1 U1135 ( .A(n1622), .Y(n4807) );
  INVX1 U1137 ( .A(n4810), .Y(n4808) );
  INVX1 U1139 ( .A(n4808), .Y(n4809) );
  AND2X1 U1141 ( .A(n8900), .B(n1619), .Y(n1621) );
  INVX1 U1143 ( .A(n1621), .Y(n4810) );
  INVX1 U1144 ( .A(n4813), .Y(n4811) );
  INVX1 U1146 ( .A(n4811), .Y(n4812) );
  AND2X1 U1148 ( .A(n8903), .B(n1619), .Y(n1620) );
  INVX1 U1150 ( .A(n1620), .Y(n4813) );
  INVX1 U1152 ( .A(n4816), .Y(n4814) );
  INVX1 U1154 ( .A(n4814), .Y(n4815) );
  AND2X1 U1156 ( .A(n10930), .B(n1576), .Y(n1618) );
  INVX1 U1158 ( .A(n1618), .Y(n4816) );
  INVX1 U1160 ( .A(n4819), .Y(n4817) );
  INVX1 U1162 ( .A(n4817), .Y(n4818) );
  AND2X1 U1164 ( .A(n10933), .B(n1576), .Y(n1617) );
  INVX1 U1166 ( .A(n1617), .Y(n4819) );
  INVX1 U1168 ( .A(n4822), .Y(n4820) );
  INVX1 U1170 ( .A(n4820), .Y(n4821) );
  AND2X1 U1172 ( .A(n10936), .B(n1576), .Y(n1616) );
  INVX1 U1174 ( .A(n1616), .Y(n4822) );
  INVX1 U1176 ( .A(n4825), .Y(n4823) );
  INVX1 U1178 ( .A(n4823), .Y(n4824) );
  AND2X1 U1180 ( .A(n10939), .B(n1576), .Y(n1615) );
  INVX1 U1182 ( .A(n1615), .Y(n4825) );
  INVX1 U1184 ( .A(n4828), .Y(n4826) );
  INVX1 U1186 ( .A(n4826), .Y(n4827) );
  AND2X1 U1188 ( .A(n10942), .B(n1576), .Y(n1614) );
  INVX1 U1190 ( .A(n1614), .Y(n4828) );
  INVX1 U1192 ( .A(n4831), .Y(n4829) );
  INVX1 U1194 ( .A(n4829), .Y(n4830) );
  AND2X1 U1196 ( .A(n10945), .B(n1576), .Y(n1613) );
  INVX1 U1198 ( .A(n1613), .Y(n4831) );
  INVX1 U1200 ( .A(n4834), .Y(n4832) );
  INVX1 U1202 ( .A(n4832), .Y(n4833) );
  AND2X1 U1204 ( .A(n10948), .B(n1576), .Y(n1612) );
  INVX1 U1206 ( .A(n1612), .Y(n4834) );
  INVX1 U1208 ( .A(n4837), .Y(n4835) );
  INVX1 U1210 ( .A(n4835), .Y(n4836) );
  AND2X1 U1212 ( .A(n10951), .B(n1576), .Y(n1611) );
  INVX1 U1214 ( .A(n1611), .Y(n4837) );
  INVX1 U1216 ( .A(n4840), .Y(n4838) );
  INVX1 U1218 ( .A(n4838), .Y(n4839) );
  AND2X1 U1220 ( .A(n10954), .B(n1576), .Y(n1610) );
  INVX1 U1222 ( .A(n1610), .Y(n4840) );
  INVX1 U1224 ( .A(n4843), .Y(n4841) );
  INVX1 U1226 ( .A(n4841), .Y(n4842) );
  AND2X1 U1228 ( .A(n10957), .B(n1576), .Y(n1609) );
  INVX1 U1229 ( .A(n1609), .Y(n4843) );
  INVX1 U1231 ( .A(n4846), .Y(n4844) );
  INVX1 U1233 ( .A(n4844), .Y(n4845) );
  AND2X1 U1235 ( .A(n10960), .B(n1576), .Y(n1608) );
  INVX1 U1237 ( .A(n1608), .Y(n4846) );
  INVX1 U1239 ( .A(n4849), .Y(n4847) );
  INVX1 U1241 ( .A(n4847), .Y(n4848) );
  AND2X1 U1243 ( .A(n10963), .B(n1576), .Y(n1607) );
  INVX1 U1245 ( .A(n1607), .Y(n4849) );
  INVX1 U1247 ( .A(n4852), .Y(n4850) );
  INVX1 U1249 ( .A(n4850), .Y(n4851) );
  AND2X1 U1251 ( .A(n10966), .B(n1576), .Y(n1606) );
  INVX1 U1253 ( .A(n1606), .Y(n4852) );
  INVX1 U1255 ( .A(n4855), .Y(n4853) );
  INVX1 U1257 ( .A(n4853), .Y(n4854) );
  AND2X1 U1259 ( .A(n10969), .B(n1576), .Y(n1605) );
  INVX1 U1261 ( .A(n1605), .Y(n4855) );
  INVX1 U1263 ( .A(n4858), .Y(n4856) );
  INVX1 U1265 ( .A(n4856), .Y(n4857) );
  AND2X1 U1267 ( .A(n10972), .B(n1576), .Y(n1604) );
  INVX1 U1269 ( .A(n1604), .Y(n4858) );
  INVX1 U1271 ( .A(n4861), .Y(n4859) );
  INVX1 U1273 ( .A(n4859), .Y(n4860) );
  AND2X1 U1275 ( .A(n10975), .B(n1576), .Y(n1603) );
  INVX1 U1277 ( .A(n1603), .Y(n4861) );
  INVX1 U1279 ( .A(n4864), .Y(n4862) );
  INVX1 U1281 ( .A(n4862), .Y(n4863) );
  AND2X1 U1283 ( .A(n10978), .B(n1576), .Y(n1602) );
  INVX1 U1285 ( .A(n1602), .Y(n4864) );
  INVX1 U1287 ( .A(n4867), .Y(n4865) );
  INVX1 U1289 ( .A(n4865), .Y(n4866) );
  AND2X1 U1291 ( .A(n10981), .B(n1576), .Y(n1601) );
  INVX1 U1293 ( .A(n1601), .Y(n4867) );
  INVX1 U1295 ( .A(n4870), .Y(n4868) );
  INVX1 U1297 ( .A(n4868), .Y(n4869) );
  AND2X1 U1299 ( .A(n10984), .B(n1576), .Y(n1600) );
  INVX1 U1301 ( .A(n1600), .Y(n4870) );
  INVX1 U1303 ( .A(n4873), .Y(n4871) );
  INVX1 U1305 ( .A(n4871), .Y(n4872) );
  AND2X1 U1307 ( .A(n10987), .B(n1576), .Y(n1599) );
  INVX1 U1309 ( .A(n1599), .Y(n4873) );
  INVX1 U1311 ( .A(n4876), .Y(n4874) );
  INVX1 U1313 ( .A(n4874), .Y(n4875) );
  AND2X1 U1314 ( .A(n10990), .B(n1576), .Y(n1598) );
  INVX1 U1316 ( .A(n1598), .Y(n4876) );
  INVX1 U1318 ( .A(n4879), .Y(n4877) );
  INVX1 U1320 ( .A(n4877), .Y(n4878) );
  AND2X1 U1322 ( .A(n10993), .B(n1576), .Y(n1597) );
  INVX1 U1324 ( .A(n1597), .Y(n4879) );
  INVX1 U1326 ( .A(n4882), .Y(n4880) );
  INVX1 U1328 ( .A(n4880), .Y(n4881) );
  AND2X1 U1330 ( .A(n10996), .B(n1576), .Y(n1596) );
  INVX1 U1332 ( .A(n1596), .Y(n4882) );
  INVX1 U1334 ( .A(n4885), .Y(n4883) );
  INVX1 U1336 ( .A(n4883), .Y(n4884) );
  AND2X1 U1338 ( .A(n10999), .B(n1576), .Y(n1595) );
  INVX1 U1340 ( .A(n1595), .Y(n4885) );
  INVX1 U1342 ( .A(n4888), .Y(n4886) );
  INVX1 U1344 ( .A(n4886), .Y(n4887) );
  AND2X1 U1346 ( .A(n11002), .B(n1576), .Y(n1594) );
  INVX1 U1348 ( .A(n1594), .Y(n4888) );
  INVX1 U1350 ( .A(n4891), .Y(n4889) );
  INVX1 U1352 ( .A(n4889), .Y(n4890) );
  AND2X1 U1354 ( .A(n11005), .B(n1576), .Y(n1593) );
  INVX1 U1356 ( .A(n1593), .Y(n4891) );
  INVX1 U1358 ( .A(n4894), .Y(n4892) );
  INVX1 U1360 ( .A(n4892), .Y(n4893) );
  AND2X1 U1362 ( .A(n11008), .B(n1576), .Y(n1592) );
  INVX1 U1364 ( .A(n1592), .Y(n4894) );
  INVX1 U1366 ( .A(n4897), .Y(n4895) );
  INVX1 U1368 ( .A(n4895), .Y(n4896) );
  AND2X1 U1370 ( .A(n11011), .B(n1576), .Y(n1591) );
  INVX1 U1372 ( .A(n1591), .Y(n4897) );
  INVX1 U1374 ( .A(n4900), .Y(n4898) );
  INVX1 U1376 ( .A(n4898), .Y(n4899) );
  AND2X1 U1378 ( .A(n11014), .B(n1576), .Y(n1590) );
  INVX1 U1380 ( .A(n1590), .Y(n4900) );
  INVX1 U1382 ( .A(n4903), .Y(n4901) );
  INVX1 U1384 ( .A(n4901), .Y(n4902) );
  AND2X1 U1386 ( .A(n11017), .B(n1576), .Y(n1589) );
  INVX1 U1388 ( .A(n1589), .Y(n4903) );
  INVX1 U1390 ( .A(n4906), .Y(n4904) );
  INVX1 U1392 ( .A(n4904), .Y(n4905) );
  AND2X1 U1394 ( .A(n11020), .B(n1576), .Y(n1588) );
  INVX1 U1396 ( .A(n1588), .Y(n4906) );
  INVX1 U1398 ( .A(n4909), .Y(n4907) );
  INVX1 U1399 ( .A(n4907), .Y(n4908) );
  AND2X1 U1401 ( .A(n11023), .B(n1576), .Y(n1587) );
  INVX1 U1403 ( .A(n1587), .Y(n4909) );
  INVX1 U1405 ( .A(n4912), .Y(n4910) );
  INVX1 U1407 ( .A(n4910), .Y(n4911) );
  AND2X1 U1409 ( .A(n11026), .B(n1576), .Y(n1586) );
  INVX1 U1411 ( .A(n1586), .Y(n4912) );
  INVX1 U1413 ( .A(n4915), .Y(n4913) );
  INVX1 U1415 ( .A(n4913), .Y(n4914) );
  AND2X1 U1417 ( .A(n11029), .B(n1576), .Y(n1585) );
  INVX1 U1419 ( .A(n1585), .Y(n4915) );
  INVX1 U1421 ( .A(n4918), .Y(n4916) );
  INVX1 U1423 ( .A(n4916), .Y(n4917) );
  AND2X1 U1425 ( .A(n11032), .B(n1576), .Y(n1584) );
  INVX1 U1427 ( .A(n1584), .Y(n4918) );
  INVX1 U1429 ( .A(n4921), .Y(n4919) );
  INVX1 U1431 ( .A(n4919), .Y(n4920) );
  AND2X1 U1433 ( .A(n11035), .B(n1576), .Y(n1583) );
  INVX1 U1435 ( .A(n1583), .Y(n4921) );
  INVX1 U1437 ( .A(n4924), .Y(n4922) );
  INVX1 U1439 ( .A(n4922), .Y(n4923) );
  AND2X1 U1441 ( .A(n11038), .B(n1576), .Y(n1582) );
  INVX1 U1443 ( .A(n1582), .Y(n4924) );
  INVX1 U1445 ( .A(n4927), .Y(n4925) );
  INVX1 U1447 ( .A(n4925), .Y(n4926) );
  AND2X1 U1449 ( .A(n11041), .B(n1576), .Y(n1581) );
  INVX1 U1451 ( .A(n1581), .Y(n4927) );
  INVX1 U1453 ( .A(n4930), .Y(n4928) );
  INVX1 U1455 ( .A(n4928), .Y(n4929) );
  AND2X1 U1457 ( .A(n11044), .B(n1576), .Y(n1580) );
  INVX1 U1459 ( .A(n1580), .Y(n4930) );
  INVX1 U1461 ( .A(n4933), .Y(n4931) );
  INVX1 U1463 ( .A(n4931), .Y(n4932) );
  AND2X1 U1465 ( .A(n11047), .B(n1576), .Y(n1579) );
  INVX1 U1467 ( .A(n1579), .Y(n4933) );
  INVX1 U1469 ( .A(n4936), .Y(n4934) );
  INVX1 U1471 ( .A(n4934), .Y(n4935) );
  AND2X1 U1473 ( .A(n11050), .B(n1576), .Y(n1578) );
  INVX1 U1475 ( .A(n1578), .Y(n4936) );
  INVX1 U1477 ( .A(n4939), .Y(n4937) );
  INVX1 U1479 ( .A(n4937), .Y(n4938) );
  AND2X1 U1481 ( .A(n11053), .B(n1576), .Y(n1577) );
  INVX1 U1483 ( .A(n1577), .Y(n4939) );
  INVX1 U1484 ( .A(n4942), .Y(n4940) );
  INVX1 U1485 ( .A(n4940), .Y(n4941) );
  AND2X1 U1489 ( .A(n8906), .B(n13045), .Y(n1574) );
  INVX1 U1491 ( .A(n1574), .Y(n4942) );
  INVX1 U1493 ( .A(n4945), .Y(n4943) );
  INVX1 U1495 ( .A(n4943), .Y(n4944) );
  AND2X1 U1497 ( .A(n8909), .B(n12992), .Y(n1573) );
  INVX1 U1499 ( .A(n1573), .Y(n4945) );
  INVX1 U1501 ( .A(n4948), .Y(n4946) );
  INVX1 U1503 ( .A(n4946), .Y(n4947) );
  AND2X1 U1505 ( .A(n8912), .B(n13045), .Y(n1572) );
  INVX1 U1507 ( .A(n1572), .Y(n4948) );
  INVX1 U1509 ( .A(n4951), .Y(n4949) );
  INVX1 U1511 ( .A(n4949), .Y(n4950) );
  AND2X1 U1513 ( .A(n8915), .B(n12969), .Y(n1571) );
  INVX1 U1515 ( .A(n1571), .Y(n4951) );
  INVX1 U1517 ( .A(n4954), .Y(n4952) );
  INVX1 U1519 ( .A(n4952), .Y(n4953) );
  AND2X1 U1521 ( .A(n8918), .B(n13045), .Y(n1570) );
  INVX1 U1523 ( .A(n1570), .Y(n4954) );
  INVX1 U1525 ( .A(n4957), .Y(n4955) );
  INVX1 U1527 ( .A(n4955), .Y(n4956) );
  AND2X1 U1529 ( .A(n8921), .B(n13032), .Y(n1569) );
  INVX1 U1531 ( .A(n1569), .Y(n4957) );
  INVX1 U1533 ( .A(n4960), .Y(n4958) );
  INVX1 U1535 ( .A(n4958), .Y(n4959) );
  AND2X1 U1537 ( .A(n8924), .B(n13045), .Y(n1568) );
  INVX1 U1539 ( .A(n1568), .Y(n4960) );
  INVX1 U1541 ( .A(n4963), .Y(n4961) );
  INVX1 U1543 ( .A(n4961), .Y(n4962) );
  AND2X1 U1545 ( .A(n8927), .B(n12990), .Y(n1567) );
  INVX1 U1547 ( .A(n1567), .Y(n4963) );
  INVX1 U1549 ( .A(n4966), .Y(n4964) );
  INVX1 U1551 ( .A(n4964), .Y(n4965) );
  AND2X1 U1553 ( .A(n8930), .B(n13045), .Y(n1566) );
  INVX1 U1555 ( .A(n1566), .Y(n4966) );
  INVX1 U1557 ( .A(n4969), .Y(n4967) );
  INVX1 U1559 ( .A(n4967), .Y(n4968) );
  AND2X1 U1561 ( .A(n8933), .B(n12967), .Y(n1565) );
  INVX1 U1563 ( .A(n1565), .Y(n4969) );
  INVX1 U1565 ( .A(n4972), .Y(n4970) );
  INVX1 U1567 ( .A(n4970), .Y(n4971) );
  AND2X1 U1569 ( .A(n8936), .B(n13045), .Y(n1564) );
  INVX1 U1571 ( .A(n1564), .Y(n4972) );
  INVX1 U1572 ( .A(n4975), .Y(n4973) );
  INVX1 U1574 ( .A(n4973), .Y(n4974) );
  AND2X1 U1576 ( .A(n8939), .B(n13032), .Y(n1563) );
  INVX1 U1578 ( .A(n1563), .Y(n4975) );
  INVX1 U1580 ( .A(n4978), .Y(n4976) );
  INVX1 U1582 ( .A(n4976), .Y(n4977) );
  AND2X1 U1584 ( .A(n8942), .B(n13045), .Y(n1562) );
  INVX1 U1586 ( .A(n1562), .Y(n4978) );
  INVX1 U1588 ( .A(n4981), .Y(n4979) );
  INVX1 U1590 ( .A(n4979), .Y(n4980) );
  AND2X1 U1592 ( .A(n8945), .B(n10796), .Y(n1561) );
  INVX1 U1594 ( .A(n1561), .Y(n4981) );
  INVX1 U1596 ( .A(n4984), .Y(n4982) );
  INVX1 U1598 ( .A(n4982), .Y(n4983) );
  AND2X1 U1600 ( .A(n8948), .B(n13045), .Y(n1560) );
  INVX1 U1602 ( .A(n1560), .Y(n4984) );
  INVX1 U1604 ( .A(n4987), .Y(n4985) );
  INVX1 U1606 ( .A(n4985), .Y(n4986) );
  AND2X1 U1608 ( .A(n8951), .B(n12992), .Y(n1559) );
  INVX1 U1610 ( .A(n1559), .Y(n4987) );
  INVX1 U1612 ( .A(n4990), .Y(n4988) );
  INVX1 U1614 ( .A(n4988), .Y(n4989) );
  AND2X1 U1616 ( .A(n8954), .B(n13045), .Y(n1558) );
  INVX1 U1618 ( .A(n1558), .Y(n4990) );
  INVX1 U1620 ( .A(n4993), .Y(n4991) );
  INVX1 U1622 ( .A(n4991), .Y(n4992) );
  AND2X1 U1624 ( .A(n8957), .B(n13032), .Y(n1557) );
  INVX1 U1626 ( .A(n1557), .Y(n4993) );
  INVX1 U1628 ( .A(n4996), .Y(n4994) );
  INVX1 U1630 ( .A(n4994), .Y(n4995) );
  AND2X1 U1632 ( .A(n8960), .B(n13045), .Y(n1556) );
  INVX1 U1634 ( .A(n1556), .Y(n4996) );
  INVX1 U1636 ( .A(n4999), .Y(n4997) );
  INVX1 U1638 ( .A(n4997), .Y(n4998) );
  AND2X1 U1640 ( .A(n8963), .B(n12967), .Y(n1555) );
  INVX1 U1642 ( .A(n1555), .Y(n4999) );
  INVX1 U1644 ( .A(n5002), .Y(n5000) );
  INVX1 U1646 ( .A(n5000), .Y(n5001) );
  AND2X1 U1648 ( .A(n8966), .B(n13045), .Y(n1554) );
  INVX1 U1650 ( .A(n1554), .Y(n5002) );
  INVX1 U1652 ( .A(n5005), .Y(n5003) );
  INVX1 U1654 ( .A(n5003), .Y(n5004) );
  AND2X1 U1656 ( .A(n8969), .B(n12969), .Y(n1553) );
  INVX1 U1657 ( .A(n1553), .Y(n5005) );
  INVX1 U1659 ( .A(n5008), .Y(n5006) );
  INVX1 U1661 ( .A(n5006), .Y(n5007) );
  AND2X1 U1663 ( .A(n8972), .B(n13045), .Y(n1552) );
  INVX1 U1665 ( .A(n1552), .Y(n5008) );
  INVX1 U1667 ( .A(n5011), .Y(n5009) );
  INVX1 U1669 ( .A(n5009), .Y(n5010) );
  AND2X1 U1671 ( .A(n8975), .B(n13032), .Y(n1551) );
  INVX1 U1673 ( .A(n1551), .Y(n5011) );
  INVX1 U1675 ( .A(n5014), .Y(n5012) );
  INVX1 U1677 ( .A(n5012), .Y(n5013) );
  AND2X1 U1679 ( .A(n8978), .B(n13045), .Y(n1550) );
  INVX1 U1681 ( .A(n1550), .Y(n5014) );
  INVX1 U1683 ( .A(n5017), .Y(n5015) );
  INVX1 U1685 ( .A(n5015), .Y(n5016) );
  AND2X1 U1687 ( .A(n8981), .B(n12990), .Y(n1549) );
  INVX1 U1689 ( .A(n1549), .Y(n5017) );
  INVX1 U1691 ( .A(n5020), .Y(n5018) );
  INVX1 U1693 ( .A(n5018), .Y(n5019) );
  AND2X1 U1695 ( .A(n8984), .B(n13045), .Y(n1548) );
  INVX1 U1697 ( .A(n1548), .Y(n5020) );
  INVX1 U1699 ( .A(n5023), .Y(n5021) );
  INVX1 U1701 ( .A(n5021), .Y(n5022) );
  AND2X1 U1703 ( .A(n8987), .B(n8762), .Y(n1547) );
  INVX1 U1705 ( .A(n1547), .Y(n5023) );
  INVX1 U1707 ( .A(n5026), .Y(n5024) );
  INVX1 U1709 ( .A(n5024), .Y(n5025) );
  AND2X1 U1711 ( .A(n8990), .B(n13045), .Y(n1546) );
  INVX1 U1713 ( .A(n1546), .Y(n5026) );
  INVX1 U1715 ( .A(n5029), .Y(n5027) );
  INVX1 U1717 ( .A(n5027), .Y(n5028) );
  AND2X1 U1719 ( .A(n8993), .B(n13032), .Y(n1545) );
  INVX1 U1721 ( .A(n1545), .Y(n5029) );
  INVX1 U1723 ( .A(n5032), .Y(n5030) );
  INVX1 U1725 ( .A(n5030), .Y(n5031) );
  AND2X1 U1727 ( .A(n8996), .B(n13045), .Y(n1544) );
  INVX1 U1729 ( .A(n1544), .Y(n5032) );
  INVX1 U1731 ( .A(n5035), .Y(n5033) );
  INVX1 U1733 ( .A(n5033), .Y(n5034) );
  AND2X1 U1735 ( .A(n8999), .B(n12990), .Y(n1543) );
  INVX1 U1737 ( .A(n1543), .Y(n5035) );
  INVX1 U1739 ( .A(n5038), .Y(n5036) );
  INVX1 U1741 ( .A(n5036), .Y(n5037) );
  AND2X1 U1742 ( .A(n9002), .B(n13045), .Y(n1542) );
  INVX1 U1744 ( .A(n1542), .Y(n5038) );
  INVX1 U1746 ( .A(n5041), .Y(n5039) );
  INVX1 U1748 ( .A(n5039), .Y(n5040) );
  AND2X1 U1750 ( .A(n9005), .B(n12969), .Y(n1541) );
  INVX1 U1752 ( .A(n1541), .Y(n5041) );
  INVX1 U1754 ( .A(n5044), .Y(n5042) );
  INVX1 U1756 ( .A(n5042), .Y(n5043) );
  AND2X1 U1758 ( .A(n9008), .B(n13045), .Y(n1540) );
  INVX1 U1760 ( .A(n1540), .Y(n5044) );
  INVX1 U1762 ( .A(n5047), .Y(n5045) );
  INVX1 U1764 ( .A(n5045), .Y(n5046) );
  AND2X1 U1766 ( .A(n9011), .B(n13032), .Y(n1539) );
  INVX1 U1768 ( .A(n1539), .Y(n5047) );
  INVX1 U1770 ( .A(n5050), .Y(n5048) );
  INVX1 U1772 ( .A(n5048), .Y(n5049) );
  AND2X1 U1774 ( .A(n9014), .B(n13045), .Y(n1538) );
  INVX1 U1776 ( .A(n1538), .Y(n5050) );
  INVX1 U1778 ( .A(n5053), .Y(n5051) );
  INVX1 U1780 ( .A(n5051), .Y(n5052) );
  AND2X1 U1782 ( .A(n9017), .B(n8662), .Y(n1537) );
  INVX1 U1784 ( .A(n1537), .Y(n5053) );
  INVX1 U1786 ( .A(n5056), .Y(n5054) );
  INVX1 U1788 ( .A(n5054), .Y(n5055) );
  AND2X1 U1790 ( .A(n9020), .B(n13045), .Y(n1536) );
  INVX1 U1792 ( .A(n1536), .Y(n5056) );
  INVX1 U1794 ( .A(n5059), .Y(n5057) );
  INVX1 U1796 ( .A(n5057), .Y(n5058) );
  AND2X1 U1798 ( .A(n9023), .B(n12992), .Y(n1535) );
  INVX1 U1800 ( .A(n1535), .Y(n5059) );
  INVX1 U1802 ( .A(n5062), .Y(n5060) );
  INVX1 U1804 ( .A(n5060), .Y(n5061) );
  AND2X1 U1806 ( .A(n9026), .B(n13045), .Y(n1534) );
  INVX1 U1808 ( .A(n1534), .Y(n5062) );
  INVX1 U1810 ( .A(n5065), .Y(n5063) );
  INVX1 U1812 ( .A(n5063), .Y(n5064) );
  AND2X1 U1814 ( .A(n9029), .B(n13032), .Y(n1533) );
  INVX1 U1816 ( .A(n1533), .Y(n5065) );
  INVX1 U1818 ( .A(n5068), .Y(n5066) );
  INVX1 U1820 ( .A(n5066), .Y(n5067) );
  AND2X1 U1822 ( .A(n11056), .B(n1489), .Y(n1531) );
  INVX1 U1824 ( .A(n1531), .Y(n5068) );
  INVX1 U1826 ( .A(n5071), .Y(n5069) );
  INVX1 U1827 ( .A(n5069), .Y(n5070) );
  AND2X1 U1829 ( .A(n11059), .B(n1489), .Y(n1530) );
  INVX1 U1831 ( .A(n1530), .Y(n5071) );
  INVX1 U1833 ( .A(n5074), .Y(n5072) );
  INVX1 U1835 ( .A(n5072), .Y(n5073) );
  AND2X1 U1837 ( .A(n11062), .B(n1489), .Y(n1529) );
  INVX1 U1839 ( .A(n1529), .Y(n5074) );
  INVX1 U1841 ( .A(n5077), .Y(n5075) );
  INVX1 U1843 ( .A(n5075), .Y(n5076) );
  AND2X1 U1845 ( .A(n11065), .B(n1489), .Y(n1528) );
  INVX1 U1847 ( .A(n1528), .Y(n5077) );
  INVX1 U1849 ( .A(n5080), .Y(n5078) );
  INVX1 U1851 ( .A(n5078), .Y(n5079) );
  AND2X1 U1853 ( .A(n11068), .B(n1489), .Y(n1527) );
  INVX1 U1855 ( .A(n1527), .Y(n5080) );
  INVX1 U1857 ( .A(n5083), .Y(n5081) );
  INVX1 U1859 ( .A(n5081), .Y(n5082) );
  AND2X1 U1861 ( .A(n11071), .B(n1489), .Y(n1526) );
  INVX1 U1863 ( .A(n1526), .Y(n5083) );
  INVX1 U1865 ( .A(n5086), .Y(n5084) );
  INVX1 U1867 ( .A(n5084), .Y(n5085) );
  AND2X1 U1869 ( .A(n11074), .B(n1489), .Y(n1525) );
  INVX1 U1871 ( .A(n1525), .Y(n5086) );
  INVX1 U1873 ( .A(n5089), .Y(n5087) );
  INVX1 U1875 ( .A(n5087), .Y(n5088) );
  AND2X1 U1877 ( .A(n11077), .B(n1489), .Y(n1524) );
  INVX1 U1879 ( .A(n1524), .Y(n5089) );
  INVX1 U1881 ( .A(n5092), .Y(n5090) );
  INVX1 U1883 ( .A(n5090), .Y(n5091) );
  AND2X1 U1885 ( .A(n11080), .B(n1489), .Y(n1523) );
  INVX1 U1887 ( .A(n1523), .Y(n5092) );
  INVX1 U1889 ( .A(n5095), .Y(n5093) );
  INVX1 U1891 ( .A(n5093), .Y(n5094) );
  AND2X1 U1893 ( .A(n11083), .B(n1489), .Y(n1522) );
  INVX1 U1895 ( .A(n1522), .Y(n5095) );
  INVX1 U1897 ( .A(n5098), .Y(n5096) );
  INVX1 U1899 ( .A(n5096), .Y(n5097) );
  AND2X1 U1901 ( .A(n11086), .B(n1489), .Y(n1521) );
  INVX1 U1903 ( .A(n1521), .Y(n5098) );
  INVX1 U1905 ( .A(n5101), .Y(n5099) );
  INVX1 U1907 ( .A(n5099), .Y(n5100) );
  AND2X1 U1909 ( .A(n11089), .B(n1489), .Y(n1520) );
  INVX1 U1911 ( .A(n1520), .Y(n5101) );
  INVX1 U1912 ( .A(n5104), .Y(n5102) );
  INVX1 U1914 ( .A(n5102), .Y(n5103) );
  AND2X1 U1916 ( .A(n11092), .B(n1489), .Y(n1519) );
  INVX1 U1918 ( .A(n1519), .Y(n5104) );
  INVX1 U1920 ( .A(n5107), .Y(n5105) );
  INVX1 U1922 ( .A(n5105), .Y(n5106) );
  AND2X1 U1924 ( .A(n11095), .B(n1489), .Y(n1518) );
  INVX1 U1926 ( .A(n1518), .Y(n5107) );
  INVX1 U1928 ( .A(n5110), .Y(n5108) );
  INVX1 U1930 ( .A(n5108), .Y(n5109) );
  AND2X1 U1932 ( .A(n11098), .B(n1489), .Y(n1517) );
  INVX1 U1934 ( .A(n1517), .Y(n5110) );
  INVX1 U1936 ( .A(n5113), .Y(n5111) );
  INVX1 U1938 ( .A(n5111), .Y(n5112) );
  AND2X1 U1940 ( .A(n11101), .B(n1489), .Y(n1516) );
  INVX1 U1942 ( .A(n1516), .Y(n5113) );
  INVX1 U1944 ( .A(n5116), .Y(n5114) );
  INVX1 U1946 ( .A(n5114), .Y(n5115) );
  AND2X1 U1948 ( .A(n11104), .B(n1489), .Y(n1515) );
  INVX1 U1950 ( .A(n1515), .Y(n5116) );
  INVX1 U1952 ( .A(n5119), .Y(n5117) );
  INVX1 U1954 ( .A(n5117), .Y(n5118) );
  AND2X1 U1956 ( .A(n11107), .B(n1489), .Y(n1514) );
  INVX1 U1958 ( .A(n1514), .Y(n5119) );
  INVX1 U1960 ( .A(n5122), .Y(n5120) );
  INVX1 U1962 ( .A(n5120), .Y(n5121) );
  AND2X1 U1964 ( .A(n11110), .B(n1489), .Y(n1513) );
  INVX1 U1966 ( .A(n1513), .Y(n5122) );
  INVX1 U1968 ( .A(n5125), .Y(n5123) );
  INVX1 U1970 ( .A(n5123), .Y(n5124) );
  AND2X1 U1972 ( .A(n11113), .B(n1489), .Y(n1512) );
  INVX1 U1974 ( .A(n1512), .Y(n5125) );
  INVX1 U1976 ( .A(n5128), .Y(n5126) );
  INVX1 U1978 ( .A(n5126), .Y(n5127) );
  AND2X1 U1980 ( .A(n11116), .B(n1489), .Y(n1511) );
  INVX1 U1982 ( .A(n1511), .Y(n5128) );
  INVX1 U1984 ( .A(n5131), .Y(n5129) );
  INVX1 U1986 ( .A(n5129), .Y(n5130) );
  AND2X1 U1988 ( .A(n11119), .B(n1489), .Y(n1510) );
  INVX1 U1990 ( .A(n1510), .Y(n5131) );
  INVX1 U1992 ( .A(n5134), .Y(n5132) );
  INVX1 U1994 ( .A(n5132), .Y(n5133) );
  AND2X1 U1996 ( .A(n11122), .B(n1489), .Y(n1509) );
  INVX1 U1997 ( .A(n1509), .Y(n5134) );
  INVX1 U1999 ( .A(n5137), .Y(n5135) );
  INVX1 U2001 ( .A(n5135), .Y(n5136) );
  AND2X1 U2003 ( .A(n11125), .B(n1489), .Y(n1508) );
  INVX1 U2005 ( .A(n1508), .Y(n5137) );
  INVX1 U2007 ( .A(n5140), .Y(n5138) );
  INVX1 U2009 ( .A(n5138), .Y(n5139) );
  AND2X1 U2011 ( .A(n11128), .B(n1489), .Y(n1507) );
  INVX1 U2013 ( .A(n1507), .Y(n5140) );
  INVX1 U2015 ( .A(n5143), .Y(n5141) );
  INVX1 U2017 ( .A(n5141), .Y(n5142) );
  AND2X1 U2019 ( .A(n11131), .B(n1489), .Y(n1506) );
  INVX1 U2021 ( .A(n1506), .Y(n5143) );
  INVX1 U2023 ( .A(n5146), .Y(n5144) );
  INVX1 U2025 ( .A(n5144), .Y(n5145) );
  AND2X1 U2027 ( .A(n11134), .B(n1489), .Y(n1505) );
  INVX1 U2029 ( .A(n1505), .Y(n5146) );
  INVX1 U2031 ( .A(n5149), .Y(n5147) );
  INVX1 U2033 ( .A(n5147), .Y(n5148) );
  AND2X1 U2035 ( .A(n11137), .B(n1489), .Y(n1504) );
  INVX1 U2037 ( .A(n1504), .Y(n5149) );
  INVX1 U2039 ( .A(n5152), .Y(n5150) );
  INVX1 U2041 ( .A(n5150), .Y(n5151) );
  AND2X1 U2043 ( .A(n11140), .B(n1489), .Y(n1503) );
  INVX1 U2045 ( .A(n1503), .Y(n5152) );
  INVX1 U2047 ( .A(n5155), .Y(n5153) );
  INVX1 U2049 ( .A(n5153), .Y(n5154) );
  AND2X1 U2051 ( .A(n11143), .B(n1489), .Y(n1502) );
  INVX1 U2053 ( .A(n1502), .Y(n5155) );
  INVX1 U2055 ( .A(n5158), .Y(n5156) );
  INVX1 U2057 ( .A(n5156), .Y(n5157) );
  AND2X1 U2059 ( .A(n11146), .B(n1489), .Y(n1501) );
  INVX1 U2061 ( .A(n1501), .Y(n5158) );
  INVX1 U2063 ( .A(n5161), .Y(n5159) );
  INVX1 U2065 ( .A(n5159), .Y(n5160) );
  AND2X1 U2067 ( .A(n11149), .B(n1489), .Y(n1500) );
  INVX1 U2069 ( .A(n1500), .Y(n5161) );
  INVX1 U2071 ( .A(n5164), .Y(n5162) );
  INVX1 U2073 ( .A(n5162), .Y(n5163) );
  AND2X1 U2075 ( .A(n11152), .B(n1489), .Y(n1499) );
  INVX1 U2077 ( .A(n1499), .Y(n5164) );
  INVX1 U2079 ( .A(n5167), .Y(n5165) );
  INVX1 U2081 ( .A(n5165), .Y(n5166) );
  AND2X1 U2082 ( .A(n11155), .B(n1489), .Y(n1498) );
  INVX1 U2084 ( .A(n1498), .Y(n5167) );
  INVX1 U2086 ( .A(n5170), .Y(n5168) );
  INVX1 U2088 ( .A(n5168), .Y(n5169) );
  AND2X1 U2090 ( .A(n11158), .B(n1489), .Y(n1497) );
  INVX1 U2092 ( .A(n1497), .Y(n5170) );
  INVX1 U2094 ( .A(n5173), .Y(n5171) );
  INVX1 U2096 ( .A(n5171), .Y(n5172) );
  AND2X1 U2098 ( .A(n11161), .B(n1489), .Y(n1496) );
  INVX1 U2100 ( .A(n1496), .Y(n5173) );
  INVX1 U2102 ( .A(n5176), .Y(n5174) );
  INVX1 U2104 ( .A(n5174), .Y(n5175) );
  AND2X1 U2106 ( .A(n11164), .B(n1489), .Y(n1495) );
  INVX1 U2108 ( .A(n1495), .Y(n5176) );
  INVX1 U2110 ( .A(n5179), .Y(n5177) );
  INVX1 U2112 ( .A(n5177), .Y(n5178) );
  AND2X1 U2114 ( .A(n11167), .B(n1489), .Y(n1494) );
  INVX1 U2116 ( .A(n1494), .Y(n5179) );
  INVX1 U2118 ( .A(n5182), .Y(n5180) );
  INVX1 U2120 ( .A(n5180), .Y(n5181) );
  AND2X1 U2122 ( .A(n11170), .B(n1489), .Y(n1493) );
  INVX1 U2124 ( .A(n1493), .Y(n5182) );
  INVX1 U2126 ( .A(n5185), .Y(n5183) );
  INVX1 U2128 ( .A(n5183), .Y(n5184) );
  AND2X1 U2130 ( .A(n11173), .B(n1489), .Y(n1492) );
  INVX1 U2132 ( .A(n1492), .Y(n5185) );
  INVX1 U2134 ( .A(n5188), .Y(n5186) );
  INVX1 U2136 ( .A(n5186), .Y(n5187) );
  AND2X1 U2138 ( .A(n11176), .B(n1489), .Y(n1491) );
  INVX1 U2140 ( .A(n1491), .Y(n5188) );
  INVX1 U2142 ( .A(n5191), .Y(n5189) );
  INVX1 U2144 ( .A(n5189), .Y(n5190) );
  AND2X1 U2146 ( .A(n11179), .B(n1489), .Y(n1490) );
  INVX1 U2148 ( .A(n1490), .Y(n5191) );
  INVX1 U2150 ( .A(n5194), .Y(n5192) );
  INVX1 U2152 ( .A(n5192), .Y(n5193) );
  AND2X1 U2154 ( .A(n9032), .B(n1445), .Y(n1487) );
  INVX1 U2156 ( .A(n1487), .Y(n5194) );
  INVX1 U2158 ( .A(n5197), .Y(n5195) );
  INVX1 U2160 ( .A(n5195), .Y(n5196) );
  AND2X1 U2162 ( .A(n9035), .B(n1445), .Y(n1486) );
  INVX1 U2164 ( .A(n1486), .Y(n5197) );
  INVX1 U2166 ( .A(n5200), .Y(n5198) );
  INVX1 U2167 ( .A(n5198), .Y(n5199) );
  AND2X1 U2168 ( .A(n9038), .B(n1445), .Y(n1485) );
  INVX1 U2172 ( .A(n1485), .Y(n5200) );
  INVX1 U2174 ( .A(n5203), .Y(n5201) );
  INVX1 U2176 ( .A(n5201), .Y(n5202) );
  AND2X1 U2178 ( .A(n9041), .B(n1445), .Y(n1484) );
  INVX1 U2180 ( .A(n1484), .Y(n5203) );
  INVX1 U2182 ( .A(n5206), .Y(n5204) );
  INVX1 U2184 ( .A(n5204), .Y(n5205) );
  AND2X1 U2186 ( .A(n9044), .B(n1445), .Y(n1483) );
  INVX1 U2188 ( .A(n1483), .Y(n5206) );
  INVX1 U2190 ( .A(n5209), .Y(n5207) );
  INVX1 U2192 ( .A(n5207), .Y(n5208) );
  AND2X1 U2194 ( .A(n9047), .B(n1445), .Y(n1482) );
  INVX1 U2196 ( .A(n1482), .Y(n5209) );
  INVX1 U2198 ( .A(n5212), .Y(n5210) );
  INVX1 U2200 ( .A(n5210), .Y(n5211) );
  AND2X1 U2202 ( .A(n9050), .B(n1445), .Y(n1481) );
  INVX1 U2204 ( .A(n1481), .Y(n5212) );
  INVX1 U2206 ( .A(n5215), .Y(n5213) );
  INVX1 U2208 ( .A(n5213), .Y(n5214) );
  AND2X1 U2210 ( .A(n9053), .B(n1445), .Y(n1480) );
  INVX1 U2212 ( .A(n1480), .Y(n5215) );
  INVX1 U2214 ( .A(n5218), .Y(n5216) );
  INVX1 U2216 ( .A(n5216), .Y(n5217) );
  AND2X1 U2218 ( .A(n9056), .B(n1445), .Y(n1479) );
  INVX1 U2220 ( .A(n1479), .Y(n5218) );
  INVX1 U2222 ( .A(n5221), .Y(n5219) );
  INVX1 U2224 ( .A(n5219), .Y(n5220) );
  AND2X1 U2226 ( .A(n9059), .B(n1445), .Y(n1478) );
  INVX1 U2228 ( .A(n1478), .Y(n5221) );
  INVX1 U2230 ( .A(n5224), .Y(n5222) );
  INVX1 U2232 ( .A(n5222), .Y(n5223) );
  AND2X1 U2234 ( .A(n9062), .B(n1445), .Y(n1477) );
  INVX1 U2236 ( .A(n1477), .Y(n5224) );
  INVX1 U2238 ( .A(n5227), .Y(n5225) );
  INVX1 U2240 ( .A(n5225), .Y(n5226) );
  AND2X1 U2242 ( .A(n9065), .B(n1445), .Y(n1476) );
  INVX1 U2244 ( .A(n1476), .Y(n5227) );
  INVX1 U2246 ( .A(n5230), .Y(n5228) );
  INVX1 U2248 ( .A(n5228), .Y(n5229) );
  AND2X1 U2250 ( .A(n9068), .B(n1445), .Y(n1475) );
  INVX1 U2252 ( .A(n1475), .Y(n5230) );
  INVX1 U2254 ( .A(n5233), .Y(n5231) );
  INVX1 U2255 ( .A(n5231), .Y(n5232) );
  AND2X1 U2258 ( .A(n9071), .B(n1445), .Y(n1474) );
  INVX1 U2260 ( .A(n1474), .Y(n5233) );
  INVX1 U2262 ( .A(n5236), .Y(n5234) );
  INVX1 U2264 ( .A(n5234), .Y(n5235) );
  AND2X1 U2266 ( .A(n9074), .B(n1445), .Y(n1473) );
  INVX1 U2268 ( .A(n1473), .Y(n5236) );
  INVX1 U2270 ( .A(n5239), .Y(n5237) );
  INVX1 U2272 ( .A(n5237), .Y(n5238) );
  AND2X1 U2274 ( .A(n9077), .B(n1445), .Y(n1472) );
  INVX1 U2276 ( .A(n1472), .Y(n5239) );
  INVX1 U2278 ( .A(n5242), .Y(n5240) );
  INVX1 U2280 ( .A(n5240), .Y(n5241) );
  AND2X1 U2282 ( .A(n9080), .B(n1445), .Y(n1471) );
  INVX1 U2284 ( .A(n1471), .Y(n5242) );
  INVX1 U2286 ( .A(n5245), .Y(n5243) );
  INVX1 U2288 ( .A(n5243), .Y(n5244) );
  AND2X1 U2290 ( .A(n9083), .B(n1445), .Y(n1470) );
  INVX1 U2292 ( .A(n1470), .Y(n5245) );
  INVX1 U2294 ( .A(n5248), .Y(n5246) );
  INVX1 U2296 ( .A(n5246), .Y(n5247) );
  AND2X1 U2298 ( .A(n9086), .B(n1445), .Y(n1469) );
  INVX1 U2300 ( .A(n1469), .Y(n5248) );
  INVX1 U2302 ( .A(n5251), .Y(n5249) );
  INVX1 U2304 ( .A(n5249), .Y(n5250) );
  AND2X1 U2306 ( .A(n9089), .B(n1445), .Y(n1468) );
  INVX1 U2308 ( .A(n1468), .Y(n5251) );
  INVX1 U2310 ( .A(n5254), .Y(n5252) );
  INVX1 U2312 ( .A(n5252), .Y(n5253) );
  AND2X1 U2314 ( .A(n9092), .B(n1445), .Y(n1467) );
  INVX1 U2316 ( .A(n1467), .Y(n5254) );
  INVX1 U2318 ( .A(n5257), .Y(n5255) );
  INVX1 U2320 ( .A(n5255), .Y(n5256) );
  AND2X1 U2322 ( .A(n9095), .B(n1445), .Y(n1466) );
  INVX1 U2324 ( .A(n1466), .Y(n5257) );
  INVX1 U2326 ( .A(n5260), .Y(n5258) );
  INVX1 U2328 ( .A(n5258), .Y(n5259) );
  AND2X1 U2330 ( .A(n9098), .B(n1445), .Y(n1465) );
  INVX1 U2332 ( .A(n1465), .Y(n5260) );
  INVX1 U2334 ( .A(n5263), .Y(n5261) );
  INVX1 U2336 ( .A(n5261), .Y(n5262) );
  AND2X1 U2338 ( .A(n9101), .B(n1445), .Y(n1464) );
  INVX1 U2340 ( .A(n1464), .Y(n5263) );
  INVX1 U2341 ( .A(n5266), .Y(n5264) );
  INVX1 U2344 ( .A(n5264), .Y(n5265) );
  AND2X1 U2346 ( .A(n9104), .B(n1445), .Y(n1463) );
  INVX1 U2348 ( .A(n1463), .Y(n5266) );
  INVX1 U2350 ( .A(n5269), .Y(n5267) );
  INVX1 U2352 ( .A(n5267), .Y(n5268) );
  AND2X1 U2354 ( .A(n9107), .B(n1445), .Y(n1462) );
  INVX1 U2356 ( .A(n1462), .Y(n5269) );
  INVX1 U2358 ( .A(n5272), .Y(n5270) );
  INVX1 U2360 ( .A(n5270), .Y(n5271) );
  AND2X1 U2362 ( .A(n9110), .B(n1445), .Y(n1461) );
  INVX1 U2364 ( .A(n1461), .Y(n5272) );
  INVX1 U2366 ( .A(n5275), .Y(n5273) );
  INVX1 U2368 ( .A(n5273), .Y(n5274) );
  AND2X1 U2370 ( .A(n9113), .B(n1445), .Y(n1460) );
  INVX1 U2372 ( .A(n1460), .Y(n5275) );
  INVX1 U2374 ( .A(n5278), .Y(n5276) );
  INVX1 U2376 ( .A(n5276), .Y(n5277) );
  AND2X1 U2378 ( .A(n9116), .B(n1445), .Y(n1459) );
  INVX1 U2380 ( .A(n1459), .Y(n5278) );
  INVX1 U2382 ( .A(n5281), .Y(n5279) );
  INVX1 U2384 ( .A(n5279), .Y(n5280) );
  AND2X1 U2386 ( .A(n9119), .B(n1445), .Y(n1458) );
  INVX1 U2388 ( .A(n1458), .Y(n5281) );
  INVX1 U2390 ( .A(n5284), .Y(n5282) );
  INVX1 U2392 ( .A(n5282), .Y(n5283) );
  AND2X1 U2394 ( .A(n9122), .B(n1445), .Y(n1457) );
  INVX1 U2396 ( .A(n1457), .Y(n5284) );
  INVX1 U2398 ( .A(n5287), .Y(n5285) );
  INVX1 U2400 ( .A(n5285), .Y(n5286) );
  AND2X1 U2402 ( .A(n9125), .B(n1445), .Y(n1456) );
  INVX1 U2404 ( .A(n1456), .Y(n5287) );
  INVX1 U2406 ( .A(n5290), .Y(n5288) );
  INVX1 U2408 ( .A(n5288), .Y(n5289) );
  AND2X1 U2410 ( .A(n9128), .B(n1445), .Y(n1455) );
  INVX1 U2412 ( .A(n1455), .Y(n5290) );
  INVX1 U2414 ( .A(n5293), .Y(n5291) );
  INVX1 U2416 ( .A(n5291), .Y(n5292) );
  AND2X1 U2418 ( .A(n9131), .B(n1445), .Y(n1454) );
  INVX1 U2420 ( .A(n1454), .Y(n5293) );
  INVX1 U2422 ( .A(n5296), .Y(n5294) );
  INVX1 U2424 ( .A(n5294), .Y(n5295) );
  AND2X1 U2426 ( .A(n9134), .B(n1445), .Y(n1453) );
  INVX1 U2427 ( .A(n1453), .Y(n5296) );
  INVX1 U2428 ( .A(n5299), .Y(n5297) );
  INVX1 U2430 ( .A(n5297), .Y(n5298) );
  AND2X1 U2432 ( .A(n9137), .B(n1445), .Y(n1452) );
  INVX1 U2434 ( .A(n1452), .Y(n5299) );
  INVX1 U2436 ( .A(n5302), .Y(n5300) );
  INVX1 U2438 ( .A(n5300), .Y(n5301) );
  AND2X1 U2440 ( .A(n9140), .B(n1445), .Y(n1451) );
  INVX1 U2442 ( .A(n1451), .Y(n5302) );
  INVX1 U2444 ( .A(n5305), .Y(n5303) );
  INVX1 U2446 ( .A(n5303), .Y(n5304) );
  AND2X1 U2448 ( .A(n9143), .B(n1445), .Y(n1450) );
  INVX1 U2450 ( .A(n1450), .Y(n5305) );
  INVX1 U2452 ( .A(n5308), .Y(n5306) );
  INVX1 U2454 ( .A(n5306), .Y(n5307) );
  AND2X1 U2456 ( .A(n9146), .B(n1445), .Y(n1449) );
  INVX1 U2458 ( .A(n1449), .Y(n5308) );
  INVX1 U2460 ( .A(n5311), .Y(n5309) );
  INVX1 U2462 ( .A(n5309), .Y(n5310) );
  AND2X1 U2464 ( .A(n9149), .B(n1445), .Y(n1448) );
  INVX1 U2466 ( .A(n1448), .Y(n5311) );
  INVX1 U2468 ( .A(n5314), .Y(n5312) );
  INVX1 U2470 ( .A(n5312), .Y(n5313) );
  AND2X1 U2472 ( .A(n9152), .B(n1445), .Y(n1447) );
  INVX1 U2474 ( .A(n1447), .Y(n5314) );
  INVX1 U2476 ( .A(n5317), .Y(n5315) );
  INVX1 U2478 ( .A(n5315), .Y(n5316) );
  AND2X1 U2480 ( .A(n9155), .B(n1445), .Y(n1446) );
  INVX1 U2482 ( .A(n1446), .Y(n5317) );
  INVX1 U2484 ( .A(n5320), .Y(n5318) );
  INVX1 U2486 ( .A(n5318), .Y(n5319) );
  AND2X1 U2488 ( .A(n11182), .B(n1402), .Y(n1444) );
  INVX1 U2490 ( .A(n1444), .Y(n5320) );
  INVX1 U2492 ( .A(n5323), .Y(n5321) );
  INVX1 U2494 ( .A(n5321), .Y(n5322) );
  AND2X1 U2496 ( .A(n11185), .B(n1402), .Y(n1443) );
  INVX1 U2498 ( .A(n1443), .Y(n5323) );
  INVX1 U2500 ( .A(n5326), .Y(n5324) );
  INVX1 U2502 ( .A(n5324), .Y(n5325) );
  AND2X1 U2504 ( .A(n11188), .B(n1402), .Y(n1442) );
  INVX1 U2506 ( .A(n1442), .Y(n5326) );
  INVX1 U2508 ( .A(n5329), .Y(n5327) );
  INVX1 U2510 ( .A(n5327), .Y(n5328) );
  AND2X1 U2512 ( .A(n11191), .B(n1402), .Y(n1441) );
  INVX1 U2513 ( .A(n1441), .Y(n5329) );
  INVX1 U2514 ( .A(n5332), .Y(n5330) );
  INVX1 U2516 ( .A(n5330), .Y(n5331) );
  AND2X1 U2518 ( .A(n11194), .B(n1402), .Y(n1440) );
  INVX1 U2520 ( .A(n1440), .Y(n5332) );
  INVX1 U2522 ( .A(n5335), .Y(n5333) );
  INVX1 U2524 ( .A(n5333), .Y(n5334) );
  AND2X1 U2526 ( .A(n11197), .B(n1402), .Y(n1439) );
  INVX1 U2528 ( .A(n1439), .Y(n5335) );
  INVX1 U2530 ( .A(n5338), .Y(n5336) );
  INVX1 U2532 ( .A(n5336), .Y(n5337) );
  AND2X1 U2534 ( .A(n11200), .B(n1402), .Y(n1438) );
  INVX1 U2536 ( .A(n1438), .Y(n5338) );
  INVX1 U2538 ( .A(n5341), .Y(n5339) );
  INVX1 U2540 ( .A(n5339), .Y(n5340) );
  AND2X1 U2542 ( .A(n11203), .B(n1402), .Y(n1437) );
  INVX1 U2544 ( .A(n1437), .Y(n5341) );
  INVX1 U2546 ( .A(n5344), .Y(n5342) );
  INVX1 U2548 ( .A(n5342), .Y(n5343) );
  AND2X1 U2550 ( .A(n11206), .B(n1402), .Y(n1436) );
  INVX1 U2552 ( .A(n1436), .Y(n5344) );
  INVX1 U2554 ( .A(n5347), .Y(n5345) );
  INVX1 U2556 ( .A(n5345), .Y(n5346) );
  AND2X1 U2558 ( .A(n11209), .B(n1402), .Y(n1435) );
  INVX1 U2560 ( .A(n1435), .Y(n5347) );
  INVX1 U2562 ( .A(n5350), .Y(n5348) );
  INVX1 U2564 ( .A(n5348), .Y(n5349) );
  AND2X1 U2566 ( .A(n11212), .B(n1402), .Y(n1434) );
  INVX1 U2568 ( .A(n1434), .Y(n5350) );
  INVX1 U2570 ( .A(n5353), .Y(n5351) );
  INVX1 U2572 ( .A(n5351), .Y(n5352) );
  AND2X1 U2574 ( .A(n11215), .B(n1402), .Y(n1433) );
  INVX1 U2576 ( .A(n1433), .Y(n5353) );
  INVX1 U2578 ( .A(n5356), .Y(n5354) );
  INVX1 U2580 ( .A(n5354), .Y(n5355) );
  AND2X1 U2582 ( .A(n11218), .B(n1402), .Y(n1432) );
  INVX1 U2584 ( .A(n1432), .Y(n5356) );
  INVX1 U2586 ( .A(n5359), .Y(n5357) );
  INVX1 U2588 ( .A(n5357), .Y(n5358) );
  AND2X1 U2590 ( .A(n11221), .B(n1402), .Y(n1431) );
  INVX1 U2592 ( .A(n1431), .Y(n5359) );
  INVX1 U2594 ( .A(n5362), .Y(n5360) );
  INVX1 U2596 ( .A(n5360), .Y(n5361) );
  AND2X1 U2598 ( .A(n11224), .B(n1402), .Y(n1430) );
  INVX1 U2599 ( .A(n1430), .Y(n5362) );
  INVX1 U2600 ( .A(n5365), .Y(n5363) );
  INVX1 U2602 ( .A(n5363), .Y(n5364) );
  AND2X1 U2604 ( .A(n11227), .B(n1402), .Y(n1429) );
  INVX1 U2606 ( .A(n1429), .Y(n5365) );
  INVX1 U2608 ( .A(n5368), .Y(n5366) );
  INVX1 U2610 ( .A(n5366), .Y(n5367) );
  AND2X1 U2612 ( .A(n11230), .B(n1402), .Y(n1428) );
  INVX1 U2614 ( .A(n1428), .Y(n5368) );
  INVX1 U2616 ( .A(n5371), .Y(n5369) );
  INVX1 U2618 ( .A(n5369), .Y(n5370) );
  AND2X1 U2620 ( .A(n11233), .B(n1402), .Y(n1427) );
  INVX1 U2622 ( .A(n1427), .Y(n5371) );
  INVX1 U2624 ( .A(n5374), .Y(n5372) );
  INVX1 U2626 ( .A(n5372), .Y(n5373) );
  AND2X1 U2628 ( .A(n11236), .B(n1402), .Y(n1426) );
  INVX1 U2630 ( .A(n1426), .Y(n5374) );
  INVX1 U2632 ( .A(n5377), .Y(n5375) );
  INVX1 U2634 ( .A(n5375), .Y(n5376) );
  AND2X1 U2636 ( .A(n11239), .B(n1402), .Y(n1425) );
  INVX1 U2638 ( .A(n1425), .Y(n5377) );
  INVX1 U2640 ( .A(n5380), .Y(n5378) );
  INVX1 U2642 ( .A(n5378), .Y(n5379) );
  AND2X1 U2644 ( .A(n11242), .B(n1402), .Y(n1424) );
  INVX1 U2646 ( .A(n1424), .Y(n5380) );
  INVX1 U2648 ( .A(n5383), .Y(n5381) );
  INVX1 U2650 ( .A(n5381), .Y(n5382) );
  AND2X1 U2652 ( .A(n11245), .B(n1402), .Y(n1423) );
  INVX1 U2654 ( .A(n1423), .Y(n5383) );
  INVX1 U2656 ( .A(n5386), .Y(n5384) );
  INVX1 U2658 ( .A(n5384), .Y(n5385) );
  AND2X1 U2660 ( .A(n11248), .B(n1402), .Y(n1422) );
  INVX1 U2662 ( .A(n1422), .Y(n5386) );
  INVX1 U2664 ( .A(n5389), .Y(n5387) );
  INVX1 U2666 ( .A(n5387), .Y(n5388) );
  AND2X1 U2668 ( .A(n11251), .B(n1402), .Y(n1421) );
  INVX1 U2670 ( .A(n1421), .Y(n5389) );
  INVX1 U2672 ( .A(n5392), .Y(n5390) );
  INVX1 U2674 ( .A(n5390), .Y(n5391) );
  AND2X1 U2676 ( .A(n11254), .B(n1402), .Y(n1420) );
  INVX1 U2678 ( .A(n1420), .Y(n5392) );
  INVX1 U2680 ( .A(n5395), .Y(n5393) );
  INVX1 U2682 ( .A(n5393), .Y(n5394) );
  AND2X1 U2684 ( .A(n11257), .B(n1402), .Y(n1419) );
  INVX1 U2685 ( .A(n1419), .Y(n5395) );
  INVX1 U2686 ( .A(n5398), .Y(n5396) );
  INVX1 U2688 ( .A(n5396), .Y(n5397) );
  AND2X1 U2690 ( .A(n11260), .B(n1402), .Y(n1418) );
  INVX1 U2692 ( .A(n1418), .Y(n5398) );
  INVX1 U2694 ( .A(n5401), .Y(n5399) );
  INVX1 U2696 ( .A(n5399), .Y(n5400) );
  AND2X1 U2698 ( .A(n11263), .B(n1402), .Y(n1417) );
  INVX1 U2700 ( .A(n1417), .Y(n5401) );
  INVX1 U2702 ( .A(n5404), .Y(n5402) );
  INVX1 U2704 ( .A(n5402), .Y(n5403) );
  AND2X1 U2706 ( .A(n11266), .B(n1402), .Y(n1416) );
  INVX1 U2708 ( .A(n1416), .Y(n5404) );
  INVX1 U2710 ( .A(n5407), .Y(n5405) );
  INVX1 U2712 ( .A(n5405), .Y(n5406) );
  AND2X1 U2714 ( .A(n11269), .B(n1402), .Y(n1415) );
  INVX1 U2716 ( .A(n1415), .Y(n5407) );
  INVX1 U2718 ( .A(n5410), .Y(n5408) );
  INVX1 U2720 ( .A(n5408), .Y(n5409) );
  AND2X1 U2722 ( .A(n11272), .B(n1402), .Y(n1414) );
  INVX1 U2724 ( .A(n1414), .Y(n5410) );
  INVX1 U2726 ( .A(n5413), .Y(n5411) );
  INVX1 U2728 ( .A(n5411), .Y(n5412) );
  AND2X1 U2730 ( .A(n11275), .B(n1402), .Y(n1413) );
  INVX1 U2732 ( .A(n1413), .Y(n5413) );
  INVX1 U2734 ( .A(n5416), .Y(n5414) );
  INVX1 U2736 ( .A(n5414), .Y(n5415) );
  AND2X1 U2738 ( .A(n11278), .B(n1402), .Y(n1412) );
  INVX1 U2740 ( .A(n1412), .Y(n5416) );
  INVX1 U2742 ( .A(n5419), .Y(n5417) );
  INVX1 U2744 ( .A(n5417), .Y(n5418) );
  AND2X1 U2746 ( .A(n11281), .B(n1402), .Y(n1411) );
  INVX1 U2748 ( .A(n1411), .Y(n5419) );
  INVX1 U2750 ( .A(n5422), .Y(n5420) );
  INVX1 U2752 ( .A(n5420), .Y(n5421) );
  AND2X1 U2754 ( .A(n11284), .B(n1402), .Y(n1410) );
  INVX1 U2756 ( .A(n1410), .Y(n5422) );
  INVX1 U2758 ( .A(n5425), .Y(n5423) );
  INVX1 U2760 ( .A(n5423), .Y(n5424) );
  AND2X1 U2762 ( .A(n11287), .B(n1402), .Y(n1409) );
  INVX1 U2764 ( .A(n1409), .Y(n5425) );
  INVX1 U2766 ( .A(n5428), .Y(n5426) );
  INVX1 U2768 ( .A(n5426), .Y(n5427) );
  AND2X1 U2770 ( .A(n11290), .B(n1402), .Y(n1408) );
  INVX1 U2771 ( .A(n1408), .Y(n5428) );
  INVX1 U2774 ( .A(n5431), .Y(n5429) );
  INVX1 U2777 ( .A(n5429), .Y(n5430) );
  AND2X1 U2780 ( .A(n11293), .B(n1402), .Y(n1407) );
  INVX1 U2783 ( .A(n1407), .Y(n5431) );
  INVX1 U2786 ( .A(n5434), .Y(n5432) );
  INVX1 U2789 ( .A(n5432), .Y(n5433) );
  AND2X1 U2792 ( .A(n11296), .B(n1402), .Y(n1406) );
  INVX1 U2795 ( .A(n1406), .Y(n5434) );
  INVX1 U2798 ( .A(n5437), .Y(n5435) );
  INVX1 U2801 ( .A(n5435), .Y(n5436) );
  AND2X1 U2804 ( .A(n11299), .B(n1402), .Y(n1405) );
  INVX1 U2807 ( .A(n1405), .Y(n5437) );
  INVX1 U2810 ( .A(n5440), .Y(n5438) );
  INVX1 U2813 ( .A(n5438), .Y(n5439) );
  AND2X1 U2816 ( .A(n11302), .B(n1402), .Y(n1404) );
  INVX1 U2819 ( .A(n1404), .Y(n5440) );
  INVX1 U2822 ( .A(n5443), .Y(n5441) );
  INVX1 U2825 ( .A(n5441), .Y(n5442) );
  AND2X1 U2828 ( .A(n11305), .B(n1402), .Y(n1403) );
  INVX1 U2831 ( .A(n1403), .Y(n5443) );
  INVX1 U2834 ( .A(n5446), .Y(n5444) );
  INVX1 U2837 ( .A(n5444), .Y(n5445) );
  AND2X1 U2840 ( .A(n9158), .B(n1358), .Y(n1400) );
  INVX1 U2843 ( .A(n1400), .Y(n5446) );
  INVX1 U2846 ( .A(n5449), .Y(n5447) );
  INVX1 U2849 ( .A(n5447), .Y(n5448) );
  AND2X1 U2852 ( .A(n9161), .B(n1358), .Y(n1399) );
  INVX1 U2855 ( .A(n1399), .Y(n5449) );
  INVX1 U2858 ( .A(n5452), .Y(n5450) );
  INVX1 U2861 ( .A(n5450), .Y(n5451) );
  AND2X1 U2864 ( .A(n9164), .B(n1358), .Y(n1398) );
  INVX1 U2867 ( .A(n1398), .Y(n5452) );
  INVX1 U2870 ( .A(n5455), .Y(n5453) );
  INVX1 U2873 ( .A(n5453), .Y(n5454) );
  AND2X1 U2876 ( .A(n9167), .B(n1358), .Y(n1397) );
  INVX1 U2879 ( .A(n1397), .Y(n5455) );
  INVX1 U2882 ( .A(n5458), .Y(n5456) );
  INVX1 U2885 ( .A(n5456), .Y(n5457) );
  AND2X1 U2888 ( .A(n9170), .B(n1358), .Y(n1396) );
  INVX1 U2891 ( .A(n1396), .Y(n5458) );
  INVX1 U2894 ( .A(n5461), .Y(n5459) );
  INVX1 U2897 ( .A(n5459), .Y(n5460) );
  AND2X1 U2898 ( .A(n9173), .B(n1358), .Y(n1395) );
  INVX1 U2901 ( .A(n1395), .Y(n5461) );
  INVX1 U2903 ( .A(n5464), .Y(n5462) );
  INVX1 U2906 ( .A(n5462), .Y(n5463) );
  AND2X1 U2907 ( .A(n9176), .B(n1358), .Y(n1394) );
  INVX1 U2909 ( .A(n1394), .Y(n5464) );
  INVX1 U2919 ( .A(n5467), .Y(n5465) );
  INVX1 U2920 ( .A(n5465), .Y(n5466) );
  AND2X1 U2921 ( .A(n9179), .B(n1358), .Y(n1393) );
  INVX1 U2923 ( .A(n1393), .Y(n5467) );
  INVX1 U2931 ( .A(n5470), .Y(n5468) );
  INVX1 U2932 ( .A(n5468), .Y(n5469) );
  AND2X1 U2934 ( .A(n9182), .B(n1358), .Y(n1392) );
  INVX1 U4377 ( .A(n1392), .Y(n5470) );
  INVX1 U4378 ( .A(n5473), .Y(n5471) );
  INVX1 U4379 ( .A(n5471), .Y(n5472) );
  AND2X1 U4380 ( .A(n9185), .B(n1358), .Y(n1391) );
  INVX1 U4381 ( .A(n1391), .Y(n5473) );
  INVX1 U4382 ( .A(n5476), .Y(n5474) );
  INVX1 U4383 ( .A(n5474), .Y(n5475) );
  AND2X1 U4384 ( .A(n9188), .B(n1358), .Y(n1390) );
  INVX1 U4385 ( .A(n1390), .Y(n5476) );
  INVX1 U4386 ( .A(n5479), .Y(n5477) );
  INVX1 U4387 ( .A(n5477), .Y(n5478) );
  AND2X1 U4388 ( .A(n9191), .B(n1358), .Y(n1389) );
  INVX1 U4389 ( .A(n1389), .Y(n5479) );
  INVX1 U4390 ( .A(n5482), .Y(n5480) );
  INVX1 U4391 ( .A(n5480), .Y(n5481) );
  AND2X1 U4392 ( .A(n9194), .B(n1358), .Y(n1388) );
  INVX1 U4393 ( .A(n1388), .Y(n5482) );
  INVX1 U4394 ( .A(n5485), .Y(n5483) );
  INVX1 U4395 ( .A(n5483), .Y(n5484) );
  AND2X1 U4396 ( .A(n9197), .B(n1358), .Y(n1387) );
  INVX1 U4397 ( .A(n1387), .Y(n5485) );
  INVX1 U4398 ( .A(n5488), .Y(n5486) );
  INVX1 U4399 ( .A(n5486), .Y(n5487) );
  AND2X1 U4400 ( .A(n9200), .B(n1358), .Y(n1386) );
  INVX1 U4401 ( .A(n1386), .Y(n5488) );
  INVX1 U4402 ( .A(n5491), .Y(n5489) );
  INVX1 U4403 ( .A(n5489), .Y(n5490) );
  AND2X1 U4404 ( .A(n9203), .B(n1358), .Y(n1385) );
  INVX1 U4405 ( .A(n1385), .Y(n5491) );
  INVX1 U4406 ( .A(n5494), .Y(n5492) );
  INVX1 U4407 ( .A(n5492), .Y(n5493) );
  AND2X1 U4408 ( .A(n9206), .B(n1358), .Y(n1384) );
  INVX1 U4409 ( .A(n1384), .Y(n5494) );
  INVX1 U4410 ( .A(n5497), .Y(n5495) );
  INVX1 U4411 ( .A(n5495), .Y(n5496) );
  AND2X1 U4412 ( .A(n9209), .B(n1358), .Y(n1383) );
  INVX1 U4413 ( .A(n1383), .Y(n5497) );
  INVX1 U4414 ( .A(n5500), .Y(n5498) );
  INVX1 U4415 ( .A(n5498), .Y(n5499) );
  AND2X1 U4416 ( .A(n9212), .B(n1358), .Y(n1382) );
  INVX1 U4417 ( .A(n1382), .Y(n5500) );
  INVX1 U4418 ( .A(n5503), .Y(n5501) );
  INVX1 U4419 ( .A(n5501), .Y(n5502) );
  AND2X1 U4420 ( .A(n9215), .B(n1358), .Y(n1381) );
  INVX1 U4421 ( .A(n1381), .Y(n5503) );
  INVX1 U4422 ( .A(n5506), .Y(n5504) );
  INVX1 U4423 ( .A(n5504), .Y(n5505) );
  AND2X1 U4424 ( .A(n9218), .B(n1358), .Y(n1380) );
  INVX1 U4425 ( .A(n1380), .Y(n5506) );
  INVX1 U4426 ( .A(n5509), .Y(n5507) );
  INVX1 U4427 ( .A(n5507), .Y(n5508) );
  AND2X1 U4428 ( .A(n9221), .B(n1358), .Y(n1379) );
  INVX1 U4429 ( .A(n1379), .Y(n5509) );
  INVX1 U4430 ( .A(n5512), .Y(n5510) );
  INVX1 U4431 ( .A(n5510), .Y(n5511) );
  AND2X1 U4432 ( .A(n9224), .B(n1358), .Y(n1378) );
  INVX1 U4433 ( .A(n1378), .Y(n5512) );
  INVX1 U4434 ( .A(n5515), .Y(n5513) );
  INVX1 U4435 ( .A(n5513), .Y(n5514) );
  AND2X1 U4436 ( .A(n9227), .B(n1358), .Y(n1377) );
  INVX1 U4437 ( .A(n1377), .Y(n5515) );
  INVX1 U4438 ( .A(n5518), .Y(n5516) );
  INVX1 U4439 ( .A(n5516), .Y(n5517) );
  AND2X1 U4440 ( .A(n9230), .B(n1358), .Y(n1376) );
  INVX1 U4441 ( .A(n1376), .Y(n5518) );
  INVX1 U4442 ( .A(n5521), .Y(n5519) );
  INVX1 U4443 ( .A(n5519), .Y(n5520) );
  AND2X1 U4444 ( .A(n9233), .B(n1358), .Y(n1375) );
  INVX1 U4445 ( .A(n1375), .Y(n5521) );
  INVX1 U4446 ( .A(n5524), .Y(n5522) );
  INVX1 U4447 ( .A(n5522), .Y(n5523) );
  AND2X1 U4448 ( .A(n9236), .B(n1358), .Y(n1374) );
  INVX1 U4449 ( .A(n1374), .Y(n5524) );
  INVX1 U4450 ( .A(n5527), .Y(n5525) );
  INVX1 U4451 ( .A(n5525), .Y(n5526) );
  AND2X1 U4452 ( .A(n9239), .B(n1358), .Y(n1373) );
  INVX1 U4453 ( .A(n1373), .Y(n5527) );
  INVX1 U4454 ( .A(n5530), .Y(n5528) );
  INVX1 U4455 ( .A(n5528), .Y(n5529) );
  AND2X1 U4456 ( .A(n9242), .B(n1358), .Y(n1372) );
  INVX1 U4457 ( .A(n1372), .Y(n5530) );
  INVX1 U4458 ( .A(n5533), .Y(n5531) );
  INVX1 U4459 ( .A(n5531), .Y(n5532) );
  AND2X1 U4460 ( .A(n9245), .B(n1358), .Y(n1371) );
  INVX1 U4461 ( .A(n1371), .Y(n5533) );
  INVX1 U4462 ( .A(n5536), .Y(n5534) );
  INVX1 U4463 ( .A(n5534), .Y(n5535) );
  AND2X1 U4464 ( .A(n9248), .B(n1358), .Y(n1370) );
  INVX1 U4465 ( .A(n1370), .Y(n5536) );
  INVX1 U4466 ( .A(n5539), .Y(n5537) );
  INVX1 U4467 ( .A(n5537), .Y(n5538) );
  AND2X1 U4468 ( .A(n9251), .B(n1358), .Y(n1369) );
  INVX1 U4469 ( .A(n1369), .Y(n5539) );
  INVX1 U4470 ( .A(n5542), .Y(n5540) );
  INVX1 U4471 ( .A(n5540), .Y(n5541) );
  AND2X1 U4472 ( .A(n9254), .B(n1358), .Y(n1368) );
  INVX1 U4473 ( .A(n1368), .Y(n5542) );
  INVX1 U4474 ( .A(n5545), .Y(n5543) );
  INVX1 U4475 ( .A(n5543), .Y(n5544) );
  AND2X1 U4476 ( .A(n9257), .B(n1358), .Y(n1367) );
  INVX1 U4477 ( .A(n1367), .Y(n5545) );
  INVX1 U4478 ( .A(n5548), .Y(n5546) );
  INVX1 U4479 ( .A(n5546), .Y(n5547) );
  AND2X1 U4480 ( .A(n9260), .B(n1358), .Y(n1366) );
  INVX1 U4481 ( .A(n1366), .Y(n5548) );
  INVX1 U4482 ( .A(n5551), .Y(n5549) );
  INVX1 U4483 ( .A(n5549), .Y(n5550) );
  AND2X1 U4484 ( .A(n9263), .B(n1358), .Y(n1365) );
  INVX1 U4485 ( .A(n1365), .Y(n5551) );
  INVX1 U4486 ( .A(n5554), .Y(n5552) );
  INVX1 U4487 ( .A(n5552), .Y(n5553) );
  AND2X1 U4488 ( .A(n9266), .B(n1358), .Y(n1364) );
  INVX1 U4489 ( .A(n1364), .Y(n5554) );
  INVX1 U4490 ( .A(n5557), .Y(n5555) );
  INVX1 U4491 ( .A(n5555), .Y(n5556) );
  AND2X1 U4492 ( .A(n9269), .B(n1358), .Y(n1363) );
  INVX1 U4493 ( .A(n1363), .Y(n5557) );
  INVX1 U4494 ( .A(n5560), .Y(n5558) );
  INVX1 U4495 ( .A(n5558), .Y(n5559) );
  AND2X1 U4496 ( .A(n9272), .B(n1358), .Y(n1362) );
  INVX1 U4497 ( .A(n1362), .Y(n5560) );
  INVX1 U4498 ( .A(n5563), .Y(n5561) );
  INVX1 U4499 ( .A(n5561), .Y(n5562) );
  AND2X1 U4500 ( .A(n9275), .B(n1358), .Y(n1361) );
  INVX1 U4501 ( .A(n1361), .Y(n5563) );
  INVX1 U4502 ( .A(n5566), .Y(n5564) );
  INVX1 U4503 ( .A(n5564), .Y(n5565) );
  AND2X1 U4504 ( .A(n9278), .B(n1358), .Y(n1360) );
  INVX1 U4505 ( .A(n1360), .Y(n5566) );
  INVX1 U4506 ( .A(n5569), .Y(n5567) );
  INVX1 U4507 ( .A(n5567), .Y(n5568) );
  AND2X1 U4508 ( .A(n9281), .B(n1358), .Y(n1359) );
  INVX1 U4509 ( .A(n1359), .Y(n5569) );
  INVX1 U4510 ( .A(n5572), .Y(n5570) );
  INVX1 U4511 ( .A(n5570), .Y(n5571) );
  AND2X1 U4512 ( .A(n11308), .B(n1314), .Y(n1356) );
  INVX1 U4513 ( .A(n1356), .Y(n5572) );
  INVX1 U4514 ( .A(n5575), .Y(n5573) );
  INVX1 U4515 ( .A(n5573), .Y(n5574) );
  AND2X1 U4516 ( .A(n11311), .B(n1314), .Y(n1355) );
  INVX1 U4517 ( .A(n1355), .Y(n5575) );
  INVX1 U4518 ( .A(n5578), .Y(n5576) );
  INVX1 U4519 ( .A(n5576), .Y(n5577) );
  AND2X1 U4520 ( .A(n11314), .B(n1314), .Y(n1354) );
  INVX1 U4521 ( .A(n1354), .Y(n5578) );
  INVX1 U4522 ( .A(n5581), .Y(n5579) );
  INVX1 U4523 ( .A(n5579), .Y(n5580) );
  AND2X1 U4524 ( .A(n11317), .B(n1314), .Y(n1353) );
  INVX1 U4525 ( .A(n1353), .Y(n5581) );
  INVX1 U4526 ( .A(n5584), .Y(n5582) );
  INVX1 U4527 ( .A(n5582), .Y(n5583) );
  AND2X1 U4528 ( .A(n11320), .B(n1314), .Y(n1352) );
  INVX1 U4529 ( .A(n1352), .Y(n5584) );
  INVX1 U4530 ( .A(n5587), .Y(n5585) );
  INVX1 U4531 ( .A(n5585), .Y(n5586) );
  AND2X1 U4532 ( .A(n11323), .B(n1314), .Y(n1351) );
  INVX1 U4533 ( .A(n1351), .Y(n5587) );
  INVX1 U4534 ( .A(n5590), .Y(n5588) );
  INVX1 U4535 ( .A(n5588), .Y(n5589) );
  AND2X1 U4536 ( .A(n11326), .B(n1314), .Y(n1350) );
  INVX1 U4537 ( .A(n1350), .Y(n5590) );
  INVX1 U4538 ( .A(n5593), .Y(n5591) );
  INVX1 U4539 ( .A(n5591), .Y(n5592) );
  AND2X1 U4540 ( .A(n11329), .B(n1314), .Y(n1349) );
  INVX1 U4541 ( .A(n1349), .Y(n5593) );
  INVX1 U4542 ( .A(n5596), .Y(n5594) );
  INVX1 U4543 ( .A(n5594), .Y(n5595) );
  AND2X1 U4544 ( .A(n11332), .B(n1314), .Y(n1348) );
  INVX1 U4545 ( .A(n1348), .Y(n5596) );
  INVX1 U4546 ( .A(n5599), .Y(n5597) );
  INVX1 U4547 ( .A(n5597), .Y(n5598) );
  AND2X1 U4548 ( .A(n11335), .B(n1314), .Y(n1347) );
  INVX1 U4549 ( .A(n1347), .Y(n5599) );
  INVX1 U4550 ( .A(n5602), .Y(n5600) );
  INVX1 U4551 ( .A(n5600), .Y(n5601) );
  AND2X1 U4552 ( .A(n11338), .B(n1314), .Y(n1346) );
  INVX1 U4553 ( .A(n1346), .Y(n5602) );
  INVX1 U4554 ( .A(n5605), .Y(n5603) );
  INVX1 U4555 ( .A(n5603), .Y(n5604) );
  AND2X1 U4556 ( .A(n11341), .B(n1314), .Y(n1345) );
  INVX1 U4557 ( .A(n1345), .Y(n5605) );
  INVX1 U4558 ( .A(n5608), .Y(n5606) );
  INVX1 U4559 ( .A(n5606), .Y(n5607) );
  AND2X1 U4560 ( .A(n11344), .B(n1314), .Y(n1344) );
  INVX1 U4561 ( .A(n1344), .Y(n5608) );
  INVX1 U4562 ( .A(n5611), .Y(n5609) );
  INVX1 U4563 ( .A(n5609), .Y(n5610) );
  AND2X1 U4564 ( .A(n11347), .B(n1314), .Y(n1343) );
  INVX1 U4565 ( .A(n1343), .Y(n5611) );
  INVX1 U4566 ( .A(n5614), .Y(n5612) );
  INVX1 U4567 ( .A(n5612), .Y(n5613) );
  AND2X1 U4568 ( .A(n11350), .B(n1314), .Y(n1342) );
  INVX1 U4569 ( .A(n1342), .Y(n5614) );
  INVX1 U4570 ( .A(n5617), .Y(n5615) );
  INVX1 U4571 ( .A(n5615), .Y(n5616) );
  AND2X1 U4572 ( .A(n11353), .B(n1314), .Y(n1341) );
  INVX1 U4573 ( .A(n1341), .Y(n5617) );
  INVX1 U4574 ( .A(n5620), .Y(n5618) );
  INVX1 U4575 ( .A(n5618), .Y(n5619) );
  AND2X1 U4576 ( .A(n11356), .B(n1314), .Y(n1340) );
  INVX1 U4577 ( .A(n1340), .Y(n5620) );
  INVX1 U4578 ( .A(n5623), .Y(n5621) );
  INVX1 U4579 ( .A(n5621), .Y(n5622) );
  AND2X1 U4580 ( .A(n11359), .B(n1314), .Y(n1339) );
  INVX1 U4581 ( .A(n1339), .Y(n5623) );
  INVX1 U4582 ( .A(n5626), .Y(n5624) );
  INVX1 U4583 ( .A(n5624), .Y(n5625) );
  AND2X1 U4584 ( .A(n11362), .B(n1314), .Y(n1338) );
  INVX1 U4585 ( .A(n1338), .Y(n5626) );
  INVX1 U4586 ( .A(n5629), .Y(n5627) );
  INVX1 U4587 ( .A(n5627), .Y(n5628) );
  AND2X1 U4588 ( .A(n11365), .B(n1314), .Y(n1337) );
  INVX1 U4589 ( .A(n1337), .Y(n5629) );
  INVX1 U4590 ( .A(n5632), .Y(n5630) );
  INVX1 U4591 ( .A(n5630), .Y(n5631) );
  AND2X1 U4592 ( .A(n11368), .B(n1314), .Y(n1336) );
  INVX1 U4593 ( .A(n1336), .Y(n5632) );
  INVX1 U4594 ( .A(n5635), .Y(n5633) );
  INVX1 U4595 ( .A(n5633), .Y(n5634) );
  AND2X1 U4596 ( .A(n11371), .B(n1314), .Y(n1335) );
  INVX1 U4597 ( .A(n1335), .Y(n5635) );
  INVX1 U4598 ( .A(n5638), .Y(n5636) );
  INVX1 U4599 ( .A(n5636), .Y(n5637) );
  AND2X1 U4600 ( .A(n11374), .B(n1314), .Y(n1334) );
  INVX1 U4601 ( .A(n1334), .Y(n5638) );
  INVX1 U4602 ( .A(n5641), .Y(n5639) );
  INVX1 U4603 ( .A(n5639), .Y(n5640) );
  AND2X1 U4604 ( .A(n11377), .B(n1314), .Y(n1333) );
  INVX1 U4605 ( .A(n1333), .Y(n5641) );
  INVX1 U4606 ( .A(n5644), .Y(n5642) );
  INVX1 U4607 ( .A(n5642), .Y(n5643) );
  AND2X1 U4608 ( .A(n11380), .B(n1314), .Y(n1332) );
  INVX1 U4609 ( .A(n1332), .Y(n5644) );
  INVX1 U4610 ( .A(n5647), .Y(n5645) );
  INVX1 U4611 ( .A(n5645), .Y(n5646) );
  AND2X1 U4612 ( .A(n11383), .B(n1314), .Y(n1331) );
  INVX1 U4613 ( .A(n1331), .Y(n5647) );
  INVX1 U4614 ( .A(n5650), .Y(n5648) );
  INVX1 U4615 ( .A(n5648), .Y(n5649) );
  AND2X1 U4616 ( .A(n11386), .B(n1314), .Y(n1330) );
  INVX1 U4617 ( .A(n1330), .Y(n5650) );
  INVX1 U4618 ( .A(n5653), .Y(n5651) );
  INVX1 U4619 ( .A(n5651), .Y(n5652) );
  AND2X1 U4620 ( .A(n11389), .B(n1314), .Y(n1329) );
  INVX1 U4621 ( .A(n1329), .Y(n5653) );
  INVX1 U4622 ( .A(n5656), .Y(n5654) );
  INVX1 U4623 ( .A(n5654), .Y(n5655) );
  AND2X1 U4624 ( .A(n11392), .B(n1314), .Y(n1328) );
  INVX1 U4625 ( .A(n1328), .Y(n5656) );
  INVX1 U4626 ( .A(n5659), .Y(n5657) );
  INVX1 U4627 ( .A(n5657), .Y(n5658) );
  AND2X1 U4628 ( .A(n11395), .B(n1314), .Y(n1327) );
  INVX1 U4629 ( .A(n1327), .Y(n5659) );
  INVX1 U4630 ( .A(n5662), .Y(n5660) );
  INVX1 U4631 ( .A(n5660), .Y(n5661) );
  AND2X1 U4632 ( .A(n11398), .B(n1314), .Y(n1326) );
  INVX1 U4633 ( .A(n1326), .Y(n5662) );
  INVX1 U4634 ( .A(n5665), .Y(n5663) );
  INVX1 U4635 ( .A(n5663), .Y(n5664) );
  AND2X1 U4636 ( .A(n11401), .B(n1314), .Y(n1325) );
  INVX1 U4637 ( .A(n1325), .Y(n5665) );
  INVX1 U4638 ( .A(n5668), .Y(n5666) );
  INVX1 U4639 ( .A(n5666), .Y(n5667) );
  AND2X1 U4640 ( .A(n11404), .B(n1314), .Y(n1324) );
  INVX1 U4641 ( .A(n1324), .Y(n5668) );
  INVX1 U4642 ( .A(n5671), .Y(n5669) );
  INVX1 U4643 ( .A(n5669), .Y(n5670) );
  AND2X1 U4644 ( .A(n11407), .B(n1314), .Y(n1323) );
  INVX1 U4645 ( .A(n1323), .Y(n5671) );
  INVX1 U4646 ( .A(n5674), .Y(n5672) );
  INVX1 U4647 ( .A(n5672), .Y(n5673) );
  AND2X1 U4648 ( .A(n11410), .B(n1314), .Y(n1322) );
  INVX1 U4649 ( .A(n1322), .Y(n5674) );
  INVX1 U4650 ( .A(n5677), .Y(n5675) );
  INVX1 U4651 ( .A(n5675), .Y(n5676) );
  AND2X1 U4652 ( .A(n11413), .B(n1314), .Y(n1321) );
  INVX1 U4653 ( .A(n1321), .Y(n5677) );
  INVX1 U4654 ( .A(n5680), .Y(n5678) );
  INVX1 U4655 ( .A(n5678), .Y(n5679) );
  AND2X1 U4656 ( .A(n11416), .B(n1314), .Y(n1320) );
  INVX1 U4657 ( .A(n1320), .Y(n5680) );
  INVX1 U4658 ( .A(n5683), .Y(n5681) );
  INVX1 U4659 ( .A(n5681), .Y(n5682) );
  AND2X1 U4660 ( .A(n11419), .B(n1314), .Y(n1319) );
  INVX1 U4661 ( .A(n1319), .Y(n5683) );
  INVX1 U4662 ( .A(n5686), .Y(n5684) );
  INVX1 U4663 ( .A(n5684), .Y(n5685) );
  AND2X1 U4664 ( .A(n11422), .B(n1314), .Y(n1318) );
  INVX1 U4665 ( .A(n1318), .Y(n5686) );
  INVX1 U4666 ( .A(n5689), .Y(n5687) );
  INVX1 U4667 ( .A(n5687), .Y(n5688) );
  AND2X1 U4668 ( .A(n11425), .B(n1314), .Y(n1317) );
  INVX1 U4669 ( .A(n1317), .Y(n5689) );
  INVX1 U4670 ( .A(n5692), .Y(n5690) );
  INVX1 U4671 ( .A(n5690), .Y(n5691) );
  AND2X1 U4672 ( .A(n11428), .B(n1314), .Y(n1316) );
  INVX1 U4673 ( .A(n1316), .Y(n5692) );
  INVX1 U4674 ( .A(n5695), .Y(n5693) );
  INVX1 U4675 ( .A(n5693), .Y(n5694) );
  AND2X1 U4676 ( .A(n11431), .B(n1314), .Y(n1315) );
  INVX1 U4677 ( .A(n1315), .Y(n5695) );
  INVX1 U4678 ( .A(n5698), .Y(n5696) );
  INVX1 U4679 ( .A(n5696), .Y(n5697) );
  AND2X1 U4680 ( .A(n9284), .B(n1271), .Y(n1313) );
  INVX1 U4681 ( .A(n1313), .Y(n5698) );
  INVX1 U4682 ( .A(n5701), .Y(n5699) );
  INVX1 U4683 ( .A(n5699), .Y(n5700) );
  AND2X1 U4684 ( .A(n9287), .B(n1271), .Y(n1312) );
  INVX1 U4685 ( .A(n1312), .Y(n5701) );
  INVX1 U4686 ( .A(n5704), .Y(n5702) );
  INVX1 U4687 ( .A(n5702), .Y(n5703) );
  AND2X1 U4688 ( .A(n9290), .B(n1271), .Y(n1311) );
  INVX1 U4689 ( .A(n1311), .Y(n5704) );
  INVX1 U4690 ( .A(n5707), .Y(n5705) );
  INVX1 U4691 ( .A(n5705), .Y(n5706) );
  AND2X1 U4692 ( .A(n9293), .B(n1271), .Y(n1310) );
  INVX1 U4693 ( .A(n1310), .Y(n5707) );
  INVX1 U4694 ( .A(n5710), .Y(n5708) );
  INVX1 U4695 ( .A(n5708), .Y(n5709) );
  AND2X1 U4696 ( .A(n9296), .B(n1271), .Y(n1309) );
  INVX1 U4697 ( .A(n1309), .Y(n5710) );
  INVX1 U4698 ( .A(n5713), .Y(n5711) );
  INVX1 U4699 ( .A(n5711), .Y(n5712) );
  AND2X1 U4700 ( .A(n9299), .B(n1271), .Y(n1308) );
  INVX1 U4701 ( .A(n1308), .Y(n5713) );
  INVX1 U4702 ( .A(n5716), .Y(n5714) );
  INVX1 U4703 ( .A(n5714), .Y(n5715) );
  AND2X1 U4704 ( .A(n9302), .B(n1271), .Y(n1307) );
  INVX1 U4705 ( .A(n1307), .Y(n5716) );
  INVX1 U4706 ( .A(n5719), .Y(n5717) );
  INVX1 U4707 ( .A(n5717), .Y(n5718) );
  AND2X1 U4708 ( .A(n9305), .B(n1271), .Y(n1306) );
  INVX1 U4709 ( .A(n1306), .Y(n5719) );
  INVX1 U4710 ( .A(n5722), .Y(n5720) );
  INVX1 U4711 ( .A(n5720), .Y(n5721) );
  AND2X1 U4712 ( .A(n9308), .B(n1271), .Y(n1305) );
  INVX1 U4713 ( .A(n1305), .Y(n5722) );
  INVX1 U4714 ( .A(n5725), .Y(n5723) );
  INVX1 U4715 ( .A(n5723), .Y(n5724) );
  AND2X1 U4716 ( .A(n9311), .B(n1271), .Y(n1304) );
  INVX1 U4717 ( .A(n1304), .Y(n5725) );
  INVX1 U4718 ( .A(n5728), .Y(n5726) );
  INVX1 U4719 ( .A(n5726), .Y(n5727) );
  AND2X1 U4720 ( .A(n9314), .B(n1271), .Y(n1303) );
  INVX1 U4721 ( .A(n1303), .Y(n5728) );
  INVX1 U4722 ( .A(n5731), .Y(n5729) );
  INVX1 U4723 ( .A(n5729), .Y(n5730) );
  AND2X1 U4724 ( .A(n9317), .B(n1271), .Y(n1302) );
  INVX1 U4725 ( .A(n1302), .Y(n5731) );
  INVX1 U4726 ( .A(n5734), .Y(n5732) );
  INVX1 U4727 ( .A(n5732), .Y(n5733) );
  AND2X1 U4728 ( .A(n9320), .B(n1271), .Y(n1301) );
  INVX1 U4729 ( .A(n1301), .Y(n5734) );
  INVX1 U4730 ( .A(n5737), .Y(n5735) );
  INVX1 U4731 ( .A(n5735), .Y(n5736) );
  AND2X1 U4732 ( .A(n9323), .B(n1271), .Y(n1300) );
  INVX1 U4733 ( .A(n1300), .Y(n5737) );
  INVX1 U4734 ( .A(n5740), .Y(n5738) );
  INVX1 U4735 ( .A(n5738), .Y(n5739) );
  AND2X1 U4736 ( .A(n9326), .B(n1271), .Y(n1299) );
  INVX1 U4737 ( .A(n1299), .Y(n5740) );
  INVX1 U4738 ( .A(n5743), .Y(n5741) );
  INVX1 U4739 ( .A(n5741), .Y(n5742) );
  AND2X1 U4740 ( .A(n9329), .B(n1271), .Y(n1298) );
  INVX1 U4741 ( .A(n1298), .Y(n5743) );
  INVX1 U4742 ( .A(n5746), .Y(n5744) );
  INVX1 U4743 ( .A(n5744), .Y(n5745) );
  AND2X1 U4744 ( .A(n9332), .B(n1271), .Y(n1297) );
  INVX1 U4745 ( .A(n1297), .Y(n5746) );
  INVX1 U4746 ( .A(n5749), .Y(n5747) );
  INVX1 U4747 ( .A(n5747), .Y(n5748) );
  AND2X1 U4748 ( .A(n9335), .B(n1271), .Y(n1296) );
  INVX1 U4749 ( .A(n1296), .Y(n5749) );
  INVX1 U4750 ( .A(n5752), .Y(n5750) );
  INVX1 U4751 ( .A(n5750), .Y(n5751) );
  AND2X1 U4752 ( .A(n9338), .B(n1271), .Y(n1295) );
  INVX1 U4753 ( .A(n1295), .Y(n5752) );
  INVX1 U4754 ( .A(n5755), .Y(n5753) );
  INVX1 U4755 ( .A(n5753), .Y(n5754) );
  AND2X1 U4756 ( .A(n9341), .B(n1271), .Y(n1294) );
  INVX1 U4757 ( .A(n1294), .Y(n5755) );
  INVX1 U4758 ( .A(n5758), .Y(n5756) );
  INVX1 U4759 ( .A(n5756), .Y(n5757) );
  AND2X1 U4760 ( .A(n9344), .B(n1271), .Y(n1293) );
  INVX1 U4761 ( .A(n1293), .Y(n5758) );
  INVX1 U4762 ( .A(n5761), .Y(n5759) );
  INVX1 U4763 ( .A(n5759), .Y(n5760) );
  AND2X1 U4764 ( .A(n9347), .B(n1271), .Y(n1292) );
  INVX1 U4765 ( .A(n1292), .Y(n5761) );
  INVX1 U4766 ( .A(n5764), .Y(n5762) );
  INVX1 U4767 ( .A(n5762), .Y(n5763) );
  AND2X1 U4768 ( .A(n9350), .B(n1271), .Y(n1291) );
  INVX1 U4769 ( .A(n1291), .Y(n5764) );
  INVX1 U4770 ( .A(n5767), .Y(n5765) );
  INVX1 U4771 ( .A(n5765), .Y(n5766) );
  AND2X1 U4772 ( .A(n9353), .B(n1271), .Y(n1290) );
  INVX1 U4773 ( .A(n1290), .Y(n5767) );
  INVX1 U4774 ( .A(n5770), .Y(n5768) );
  INVX1 U4775 ( .A(n5768), .Y(n5769) );
  AND2X1 U4776 ( .A(n9356), .B(n1271), .Y(n1289) );
  INVX1 U4777 ( .A(n1289), .Y(n5770) );
  INVX1 U4778 ( .A(n5773), .Y(n5771) );
  INVX1 U4779 ( .A(n5771), .Y(n5772) );
  AND2X1 U4780 ( .A(n9359), .B(n1271), .Y(n1288) );
  INVX1 U4781 ( .A(n1288), .Y(n5773) );
  INVX1 U4782 ( .A(n5776), .Y(n5774) );
  INVX1 U4783 ( .A(n5774), .Y(n5775) );
  AND2X1 U4784 ( .A(n9362), .B(n1271), .Y(n1287) );
  INVX1 U4785 ( .A(n1287), .Y(n5776) );
  INVX1 U4786 ( .A(n5779), .Y(n5777) );
  INVX1 U4787 ( .A(n5777), .Y(n5778) );
  AND2X1 U4788 ( .A(n9365), .B(n1271), .Y(n1286) );
  INVX1 U4789 ( .A(n1286), .Y(n5779) );
  INVX1 U4790 ( .A(n5782), .Y(n5780) );
  INVX1 U4791 ( .A(n5780), .Y(n5781) );
  AND2X1 U4792 ( .A(n9368), .B(n1271), .Y(n1285) );
  INVX1 U4793 ( .A(n1285), .Y(n5782) );
  INVX1 U4794 ( .A(n5785), .Y(n5783) );
  INVX1 U4795 ( .A(n5783), .Y(n5784) );
  AND2X1 U4796 ( .A(n9371), .B(n1271), .Y(n1284) );
  INVX1 U4797 ( .A(n1284), .Y(n5785) );
  INVX1 U4798 ( .A(n5788), .Y(n5786) );
  INVX1 U4799 ( .A(n5786), .Y(n5787) );
  AND2X1 U4800 ( .A(n9374), .B(n1271), .Y(n1283) );
  INVX1 U4801 ( .A(n1283), .Y(n5788) );
  INVX1 U4802 ( .A(n5791), .Y(n5789) );
  INVX1 U4803 ( .A(n5789), .Y(n5790) );
  AND2X1 U4804 ( .A(n9377), .B(n1271), .Y(n1282) );
  INVX1 U4805 ( .A(n1282), .Y(n5791) );
  INVX1 U4806 ( .A(n5794), .Y(n5792) );
  INVX1 U4807 ( .A(n5792), .Y(n5793) );
  AND2X1 U4808 ( .A(n9380), .B(n1271), .Y(n1281) );
  INVX1 U4809 ( .A(n1281), .Y(n5794) );
  INVX1 U4810 ( .A(n5797), .Y(n5795) );
  INVX1 U4811 ( .A(n5795), .Y(n5796) );
  AND2X1 U4812 ( .A(n9383), .B(n1271), .Y(n1280) );
  INVX1 U4813 ( .A(n1280), .Y(n5797) );
  INVX1 U4814 ( .A(n5800), .Y(n5798) );
  INVX1 U4815 ( .A(n5798), .Y(n5799) );
  AND2X1 U4816 ( .A(n9386), .B(n1271), .Y(n1279) );
  INVX1 U4817 ( .A(n1279), .Y(n5800) );
  INVX1 U4818 ( .A(n5803), .Y(n5801) );
  INVX1 U4819 ( .A(n5801), .Y(n5802) );
  AND2X1 U4820 ( .A(n9389), .B(n1271), .Y(n1278) );
  INVX1 U4821 ( .A(n1278), .Y(n5803) );
  INVX1 U4822 ( .A(n5806), .Y(n5804) );
  INVX1 U4823 ( .A(n5804), .Y(n5805) );
  AND2X1 U4824 ( .A(n9392), .B(n1271), .Y(n1277) );
  INVX1 U4825 ( .A(n1277), .Y(n5806) );
  INVX1 U4826 ( .A(n5809), .Y(n5807) );
  INVX1 U4827 ( .A(n5807), .Y(n5808) );
  AND2X1 U4828 ( .A(n9395), .B(n1271), .Y(n1276) );
  INVX1 U4829 ( .A(n1276), .Y(n5809) );
  INVX1 U4830 ( .A(n5812), .Y(n5810) );
  INVX1 U4831 ( .A(n5810), .Y(n5811) );
  AND2X1 U4832 ( .A(n9398), .B(n1271), .Y(n1275) );
  INVX1 U4833 ( .A(n1275), .Y(n5812) );
  INVX1 U4834 ( .A(n5815), .Y(n5813) );
  INVX1 U4835 ( .A(n5813), .Y(n5814) );
  AND2X1 U4836 ( .A(n9401), .B(n1271), .Y(n1274) );
  INVX1 U4837 ( .A(n1274), .Y(n5815) );
  INVX1 U4838 ( .A(n5818), .Y(n5816) );
  INVX1 U4839 ( .A(n5816), .Y(n5817) );
  AND2X1 U4840 ( .A(n9404), .B(n1271), .Y(n1273) );
  INVX1 U4841 ( .A(n1273), .Y(n5818) );
  INVX1 U4842 ( .A(n5821), .Y(n5819) );
  INVX1 U4843 ( .A(n5819), .Y(n5820) );
  AND2X1 U4844 ( .A(n9407), .B(n1271), .Y(n1272) );
  INVX1 U4845 ( .A(n1272), .Y(n5821) );
  INVX1 U4846 ( .A(n5824), .Y(n5822) );
  INVX1 U4847 ( .A(n5822), .Y(n5823) );
  AND2X1 U4848 ( .A(n11434), .B(n13034), .Y(n1270) );
  INVX1 U4849 ( .A(n1270), .Y(n5824) );
  INVX1 U4850 ( .A(n5827), .Y(n5825) );
  INVX1 U4851 ( .A(n5825), .Y(n5826) );
  AND2X1 U4852 ( .A(n11437), .B(n13035), .Y(n1269) );
  INVX1 U4853 ( .A(n1269), .Y(n5827) );
  INVX1 U4854 ( .A(n5830), .Y(n5828) );
  INVX1 U4855 ( .A(n5828), .Y(n5829) );
  AND2X1 U4856 ( .A(n11440), .B(n13036), .Y(n1268) );
  INVX1 U4857 ( .A(n1268), .Y(n5830) );
  INVX1 U4858 ( .A(n5833), .Y(n5831) );
  INVX1 U4859 ( .A(n5831), .Y(n5832) );
  AND2X1 U4860 ( .A(n11443), .B(n13034), .Y(n1267) );
  INVX1 U4861 ( .A(n1267), .Y(n5833) );
  INVX1 U4862 ( .A(n5836), .Y(n5834) );
  INVX1 U4863 ( .A(n5834), .Y(n5835) );
  AND2X1 U4864 ( .A(n11446), .B(n8654), .Y(n1266) );
  INVX1 U4865 ( .A(n1266), .Y(n5836) );
  INVX1 U4866 ( .A(n5839), .Y(n5837) );
  INVX1 U4867 ( .A(n5837), .Y(n5838) );
  AND2X1 U4868 ( .A(n11449), .B(n8768), .Y(n1265) );
  INVX1 U4869 ( .A(n1265), .Y(n5839) );
  INVX1 U4870 ( .A(n5842), .Y(n5840) );
  INVX1 U4871 ( .A(n5840), .Y(n5841) );
  AND2X1 U4872 ( .A(n11452), .B(n13034), .Y(n1264) );
  INVX1 U4873 ( .A(n1264), .Y(n5842) );
  INVX1 U4874 ( .A(n5845), .Y(n5843) );
  INVX1 U4875 ( .A(n5843), .Y(n5844) );
  AND2X1 U4876 ( .A(n11455), .B(n8754), .Y(n1263) );
  INVX1 U4877 ( .A(n1263), .Y(n5845) );
  INVX1 U4878 ( .A(n5848), .Y(n5846) );
  INVX1 U4879 ( .A(n5846), .Y(n5847) );
  AND2X1 U4880 ( .A(n11458), .B(n8642), .Y(n1262) );
  INVX1 U4881 ( .A(n1262), .Y(n5848) );
  INVX1 U4882 ( .A(n5851), .Y(n5849) );
  INVX1 U4883 ( .A(n5849), .Y(n5850) );
  AND2X1 U4884 ( .A(n11461), .B(n13034), .Y(n1261) );
  INVX1 U4885 ( .A(n1261), .Y(n5851) );
  INVX1 U4886 ( .A(n5854), .Y(n5852) );
  INVX1 U4887 ( .A(n5852), .Y(n5853) );
  AND2X1 U4888 ( .A(n11464), .B(n8630), .Y(n1260) );
  INVX1 U4889 ( .A(n1260), .Y(n5854) );
  INVX1 U4890 ( .A(n5857), .Y(n5855) );
  INVX1 U4891 ( .A(n5855), .Y(n5856) );
  AND2X1 U4892 ( .A(n11467), .B(n8768), .Y(n1259) );
  INVX1 U4893 ( .A(n1259), .Y(n5857) );
  INVX1 U4894 ( .A(n5860), .Y(n5858) );
  INVX1 U4895 ( .A(n5858), .Y(n5859) );
  AND2X1 U4896 ( .A(n11470), .B(n13034), .Y(n1258) );
  INVX1 U4897 ( .A(n1258), .Y(n5860) );
  INVX1 U4898 ( .A(n5863), .Y(n5861) );
  INVX1 U4899 ( .A(n5861), .Y(n5862) );
  AND2X1 U4900 ( .A(n11473), .B(n13026), .Y(n1257) );
  INVX1 U4901 ( .A(n1257), .Y(n5863) );
  INVX1 U4902 ( .A(n5866), .Y(n5864) );
  INVX1 U4903 ( .A(n5864), .Y(n5865) );
  AND2X1 U4904 ( .A(n11476), .B(n13026), .Y(n1256) );
  INVX1 U4905 ( .A(n1256), .Y(n5866) );
  INVX1 U4906 ( .A(n5869), .Y(n5867) );
  INVX1 U4907 ( .A(n5867), .Y(n5868) );
  AND2X1 U4908 ( .A(n11479), .B(n13034), .Y(n1255) );
  INVX1 U4909 ( .A(n1255), .Y(n5869) );
  INVX1 U4910 ( .A(n5872), .Y(n5870) );
  INVX1 U4911 ( .A(n5870), .Y(n5871) );
  AND2X1 U4912 ( .A(n11482), .B(n13035), .Y(n1254) );
  INVX1 U4913 ( .A(n1254), .Y(n5872) );
  INVX1 U4914 ( .A(n5875), .Y(n5873) );
  INVX1 U4915 ( .A(n5873), .Y(n5874) );
  AND2X1 U4916 ( .A(n11485), .B(n8636), .Y(n1253) );
  INVX1 U4917 ( .A(n1253), .Y(n5875) );
  INVX1 U4918 ( .A(n5878), .Y(n5876) );
  INVX1 U4919 ( .A(n5876), .Y(n5877) );
  AND2X1 U4920 ( .A(n11488), .B(n13034), .Y(n1252) );
  INVX1 U4921 ( .A(n1252), .Y(n5878) );
  INVX1 U4922 ( .A(n5881), .Y(n5879) );
  INVX1 U4923 ( .A(n5879), .Y(n5880) );
  AND2X1 U4924 ( .A(n11491), .B(n8760), .Y(n1251) );
  INVX1 U4925 ( .A(n1251), .Y(n5881) );
  INVX1 U4926 ( .A(n5884), .Y(n5882) );
  INVX1 U4927 ( .A(n5882), .Y(n5883) );
  AND2X1 U4928 ( .A(n11494), .B(n10802), .Y(n1250) );
  INVX1 U4929 ( .A(n1250), .Y(n5884) );
  INVX1 U4930 ( .A(n5887), .Y(n5885) );
  INVX1 U4931 ( .A(n5885), .Y(n5886) );
  AND2X1 U4932 ( .A(n11497), .B(n13034), .Y(n1249) );
  INVX1 U4933 ( .A(n1249), .Y(n5887) );
  INVX1 U4934 ( .A(n5890), .Y(n5888) );
  INVX1 U4935 ( .A(n5888), .Y(n5889) );
  AND2X1 U4936 ( .A(n11500), .B(n12975), .Y(n1248) );
  INVX1 U4937 ( .A(n1248), .Y(n5890) );
  INVX1 U4938 ( .A(n5893), .Y(n5891) );
  INVX1 U4939 ( .A(n5891), .Y(n5892) );
  AND2X1 U4940 ( .A(n11503), .B(n13026), .Y(n1247) );
  INVX1 U4941 ( .A(n1247), .Y(n5893) );
  INVX1 U4942 ( .A(n5896), .Y(n5894) );
  INVX1 U4943 ( .A(n5894), .Y(n5895) );
  AND2X1 U4944 ( .A(n11506), .B(n13034), .Y(n1246) );
  INVX1 U4945 ( .A(n1246), .Y(n5896) );
  INVX1 U4946 ( .A(n5899), .Y(n5897) );
  INVX1 U4947 ( .A(n5897), .Y(n5898) );
  AND2X1 U4948 ( .A(n11509), .B(n8656), .Y(n1245) );
  INVX1 U4949 ( .A(n1245), .Y(n5899) );
  INVX1 U4950 ( .A(n5902), .Y(n5900) );
  INVX1 U4951 ( .A(n5900), .Y(n5901) );
  AND2X1 U4952 ( .A(n11512), .B(n12984), .Y(n1244) );
  INVX1 U4953 ( .A(n1244), .Y(n5902) );
  INVX1 U4954 ( .A(n5905), .Y(n5903) );
  INVX1 U4955 ( .A(n5903), .Y(n5904) );
  AND2X1 U4956 ( .A(n11515), .B(n13034), .Y(n1243) );
  INVX1 U4957 ( .A(n1243), .Y(n5905) );
  INVX1 U4958 ( .A(n5908), .Y(n5906) );
  INVX1 U4959 ( .A(n5906), .Y(n5907) );
  AND2X1 U4960 ( .A(n11518), .B(n12962), .Y(n1242) );
  INVX1 U4961 ( .A(n1242), .Y(n5908) );
  INVX1 U4962 ( .A(n5911), .Y(n5909) );
  INVX1 U4963 ( .A(n5909), .Y(n5910) );
  AND2X1 U4964 ( .A(n11521), .B(n12962), .Y(n1241) );
  INVX1 U4965 ( .A(n1241), .Y(n5911) );
  INVX1 U4966 ( .A(n5914), .Y(n5912) );
  INVX1 U4967 ( .A(n5912), .Y(n5913) );
  AND2X1 U4968 ( .A(n11524), .B(n13034), .Y(n1240) );
  INVX1 U4969 ( .A(n1240), .Y(n5914) );
  INVX1 U4970 ( .A(n5917), .Y(n5915) );
  INVX1 U4971 ( .A(n5915), .Y(n5916) );
  AND2X1 U4972 ( .A(n11527), .B(n12975), .Y(n1239) );
  INVX1 U4973 ( .A(n1239), .Y(n5917) );
  INVX1 U4974 ( .A(n5920), .Y(n5918) );
  INVX1 U4975 ( .A(n5918), .Y(n5919) );
  AND2X1 U4976 ( .A(n11530), .B(n13026), .Y(n1238) );
  INVX1 U4977 ( .A(n1238), .Y(n5920) );
  INVX1 U4978 ( .A(n5923), .Y(n5921) );
  INVX1 U4979 ( .A(n5921), .Y(n5922) );
  AND2X1 U4980 ( .A(n11533), .B(n13034), .Y(n1237) );
  INVX1 U4981 ( .A(n1237), .Y(n5923) );
  INVX1 U4982 ( .A(n5926), .Y(n5924) );
  INVX1 U4983 ( .A(n5924), .Y(n5925) );
  AND2X1 U4984 ( .A(n11536), .B(n12984), .Y(n1236) );
  INVX1 U4985 ( .A(n1236), .Y(n5926) );
  INVX1 U4986 ( .A(n5929), .Y(n5927) );
  INVX1 U4987 ( .A(n5927), .Y(n5928) );
  AND2X1 U4988 ( .A(n11539), .B(n13036), .Y(n1235) );
  INVX1 U4989 ( .A(n1235), .Y(n5929) );
  INVX1 U4990 ( .A(n5932), .Y(n5930) );
  INVX1 U4991 ( .A(n5930), .Y(n5931) );
  AND2X1 U4992 ( .A(n11542), .B(n13034), .Y(n1234) );
  INVX1 U4993 ( .A(n1234), .Y(n5932) );
  INVX1 U4994 ( .A(n5935), .Y(n5933) );
  INVX1 U4995 ( .A(n5933), .Y(n5934) );
  AND2X1 U4996 ( .A(n11545), .B(n13026), .Y(n1233) );
  INVX1 U4997 ( .A(n1233), .Y(n5935) );
  INVX1 U4998 ( .A(n5938), .Y(n5936) );
  INVX1 U4999 ( .A(n5936), .Y(n5937) );
  AND2X1 U5000 ( .A(n11548), .B(n8668), .Y(n1232) );
  INVX1 U5001 ( .A(n1232), .Y(n5938) );
  INVX1 U5002 ( .A(n5941), .Y(n5939) );
  INVX1 U5003 ( .A(n5939), .Y(n5940) );
  AND2X1 U5004 ( .A(n11551), .B(n13034), .Y(n1231) );
  INVX1 U5005 ( .A(n1231), .Y(n5941) );
  INVX1 U5006 ( .A(n5944), .Y(n5942) );
  INVX1 U5007 ( .A(n5942), .Y(n5943) );
  AND2X1 U5008 ( .A(n11554), .B(n13035), .Y(n1230) );
  INVX1 U5009 ( .A(n1230), .Y(n5944) );
  INVX1 U5010 ( .A(n5947), .Y(n5945) );
  INVX1 U5011 ( .A(n5945), .Y(n5946) );
  AND2X1 U5012 ( .A(n11557), .B(n13026), .Y(n1229) );
  INVX1 U5013 ( .A(n1229), .Y(n5947) );
  INVX1 U5014 ( .A(n5950), .Y(n5948) );
  INVX1 U5015 ( .A(n5948), .Y(n5949) );
  AND2X1 U5016 ( .A(n9410), .B(n1185), .Y(n1227) );
  INVX1 U5017 ( .A(n1227), .Y(n5950) );
  INVX1 U5018 ( .A(n5953), .Y(n5951) );
  INVX1 U5019 ( .A(n5951), .Y(n5952) );
  AND2X1 U5020 ( .A(n9413), .B(n1185), .Y(n1226) );
  INVX1 U5021 ( .A(n1226), .Y(n5953) );
  INVX1 U5022 ( .A(n5956), .Y(n5954) );
  INVX1 U5023 ( .A(n5954), .Y(n5955) );
  AND2X1 U5024 ( .A(n9416), .B(n1185), .Y(n1225) );
  INVX1 U5025 ( .A(n1225), .Y(n5956) );
  INVX1 U5026 ( .A(n5959), .Y(n5957) );
  INVX1 U5027 ( .A(n5957), .Y(n5958) );
  AND2X1 U5028 ( .A(n9419), .B(n1185), .Y(n1224) );
  INVX1 U5029 ( .A(n1224), .Y(n5959) );
  INVX1 U5030 ( .A(n5962), .Y(n5960) );
  INVX1 U5031 ( .A(n5960), .Y(n5961) );
  AND2X1 U5032 ( .A(n9422), .B(n1185), .Y(n1223) );
  INVX1 U5033 ( .A(n1223), .Y(n5962) );
  INVX1 U5034 ( .A(n5965), .Y(n5963) );
  INVX1 U5035 ( .A(n5963), .Y(n5964) );
  AND2X1 U5036 ( .A(n9425), .B(n1185), .Y(n1222) );
  INVX1 U5037 ( .A(n1222), .Y(n5965) );
  INVX1 U5038 ( .A(n5968), .Y(n5966) );
  INVX1 U5039 ( .A(n5966), .Y(n5967) );
  AND2X1 U5040 ( .A(n9428), .B(n1185), .Y(n1221) );
  INVX1 U5041 ( .A(n1221), .Y(n5968) );
  INVX1 U5042 ( .A(n5971), .Y(n5969) );
  INVX1 U5043 ( .A(n5969), .Y(n5970) );
  AND2X1 U5044 ( .A(n9431), .B(n1185), .Y(n1220) );
  INVX1 U5045 ( .A(n1220), .Y(n5971) );
  INVX1 U5046 ( .A(n5974), .Y(n5972) );
  INVX1 U5047 ( .A(n5972), .Y(n5973) );
  AND2X1 U5048 ( .A(n9434), .B(n1185), .Y(n1219) );
  INVX1 U5049 ( .A(n1219), .Y(n5974) );
  INVX1 U5050 ( .A(n5977), .Y(n5975) );
  INVX1 U5051 ( .A(n5975), .Y(n5976) );
  AND2X1 U5052 ( .A(n9437), .B(n1185), .Y(n1218) );
  INVX1 U5053 ( .A(n1218), .Y(n5977) );
  INVX1 U5054 ( .A(n5980), .Y(n5978) );
  INVX1 U5055 ( .A(n5978), .Y(n5979) );
  AND2X1 U5056 ( .A(n9440), .B(n1185), .Y(n1217) );
  INVX1 U5057 ( .A(n1217), .Y(n5980) );
  INVX1 U5058 ( .A(n5983), .Y(n5981) );
  INVX1 U5059 ( .A(n5981), .Y(n5982) );
  AND2X1 U5060 ( .A(n9443), .B(n1185), .Y(n1216) );
  INVX1 U5061 ( .A(n1216), .Y(n5983) );
  INVX1 U5062 ( .A(n5986), .Y(n5984) );
  INVX1 U5063 ( .A(n5984), .Y(n5985) );
  AND2X1 U5064 ( .A(n9446), .B(n1185), .Y(n1215) );
  INVX1 U5065 ( .A(n1215), .Y(n5986) );
  INVX1 U5066 ( .A(n5989), .Y(n5987) );
  INVX1 U5067 ( .A(n5987), .Y(n5988) );
  AND2X1 U5068 ( .A(n9449), .B(n1185), .Y(n1214) );
  INVX1 U5069 ( .A(n1214), .Y(n5989) );
  INVX1 U5070 ( .A(n5992), .Y(n5990) );
  INVX1 U5071 ( .A(n5990), .Y(n5991) );
  AND2X1 U5072 ( .A(n9452), .B(n1185), .Y(n1213) );
  INVX1 U5073 ( .A(n1213), .Y(n5992) );
  INVX1 U5074 ( .A(n5995), .Y(n5993) );
  INVX1 U5075 ( .A(n5993), .Y(n5994) );
  AND2X1 U5076 ( .A(n9455), .B(n1185), .Y(n1212) );
  INVX1 U5077 ( .A(n1212), .Y(n5995) );
  INVX1 U5078 ( .A(n5998), .Y(n5996) );
  INVX1 U5079 ( .A(n5996), .Y(n5997) );
  AND2X1 U5080 ( .A(n9458), .B(n1185), .Y(n1211) );
  INVX1 U5081 ( .A(n1211), .Y(n5998) );
  INVX1 U5082 ( .A(n6001), .Y(n5999) );
  INVX1 U5083 ( .A(n5999), .Y(n6000) );
  AND2X1 U5084 ( .A(n9461), .B(n1185), .Y(n1210) );
  INVX1 U5085 ( .A(n1210), .Y(n6001) );
  INVX1 U5086 ( .A(n6004), .Y(n6002) );
  INVX1 U5087 ( .A(n6002), .Y(n6003) );
  AND2X1 U5088 ( .A(n9464), .B(n1185), .Y(n1209) );
  INVX1 U5089 ( .A(n1209), .Y(n6004) );
  INVX1 U5090 ( .A(n6007), .Y(n6005) );
  INVX1 U5091 ( .A(n6005), .Y(n6006) );
  AND2X1 U5092 ( .A(n9467), .B(n1185), .Y(n1208) );
  INVX1 U5093 ( .A(n1208), .Y(n6007) );
  INVX1 U5094 ( .A(n6010), .Y(n6008) );
  INVX1 U5095 ( .A(n6008), .Y(n6009) );
  AND2X1 U5096 ( .A(n9470), .B(n1185), .Y(n1207) );
  INVX1 U5097 ( .A(n1207), .Y(n6010) );
  INVX1 U5098 ( .A(n6013), .Y(n6011) );
  INVX1 U5099 ( .A(n6011), .Y(n6012) );
  AND2X1 U5100 ( .A(n9473), .B(n1185), .Y(n1206) );
  INVX1 U5101 ( .A(n1206), .Y(n6013) );
  INVX1 U5102 ( .A(n6016), .Y(n6014) );
  INVX1 U5103 ( .A(n6014), .Y(n6015) );
  AND2X1 U5104 ( .A(n9476), .B(n1185), .Y(n1205) );
  INVX1 U5105 ( .A(n1205), .Y(n6016) );
  INVX1 U5106 ( .A(n6019), .Y(n6017) );
  INVX1 U5107 ( .A(n6017), .Y(n6018) );
  AND2X1 U5108 ( .A(n9479), .B(n1185), .Y(n1204) );
  INVX1 U5109 ( .A(n1204), .Y(n6019) );
  INVX1 U5110 ( .A(n6022), .Y(n6020) );
  INVX1 U5111 ( .A(n6020), .Y(n6021) );
  AND2X1 U5112 ( .A(n9482), .B(n1185), .Y(n1203) );
  INVX1 U5113 ( .A(n1203), .Y(n6022) );
  INVX1 U5114 ( .A(n6025), .Y(n6023) );
  INVX1 U5115 ( .A(n6023), .Y(n6024) );
  AND2X1 U5116 ( .A(n9485), .B(n1185), .Y(n1202) );
  INVX1 U5117 ( .A(n1202), .Y(n6025) );
  INVX1 U5118 ( .A(n6028), .Y(n6026) );
  INVX1 U5119 ( .A(n6026), .Y(n6027) );
  AND2X1 U5120 ( .A(n9488), .B(n1185), .Y(n1201) );
  INVX1 U5121 ( .A(n1201), .Y(n6028) );
  INVX1 U5122 ( .A(n6031), .Y(n6029) );
  INVX1 U5123 ( .A(n6029), .Y(n6030) );
  AND2X1 U5124 ( .A(n9491), .B(n1185), .Y(n1200) );
  INVX1 U5125 ( .A(n1200), .Y(n6031) );
  INVX1 U5126 ( .A(n6034), .Y(n6032) );
  INVX1 U5127 ( .A(n6032), .Y(n6033) );
  AND2X1 U5128 ( .A(n9494), .B(n1185), .Y(n1199) );
  INVX1 U5129 ( .A(n1199), .Y(n6034) );
  INVX1 U5130 ( .A(n6037), .Y(n6035) );
  INVX1 U5131 ( .A(n6035), .Y(n6036) );
  AND2X1 U5132 ( .A(n9497), .B(n1185), .Y(n1198) );
  INVX1 U5133 ( .A(n1198), .Y(n6037) );
  INVX1 U5134 ( .A(n6040), .Y(n6038) );
  INVX1 U5135 ( .A(n6038), .Y(n6039) );
  AND2X1 U5136 ( .A(n9500), .B(n1185), .Y(n1197) );
  INVX1 U5137 ( .A(n1197), .Y(n6040) );
  INVX1 U5138 ( .A(n6043), .Y(n6041) );
  INVX1 U5139 ( .A(n6041), .Y(n6042) );
  AND2X1 U5140 ( .A(n9503), .B(n1185), .Y(n1196) );
  INVX1 U5141 ( .A(n1196), .Y(n6043) );
  INVX1 U5142 ( .A(n6046), .Y(n6044) );
  INVX1 U5143 ( .A(n6044), .Y(n6045) );
  AND2X1 U5144 ( .A(n9506), .B(n1185), .Y(n1195) );
  INVX1 U5145 ( .A(n1195), .Y(n6046) );
  INVX1 U5146 ( .A(n6049), .Y(n6047) );
  INVX1 U5147 ( .A(n6047), .Y(n6048) );
  AND2X1 U5148 ( .A(n9509), .B(n1185), .Y(n1194) );
  INVX1 U5149 ( .A(n1194), .Y(n6049) );
  INVX1 U5150 ( .A(n6052), .Y(n6050) );
  INVX1 U5151 ( .A(n6050), .Y(n6051) );
  AND2X1 U5152 ( .A(n9512), .B(n1185), .Y(n1193) );
  INVX1 U5153 ( .A(n1193), .Y(n6052) );
  INVX1 U5154 ( .A(n6055), .Y(n6053) );
  INVX1 U5155 ( .A(n6053), .Y(n6054) );
  AND2X1 U5156 ( .A(n9515), .B(n1185), .Y(n1192) );
  INVX1 U5157 ( .A(n1192), .Y(n6055) );
  INVX1 U5158 ( .A(n6058), .Y(n6056) );
  INVX1 U5159 ( .A(n6056), .Y(n6057) );
  AND2X1 U5160 ( .A(n9518), .B(n1185), .Y(n1191) );
  INVX1 U5161 ( .A(n1191), .Y(n6058) );
  INVX1 U5162 ( .A(n6061), .Y(n6059) );
  INVX1 U5163 ( .A(n6059), .Y(n6060) );
  AND2X1 U5164 ( .A(n9521), .B(n1185), .Y(n1190) );
  INVX1 U5165 ( .A(n1190), .Y(n6061) );
  INVX1 U5166 ( .A(n6064), .Y(n6062) );
  INVX1 U5167 ( .A(n6062), .Y(n6063) );
  AND2X1 U5168 ( .A(n9524), .B(n1185), .Y(n1189) );
  INVX1 U5169 ( .A(n1189), .Y(n6064) );
  INVX1 U5170 ( .A(n6067), .Y(n6065) );
  INVX1 U5171 ( .A(n6065), .Y(n6066) );
  AND2X1 U5172 ( .A(n9527), .B(n1185), .Y(n1188) );
  INVX1 U5173 ( .A(n1188), .Y(n6067) );
  INVX1 U5174 ( .A(n6070), .Y(n6068) );
  INVX1 U5175 ( .A(n6068), .Y(n6069) );
  AND2X1 U5176 ( .A(n9530), .B(n1185), .Y(n1187) );
  INVX1 U5177 ( .A(n1187), .Y(n6070) );
  INVX1 U5178 ( .A(n6073), .Y(n6071) );
  INVX1 U5179 ( .A(n6071), .Y(n6072) );
  AND2X1 U5180 ( .A(n9533), .B(n1185), .Y(n1186) );
  INVX1 U5181 ( .A(n1186), .Y(n6073) );
  INVX1 U5182 ( .A(n6076), .Y(n6074) );
  INVX1 U5183 ( .A(n6074), .Y(n6075) );
  AND2X1 U5184 ( .A(n11560), .B(n1142), .Y(n1184) );
  INVX1 U5185 ( .A(n1184), .Y(n6076) );
  INVX1 U5186 ( .A(n6079), .Y(n6077) );
  INVX1 U5187 ( .A(n6077), .Y(n6078) );
  AND2X1 U5188 ( .A(n11563), .B(n1142), .Y(n1183) );
  INVX1 U5189 ( .A(n1183), .Y(n6079) );
  INVX1 U5190 ( .A(n6082), .Y(n6080) );
  INVX1 U5191 ( .A(n6080), .Y(n6081) );
  AND2X1 U5192 ( .A(n11566), .B(n1142), .Y(n1182) );
  INVX1 U5193 ( .A(n1182), .Y(n6082) );
  INVX1 U5194 ( .A(n6085), .Y(n6083) );
  INVX1 U5195 ( .A(n6083), .Y(n6084) );
  AND2X1 U5196 ( .A(n11569), .B(n1142), .Y(n1181) );
  INVX1 U5197 ( .A(n1181), .Y(n6085) );
  INVX1 U5198 ( .A(n6088), .Y(n6086) );
  INVX1 U5199 ( .A(n6086), .Y(n6087) );
  AND2X1 U5200 ( .A(n11572), .B(n1142), .Y(n1180) );
  INVX1 U5201 ( .A(n1180), .Y(n6088) );
  INVX1 U5202 ( .A(n6091), .Y(n6089) );
  INVX1 U5203 ( .A(n6089), .Y(n6090) );
  AND2X1 U5204 ( .A(n11575), .B(n1142), .Y(n1179) );
  INVX1 U5205 ( .A(n1179), .Y(n6091) );
  INVX1 U5206 ( .A(n6094), .Y(n6092) );
  INVX1 U5207 ( .A(n6092), .Y(n6093) );
  AND2X1 U5208 ( .A(n11578), .B(n1142), .Y(n1178) );
  INVX1 U5209 ( .A(n1178), .Y(n6094) );
  INVX1 U5210 ( .A(n6097), .Y(n6095) );
  INVX1 U5211 ( .A(n6095), .Y(n6096) );
  AND2X1 U5212 ( .A(n11581), .B(n1142), .Y(n1177) );
  INVX1 U5213 ( .A(n1177), .Y(n6097) );
  INVX1 U5214 ( .A(n6100), .Y(n6098) );
  INVX1 U5215 ( .A(n6098), .Y(n6099) );
  AND2X1 U5216 ( .A(n11584), .B(n1142), .Y(n1176) );
  INVX1 U5217 ( .A(n1176), .Y(n6100) );
  INVX1 U5218 ( .A(n6103), .Y(n6101) );
  INVX1 U5219 ( .A(n6101), .Y(n6102) );
  AND2X1 U5220 ( .A(n11587), .B(n1142), .Y(n1175) );
  INVX1 U5221 ( .A(n1175), .Y(n6103) );
  INVX1 U5222 ( .A(n6106), .Y(n6104) );
  INVX1 U5223 ( .A(n6104), .Y(n6105) );
  AND2X1 U5224 ( .A(n11590), .B(n1142), .Y(n1174) );
  INVX1 U5225 ( .A(n1174), .Y(n6106) );
  INVX1 U5226 ( .A(n6109), .Y(n6107) );
  INVX1 U5227 ( .A(n6107), .Y(n6108) );
  AND2X1 U5228 ( .A(n11593), .B(n1142), .Y(n1173) );
  INVX1 U5229 ( .A(n1173), .Y(n6109) );
  INVX1 U5230 ( .A(n6112), .Y(n6110) );
  INVX1 U5231 ( .A(n6110), .Y(n6111) );
  AND2X1 U5232 ( .A(n11596), .B(n1142), .Y(n1172) );
  INVX1 U5233 ( .A(n1172), .Y(n6112) );
  INVX1 U5234 ( .A(n6115), .Y(n6113) );
  INVX1 U5235 ( .A(n6113), .Y(n6114) );
  AND2X1 U5236 ( .A(n11599), .B(n1142), .Y(n1171) );
  INVX1 U5237 ( .A(n1171), .Y(n6115) );
  INVX1 U5238 ( .A(n6118), .Y(n6116) );
  INVX1 U5239 ( .A(n6116), .Y(n6117) );
  AND2X1 U5240 ( .A(n11602), .B(n1142), .Y(n1170) );
  INVX1 U5241 ( .A(n1170), .Y(n6118) );
  INVX1 U5242 ( .A(n6121), .Y(n6119) );
  INVX1 U5243 ( .A(n6119), .Y(n6120) );
  AND2X1 U5244 ( .A(n11605), .B(n1142), .Y(n1169) );
  INVX1 U5245 ( .A(n1169), .Y(n6121) );
  INVX1 U5246 ( .A(n6124), .Y(n6122) );
  INVX1 U5247 ( .A(n6122), .Y(n6123) );
  AND2X1 U5248 ( .A(n11608), .B(n1142), .Y(n1168) );
  INVX1 U5249 ( .A(n1168), .Y(n6124) );
  INVX1 U5250 ( .A(n6127), .Y(n6125) );
  INVX1 U5251 ( .A(n6125), .Y(n6126) );
  AND2X1 U5252 ( .A(n11611), .B(n1142), .Y(n1167) );
  INVX1 U5253 ( .A(n1167), .Y(n6127) );
  INVX1 U5254 ( .A(n6130), .Y(n6128) );
  INVX1 U5255 ( .A(n6128), .Y(n6129) );
  AND2X1 U5256 ( .A(n11614), .B(n1142), .Y(n1166) );
  INVX1 U5257 ( .A(n1166), .Y(n6130) );
  INVX1 U5258 ( .A(n6133), .Y(n6131) );
  INVX1 U5259 ( .A(n6131), .Y(n6132) );
  AND2X1 U5260 ( .A(n11617), .B(n1142), .Y(n1165) );
  INVX1 U5261 ( .A(n1165), .Y(n6133) );
  INVX1 U5262 ( .A(n6136), .Y(n6134) );
  INVX1 U5263 ( .A(n6134), .Y(n6135) );
  AND2X1 U5264 ( .A(n11620), .B(n1142), .Y(n1164) );
  INVX1 U5265 ( .A(n1164), .Y(n6136) );
  INVX1 U5266 ( .A(n6139), .Y(n6137) );
  INVX1 U5267 ( .A(n6137), .Y(n6138) );
  AND2X1 U5268 ( .A(n11623), .B(n1142), .Y(n1163) );
  INVX1 U5269 ( .A(n1163), .Y(n6139) );
  INVX1 U5270 ( .A(n6142), .Y(n6140) );
  INVX1 U5271 ( .A(n6140), .Y(n6141) );
  AND2X1 U5272 ( .A(n11626), .B(n1142), .Y(n1162) );
  INVX1 U5273 ( .A(n1162), .Y(n6142) );
  INVX1 U5274 ( .A(n6145), .Y(n6143) );
  INVX1 U5275 ( .A(n6143), .Y(n6144) );
  AND2X1 U5276 ( .A(n11629), .B(n1142), .Y(n1161) );
  INVX1 U5277 ( .A(n1161), .Y(n6145) );
  INVX1 U5278 ( .A(n6148), .Y(n6146) );
  INVX1 U5279 ( .A(n6146), .Y(n6147) );
  AND2X1 U5280 ( .A(n11632), .B(n1142), .Y(n1160) );
  INVX1 U5281 ( .A(n1160), .Y(n6148) );
  INVX1 U5282 ( .A(n6151), .Y(n6149) );
  INVX1 U5283 ( .A(n6149), .Y(n6150) );
  AND2X1 U5284 ( .A(n11635), .B(n1142), .Y(n1159) );
  INVX1 U5285 ( .A(n1159), .Y(n6151) );
  INVX1 U5286 ( .A(n6154), .Y(n6152) );
  INVX1 U5287 ( .A(n6152), .Y(n6153) );
  AND2X1 U5288 ( .A(n11638), .B(n1142), .Y(n1158) );
  INVX1 U5289 ( .A(n1158), .Y(n6154) );
  INVX1 U5290 ( .A(n6157), .Y(n6155) );
  INVX1 U5291 ( .A(n6155), .Y(n6156) );
  AND2X1 U5292 ( .A(n11641), .B(n1142), .Y(n1157) );
  INVX1 U5293 ( .A(n1157), .Y(n6157) );
  INVX1 U5294 ( .A(n6160), .Y(n6158) );
  INVX1 U5295 ( .A(n6158), .Y(n6159) );
  AND2X1 U5296 ( .A(n11644), .B(n1142), .Y(n1156) );
  INVX1 U5297 ( .A(n1156), .Y(n6160) );
  INVX1 U5298 ( .A(n6163), .Y(n6161) );
  INVX1 U5299 ( .A(n6161), .Y(n6162) );
  AND2X1 U5300 ( .A(n11647), .B(n1142), .Y(n1155) );
  INVX1 U5301 ( .A(n1155), .Y(n6163) );
  INVX1 U5302 ( .A(n6166), .Y(n6164) );
  INVX1 U5303 ( .A(n6164), .Y(n6165) );
  AND2X1 U5304 ( .A(n11650), .B(n1142), .Y(n1154) );
  INVX1 U5305 ( .A(n1154), .Y(n6166) );
  INVX1 U5306 ( .A(n6169), .Y(n6167) );
  INVX1 U5307 ( .A(n6167), .Y(n6168) );
  AND2X1 U5308 ( .A(n11653), .B(n1142), .Y(n1153) );
  INVX1 U5309 ( .A(n1153), .Y(n6169) );
  INVX1 U5310 ( .A(n6172), .Y(n6170) );
  INVX1 U5311 ( .A(n6170), .Y(n6171) );
  AND2X1 U5312 ( .A(n11656), .B(n1142), .Y(n1152) );
  INVX1 U5313 ( .A(n1152), .Y(n6172) );
  INVX1 U5314 ( .A(n6175), .Y(n6173) );
  INVX1 U5315 ( .A(n6173), .Y(n6174) );
  AND2X1 U5316 ( .A(n11659), .B(n1142), .Y(n1151) );
  INVX1 U5317 ( .A(n1151), .Y(n6175) );
  INVX1 U5318 ( .A(n6178), .Y(n6176) );
  INVX1 U5319 ( .A(n6176), .Y(n6177) );
  AND2X1 U5320 ( .A(n11662), .B(n1142), .Y(n1150) );
  INVX1 U5321 ( .A(n1150), .Y(n6178) );
  INVX1 U5322 ( .A(n6181), .Y(n6179) );
  INVX1 U5323 ( .A(n6179), .Y(n6180) );
  AND2X1 U5324 ( .A(n11665), .B(n1142), .Y(n1149) );
  INVX1 U5325 ( .A(n1149), .Y(n6181) );
  INVX1 U5326 ( .A(n6184), .Y(n6182) );
  INVX1 U5327 ( .A(n6182), .Y(n6183) );
  AND2X1 U5328 ( .A(n11668), .B(n1142), .Y(n1148) );
  INVX1 U5329 ( .A(n1148), .Y(n6184) );
  INVX1 U5330 ( .A(n6187), .Y(n6185) );
  INVX1 U5331 ( .A(n6185), .Y(n6186) );
  AND2X1 U5332 ( .A(n11671), .B(n1142), .Y(n1147) );
  INVX1 U5333 ( .A(n1147), .Y(n6187) );
  INVX1 U5334 ( .A(n6190), .Y(n6188) );
  INVX1 U5335 ( .A(n6188), .Y(n6189) );
  AND2X1 U5336 ( .A(n11674), .B(n1142), .Y(n1146) );
  INVX1 U5337 ( .A(n1146), .Y(n6190) );
  INVX1 U5338 ( .A(n6193), .Y(n6191) );
  INVX1 U5339 ( .A(n6191), .Y(n6192) );
  AND2X1 U5340 ( .A(n11677), .B(n1142), .Y(n1145) );
  INVX1 U5341 ( .A(n1145), .Y(n6193) );
  INVX1 U5342 ( .A(n6196), .Y(n6194) );
  INVX1 U5343 ( .A(n6194), .Y(n6195) );
  AND2X1 U5344 ( .A(n11680), .B(n1142), .Y(n1144) );
  INVX1 U5345 ( .A(n1144), .Y(n6196) );
  INVX1 U5346 ( .A(n6199), .Y(n6197) );
  INVX1 U5347 ( .A(n6197), .Y(n6198) );
  AND2X1 U5348 ( .A(n11683), .B(n1142), .Y(n1143) );
  INVX1 U5349 ( .A(n1143), .Y(n6199) );
  INVX1 U5350 ( .A(n6202), .Y(n6200) );
  INVX1 U5351 ( .A(n6200), .Y(n6201) );
  AND2X1 U5352 ( .A(n9536), .B(n1099), .Y(n1141) );
  INVX1 U5353 ( .A(n1141), .Y(n6202) );
  INVX1 U5354 ( .A(n6205), .Y(n6203) );
  INVX1 U5355 ( .A(n6203), .Y(n6204) );
  AND2X1 U5356 ( .A(n9539), .B(n1099), .Y(n1140) );
  INVX1 U5357 ( .A(n1140), .Y(n6205) );
  INVX1 U5358 ( .A(n6208), .Y(n6206) );
  INVX1 U5359 ( .A(n6206), .Y(n6207) );
  AND2X1 U5360 ( .A(n9542), .B(n1099), .Y(n1139) );
  INVX1 U5361 ( .A(n1139), .Y(n6208) );
  INVX1 U5362 ( .A(n6211), .Y(n6209) );
  INVX1 U5363 ( .A(n6209), .Y(n6210) );
  AND2X1 U5364 ( .A(n9545), .B(n1099), .Y(n1138) );
  INVX1 U5365 ( .A(n1138), .Y(n6211) );
  INVX1 U5366 ( .A(n6214), .Y(n6212) );
  INVX1 U5367 ( .A(n6212), .Y(n6213) );
  AND2X1 U5368 ( .A(n9548), .B(n1099), .Y(n1137) );
  INVX1 U5369 ( .A(n1137), .Y(n6214) );
  INVX1 U5370 ( .A(n6217), .Y(n6215) );
  INVX1 U5371 ( .A(n6215), .Y(n6216) );
  AND2X1 U5372 ( .A(n9551), .B(n1099), .Y(n1136) );
  INVX1 U5373 ( .A(n1136), .Y(n6217) );
  INVX1 U5374 ( .A(n6220), .Y(n6218) );
  INVX1 U5375 ( .A(n6218), .Y(n6219) );
  AND2X1 U5376 ( .A(n9554), .B(n1099), .Y(n1135) );
  INVX1 U5377 ( .A(n1135), .Y(n6220) );
  INVX1 U5378 ( .A(n6223), .Y(n6221) );
  INVX1 U5379 ( .A(n6221), .Y(n6222) );
  AND2X1 U5380 ( .A(n9557), .B(n1099), .Y(n1134) );
  INVX1 U5381 ( .A(n1134), .Y(n6223) );
  INVX1 U5382 ( .A(n6226), .Y(n6224) );
  INVX1 U5383 ( .A(n6224), .Y(n6225) );
  AND2X1 U5384 ( .A(n9560), .B(n1099), .Y(n1133) );
  INVX1 U5385 ( .A(n1133), .Y(n6226) );
  INVX1 U5386 ( .A(n6229), .Y(n6227) );
  INVX1 U5387 ( .A(n6227), .Y(n6228) );
  AND2X1 U5388 ( .A(n9563), .B(n1099), .Y(n1132) );
  INVX1 U5389 ( .A(n1132), .Y(n6229) );
  INVX1 U5390 ( .A(n6232), .Y(n6230) );
  INVX1 U5391 ( .A(n6230), .Y(n6231) );
  AND2X1 U5392 ( .A(n9566), .B(n1099), .Y(n1131) );
  INVX1 U5393 ( .A(n1131), .Y(n6232) );
  INVX1 U5394 ( .A(n6235), .Y(n6233) );
  INVX1 U5395 ( .A(n6233), .Y(n6234) );
  AND2X1 U5396 ( .A(n9569), .B(n1099), .Y(n1130) );
  INVX1 U5397 ( .A(n1130), .Y(n6235) );
  INVX1 U5398 ( .A(n6238), .Y(n6236) );
  INVX1 U5399 ( .A(n6236), .Y(n6237) );
  AND2X1 U5400 ( .A(n9572), .B(n1099), .Y(n1129) );
  INVX1 U5401 ( .A(n1129), .Y(n6238) );
  INVX1 U5402 ( .A(n6241), .Y(n6239) );
  INVX1 U5403 ( .A(n6239), .Y(n6240) );
  AND2X1 U5404 ( .A(n9575), .B(n1099), .Y(n1128) );
  INVX1 U5405 ( .A(n1128), .Y(n6241) );
  INVX1 U5406 ( .A(n6244), .Y(n6242) );
  INVX1 U5407 ( .A(n6242), .Y(n6243) );
  AND2X1 U5408 ( .A(n9578), .B(n1099), .Y(n1127) );
  INVX1 U5409 ( .A(n1127), .Y(n6244) );
  INVX1 U5410 ( .A(n6247), .Y(n6245) );
  INVX1 U5411 ( .A(n6245), .Y(n6246) );
  AND2X1 U5412 ( .A(n9581), .B(n1099), .Y(n1126) );
  INVX1 U5413 ( .A(n1126), .Y(n6247) );
  INVX1 U5414 ( .A(n6250), .Y(n6248) );
  INVX1 U5415 ( .A(n6248), .Y(n6249) );
  AND2X1 U5416 ( .A(n9584), .B(n1099), .Y(n1125) );
  INVX1 U5417 ( .A(n1125), .Y(n6250) );
  INVX1 U5418 ( .A(n6253), .Y(n6251) );
  INVX1 U5419 ( .A(n6251), .Y(n6252) );
  AND2X1 U5420 ( .A(n9587), .B(n1099), .Y(n1124) );
  INVX1 U5421 ( .A(n1124), .Y(n6253) );
  INVX1 U5422 ( .A(n6256), .Y(n6254) );
  INVX1 U5423 ( .A(n6254), .Y(n6255) );
  AND2X1 U5424 ( .A(n9590), .B(n1099), .Y(n1123) );
  INVX1 U5425 ( .A(n1123), .Y(n6256) );
  INVX1 U5426 ( .A(n6259), .Y(n6257) );
  INVX1 U5427 ( .A(n6257), .Y(n6258) );
  AND2X1 U5428 ( .A(n9593), .B(n1099), .Y(n1122) );
  INVX1 U5429 ( .A(n1122), .Y(n6259) );
  INVX1 U5430 ( .A(n6262), .Y(n6260) );
  INVX1 U5431 ( .A(n6260), .Y(n6261) );
  AND2X1 U5432 ( .A(n9596), .B(n1099), .Y(n1121) );
  INVX1 U5433 ( .A(n1121), .Y(n6262) );
  INVX1 U5434 ( .A(n6265), .Y(n6263) );
  INVX1 U5435 ( .A(n6263), .Y(n6264) );
  AND2X1 U5436 ( .A(n9599), .B(n1099), .Y(n1120) );
  INVX1 U5437 ( .A(n1120), .Y(n6265) );
  INVX1 U5438 ( .A(n6268), .Y(n6266) );
  INVX1 U5439 ( .A(n6266), .Y(n6267) );
  AND2X1 U5440 ( .A(n9602), .B(n1099), .Y(n1119) );
  INVX1 U5441 ( .A(n1119), .Y(n6268) );
  INVX1 U5442 ( .A(n6271), .Y(n6269) );
  INVX1 U5443 ( .A(n6269), .Y(n6270) );
  AND2X1 U5444 ( .A(n9605), .B(n1099), .Y(n1118) );
  INVX1 U5445 ( .A(n1118), .Y(n6271) );
  INVX1 U5446 ( .A(n6274), .Y(n6272) );
  INVX1 U5447 ( .A(n6272), .Y(n6273) );
  AND2X1 U5448 ( .A(n9608), .B(n1099), .Y(n1117) );
  INVX1 U5449 ( .A(n1117), .Y(n6274) );
  INVX1 U5450 ( .A(n6277), .Y(n6275) );
  INVX1 U5451 ( .A(n6275), .Y(n6276) );
  AND2X1 U5452 ( .A(n9611), .B(n1099), .Y(n1116) );
  INVX1 U5453 ( .A(n1116), .Y(n6277) );
  INVX1 U5454 ( .A(n6280), .Y(n6278) );
  INVX1 U5455 ( .A(n6278), .Y(n6279) );
  AND2X1 U5456 ( .A(n9614), .B(n1099), .Y(n1115) );
  INVX1 U5457 ( .A(n1115), .Y(n6280) );
  INVX1 U5458 ( .A(n6283), .Y(n6281) );
  INVX1 U5459 ( .A(n6281), .Y(n6282) );
  AND2X1 U5460 ( .A(n9617), .B(n1099), .Y(n1114) );
  INVX1 U5461 ( .A(n1114), .Y(n6283) );
  INVX1 U5462 ( .A(n6286), .Y(n6284) );
  INVX1 U5463 ( .A(n6284), .Y(n6285) );
  AND2X1 U5464 ( .A(n9620), .B(n1099), .Y(n1113) );
  INVX1 U5465 ( .A(n1113), .Y(n6286) );
  INVX1 U5466 ( .A(n6289), .Y(n6287) );
  INVX1 U5467 ( .A(n6287), .Y(n6288) );
  AND2X1 U5468 ( .A(n9623), .B(n1099), .Y(n1112) );
  INVX1 U5469 ( .A(n1112), .Y(n6289) );
  INVX1 U5470 ( .A(n6292), .Y(n6290) );
  INVX1 U5471 ( .A(n6290), .Y(n6291) );
  AND2X1 U5472 ( .A(n9626), .B(n1099), .Y(n1111) );
  INVX1 U5473 ( .A(n1111), .Y(n6292) );
  INVX1 U5474 ( .A(n6295), .Y(n6293) );
  INVX1 U5475 ( .A(n6293), .Y(n6294) );
  AND2X1 U5476 ( .A(n9629), .B(n1099), .Y(n1110) );
  INVX1 U5477 ( .A(n1110), .Y(n6295) );
  INVX1 U5478 ( .A(n6298), .Y(n6296) );
  INVX1 U5479 ( .A(n6296), .Y(n6297) );
  AND2X1 U5480 ( .A(n9632), .B(n1099), .Y(n1109) );
  INVX1 U5481 ( .A(n1109), .Y(n6298) );
  INVX1 U5482 ( .A(n6301), .Y(n6299) );
  INVX1 U5483 ( .A(n6299), .Y(n6300) );
  AND2X1 U5484 ( .A(n9635), .B(n1099), .Y(n1108) );
  INVX1 U5485 ( .A(n1108), .Y(n6301) );
  INVX1 U5486 ( .A(n6304), .Y(n6302) );
  INVX1 U5487 ( .A(n6302), .Y(n6303) );
  AND2X1 U5488 ( .A(n9638), .B(n1099), .Y(n1107) );
  INVX1 U5489 ( .A(n1107), .Y(n6304) );
  INVX1 U5490 ( .A(n6307), .Y(n6305) );
  INVX1 U5491 ( .A(n6305), .Y(n6306) );
  AND2X1 U5492 ( .A(n9641), .B(n1099), .Y(n1106) );
  INVX1 U5493 ( .A(n1106), .Y(n6307) );
  INVX1 U5494 ( .A(n6310), .Y(n6308) );
  INVX1 U5495 ( .A(n6308), .Y(n6309) );
  AND2X1 U5496 ( .A(n9644), .B(n1099), .Y(n1105) );
  INVX1 U5497 ( .A(n1105), .Y(n6310) );
  INVX1 U5498 ( .A(n6313), .Y(n6311) );
  INVX1 U5499 ( .A(n6311), .Y(n6312) );
  AND2X1 U5500 ( .A(n9647), .B(n1099), .Y(n1104) );
  INVX1 U5501 ( .A(n1104), .Y(n6313) );
  INVX1 U5502 ( .A(n6316), .Y(n6314) );
  INVX1 U5503 ( .A(n6314), .Y(n6315) );
  AND2X1 U5504 ( .A(n9650), .B(n1099), .Y(n1103) );
  INVX1 U5505 ( .A(n1103), .Y(n6316) );
  INVX1 U5506 ( .A(n6319), .Y(n6317) );
  INVX1 U5507 ( .A(n6317), .Y(n6318) );
  AND2X1 U5508 ( .A(n9653), .B(n1099), .Y(n1102) );
  INVX1 U5509 ( .A(n1102), .Y(n6319) );
  INVX1 U5510 ( .A(n6322), .Y(n6320) );
  INVX1 U5511 ( .A(n6320), .Y(n6321) );
  AND2X1 U5512 ( .A(n9656), .B(n1099), .Y(n1101) );
  INVX1 U5513 ( .A(n1101), .Y(n6322) );
  INVX1 U5514 ( .A(n6325), .Y(n6323) );
  INVX1 U5515 ( .A(n6323), .Y(n6324) );
  AND2X1 U5516 ( .A(n9659), .B(n1099), .Y(n1100) );
  INVX1 U5517 ( .A(n1100), .Y(n6325) );
  INVX1 U5518 ( .A(n6328), .Y(n6326) );
  INVX1 U5519 ( .A(n6326), .Y(n6327) );
  AND2X1 U5520 ( .A(n11686), .B(n1056), .Y(n1098) );
  INVX1 U5521 ( .A(n1098), .Y(n6328) );
  INVX1 U5522 ( .A(n6331), .Y(n6329) );
  INVX1 U5523 ( .A(n6329), .Y(n6330) );
  AND2X1 U5524 ( .A(n11689), .B(n1056), .Y(n1097) );
  INVX1 U5525 ( .A(n1097), .Y(n6331) );
  INVX1 U5526 ( .A(n6334), .Y(n6332) );
  INVX1 U5527 ( .A(n6332), .Y(n6333) );
  AND2X1 U5528 ( .A(n11692), .B(n1056), .Y(n1096) );
  INVX1 U5529 ( .A(n1096), .Y(n6334) );
  INVX1 U5530 ( .A(n6337), .Y(n6335) );
  INVX1 U5531 ( .A(n6335), .Y(n6336) );
  AND2X1 U5532 ( .A(n11695), .B(n1056), .Y(n1095) );
  INVX1 U5533 ( .A(n1095), .Y(n6337) );
  INVX1 U5534 ( .A(n6340), .Y(n6338) );
  INVX1 U5535 ( .A(n6338), .Y(n6339) );
  AND2X1 U5536 ( .A(n11698), .B(n1056), .Y(n1094) );
  INVX1 U5537 ( .A(n1094), .Y(n6340) );
  INVX1 U5538 ( .A(n6343), .Y(n6341) );
  INVX1 U5539 ( .A(n6341), .Y(n6342) );
  AND2X1 U5540 ( .A(n11701), .B(n1056), .Y(n1093) );
  INVX1 U5541 ( .A(n1093), .Y(n6343) );
  INVX1 U5542 ( .A(n6346), .Y(n6344) );
  INVX1 U5543 ( .A(n6344), .Y(n6345) );
  AND2X1 U5544 ( .A(n11704), .B(n1056), .Y(n1092) );
  INVX1 U5545 ( .A(n1092), .Y(n6346) );
  INVX1 U5546 ( .A(n6349), .Y(n6347) );
  INVX1 U5547 ( .A(n6347), .Y(n6348) );
  AND2X1 U5548 ( .A(n11707), .B(n1056), .Y(n1091) );
  INVX1 U5549 ( .A(n1091), .Y(n6349) );
  INVX1 U5550 ( .A(n6352), .Y(n6350) );
  INVX1 U5551 ( .A(n6350), .Y(n6351) );
  AND2X1 U5552 ( .A(n11710), .B(n1056), .Y(n1090) );
  INVX1 U5553 ( .A(n1090), .Y(n6352) );
  INVX1 U5554 ( .A(n6355), .Y(n6353) );
  INVX1 U5555 ( .A(n6353), .Y(n6354) );
  AND2X1 U5556 ( .A(n11713), .B(n1056), .Y(n1089) );
  INVX1 U5557 ( .A(n1089), .Y(n6355) );
  INVX1 U5558 ( .A(n6358), .Y(n6356) );
  INVX1 U5559 ( .A(n6356), .Y(n6357) );
  AND2X1 U5560 ( .A(n11716), .B(n1056), .Y(n1088) );
  INVX1 U5561 ( .A(n1088), .Y(n6358) );
  INVX1 U5562 ( .A(n6361), .Y(n6359) );
  INVX1 U5563 ( .A(n6359), .Y(n6360) );
  AND2X1 U5564 ( .A(n11719), .B(n1056), .Y(n1087) );
  INVX1 U5565 ( .A(n1087), .Y(n6361) );
  INVX1 U5566 ( .A(n6364), .Y(n6362) );
  INVX1 U5567 ( .A(n6362), .Y(n6363) );
  AND2X1 U5568 ( .A(n11722), .B(n1056), .Y(n1086) );
  INVX1 U5569 ( .A(n1086), .Y(n6364) );
  INVX1 U5570 ( .A(n6367), .Y(n6365) );
  INVX1 U5571 ( .A(n6365), .Y(n6366) );
  AND2X1 U5572 ( .A(n11725), .B(n1056), .Y(n1085) );
  INVX1 U5573 ( .A(n1085), .Y(n6367) );
  INVX1 U5574 ( .A(n6370), .Y(n6368) );
  INVX1 U5575 ( .A(n6368), .Y(n6369) );
  AND2X1 U5576 ( .A(n11728), .B(n1056), .Y(n1084) );
  INVX1 U5577 ( .A(n1084), .Y(n6370) );
  INVX1 U5578 ( .A(n6373), .Y(n6371) );
  INVX1 U5579 ( .A(n6371), .Y(n6372) );
  AND2X1 U5580 ( .A(n11731), .B(n1056), .Y(n1083) );
  INVX1 U5581 ( .A(n1083), .Y(n6373) );
  INVX1 U5582 ( .A(n6376), .Y(n6374) );
  INVX1 U5583 ( .A(n6374), .Y(n6375) );
  AND2X1 U5584 ( .A(n11734), .B(n1056), .Y(n1082) );
  INVX1 U5585 ( .A(n1082), .Y(n6376) );
  INVX1 U5586 ( .A(n6379), .Y(n6377) );
  INVX1 U5587 ( .A(n6377), .Y(n6378) );
  AND2X1 U5588 ( .A(n11737), .B(n1056), .Y(n1081) );
  INVX1 U5589 ( .A(n1081), .Y(n6379) );
  INVX1 U5590 ( .A(n6382), .Y(n6380) );
  INVX1 U5591 ( .A(n6380), .Y(n6381) );
  AND2X1 U5592 ( .A(n11740), .B(n1056), .Y(n1080) );
  INVX1 U5593 ( .A(n1080), .Y(n6382) );
  INVX1 U5594 ( .A(n6385), .Y(n6383) );
  INVX1 U5595 ( .A(n6383), .Y(n6384) );
  AND2X1 U5596 ( .A(n11743), .B(n1056), .Y(n1079) );
  INVX1 U5597 ( .A(n1079), .Y(n6385) );
  INVX1 U5598 ( .A(n6388), .Y(n6386) );
  INVX1 U5599 ( .A(n6386), .Y(n6387) );
  AND2X1 U5600 ( .A(n11746), .B(n1056), .Y(n1078) );
  INVX1 U5601 ( .A(n1078), .Y(n6388) );
  INVX1 U5602 ( .A(n6391), .Y(n6389) );
  INVX1 U5603 ( .A(n6389), .Y(n6390) );
  AND2X1 U5604 ( .A(n11749), .B(n1056), .Y(n1077) );
  INVX1 U5605 ( .A(n1077), .Y(n6391) );
  INVX1 U5606 ( .A(n6394), .Y(n6392) );
  INVX1 U5607 ( .A(n6392), .Y(n6393) );
  AND2X1 U5608 ( .A(n11752), .B(n1056), .Y(n1076) );
  INVX1 U5609 ( .A(n1076), .Y(n6394) );
  INVX1 U5610 ( .A(n6397), .Y(n6395) );
  INVX1 U5611 ( .A(n6395), .Y(n6396) );
  AND2X1 U5612 ( .A(n11755), .B(n1056), .Y(n1075) );
  INVX1 U5613 ( .A(n1075), .Y(n6397) );
  INVX1 U5614 ( .A(n6400), .Y(n6398) );
  INVX1 U5615 ( .A(n6398), .Y(n6399) );
  AND2X1 U5616 ( .A(n11758), .B(n1056), .Y(n1074) );
  INVX1 U5617 ( .A(n1074), .Y(n6400) );
  INVX1 U5618 ( .A(n6403), .Y(n6401) );
  INVX1 U5619 ( .A(n6401), .Y(n6402) );
  AND2X1 U5620 ( .A(n11761), .B(n1056), .Y(n1073) );
  INVX1 U5621 ( .A(n1073), .Y(n6403) );
  INVX1 U5622 ( .A(n6406), .Y(n6404) );
  INVX1 U5623 ( .A(n6404), .Y(n6405) );
  AND2X1 U5624 ( .A(n11764), .B(n1056), .Y(n1072) );
  INVX1 U5625 ( .A(n1072), .Y(n6406) );
  INVX1 U5626 ( .A(n6409), .Y(n6407) );
  INVX1 U5627 ( .A(n6407), .Y(n6408) );
  AND2X1 U5628 ( .A(n11767), .B(n1056), .Y(n1071) );
  INVX1 U5629 ( .A(n1071), .Y(n6409) );
  INVX1 U5630 ( .A(n6412), .Y(n6410) );
  INVX1 U5631 ( .A(n6410), .Y(n6411) );
  AND2X1 U5632 ( .A(n11770), .B(n1056), .Y(n1070) );
  INVX1 U5633 ( .A(n1070), .Y(n6412) );
  INVX1 U5634 ( .A(n6415), .Y(n6413) );
  INVX1 U5635 ( .A(n6413), .Y(n6414) );
  AND2X1 U5636 ( .A(n11773), .B(n1056), .Y(n1069) );
  INVX1 U5637 ( .A(n1069), .Y(n6415) );
  INVX1 U5638 ( .A(n6418), .Y(n6416) );
  INVX1 U5639 ( .A(n6416), .Y(n6417) );
  AND2X1 U5640 ( .A(n11776), .B(n1056), .Y(n1068) );
  INVX1 U5641 ( .A(n1068), .Y(n6418) );
  INVX1 U5642 ( .A(n6421), .Y(n6419) );
  INVX1 U5643 ( .A(n6419), .Y(n6420) );
  AND2X1 U5644 ( .A(n11779), .B(n1056), .Y(n1067) );
  INVX1 U5645 ( .A(n1067), .Y(n6421) );
  INVX1 U5646 ( .A(n6424), .Y(n6422) );
  INVX1 U5647 ( .A(n6422), .Y(n6423) );
  AND2X1 U5648 ( .A(n11782), .B(n1056), .Y(n1066) );
  INVX1 U5649 ( .A(n1066), .Y(n6424) );
  INVX1 U5650 ( .A(n6427), .Y(n6425) );
  INVX1 U5651 ( .A(n6425), .Y(n6426) );
  AND2X1 U5652 ( .A(n11785), .B(n1056), .Y(n1065) );
  INVX1 U5653 ( .A(n1065), .Y(n6427) );
  INVX1 U5654 ( .A(n6430), .Y(n6428) );
  INVX1 U5655 ( .A(n6428), .Y(n6429) );
  AND2X1 U5656 ( .A(n11788), .B(n1056), .Y(n1064) );
  INVX1 U5657 ( .A(n1064), .Y(n6430) );
  INVX1 U5658 ( .A(n6433), .Y(n6431) );
  INVX1 U5659 ( .A(n6431), .Y(n6432) );
  AND2X1 U5660 ( .A(n11791), .B(n1056), .Y(n1063) );
  INVX1 U5661 ( .A(n1063), .Y(n6433) );
  INVX1 U5662 ( .A(n6436), .Y(n6434) );
  INVX1 U5663 ( .A(n6434), .Y(n6435) );
  AND2X1 U5664 ( .A(n11794), .B(n1056), .Y(n1062) );
  INVX1 U5665 ( .A(n1062), .Y(n6436) );
  INVX1 U5666 ( .A(n6439), .Y(n6437) );
  INVX1 U5667 ( .A(n6437), .Y(n6438) );
  AND2X1 U5668 ( .A(n11797), .B(n1056), .Y(n1061) );
  INVX1 U5669 ( .A(n1061), .Y(n6439) );
  INVX1 U5670 ( .A(n6442), .Y(n6440) );
  INVX1 U5671 ( .A(n6440), .Y(n6441) );
  AND2X1 U5672 ( .A(n11800), .B(n1056), .Y(n1060) );
  INVX1 U5673 ( .A(n1060), .Y(n6442) );
  INVX1 U5674 ( .A(n6445), .Y(n6443) );
  INVX1 U5675 ( .A(n6443), .Y(n6444) );
  AND2X1 U5676 ( .A(n11803), .B(n1056), .Y(n1059) );
  INVX1 U5677 ( .A(n1059), .Y(n6445) );
  INVX1 U5678 ( .A(n6448), .Y(n6446) );
  INVX1 U5679 ( .A(n6446), .Y(n6447) );
  AND2X1 U5680 ( .A(n11806), .B(n1056), .Y(n1058) );
  INVX1 U5681 ( .A(n1058), .Y(n6448) );
  INVX1 U5682 ( .A(n6451), .Y(n6449) );
  INVX1 U5683 ( .A(n6449), .Y(n6450) );
  AND2X1 U5684 ( .A(n11809), .B(n1056), .Y(n1057) );
  INVX1 U5685 ( .A(n1057), .Y(n6451) );
  INVX1 U5686 ( .A(n6454), .Y(n6452) );
  INVX1 U5687 ( .A(n6452), .Y(n6453) );
  AND2X1 U5688 ( .A(n9662), .B(n1012), .Y(n1054) );
  INVX1 U5689 ( .A(n1054), .Y(n6454) );
  INVX1 U5690 ( .A(n6457), .Y(n6455) );
  INVX1 U5691 ( .A(n6455), .Y(n6456) );
  AND2X1 U5692 ( .A(n9665), .B(n1012), .Y(n1053) );
  INVX1 U5693 ( .A(n1053), .Y(n6457) );
  INVX1 U5694 ( .A(n6460), .Y(n6458) );
  INVX1 U5695 ( .A(n6458), .Y(n6459) );
  AND2X1 U5696 ( .A(n9668), .B(n1012), .Y(n1052) );
  INVX1 U5697 ( .A(n1052), .Y(n6460) );
  INVX1 U5698 ( .A(n6463), .Y(n6461) );
  INVX1 U5699 ( .A(n6461), .Y(n6462) );
  AND2X1 U5700 ( .A(n9671), .B(n1012), .Y(n1051) );
  INVX1 U5701 ( .A(n1051), .Y(n6463) );
  INVX1 U5702 ( .A(n6466), .Y(n6464) );
  INVX1 U5703 ( .A(n6464), .Y(n6465) );
  AND2X1 U5704 ( .A(n9674), .B(n1012), .Y(n1050) );
  INVX1 U5705 ( .A(n1050), .Y(n6466) );
  INVX1 U5706 ( .A(n6469), .Y(n6467) );
  INVX1 U5707 ( .A(n6467), .Y(n6468) );
  AND2X1 U5708 ( .A(n9677), .B(n1012), .Y(n1049) );
  INVX1 U5709 ( .A(n1049), .Y(n6469) );
  INVX1 U5710 ( .A(n6472), .Y(n6470) );
  INVX1 U5711 ( .A(n6470), .Y(n6471) );
  AND2X1 U5712 ( .A(n9680), .B(n1012), .Y(n1048) );
  INVX1 U5713 ( .A(n1048), .Y(n6472) );
  INVX1 U5714 ( .A(n6475), .Y(n6473) );
  INVX1 U5715 ( .A(n6473), .Y(n6474) );
  AND2X1 U5716 ( .A(n9683), .B(n1012), .Y(n1047) );
  INVX1 U5717 ( .A(n1047), .Y(n6475) );
  INVX1 U5718 ( .A(n6478), .Y(n6476) );
  INVX1 U5719 ( .A(n6476), .Y(n6477) );
  AND2X1 U5720 ( .A(n9686), .B(n1012), .Y(n1046) );
  INVX1 U5721 ( .A(n1046), .Y(n6478) );
  INVX1 U5722 ( .A(n6481), .Y(n6479) );
  INVX1 U5723 ( .A(n6479), .Y(n6480) );
  AND2X1 U5724 ( .A(n9689), .B(n1012), .Y(n1045) );
  INVX1 U5725 ( .A(n1045), .Y(n6481) );
  INVX1 U5726 ( .A(n6484), .Y(n6482) );
  INVX1 U5727 ( .A(n6482), .Y(n6483) );
  AND2X1 U5728 ( .A(n9692), .B(n1012), .Y(n1044) );
  INVX1 U5729 ( .A(n1044), .Y(n6484) );
  INVX1 U5730 ( .A(n6487), .Y(n6485) );
  INVX1 U5731 ( .A(n6485), .Y(n6486) );
  AND2X1 U5732 ( .A(n9695), .B(n1012), .Y(n1043) );
  INVX1 U5733 ( .A(n1043), .Y(n6487) );
  INVX1 U5734 ( .A(n6490), .Y(n6488) );
  INVX1 U5735 ( .A(n6488), .Y(n6489) );
  AND2X1 U5736 ( .A(n9698), .B(n1012), .Y(n1042) );
  INVX1 U5737 ( .A(n1042), .Y(n6490) );
  INVX1 U5738 ( .A(n6493), .Y(n6491) );
  INVX1 U5739 ( .A(n6491), .Y(n6492) );
  AND2X1 U5740 ( .A(n9701), .B(n1012), .Y(n1041) );
  INVX1 U5741 ( .A(n1041), .Y(n6493) );
  INVX1 U5742 ( .A(n6496), .Y(n6494) );
  INVX1 U5743 ( .A(n6494), .Y(n6495) );
  AND2X1 U5744 ( .A(n9704), .B(n1012), .Y(n1040) );
  INVX1 U5745 ( .A(n1040), .Y(n6496) );
  INVX1 U5746 ( .A(n6499), .Y(n6497) );
  INVX1 U5747 ( .A(n6497), .Y(n6498) );
  AND2X1 U5748 ( .A(n9707), .B(n1012), .Y(n1039) );
  INVX1 U5749 ( .A(n1039), .Y(n6499) );
  INVX1 U5750 ( .A(n6502), .Y(n6500) );
  INVX1 U5751 ( .A(n6500), .Y(n6501) );
  AND2X1 U5752 ( .A(n9710), .B(n1012), .Y(n1038) );
  INVX1 U5753 ( .A(n1038), .Y(n6502) );
  INVX1 U5754 ( .A(n6505), .Y(n6503) );
  INVX1 U5755 ( .A(n6503), .Y(n6504) );
  AND2X1 U5756 ( .A(n9713), .B(n1012), .Y(n1037) );
  INVX1 U5757 ( .A(n1037), .Y(n6505) );
  INVX1 U5758 ( .A(n6508), .Y(n6506) );
  INVX1 U5759 ( .A(n6506), .Y(n6507) );
  AND2X1 U5760 ( .A(n9716), .B(n1012), .Y(n1036) );
  INVX1 U5761 ( .A(n1036), .Y(n6508) );
  INVX1 U5762 ( .A(n6511), .Y(n6509) );
  INVX1 U5763 ( .A(n6509), .Y(n6510) );
  AND2X1 U5764 ( .A(n9719), .B(n1012), .Y(n1035) );
  INVX1 U5765 ( .A(n1035), .Y(n6511) );
  INVX1 U5766 ( .A(n6514), .Y(n6512) );
  INVX1 U5767 ( .A(n6512), .Y(n6513) );
  AND2X1 U5768 ( .A(n9722), .B(n1012), .Y(n1034) );
  INVX1 U5769 ( .A(n1034), .Y(n6514) );
  INVX1 U5770 ( .A(n6517), .Y(n6515) );
  INVX1 U5771 ( .A(n6515), .Y(n6516) );
  AND2X1 U5772 ( .A(n9725), .B(n1012), .Y(n1033) );
  INVX1 U5773 ( .A(n1033), .Y(n6517) );
  INVX1 U5774 ( .A(n6520), .Y(n6518) );
  INVX1 U5775 ( .A(n6518), .Y(n6519) );
  AND2X1 U5776 ( .A(n9728), .B(n1012), .Y(n1032) );
  INVX1 U5777 ( .A(n1032), .Y(n6520) );
  INVX1 U5778 ( .A(n6523), .Y(n6521) );
  INVX1 U5779 ( .A(n6521), .Y(n6522) );
  AND2X1 U5780 ( .A(n9731), .B(n1012), .Y(n1031) );
  INVX1 U5781 ( .A(n1031), .Y(n6523) );
  INVX1 U5782 ( .A(n6526), .Y(n6524) );
  INVX1 U5783 ( .A(n6524), .Y(n6525) );
  AND2X1 U5784 ( .A(n9734), .B(n1012), .Y(n1030) );
  INVX1 U5785 ( .A(n1030), .Y(n6526) );
  INVX1 U5786 ( .A(n6529), .Y(n6527) );
  INVX1 U5787 ( .A(n6527), .Y(n6528) );
  AND2X1 U5788 ( .A(n9737), .B(n1012), .Y(n1029) );
  INVX1 U5789 ( .A(n1029), .Y(n6529) );
  INVX1 U5790 ( .A(n6532), .Y(n6530) );
  INVX1 U5791 ( .A(n6530), .Y(n6531) );
  AND2X1 U5792 ( .A(n9740), .B(n1012), .Y(n1028) );
  INVX1 U5793 ( .A(n1028), .Y(n6532) );
  INVX1 U5794 ( .A(n6535), .Y(n6533) );
  INVX1 U5795 ( .A(n6533), .Y(n6534) );
  AND2X1 U5796 ( .A(n9743), .B(n1012), .Y(n1027) );
  INVX1 U5797 ( .A(n1027), .Y(n6535) );
  INVX1 U5798 ( .A(n6538), .Y(n6536) );
  INVX1 U5799 ( .A(n6536), .Y(n6537) );
  AND2X1 U5800 ( .A(n9746), .B(n1012), .Y(n1026) );
  INVX1 U5801 ( .A(n1026), .Y(n6538) );
  INVX1 U5802 ( .A(n6541), .Y(n6539) );
  INVX1 U5803 ( .A(n6539), .Y(n6540) );
  AND2X1 U5804 ( .A(n9749), .B(n1012), .Y(n1025) );
  INVX1 U5805 ( .A(n1025), .Y(n6541) );
  INVX1 U5806 ( .A(n6544), .Y(n6542) );
  INVX1 U5807 ( .A(n6542), .Y(n6543) );
  AND2X1 U5808 ( .A(n9752), .B(n1012), .Y(n1024) );
  INVX1 U5809 ( .A(n1024), .Y(n6544) );
  INVX1 U5810 ( .A(n6547), .Y(n6545) );
  INVX1 U5811 ( .A(n6545), .Y(n6546) );
  AND2X1 U5812 ( .A(n9755), .B(n1012), .Y(n1023) );
  INVX1 U5813 ( .A(n1023), .Y(n6547) );
  INVX1 U5814 ( .A(n6550), .Y(n6548) );
  INVX1 U5815 ( .A(n6548), .Y(n6549) );
  AND2X1 U5816 ( .A(n9758), .B(n1012), .Y(n1022) );
  INVX1 U5817 ( .A(n1022), .Y(n6550) );
  INVX1 U5818 ( .A(n6553), .Y(n6551) );
  INVX1 U5819 ( .A(n6551), .Y(n6552) );
  AND2X1 U5820 ( .A(n9761), .B(n1012), .Y(n1021) );
  INVX1 U5821 ( .A(n1021), .Y(n6553) );
  INVX1 U5822 ( .A(n6556), .Y(n6554) );
  INVX1 U5823 ( .A(n6554), .Y(n6555) );
  AND2X1 U5824 ( .A(n9764), .B(n1012), .Y(n1020) );
  INVX1 U5825 ( .A(n1020), .Y(n6556) );
  INVX1 U5826 ( .A(n6559), .Y(n6557) );
  INVX1 U5827 ( .A(n6557), .Y(n6558) );
  AND2X1 U5828 ( .A(n9767), .B(n1012), .Y(n1019) );
  INVX1 U5829 ( .A(n1019), .Y(n6559) );
  INVX1 U5830 ( .A(n6562), .Y(n6560) );
  INVX1 U5831 ( .A(n6560), .Y(n6561) );
  AND2X1 U5832 ( .A(n9770), .B(n1012), .Y(n1018) );
  INVX1 U5833 ( .A(n1018), .Y(n6562) );
  INVX1 U5834 ( .A(n6565), .Y(n6563) );
  INVX1 U5835 ( .A(n6563), .Y(n6564) );
  AND2X1 U5836 ( .A(n9773), .B(n1012), .Y(n1017) );
  INVX1 U5837 ( .A(n1017), .Y(n6565) );
  INVX1 U5838 ( .A(n6568), .Y(n6566) );
  INVX1 U5839 ( .A(n6566), .Y(n6567) );
  AND2X1 U5840 ( .A(n9776), .B(n1012), .Y(n1016) );
  INVX1 U5841 ( .A(n1016), .Y(n6568) );
  INVX1 U5842 ( .A(n6571), .Y(n6569) );
  INVX1 U5843 ( .A(n6569), .Y(n6570) );
  AND2X1 U5844 ( .A(n9779), .B(n1012), .Y(n1015) );
  INVX1 U5845 ( .A(n1015), .Y(n6571) );
  INVX1 U5846 ( .A(n6574), .Y(n6572) );
  INVX1 U5847 ( .A(n6572), .Y(n6573) );
  AND2X1 U5848 ( .A(n9782), .B(n1012), .Y(n1014) );
  INVX1 U5849 ( .A(n1014), .Y(n6574) );
  INVX1 U5850 ( .A(n6577), .Y(n6575) );
  INVX1 U5851 ( .A(n6575), .Y(n6576) );
  AND2X1 U5852 ( .A(n9785), .B(n1012), .Y(n1013) );
  INVX1 U5853 ( .A(n1013), .Y(n6577) );
  INVX1 U5854 ( .A(n6580), .Y(n6578) );
  INVX1 U5855 ( .A(n6578), .Y(n6579) );
  AND2X1 U5856 ( .A(n11812), .B(n968), .Y(n1010) );
  INVX1 U5857 ( .A(n1010), .Y(n6580) );
  INVX1 U5858 ( .A(n6583), .Y(n6581) );
  INVX1 U5859 ( .A(n6581), .Y(n6582) );
  AND2X1 U5860 ( .A(n11815), .B(n968), .Y(n1009) );
  INVX1 U5861 ( .A(n1009), .Y(n6583) );
  INVX1 U5862 ( .A(n6586), .Y(n6584) );
  INVX1 U5863 ( .A(n6584), .Y(n6585) );
  AND2X1 U5864 ( .A(n11818), .B(n968), .Y(n1008) );
  INVX1 U5865 ( .A(n1008), .Y(n6586) );
  INVX1 U5866 ( .A(n6589), .Y(n6587) );
  INVX1 U5867 ( .A(n6587), .Y(n6588) );
  AND2X1 U5868 ( .A(n11821), .B(n968), .Y(n1007) );
  INVX1 U5869 ( .A(n1007), .Y(n6589) );
  INVX1 U5870 ( .A(n6592), .Y(n6590) );
  INVX1 U5871 ( .A(n6590), .Y(n6591) );
  AND2X1 U5872 ( .A(n11824), .B(n968), .Y(n1006) );
  INVX1 U5873 ( .A(n1006), .Y(n6592) );
  INVX1 U5874 ( .A(n6595), .Y(n6593) );
  INVX1 U5875 ( .A(n6593), .Y(n6594) );
  AND2X1 U5876 ( .A(n11827), .B(n968), .Y(n1005) );
  INVX1 U5877 ( .A(n1005), .Y(n6595) );
  INVX1 U5878 ( .A(n6598), .Y(n6596) );
  INVX1 U5879 ( .A(n6596), .Y(n6597) );
  AND2X1 U5880 ( .A(n11830), .B(n968), .Y(n1004) );
  INVX1 U5881 ( .A(n1004), .Y(n6598) );
  INVX1 U5882 ( .A(n6601), .Y(n6599) );
  INVX1 U5883 ( .A(n6599), .Y(n6600) );
  AND2X1 U5884 ( .A(n11833), .B(n968), .Y(n1003) );
  INVX1 U5885 ( .A(n1003), .Y(n6601) );
  INVX1 U5886 ( .A(n6604), .Y(n6602) );
  INVX1 U5887 ( .A(n6602), .Y(n6603) );
  AND2X1 U5888 ( .A(n11836), .B(n968), .Y(n1002) );
  INVX1 U5889 ( .A(n1002), .Y(n6604) );
  INVX1 U5890 ( .A(n6607), .Y(n6605) );
  INVX1 U5891 ( .A(n6605), .Y(n6606) );
  AND2X1 U5892 ( .A(n11839), .B(n968), .Y(n1001) );
  INVX1 U5893 ( .A(n1001), .Y(n6607) );
  INVX1 U5894 ( .A(n6610), .Y(n6608) );
  INVX1 U5895 ( .A(n6608), .Y(n6609) );
  AND2X1 U5896 ( .A(n11842), .B(n968), .Y(n1000) );
  INVX1 U5897 ( .A(n1000), .Y(n6610) );
  INVX1 U5898 ( .A(n6613), .Y(n6611) );
  INVX1 U5899 ( .A(n6611), .Y(n6612) );
  AND2X1 U5900 ( .A(n11845), .B(n968), .Y(n999) );
  INVX1 U5901 ( .A(n999), .Y(n6613) );
  INVX1 U5902 ( .A(n6616), .Y(n6614) );
  INVX1 U5903 ( .A(n6614), .Y(n6615) );
  AND2X1 U5904 ( .A(n11848), .B(n968), .Y(n998) );
  INVX1 U5905 ( .A(n998), .Y(n6616) );
  INVX1 U5906 ( .A(n6619), .Y(n6617) );
  INVX1 U5907 ( .A(n6617), .Y(n6618) );
  AND2X1 U5908 ( .A(n11851), .B(n968), .Y(n997) );
  INVX1 U5909 ( .A(n997), .Y(n6619) );
  INVX1 U5910 ( .A(n6622), .Y(n6620) );
  INVX1 U5911 ( .A(n6620), .Y(n6621) );
  AND2X1 U5912 ( .A(n11854), .B(n968), .Y(n996) );
  INVX1 U5913 ( .A(n996), .Y(n6622) );
  INVX1 U5914 ( .A(n6625), .Y(n6623) );
  INVX1 U5915 ( .A(n6623), .Y(n6624) );
  AND2X1 U5916 ( .A(n11857), .B(n968), .Y(n995) );
  INVX1 U5917 ( .A(n995), .Y(n6625) );
  INVX1 U5918 ( .A(n6628), .Y(n6626) );
  INVX1 U5919 ( .A(n6626), .Y(n6627) );
  AND2X1 U5920 ( .A(n11860), .B(n968), .Y(n994) );
  INVX1 U5921 ( .A(n994), .Y(n6628) );
  INVX1 U5922 ( .A(n6631), .Y(n6629) );
  INVX1 U5923 ( .A(n6629), .Y(n6630) );
  AND2X1 U5924 ( .A(n11863), .B(n968), .Y(n993) );
  INVX1 U5925 ( .A(n993), .Y(n6631) );
  INVX1 U5926 ( .A(n6634), .Y(n6632) );
  INVX1 U5927 ( .A(n6632), .Y(n6633) );
  AND2X1 U5928 ( .A(n11866), .B(n968), .Y(n992) );
  INVX1 U5929 ( .A(n992), .Y(n6634) );
  INVX1 U5930 ( .A(n6637), .Y(n6635) );
  INVX1 U5931 ( .A(n6635), .Y(n6636) );
  AND2X1 U5932 ( .A(n11869), .B(n968), .Y(n991) );
  INVX1 U5933 ( .A(n991), .Y(n6637) );
  INVX1 U5934 ( .A(n6640), .Y(n6638) );
  INVX1 U5935 ( .A(n6638), .Y(n6639) );
  AND2X1 U5936 ( .A(n11872), .B(n968), .Y(n990) );
  INVX1 U5937 ( .A(n990), .Y(n6640) );
  INVX1 U5938 ( .A(n6643), .Y(n6641) );
  INVX1 U5939 ( .A(n6641), .Y(n6642) );
  AND2X1 U5940 ( .A(n11875), .B(n968), .Y(n989) );
  INVX1 U5941 ( .A(n989), .Y(n6643) );
  INVX1 U5942 ( .A(n6646), .Y(n6644) );
  INVX1 U5943 ( .A(n6644), .Y(n6645) );
  AND2X1 U5944 ( .A(n11878), .B(n968), .Y(n988) );
  INVX1 U5945 ( .A(n988), .Y(n6646) );
  INVX1 U5946 ( .A(n6649), .Y(n6647) );
  INVX1 U5947 ( .A(n6647), .Y(n6648) );
  AND2X1 U5948 ( .A(n11881), .B(n968), .Y(n987) );
  INVX1 U5949 ( .A(n987), .Y(n6649) );
  INVX1 U5950 ( .A(n6652), .Y(n6650) );
  INVX1 U5951 ( .A(n6650), .Y(n6651) );
  AND2X1 U5952 ( .A(n11884), .B(n968), .Y(n986) );
  INVX1 U5953 ( .A(n986), .Y(n6652) );
  INVX1 U5954 ( .A(n6655), .Y(n6653) );
  INVX1 U5955 ( .A(n6653), .Y(n6654) );
  AND2X1 U5956 ( .A(n11887), .B(n968), .Y(n985) );
  INVX1 U5957 ( .A(n985), .Y(n6655) );
  INVX1 U5958 ( .A(n6658), .Y(n6656) );
  INVX1 U5959 ( .A(n6656), .Y(n6657) );
  AND2X1 U5960 ( .A(n11890), .B(n968), .Y(n984) );
  INVX1 U5961 ( .A(n984), .Y(n6658) );
  INVX1 U5962 ( .A(n6661), .Y(n6659) );
  INVX1 U5963 ( .A(n6659), .Y(n6660) );
  AND2X1 U5964 ( .A(n11893), .B(n968), .Y(n983) );
  INVX1 U5965 ( .A(n983), .Y(n6661) );
  INVX1 U5966 ( .A(n6664), .Y(n6662) );
  INVX1 U5967 ( .A(n6662), .Y(n6663) );
  AND2X1 U5968 ( .A(n11896), .B(n968), .Y(n982) );
  INVX1 U5969 ( .A(n982), .Y(n6664) );
  INVX1 U5970 ( .A(n6667), .Y(n6665) );
  INVX1 U5971 ( .A(n6665), .Y(n6666) );
  AND2X1 U5972 ( .A(n11899), .B(n968), .Y(n981) );
  INVX1 U5973 ( .A(n981), .Y(n6667) );
  INVX1 U5974 ( .A(n6670), .Y(n6668) );
  INVX1 U5975 ( .A(n6668), .Y(n6669) );
  AND2X1 U5976 ( .A(n11902), .B(n968), .Y(n980) );
  INVX1 U5977 ( .A(n980), .Y(n6670) );
  INVX1 U5978 ( .A(n6673), .Y(n6671) );
  INVX1 U5979 ( .A(n6671), .Y(n6672) );
  AND2X1 U5980 ( .A(n11905), .B(n968), .Y(n979) );
  INVX1 U5981 ( .A(n979), .Y(n6673) );
  INVX1 U5982 ( .A(n6676), .Y(n6674) );
  INVX1 U5983 ( .A(n6674), .Y(n6675) );
  AND2X1 U5984 ( .A(n11908), .B(n968), .Y(n978) );
  INVX1 U5985 ( .A(n978), .Y(n6676) );
  INVX1 U5986 ( .A(n6679), .Y(n6677) );
  INVX1 U5987 ( .A(n6677), .Y(n6678) );
  AND2X1 U5988 ( .A(n11911), .B(n968), .Y(n977) );
  INVX1 U5989 ( .A(n977), .Y(n6679) );
  INVX1 U5990 ( .A(n6682), .Y(n6680) );
  INVX1 U5991 ( .A(n6680), .Y(n6681) );
  AND2X1 U5992 ( .A(n11914), .B(n968), .Y(n976) );
  INVX1 U5993 ( .A(n976), .Y(n6682) );
  INVX1 U5994 ( .A(n6685), .Y(n6683) );
  INVX1 U5995 ( .A(n6683), .Y(n6684) );
  AND2X1 U5996 ( .A(n11917), .B(n968), .Y(n975) );
  INVX1 U5997 ( .A(n975), .Y(n6685) );
  INVX1 U5998 ( .A(n6688), .Y(n6686) );
  INVX1 U5999 ( .A(n6686), .Y(n6687) );
  AND2X1 U6000 ( .A(n11920), .B(n968), .Y(n974) );
  INVX1 U6001 ( .A(n974), .Y(n6688) );
  INVX1 U6002 ( .A(n6691), .Y(n6689) );
  INVX1 U6003 ( .A(n6689), .Y(n6690) );
  AND2X1 U6004 ( .A(n11923), .B(n968), .Y(n973) );
  INVX1 U6005 ( .A(n973), .Y(n6691) );
  INVX1 U6006 ( .A(n6694), .Y(n6692) );
  INVX1 U6007 ( .A(n6692), .Y(n6693) );
  AND2X1 U6008 ( .A(n11926), .B(n968), .Y(n972) );
  INVX1 U6009 ( .A(n972), .Y(n6694) );
  INVX1 U6010 ( .A(n6697), .Y(n6695) );
  INVX1 U6011 ( .A(n6695), .Y(n6696) );
  AND2X1 U6012 ( .A(n11929), .B(n968), .Y(n971) );
  INVX1 U6013 ( .A(n971), .Y(n6697) );
  INVX1 U6014 ( .A(n6700), .Y(n6698) );
  INVX1 U6015 ( .A(n6698), .Y(n6699) );
  AND2X1 U6016 ( .A(n11932), .B(n968), .Y(n970) );
  INVX1 U6017 ( .A(n970), .Y(n6700) );
  INVX1 U6018 ( .A(n6703), .Y(n6701) );
  INVX1 U6019 ( .A(n6701), .Y(n6702) );
  AND2X1 U6020 ( .A(n11935), .B(n968), .Y(n969) );
  INVX1 U6021 ( .A(n969), .Y(n6703) );
  INVX1 U6022 ( .A(n6706), .Y(n6704) );
  INVX1 U6023 ( .A(n6704), .Y(n6705) );
  AND2X1 U6024 ( .A(n9788), .B(n925), .Y(n967) );
  INVX1 U6025 ( .A(n967), .Y(n6706) );
  INVX1 U6026 ( .A(n6709), .Y(n6707) );
  INVX1 U6027 ( .A(n6707), .Y(n6708) );
  AND2X1 U6028 ( .A(n9791), .B(n925), .Y(n966) );
  INVX1 U6029 ( .A(n966), .Y(n6709) );
  INVX1 U6030 ( .A(n6712), .Y(n6710) );
  INVX1 U6031 ( .A(n6710), .Y(n6711) );
  AND2X1 U6032 ( .A(n9794), .B(n925), .Y(n965) );
  INVX1 U6033 ( .A(n965), .Y(n6712) );
  INVX1 U6034 ( .A(n6715), .Y(n6713) );
  INVX1 U6035 ( .A(n6713), .Y(n6714) );
  AND2X1 U6036 ( .A(n9797), .B(n925), .Y(n964) );
  INVX1 U6037 ( .A(n964), .Y(n6715) );
  INVX1 U6038 ( .A(n6718), .Y(n6716) );
  INVX1 U6039 ( .A(n6716), .Y(n6717) );
  AND2X1 U6040 ( .A(n9800), .B(n925), .Y(n963) );
  INVX1 U6041 ( .A(n963), .Y(n6718) );
  INVX1 U6042 ( .A(n6721), .Y(n6719) );
  INVX1 U6043 ( .A(n6719), .Y(n6720) );
  AND2X1 U6044 ( .A(n9803), .B(n925), .Y(n962) );
  INVX1 U6045 ( .A(n962), .Y(n6721) );
  INVX1 U6046 ( .A(n6724), .Y(n6722) );
  INVX1 U6047 ( .A(n6722), .Y(n6723) );
  AND2X1 U6048 ( .A(n9806), .B(n925), .Y(n961) );
  INVX1 U6049 ( .A(n961), .Y(n6724) );
  INVX1 U6050 ( .A(n6727), .Y(n6725) );
  INVX1 U6051 ( .A(n6725), .Y(n6726) );
  AND2X1 U6052 ( .A(n9809), .B(n925), .Y(n960) );
  INVX1 U6053 ( .A(n960), .Y(n6727) );
  INVX1 U6054 ( .A(n6730), .Y(n6728) );
  INVX1 U6055 ( .A(n6728), .Y(n6729) );
  AND2X1 U6056 ( .A(n9812), .B(n925), .Y(n959) );
  INVX1 U6057 ( .A(n959), .Y(n6730) );
  INVX1 U6058 ( .A(n6733), .Y(n6731) );
  INVX1 U6059 ( .A(n6731), .Y(n6732) );
  AND2X1 U6060 ( .A(n9815), .B(n925), .Y(n958) );
  INVX1 U6061 ( .A(n958), .Y(n6733) );
  INVX1 U6062 ( .A(n6736), .Y(n6734) );
  INVX1 U6063 ( .A(n6734), .Y(n6735) );
  AND2X1 U6064 ( .A(n9818), .B(n925), .Y(n957) );
  INVX1 U6065 ( .A(n957), .Y(n6736) );
  INVX1 U6066 ( .A(n6739), .Y(n6737) );
  INVX1 U6067 ( .A(n6737), .Y(n6738) );
  AND2X1 U6068 ( .A(n9821), .B(n925), .Y(n956) );
  INVX1 U6069 ( .A(n956), .Y(n6739) );
  INVX1 U6070 ( .A(n6742), .Y(n6740) );
  INVX1 U6071 ( .A(n6740), .Y(n6741) );
  AND2X1 U6072 ( .A(n9824), .B(n925), .Y(n955) );
  INVX1 U6073 ( .A(n955), .Y(n6742) );
  INVX1 U6074 ( .A(n6745), .Y(n6743) );
  INVX1 U6075 ( .A(n6743), .Y(n6744) );
  AND2X1 U6076 ( .A(n9827), .B(n925), .Y(n954) );
  INVX1 U6077 ( .A(n954), .Y(n6745) );
  INVX1 U6078 ( .A(n6748), .Y(n6746) );
  INVX1 U6079 ( .A(n6746), .Y(n6747) );
  AND2X1 U6080 ( .A(n9830), .B(n925), .Y(n953) );
  INVX1 U6081 ( .A(n953), .Y(n6748) );
  INVX1 U6082 ( .A(n6751), .Y(n6749) );
  INVX1 U6083 ( .A(n6749), .Y(n6750) );
  AND2X1 U6084 ( .A(n9833), .B(n925), .Y(n952) );
  INVX1 U6085 ( .A(n952), .Y(n6751) );
  INVX1 U6086 ( .A(n6754), .Y(n6752) );
  INVX1 U6087 ( .A(n6752), .Y(n6753) );
  AND2X1 U6088 ( .A(n9836), .B(n925), .Y(n951) );
  INVX1 U6089 ( .A(n951), .Y(n6754) );
  INVX1 U6090 ( .A(n6757), .Y(n6755) );
  INVX1 U6091 ( .A(n6755), .Y(n6756) );
  AND2X1 U6092 ( .A(n9839), .B(n925), .Y(n950) );
  INVX1 U6093 ( .A(n950), .Y(n6757) );
  INVX1 U6094 ( .A(n6760), .Y(n6758) );
  INVX1 U6095 ( .A(n6758), .Y(n6759) );
  AND2X1 U6096 ( .A(n9842), .B(n925), .Y(n949) );
  INVX1 U6097 ( .A(n949), .Y(n6760) );
  INVX1 U6098 ( .A(n6763), .Y(n6761) );
  INVX1 U6099 ( .A(n6761), .Y(n6762) );
  AND2X1 U6100 ( .A(n9845), .B(n925), .Y(n948) );
  INVX1 U6101 ( .A(n948), .Y(n6763) );
  INVX1 U6102 ( .A(n6766), .Y(n6764) );
  INVX1 U6103 ( .A(n6764), .Y(n6765) );
  AND2X1 U6104 ( .A(n9848), .B(n925), .Y(n947) );
  INVX1 U6105 ( .A(n947), .Y(n6766) );
  INVX1 U6106 ( .A(n6769), .Y(n6767) );
  INVX1 U6107 ( .A(n6767), .Y(n6768) );
  AND2X1 U6108 ( .A(n9851), .B(n925), .Y(n946) );
  INVX1 U6109 ( .A(n946), .Y(n6769) );
  INVX1 U6110 ( .A(n6772), .Y(n6770) );
  INVX1 U6111 ( .A(n6770), .Y(n6771) );
  AND2X1 U6112 ( .A(n9854), .B(n925), .Y(n945) );
  INVX1 U6113 ( .A(n945), .Y(n6772) );
  INVX1 U6114 ( .A(n6775), .Y(n6773) );
  INVX1 U6115 ( .A(n6773), .Y(n6774) );
  AND2X1 U6116 ( .A(n9857), .B(n925), .Y(n944) );
  INVX1 U6117 ( .A(n944), .Y(n6775) );
  INVX1 U6118 ( .A(n6778), .Y(n6776) );
  INVX1 U6119 ( .A(n6776), .Y(n6777) );
  AND2X1 U6120 ( .A(n9860), .B(n925), .Y(n943) );
  INVX1 U6121 ( .A(n943), .Y(n6778) );
  INVX1 U6122 ( .A(n6781), .Y(n6779) );
  INVX1 U6123 ( .A(n6779), .Y(n6780) );
  AND2X1 U6124 ( .A(n9863), .B(n925), .Y(n942) );
  INVX1 U6125 ( .A(n942), .Y(n6781) );
  INVX1 U6126 ( .A(n6784), .Y(n6782) );
  INVX1 U6127 ( .A(n6782), .Y(n6783) );
  AND2X1 U6128 ( .A(n9866), .B(n925), .Y(n941) );
  INVX1 U6129 ( .A(n941), .Y(n6784) );
  INVX1 U6130 ( .A(n6787), .Y(n6785) );
  INVX1 U6131 ( .A(n6785), .Y(n6786) );
  AND2X1 U6132 ( .A(n9869), .B(n925), .Y(n940) );
  INVX1 U6133 ( .A(n940), .Y(n6787) );
  INVX1 U6134 ( .A(n6790), .Y(n6788) );
  INVX1 U6135 ( .A(n6788), .Y(n6789) );
  AND2X1 U6136 ( .A(n9872), .B(n925), .Y(n939) );
  INVX1 U6137 ( .A(n939), .Y(n6790) );
  INVX1 U6138 ( .A(n6793), .Y(n6791) );
  INVX1 U6139 ( .A(n6791), .Y(n6792) );
  AND2X1 U6140 ( .A(n9875), .B(n925), .Y(n938) );
  INVX1 U6141 ( .A(n938), .Y(n6793) );
  INVX1 U6142 ( .A(n6796), .Y(n6794) );
  INVX1 U6143 ( .A(n6794), .Y(n6795) );
  AND2X1 U6144 ( .A(n9878), .B(n925), .Y(n937) );
  INVX1 U6145 ( .A(n937), .Y(n6796) );
  INVX1 U6146 ( .A(n6799), .Y(n6797) );
  INVX1 U6147 ( .A(n6797), .Y(n6798) );
  AND2X1 U6148 ( .A(n9881), .B(n925), .Y(n936) );
  INVX1 U6149 ( .A(n936), .Y(n6799) );
  INVX1 U6150 ( .A(n6802), .Y(n6800) );
  INVX1 U6151 ( .A(n6800), .Y(n6801) );
  AND2X1 U6152 ( .A(n9884), .B(n925), .Y(n935) );
  INVX1 U6153 ( .A(n935), .Y(n6802) );
  INVX1 U6154 ( .A(n6805), .Y(n6803) );
  INVX1 U6155 ( .A(n6803), .Y(n6804) );
  AND2X1 U6156 ( .A(n9887), .B(n925), .Y(n934) );
  INVX1 U6157 ( .A(n934), .Y(n6805) );
  INVX1 U6158 ( .A(n6808), .Y(n6806) );
  INVX1 U6159 ( .A(n6806), .Y(n6807) );
  AND2X1 U6160 ( .A(n9890), .B(n925), .Y(n933) );
  INVX1 U6161 ( .A(n933), .Y(n6808) );
  INVX1 U6162 ( .A(n6811), .Y(n6809) );
  INVX1 U6163 ( .A(n6809), .Y(n6810) );
  AND2X1 U6164 ( .A(n9893), .B(n925), .Y(n932) );
  INVX1 U6165 ( .A(n932), .Y(n6811) );
  INVX1 U6166 ( .A(n6814), .Y(n6812) );
  INVX1 U6167 ( .A(n6812), .Y(n6813) );
  AND2X1 U6168 ( .A(n9896), .B(n925), .Y(n931) );
  INVX1 U6169 ( .A(n931), .Y(n6814) );
  INVX1 U6170 ( .A(n6817), .Y(n6815) );
  INVX1 U6171 ( .A(n6815), .Y(n6816) );
  AND2X1 U6172 ( .A(n9899), .B(n925), .Y(n930) );
  INVX1 U6173 ( .A(n930), .Y(n6817) );
  INVX1 U6174 ( .A(n6820), .Y(n6818) );
  INVX1 U6175 ( .A(n6818), .Y(n6819) );
  AND2X1 U6176 ( .A(n9902), .B(n925), .Y(n929) );
  INVX1 U6177 ( .A(n929), .Y(n6820) );
  INVX1 U6178 ( .A(n6823), .Y(n6821) );
  INVX1 U6179 ( .A(n6821), .Y(n6822) );
  AND2X1 U6180 ( .A(n9905), .B(n925), .Y(n928) );
  INVX1 U6181 ( .A(n928), .Y(n6823) );
  INVX1 U6182 ( .A(n6826), .Y(n6824) );
  INVX1 U6183 ( .A(n6824), .Y(n6825) );
  AND2X1 U6184 ( .A(n9908), .B(n925), .Y(n927) );
  INVX1 U6185 ( .A(n927), .Y(n6826) );
  INVX1 U6186 ( .A(n6829), .Y(n6827) );
  INVX1 U6187 ( .A(n6827), .Y(n6828) );
  AND2X1 U6188 ( .A(n9911), .B(n925), .Y(n926) );
  INVX1 U6189 ( .A(n926), .Y(n6829) );
  INVX1 U6190 ( .A(n6832), .Y(n6830) );
  INVX1 U6191 ( .A(n6830), .Y(n6831) );
  AND2X1 U6192 ( .A(n11938), .B(n882), .Y(n924) );
  INVX1 U6193 ( .A(n924), .Y(n6832) );
  INVX1 U6194 ( .A(n6835), .Y(n6833) );
  INVX1 U6195 ( .A(n6833), .Y(n6834) );
  AND2X1 U6196 ( .A(n11941), .B(n882), .Y(n923) );
  INVX1 U6197 ( .A(n923), .Y(n6835) );
  INVX1 U6198 ( .A(n6838), .Y(n6836) );
  INVX1 U6199 ( .A(n6836), .Y(n6837) );
  AND2X1 U6200 ( .A(n11944), .B(n882), .Y(n922) );
  INVX1 U6201 ( .A(n922), .Y(n6838) );
  INVX1 U6202 ( .A(n6841), .Y(n6839) );
  INVX1 U6203 ( .A(n6839), .Y(n6840) );
  AND2X1 U6204 ( .A(n11947), .B(n882), .Y(n921) );
  INVX1 U6205 ( .A(n921), .Y(n6841) );
  INVX1 U6206 ( .A(n6844), .Y(n6842) );
  INVX1 U6207 ( .A(n6842), .Y(n6843) );
  AND2X1 U6208 ( .A(n11950), .B(n882), .Y(n920) );
  INVX1 U6209 ( .A(n920), .Y(n6844) );
  INVX1 U6210 ( .A(n6847), .Y(n6845) );
  INVX1 U6211 ( .A(n6845), .Y(n6846) );
  AND2X1 U6212 ( .A(n11953), .B(n882), .Y(n919) );
  INVX1 U6213 ( .A(n919), .Y(n6847) );
  INVX1 U6214 ( .A(n6850), .Y(n6848) );
  INVX1 U6215 ( .A(n6848), .Y(n6849) );
  AND2X1 U6216 ( .A(n11956), .B(n882), .Y(n918) );
  INVX1 U6217 ( .A(n918), .Y(n6850) );
  INVX1 U6218 ( .A(n6853), .Y(n6851) );
  INVX1 U6219 ( .A(n6851), .Y(n6852) );
  AND2X1 U6220 ( .A(n11959), .B(n882), .Y(n917) );
  INVX1 U6221 ( .A(n917), .Y(n6853) );
  INVX1 U6222 ( .A(n6856), .Y(n6854) );
  INVX1 U6223 ( .A(n6854), .Y(n6855) );
  AND2X1 U6224 ( .A(n11962), .B(n882), .Y(n916) );
  INVX1 U6225 ( .A(n916), .Y(n6856) );
  INVX1 U6226 ( .A(n6859), .Y(n6857) );
  INVX1 U6227 ( .A(n6857), .Y(n6858) );
  AND2X1 U6228 ( .A(n11965), .B(n882), .Y(n915) );
  INVX1 U6229 ( .A(n915), .Y(n6859) );
  INVX1 U6230 ( .A(n6862), .Y(n6860) );
  INVX1 U6231 ( .A(n6860), .Y(n6861) );
  AND2X1 U6232 ( .A(n11968), .B(n882), .Y(n914) );
  INVX1 U6233 ( .A(n914), .Y(n6862) );
  INVX1 U6234 ( .A(n6865), .Y(n6863) );
  INVX1 U6235 ( .A(n6863), .Y(n6864) );
  AND2X1 U6236 ( .A(n11971), .B(n882), .Y(n913) );
  INVX1 U6237 ( .A(n913), .Y(n6865) );
  INVX1 U6238 ( .A(n6868), .Y(n6866) );
  INVX1 U6239 ( .A(n6866), .Y(n6867) );
  AND2X1 U6240 ( .A(n11974), .B(n882), .Y(n912) );
  INVX1 U6241 ( .A(n912), .Y(n6868) );
  INVX1 U6242 ( .A(n6871), .Y(n6869) );
  INVX1 U6243 ( .A(n6869), .Y(n6870) );
  AND2X1 U6244 ( .A(n11977), .B(n882), .Y(n911) );
  INVX1 U6245 ( .A(n911), .Y(n6871) );
  INVX1 U6246 ( .A(n6874), .Y(n6872) );
  INVX1 U6247 ( .A(n6872), .Y(n6873) );
  AND2X1 U6248 ( .A(n11980), .B(n882), .Y(n910) );
  INVX1 U6249 ( .A(n910), .Y(n6874) );
  INVX1 U6250 ( .A(n6877), .Y(n6875) );
  INVX1 U6251 ( .A(n6875), .Y(n6876) );
  AND2X1 U6252 ( .A(n11983), .B(n882), .Y(n909) );
  INVX1 U6253 ( .A(n909), .Y(n6877) );
  INVX1 U6254 ( .A(n6880), .Y(n6878) );
  INVX1 U6255 ( .A(n6878), .Y(n6879) );
  AND2X1 U6256 ( .A(n11986), .B(n882), .Y(n908) );
  INVX1 U6257 ( .A(n908), .Y(n6880) );
  INVX1 U6258 ( .A(n6883), .Y(n6881) );
  INVX1 U6259 ( .A(n6881), .Y(n6882) );
  AND2X1 U6260 ( .A(n11989), .B(n882), .Y(n907) );
  INVX1 U6261 ( .A(n907), .Y(n6883) );
  INVX1 U6262 ( .A(n6886), .Y(n6884) );
  INVX1 U6263 ( .A(n6884), .Y(n6885) );
  AND2X1 U6264 ( .A(n11992), .B(n882), .Y(n906) );
  INVX1 U6265 ( .A(n906), .Y(n6886) );
  INVX1 U6266 ( .A(n6889), .Y(n6887) );
  INVX1 U6267 ( .A(n6887), .Y(n6888) );
  AND2X1 U6268 ( .A(n11995), .B(n882), .Y(n905) );
  INVX1 U6269 ( .A(n905), .Y(n6889) );
  INVX1 U6270 ( .A(n6892), .Y(n6890) );
  INVX1 U6271 ( .A(n6890), .Y(n6891) );
  AND2X1 U6272 ( .A(n11998), .B(n882), .Y(n904) );
  INVX1 U6273 ( .A(n904), .Y(n6892) );
  INVX1 U6274 ( .A(n6895), .Y(n6893) );
  INVX1 U6275 ( .A(n6893), .Y(n6894) );
  AND2X1 U6276 ( .A(n12001), .B(n882), .Y(n903) );
  INVX1 U6277 ( .A(n903), .Y(n6895) );
  INVX1 U6278 ( .A(n6898), .Y(n6896) );
  INVX1 U6279 ( .A(n6896), .Y(n6897) );
  AND2X1 U6280 ( .A(n12004), .B(n882), .Y(n902) );
  INVX1 U6281 ( .A(n902), .Y(n6898) );
  INVX1 U6282 ( .A(n6901), .Y(n6899) );
  INVX1 U6283 ( .A(n6899), .Y(n6900) );
  AND2X1 U6284 ( .A(n12007), .B(n882), .Y(n901) );
  INVX1 U6285 ( .A(n901), .Y(n6901) );
  INVX1 U6286 ( .A(n6904), .Y(n6902) );
  INVX1 U6287 ( .A(n6902), .Y(n6903) );
  AND2X1 U6288 ( .A(n12010), .B(n882), .Y(n900) );
  INVX1 U6289 ( .A(n900), .Y(n6904) );
  INVX1 U6290 ( .A(n6907), .Y(n6905) );
  INVX1 U6291 ( .A(n6905), .Y(n6906) );
  AND2X1 U6292 ( .A(n12013), .B(n882), .Y(n899) );
  INVX1 U6293 ( .A(n899), .Y(n6907) );
  INVX1 U6294 ( .A(n6910), .Y(n6908) );
  INVX1 U6295 ( .A(n6908), .Y(n6909) );
  AND2X1 U6296 ( .A(n12016), .B(n882), .Y(n898) );
  INVX1 U6297 ( .A(n898), .Y(n6910) );
  INVX1 U6298 ( .A(n6913), .Y(n6911) );
  INVX1 U6299 ( .A(n6911), .Y(n6912) );
  AND2X1 U6300 ( .A(n12019), .B(n882), .Y(n897) );
  INVX1 U6301 ( .A(n897), .Y(n6913) );
  INVX1 U6302 ( .A(n6916), .Y(n6914) );
  INVX1 U6303 ( .A(n6914), .Y(n6915) );
  AND2X1 U6304 ( .A(n12022), .B(n882), .Y(n896) );
  INVX1 U6305 ( .A(n896), .Y(n6916) );
  INVX1 U6306 ( .A(n6919), .Y(n6917) );
  INVX1 U6307 ( .A(n6917), .Y(n6918) );
  AND2X1 U6308 ( .A(n12025), .B(n882), .Y(n895) );
  INVX1 U6309 ( .A(n895), .Y(n6919) );
  INVX1 U6310 ( .A(n6922), .Y(n6920) );
  INVX1 U6311 ( .A(n6920), .Y(n6921) );
  AND2X1 U6312 ( .A(n12028), .B(n882), .Y(n894) );
  INVX1 U6313 ( .A(n894), .Y(n6922) );
  INVX1 U6314 ( .A(n6925), .Y(n6923) );
  INVX1 U6315 ( .A(n6923), .Y(n6924) );
  AND2X1 U6316 ( .A(n12031), .B(n882), .Y(n893) );
  INVX1 U6317 ( .A(n893), .Y(n6925) );
  INVX1 U6318 ( .A(n6928), .Y(n6926) );
  INVX1 U6319 ( .A(n6926), .Y(n6927) );
  AND2X1 U6320 ( .A(n12034), .B(n882), .Y(n892) );
  INVX1 U6321 ( .A(n892), .Y(n6928) );
  INVX1 U6322 ( .A(n6931), .Y(n6929) );
  INVX1 U6323 ( .A(n6929), .Y(n6930) );
  AND2X1 U6324 ( .A(n12037), .B(n882), .Y(n891) );
  INVX1 U6325 ( .A(n891), .Y(n6931) );
  INVX1 U6326 ( .A(n6934), .Y(n6932) );
  INVX1 U6327 ( .A(n6932), .Y(n6933) );
  AND2X1 U6328 ( .A(n12040), .B(n882), .Y(n890) );
  INVX1 U6329 ( .A(n890), .Y(n6934) );
  INVX1 U6330 ( .A(n6937), .Y(n6935) );
  INVX1 U6331 ( .A(n6935), .Y(n6936) );
  AND2X1 U6332 ( .A(n12043), .B(n882), .Y(n889) );
  INVX1 U6333 ( .A(n889), .Y(n6937) );
  INVX1 U6334 ( .A(n6940), .Y(n6938) );
  INVX1 U6335 ( .A(n6938), .Y(n6939) );
  AND2X1 U6336 ( .A(n12046), .B(n882), .Y(n888) );
  INVX1 U6337 ( .A(n888), .Y(n6940) );
  INVX1 U6338 ( .A(n6943), .Y(n6941) );
  INVX1 U6339 ( .A(n6941), .Y(n6942) );
  AND2X1 U6340 ( .A(n12049), .B(n882), .Y(n887) );
  INVX1 U6341 ( .A(n887), .Y(n6943) );
  INVX1 U6342 ( .A(n6946), .Y(n6944) );
  INVX1 U6343 ( .A(n6944), .Y(n6945) );
  AND2X1 U6344 ( .A(n12052), .B(n882), .Y(n886) );
  INVX1 U6345 ( .A(n886), .Y(n6946) );
  INVX1 U6346 ( .A(n6949), .Y(n6947) );
  INVX1 U6347 ( .A(n6947), .Y(n6948) );
  AND2X1 U6348 ( .A(n12055), .B(n882), .Y(n885) );
  INVX1 U6349 ( .A(n885), .Y(n6949) );
  INVX1 U6350 ( .A(n6952), .Y(n6950) );
  INVX1 U6351 ( .A(n6950), .Y(n6951) );
  AND2X1 U6352 ( .A(n12058), .B(n882), .Y(n884) );
  INVX1 U6353 ( .A(n884), .Y(n6952) );
  INVX1 U6354 ( .A(n6955), .Y(n6953) );
  INVX1 U6355 ( .A(n6953), .Y(n6954) );
  AND2X1 U6356 ( .A(n12061), .B(n882), .Y(n883) );
  INVX1 U6357 ( .A(n883), .Y(n6955) );
  INVX1 U6358 ( .A(n6958), .Y(n6956) );
  INVX1 U6359 ( .A(n6956), .Y(n6957) );
  AND2X1 U6360 ( .A(n9914), .B(n839), .Y(n881) );
  INVX1 U6361 ( .A(n881), .Y(n6958) );
  INVX1 U6362 ( .A(n6961), .Y(n6959) );
  INVX1 U6363 ( .A(n6959), .Y(n6960) );
  AND2X1 U6364 ( .A(n9917), .B(n839), .Y(n880) );
  INVX1 U6365 ( .A(n880), .Y(n6961) );
  INVX1 U6366 ( .A(n6964), .Y(n6962) );
  INVX1 U6367 ( .A(n6962), .Y(n6963) );
  AND2X1 U6368 ( .A(n9920), .B(n839), .Y(n879) );
  INVX1 U6369 ( .A(n879), .Y(n6964) );
  INVX1 U6370 ( .A(n6967), .Y(n6965) );
  INVX1 U6371 ( .A(n6965), .Y(n6966) );
  AND2X1 U6372 ( .A(n9923), .B(n839), .Y(n878) );
  INVX1 U6373 ( .A(n878), .Y(n6967) );
  INVX1 U6374 ( .A(n6970), .Y(n6968) );
  INVX1 U6375 ( .A(n6968), .Y(n6969) );
  AND2X1 U6376 ( .A(n9926), .B(n839), .Y(n877) );
  INVX1 U6377 ( .A(n877), .Y(n6970) );
  INVX1 U6378 ( .A(n6973), .Y(n6971) );
  INVX1 U6379 ( .A(n6971), .Y(n6972) );
  AND2X1 U6380 ( .A(n9929), .B(n839), .Y(n876) );
  INVX1 U6381 ( .A(n876), .Y(n6973) );
  INVX1 U6382 ( .A(n6976), .Y(n6974) );
  INVX1 U6383 ( .A(n6974), .Y(n6975) );
  AND2X1 U6384 ( .A(n9932), .B(n839), .Y(n875) );
  INVX1 U6385 ( .A(n875), .Y(n6976) );
  INVX1 U6386 ( .A(n6979), .Y(n6977) );
  INVX1 U6387 ( .A(n6977), .Y(n6978) );
  AND2X1 U6388 ( .A(n9935), .B(n839), .Y(n874) );
  INVX1 U6389 ( .A(n874), .Y(n6979) );
  INVX1 U6390 ( .A(n6982), .Y(n6980) );
  INVX1 U6391 ( .A(n6980), .Y(n6981) );
  AND2X1 U6392 ( .A(n9938), .B(n839), .Y(n873) );
  INVX1 U6393 ( .A(n873), .Y(n6982) );
  INVX1 U6394 ( .A(n6985), .Y(n6983) );
  INVX1 U6395 ( .A(n6983), .Y(n6984) );
  AND2X1 U6396 ( .A(n9941), .B(n839), .Y(n872) );
  INVX1 U6397 ( .A(n872), .Y(n6985) );
  INVX1 U6398 ( .A(n6988), .Y(n6986) );
  INVX1 U6399 ( .A(n6986), .Y(n6987) );
  AND2X1 U6400 ( .A(n9944), .B(n839), .Y(n871) );
  INVX1 U6401 ( .A(n871), .Y(n6988) );
  INVX1 U6402 ( .A(n6991), .Y(n6989) );
  INVX1 U6403 ( .A(n6989), .Y(n6990) );
  AND2X1 U6404 ( .A(n9947), .B(n839), .Y(n870) );
  INVX1 U6405 ( .A(n870), .Y(n6991) );
  INVX1 U6406 ( .A(n6994), .Y(n6992) );
  INVX1 U6407 ( .A(n6992), .Y(n6993) );
  AND2X1 U6408 ( .A(n9950), .B(n839), .Y(n869) );
  INVX1 U6409 ( .A(n869), .Y(n6994) );
  INVX1 U6410 ( .A(n6997), .Y(n6995) );
  INVX1 U6411 ( .A(n6995), .Y(n6996) );
  AND2X1 U6412 ( .A(n9953), .B(n839), .Y(n868) );
  INVX1 U6413 ( .A(n868), .Y(n6997) );
  INVX1 U6414 ( .A(n7000), .Y(n6998) );
  INVX1 U6415 ( .A(n6998), .Y(n6999) );
  AND2X1 U6416 ( .A(n9956), .B(n839), .Y(n867) );
  INVX1 U6417 ( .A(n867), .Y(n7000) );
  INVX1 U6418 ( .A(n7003), .Y(n7001) );
  INVX1 U6419 ( .A(n7001), .Y(n7002) );
  AND2X1 U6420 ( .A(n9959), .B(n839), .Y(n866) );
  INVX1 U6421 ( .A(n866), .Y(n7003) );
  INVX1 U6422 ( .A(n7006), .Y(n7004) );
  INVX1 U6423 ( .A(n7004), .Y(n7005) );
  AND2X1 U6424 ( .A(n9962), .B(n839), .Y(n865) );
  INVX1 U6425 ( .A(n865), .Y(n7006) );
  INVX1 U6426 ( .A(n7009), .Y(n7007) );
  INVX1 U6427 ( .A(n7007), .Y(n7008) );
  AND2X1 U6428 ( .A(n9965), .B(n839), .Y(n864) );
  INVX1 U6429 ( .A(n864), .Y(n7009) );
  INVX1 U6430 ( .A(n7012), .Y(n7010) );
  INVX1 U6431 ( .A(n7010), .Y(n7011) );
  AND2X1 U6432 ( .A(n9968), .B(n839), .Y(n863) );
  INVX1 U6433 ( .A(n863), .Y(n7012) );
  INVX1 U6434 ( .A(n7015), .Y(n7013) );
  INVX1 U6435 ( .A(n7013), .Y(n7014) );
  AND2X1 U6436 ( .A(n9971), .B(n839), .Y(n862) );
  INVX1 U6437 ( .A(n862), .Y(n7015) );
  INVX1 U6438 ( .A(n7018), .Y(n7016) );
  INVX1 U6439 ( .A(n7016), .Y(n7017) );
  AND2X1 U6440 ( .A(n9974), .B(n839), .Y(n861) );
  INVX1 U6441 ( .A(n861), .Y(n7018) );
  INVX1 U6442 ( .A(n7021), .Y(n7019) );
  INVX1 U6443 ( .A(n7019), .Y(n7020) );
  AND2X1 U6444 ( .A(n9977), .B(n839), .Y(n860) );
  INVX1 U6445 ( .A(n860), .Y(n7021) );
  INVX1 U6446 ( .A(n7024), .Y(n7022) );
  INVX1 U6447 ( .A(n7022), .Y(n7023) );
  AND2X1 U6448 ( .A(n9980), .B(n839), .Y(n859) );
  INVX1 U6449 ( .A(n859), .Y(n7024) );
  INVX1 U6450 ( .A(n7027), .Y(n7025) );
  INVX1 U6451 ( .A(n7025), .Y(n7026) );
  AND2X1 U6452 ( .A(n9983), .B(n839), .Y(n858) );
  INVX1 U6453 ( .A(n858), .Y(n7027) );
  INVX1 U6454 ( .A(n7030), .Y(n7028) );
  INVX1 U6455 ( .A(n7028), .Y(n7029) );
  AND2X1 U6456 ( .A(n9986), .B(n839), .Y(n857) );
  INVX1 U6457 ( .A(n857), .Y(n7030) );
  INVX1 U6458 ( .A(n7033), .Y(n7031) );
  INVX1 U6459 ( .A(n7031), .Y(n7032) );
  AND2X1 U6460 ( .A(n9989), .B(n839), .Y(n856) );
  INVX1 U6461 ( .A(n856), .Y(n7033) );
  INVX1 U6462 ( .A(n7036), .Y(n7034) );
  INVX1 U6463 ( .A(n7034), .Y(n7035) );
  AND2X1 U6464 ( .A(n9992), .B(n839), .Y(n855) );
  INVX1 U6465 ( .A(n855), .Y(n7036) );
  INVX1 U6466 ( .A(n7039), .Y(n7037) );
  INVX1 U6467 ( .A(n7037), .Y(n7038) );
  AND2X1 U6468 ( .A(n9995), .B(n839), .Y(n854) );
  INVX1 U6469 ( .A(n854), .Y(n7039) );
  INVX1 U6470 ( .A(n7042), .Y(n7040) );
  INVX1 U6471 ( .A(n7040), .Y(n7041) );
  AND2X1 U6472 ( .A(n9998), .B(n839), .Y(n853) );
  INVX1 U6473 ( .A(n853), .Y(n7042) );
  INVX1 U6474 ( .A(n7045), .Y(n7043) );
  INVX1 U6475 ( .A(n7043), .Y(n7044) );
  AND2X1 U6476 ( .A(n10001), .B(n839), .Y(n852) );
  INVX1 U6477 ( .A(n852), .Y(n7045) );
  INVX1 U6478 ( .A(n7048), .Y(n7046) );
  INVX1 U6479 ( .A(n7046), .Y(n7047) );
  AND2X1 U6480 ( .A(n10004), .B(n839), .Y(n851) );
  INVX1 U6481 ( .A(n851), .Y(n7048) );
  INVX1 U6482 ( .A(n7051), .Y(n7049) );
  INVX1 U6483 ( .A(n7049), .Y(n7050) );
  AND2X1 U6484 ( .A(n10007), .B(n839), .Y(n850) );
  INVX1 U6485 ( .A(n850), .Y(n7051) );
  INVX1 U6486 ( .A(n7054), .Y(n7052) );
  INVX1 U6487 ( .A(n7052), .Y(n7053) );
  AND2X1 U6488 ( .A(n10010), .B(n839), .Y(n849) );
  INVX1 U6489 ( .A(n849), .Y(n7054) );
  INVX1 U6490 ( .A(n7057), .Y(n7055) );
  INVX1 U6491 ( .A(n7055), .Y(n7056) );
  AND2X1 U6492 ( .A(n10013), .B(n839), .Y(n848) );
  INVX1 U6493 ( .A(n848), .Y(n7057) );
  INVX1 U6494 ( .A(n7060), .Y(n7058) );
  INVX1 U6495 ( .A(n7058), .Y(n7059) );
  AND2X1 U6496 ( .A(n10016), .B(n839), .Y(n847) );
  INVX1 U6497 ( .A(n847), .Y(n7060) );
  INVX1 U6498 ( .A(n7063), .Y(n7061) );
  INVX1 U6499 ( .A(n7061), .Y(n7062) );
  AND2X1 U6500 ( .A(n10019), .B(n839), .Y(n846) );
  INVX1 U6501 ( .A(n846), .Y(n7063) );
  INVX1 U6502 ( .A(n7066), .Y(n7064) );
  INVX1 U6503 ( .A(n7064), .Y(n7065) );
  AND2X1 U6504 ( .A(n10022), .B(n839), .Y(n845) );
  INVX1 U6505 ( .A(n845), .Y(n7066) );
  INVX1 U6506 ( .A(n7069), .Y(n7067) );
  INVX1 U6507 ( .A(n7067), .Y(n7068) );
  AND2X1 U6508 ( .A(n10025), .B(n839), .Y(n844) );
  INVX1 U6509 ( .A(n844), .Y(n7069) );
  INVX1 U6510 ( .A(n7072), .Y(n7070) );
  INVX1 U6511 ( .A(n7070), .Y(n7071) );
  AND2X1 U6512 ( .A(n10028), .B(n839), .Y(n843) );
  INVX1 U6513 ( .A(n843), .Y(n7072) );
  INVX1 U6514 ( .A(n7075), .Y(n7073) );
  INVX1 U6515 ( .A(n7073), .Y(n7074) );
  AND2X1 U6516 ( .A(n10031), .B(n839), .Y(n842) );
  INVX1 U6517 ( .A(n842), .Y(n7075) );
  INVX1 U6518 ( .A(n7078), .Y(n7076) );
  INVX1 U6519 ( .A(n7076), .Y(n7077) );
  AND2X1 U6520 ( .A(n10034), .B(n839), .Y(n841) );
  INVX1 U6521 ( .A(n841), .Y(n7078) );
  INVX1 U6522 ( .A(n7081), .Y(n7079) );
  INVX1 U6523 ( .A(n7079), .Y(n7080) );
  AND2X1 U6524 ( .A(n10037), .B(n839), .Y(n840) );
  INVX1 U6525 ( .A(n840), .Y(n7081) );
  INVX1 U6526 ( .A(n7084), .Y(n7082) );
  INVX1 U6527 ( .A(n7082), .Y(n7083) );
  AND2X1 U6528 ( .A(n12064), .B(n13038), .Y(n838) );
  INVX1 U6529 ( .A(n838), .Y(n7084) );
  INVX1 U6530 ( .A(n7087), .Y(n7085) );
  INVX1 U6531 ( .A(n7085), .Y(n7086) );
  AND2X1 U6532 ( .A(n12067), .B(n13039), .Y(n837) );
  INVX1 U6533 ( .A(n837), .Y(n7087) );
  INVX1 U6534 ( .A(n7090), .Y(n7088) );
  INVX1 U6535 ( .A(n7088), .Y(n7089) );
  AND2X1 U6536 ( .A(n12070), .B(n13040), .Y(n836) );
  INVX1 U6537 ( .A(n836), .Y(n7090) );
  INVX1 U6538 ( .A(n7093), .Y(n7091) );
  INVX1 U6539 ( .A(n7091), .Y(n7092) );
  AND2X1 U6540 ( .A(n12073), .B(n13038), .Y(n835) );
  INVX1 U6541 ( .A(n835), .Y(n7093) );
  INVX1 U6542 ( .A(n7096), .Y(n7094) );
  INVX1 U6543 ( .A(n7094), .Y(n7095) );
  AND2X1 U6544 ( .A(n12076), .B(n8652), .Y(n834) );
  INVX1 U6545 ( .A(n834), .Y(n7096) );
  INVX1 U6546 ( .A(n7099), .Y(n7097) );
  INVX1 U6547 ( .A(n7097), .Y(n7098) );
  AND2X1 U6548 ( .A(n12079), .B(n8766), .Y(n833) );
  INVX1 U6549 ( .A(n833), .Y(n7099) );
  INVX1 U6550 ( .A(n7102), .Y(n7100) );
  INVX1 U6551 ( .A(n7100), .Y(n7101) );
  AND2X1 U6552 ( .A(n12082), .B(n13038), .Y(n832) );
  INVX1 U6553 ( .A(n832), .Y(n7102) );
  INVX1 U6554 ( .A(n7105), .Y(n7103) );
  INVX1 U6555 ( .A(n7103), .Y(n7104) );
  AND2X1 U6556 ( .A(n12085), .B(n8756), .Y(n831) );
  INVX1 U6557 ( .A(n831), .Y(n7105) );
  INVX1 U6558 ( .A(n7108), .Y(n7106) );
  INVX1 U6559 ( .A(n7106), .Y(n7107) );
  AND2X1 U6560 ( .A(n12088), .B(n8640), .Y(n830) );
  INVX1 U6561 ( .A(n830), .Y(n7108) );
  INVX1 U6562 ( .A(n7111), .Y(n7109) );
  INVX1 U6563 ( .A(n7109), .Y(n7110) );
  AND2X1 U6564 ( .A(n12091), .B(n13038), .Y(n829) );
  INVX1 U6565 ( .A(n829), .Y(n7111) );
  INVX1 U6566 ( .A(n7114), .Y(n7112) );
  INVX1 U6567 ( .A(n7112), .Y(n7113) );
  AND2X1 U6568 ( .A(n12094), .B(n8632), .Y(n828) );
  INVX1 U6569 ( .A(n828), .Y(n7114) );
  INVX1 U6570 ( .A(n7117), .Y(n7115) );
  INVX1 U6571 ( .A(n7115), .Y(n7116) );
  AND2X1 U6572 ( .A(n12097), .B(n8766), .Y(n827) );
  INVX1 U6573 ( .A(n827), .Y(n7117) );
  INVX1 U6574 ( .A(n7120), .Y(n7118) );
  INVX1 U6575 ( .A(n7118), .Y(n7119) );
  AND2X1 U6576 ( .A(n12100), .B(n13038), .Y(n826) );
  INVX1 U6577 ( .A(n826), .Y(n7120) );
  INVX1 U6578 ( .A(n7123), .Y(n7121) );
  INVX1 U6579 ( .A(n7121), .Y(n7122) );
  AND2X1 U6580 ( .A(n12103), .B(n13025), .Y(n825) );
  INVX1 U6581 ( .A(n825), .Y(n7123) );
  INVX1 U6582 ( .A(n7126), .Y(n7124) );
  INVX1 U6583 ( .A(n7124), .Y(n7125) );
  AND2X1 U6584 ( .A(n12106), .B(n13025), .Y(n824) );
  INVX1 U6585 ( .A(n824), .Y(n7126) );
  INVX1 U6586 ( .A(n7129), .Y(n7127) );
  INVX1 U6587 ( .A(n7127), .Y(n7128) );
  AND2X1 U6588 ( .A(n12109), .B(n13038), .Y(n823) );
  INVX1 U6589 ( .A(n823), .Y(n7129) );
  INVX1 U6590 ( .A(n7132), .Y(n7130) );
  INVX1 U6591 ( .A(n7130), .Y(n7131) );
  AND2X1 U6592 ( .A(n12112), .B(n13039), .Y(n822) );
  INVX1 U6593 ( .A(n822), .Y(n7132) );
  INVX1 U6594 ( .A(n7135), .Y(n7133) );
  INVX1 U6595 ( .A(n7133), .Y(n7134) );
  AND2X1 U6596 ( .A(n12115), .B(n8634), .Y(n821) );
  INVX1 U6597 ( .A(n821), .Y(n7135) );
  INVX1 U6598 ( .A(n7138), .Y(n7136) );
  INVX1 U6599 ( .A(n7136), .Y(n7137) );
  AND2X1 U6600 ( .A(n12118), .B(n13038), .Y(n820) );
  INVX1 U6601 ( .A(n820), .Y(n7138) );
  INVX1 U6602 ( .A(n7141), .Y(n7139) );
  INVX1 U6603 ( .A(n7139), .Y(n7140) );
  AND2X1 U6604 ( .A(n12121), .B(n8758), .Y(n819) );
  INVX1 U6605 ( .A(n819), .Y(n7141) );
  INVX1 U6606 ( .A(n7144), .Y(n7142) );
  INVX1 U6607 ( .A(n7142), .Y(n7143) );
  AND2X1 U6608 ( .A(n12124), .B(n10800), .Y(n818) );
  INVX1 U6609 ( .A(n818), .Y(n7144) );
  INVX1 U6610 ( .A(n7147), .Y(n7145) );
  INVX1 U6611 ( .A(n7145), .Y(n7146) );
  AND2X1 U6612 ( .A(n12127), .B(n13038), .Y(n817) );
  INVX1 U6613 ( .A(n817), .Y(n7147) );
  INVX1 U6614 ( .A(n7150), .Y(n7148) );
  INVX1 U6615 ( .A(n7148), .Y(n7149) );
  AND2X1 U6616 ( .A(n12130), .B(n12973), .Y(n816) );
  INVX1 U6617 ( .A(n816), .Y(n7150) );
  INVX1 U6618 ( .A(n7153), .Y(n7151) );
  INVX1 U6619 ( .A(n7151), .Y(n7152) );
  AND2X1 U6620 ( .A(n12133), .B(n13025), .Y(n815) );
  INVX1 U6621 ( .A(n815), .Y(n7153) );
  INVX1 U6622 ( .A(n7156), .Y(n7154) );
  INVX1 U6623 ( .A(n7154), .Y(n7155) );
  AND2X1 U6624 ( .A(n12136), .B(n13038), .Y(n814) );
  INVX1 U6625 ( .A(n814), .Y(n7156) );
  INVX1 U6626 ( .A(n7159), .Y(n7157) );
  INVX1 U6627 ( .A(n7157), .Y(n7158) );
  AND2X1 U6628 ( .A(n12139), .B(n8658), .Y(n813) );
  INVX1 U6629 ( .A(n813), .Y(n7159) );
  INVX1 U6630 ( .A(n7162), .Y(n7160) );
  INVX1 U6631 ( .A(n7160), .Y(n7161) );
  AND2X1 U6632 ( .A(n12142), .B(n12986), .Y(n812) );
  INVX1 U6633 ( .A(n812), .Y(n7162) );
  INVX1 U6634 ( .A(n7165), .Y(n7163) );
  INVX1 U6635 ( .A(n7163), .Y(n7164) );
  AND2X1 U6636 ( .A(n12145), .B(n13038), .Y(n811) );
  INVX1 U6637 ( .A(n811), .Y(n7165) );
  INVX1 U6638 ( .A(n7168), .Y(n7166) );
  INVX1 U6639 ( .A(n7166), .Y(n7167) );
  AND2X1 U6640 ( .A(n12148), .B(n12961), .Y(n810) );
  INVX1 U6641 ( .A(n810), .Y(n7168) );
  INVX1 U6642 ( .A(n7171), .Y(n7169) );
  INVX1 U6643 ( .A(n7169), .Y(n7170) );
  AND2X1 U6644 ( .A(n12151), .B(n12961), .Y(n809) );
  INVX1 U6645 ( .A(n809), .Y(n7171) );
  INVX1 U6646 ( .A(n7174), .Y(n7172) );
  INVX1 U6647 ( .A(n7172), .Y(n7173) );
  AND2X1 U6648 ( .A(n12154), .B(n13038), .Y(n808) );
  INVX1 U6649 ( .A(n808), .Y(n7174) );
  INVX1 U6650 ( .A(n7177), .Y(n7175) );
  INVX1 U6651 ( .A(n7175), .Y(n7176) );
  AND2X1 U6652 ( .A(n12157), .B(n12973), .Y(n807) );
  INVX1 U6653 ( .A(n807), .Y(n7177) );
  INVX1 U6654 ( .A(n7180), .Y(n7178) );
  INVX1 U6655 ( .A(n7178), .Y(n7179) );
  AND2X1 U6656 ( .A(n12160), .B(n13025), .Y(n806) );
  INVX1 U6657 ( .A(n806), .Y(n7180) );
  INVX1 U6658 ( .A(n7183), .Y(n7181) );
  INVX1 U6659 ( .A(n7181), .Y(n7182) );
  AND2X1 U6660 ( .A(n12163), .B(n13038), .Y(n805) );
  INVX1 U6661 ( .A(n805), .Y(n7183) );
  INVX1 U6662 ( .A(n7186), .Y(n7184) );
  INVX1 U6663 ( .A(n7184), .Y(n7185) );
  AND2X1 U6664 ( .A(n12166), .B(n12986), .Y(n804) );
  INVX1 U6665 ( .A(n804), .Y(n7186) );
  INVX1 U6666 ( .A(n7189), .Y(n7187) );
  INVX1 U6667 ( .A(n7187), .Y(n7188) );
  AND2X1 U6668 ( .A(n12169), .B(n13040), .Y(n803) );
  INVX1 U6669 ( .A(n803), .Y(n7189) );
  INVX1 U6670 ( .A(n7192), .Y(n7190) );
  INVX1 U6671 ( .A(n7190), .Y(n7191) );
  AND2X1 U6672 ( .A(n12172), .B(n13038), .Y(n802) );
  INVX1 U6673 ( .A(n802), .Y(n7192) );
  INVX1 U6674 ( .A(n7195), .Y(n7193) );
  INVX1 U6675 ( .A(n7193), .Y(n7194) );
  AND2X1 U6676 ( .A(n12175), .B(n13025), .Y(n801) );
  INVX1 U6677 ( .A(n801), .Y(n7195) );
  INVX1 U6678 ( .A(n7198), .Y(n7196) );
  INVX1 U6679 ( .A(n7196), .Y(n7197) );
  AND2X1 U6680 ( .A(n12178), .B(n8666), .Y(n800) );
  INVX1 U6681 ( .A(n800), .Y(n7198) );
  INVX1 U6682 ( .A(n7201), .Y(n7199) );
  INVX1 U6683 ( .A(n7199), .Y(n7200) );
  AND2X1 U6684 ( .A(n12181), .B(n13038), .Y(n799) );
  INVX1 U6685 ( .A(n799), .Y(n7201) );
  INVX1 U6686 ( .A(n7204), .Y(n7202) );
  INVX1 U6687 ( .A(n7202), .Y(n7203) );
  AND2X1 U6688 ( .A(n12184), .B(n13039), .Y(n798) );
  INVX1 U6689 ( .A(n798), .Y(n7204) );
  INVX1 U6690 ( .A(n7207), .Y(n7205) );
  INVX1 U6691 ( .A(n7205), .Y(n7206) );
  AND2X1 U6692 ( .A(n12187), .B(n13025), .Y(n797) );
  INVX1 U6693 ( .A(n797), .Y(n7207) );
  INVX1 U6694 ( .A(n7210), .Y(n7208) );
  INVX1 U6695 ( .A(n7208), .Y(n7209) );
  AND2X1 U6696 ( .A(n10040), .B(n753), .Y(n795) );
  INVX1 U6697 ( .A(n795), .Y(n7210) );
  INVX1 U6698 ( .A(n7213), .Y(n7211) );
  INVX1 U6699 ( .A(n7211), .Y(n7212) );
  AND2X1 U6700 ( .A(n10043), .B(n753), .Y(n794) );
  INVX1 U6701 ( .A(n794), .Y(n7213) );
  INVX1 U6702 ( .A(n7216), .Y(n7214) );
  INVX1 U6703 ( .A(n7214), .Y(n7215) );
  AND2X1 U6704 ( .A(n10046), .B(n753), .Y(n793) );
  INVX1 U6705 ( .A(n793), .Y(n7216) );
  INVX1 U6706 ( .A(n7219), .Y(n7217) );
  INVX1 U6707 ( .A(n7217), .Y(n7218) );
  AND2X1 U6708 ( .A(n10049), .B(n753), .Y(n792) );
  INVX1 U6709 ( .A(n792), .Y(n7219) );
  INVX1 U6710 ( .A(n7222), .Y(n7220) );
  INVX1 U6711 ( .A(n7220), .Y(n7221) );
  AND2X1 U6712 ( .A(n10052), .B(n753), .Y(n791) );
  INVX1 U6713 ( .A(n791), .Y(n7222) );
  INVX1 U6714 ( .A(n7225), .Y(n7223) );
  INVX1 U6715 ( .A(n7223), .Y(n7224) );
  AND2X1 U6716 ( .A(n10055), .B(n753), .Y(n790) );
  INVX1 U6717 ( .A(n790), .Y(n7225) );
  INVX1 U6718 ( .A(n7228), .Y(n7226) );
  INVX1 U6719 ( .A(n7226), .Y(n7227) );
  AND2X1 U6720 ( .A(n10058), .B(n753), .Y(n789) );
  INVX1 U6721 ( .A(n789), .Y(n7228) );
  INVX1 U6722 ( .A(n7231), .Y(n7229) );
  INVX1 U6723 ( .A(n7229), .Y(n7230) );
  AND2X1 U6724 ( .A(n10061), .B(n753), .Y(n788) );
  INVX1 U6725 ( .A(n788), .Y(n7231) );
  INVX1 U6726 ( .A(n7234), .Y(n7232) );
  INVX1 U6727 ( .A(n7232), .Y(n7233) );
  AND2X1 U6728 ( .A(n10064), .B(n753), .Y(n787) );
  INVX1 U6729 ( .A(n787), .Y(n7234) );
  INVX1 U6730 ( .A(n7237), .Y(n7235) );
  INVX1 U6731 ( .A(n7235), .Y(n7236) );
  AND2X1 U6732 ( .A(n10067), .B(n753), .Y(n786) );
  INVX1 U6733 ( .A(n786), .Y(n7237) );
  INVX1 U6734 ( .A(n7240), .Y(n7238) );
  INVX1 U6735 ( .A(n7238), .Y(n7239) );
  AND2X1 U6736 ( .A(n10070), .B(n753), .Y(n785) );
  INVX1 U6737 ( .A(n785), .Y(n7240) );
  INVX1 U6738 ( .A(n7243), .Y(n7241) );
  INVX1 U6739 ( .A(n7241), .Y(n7242) );
  AND2X1 U6740 ( .A(n10073), .B(n753), .Y(n784) );
  INVX1 U6741 ( .A(n784), .Y(n7243) );
  INVX1 U6742 ( .A(n7246), .Y(n7244) );
  INVX1 U6743 ( .A(n7244), .Y(n7245) );
  AND2X1 U6744 ( .A(n10076), .B(n753), .Y(n783) );
  INVX1 U6745 ( .A(n783), .Y(n7246) );
  INVX1 U6746 ( .A(n7249), .Y(n7247) );
  INVX1 U6747 ( .A(n7247), .Y(n7248) );
  AND2X1 U6748 ( .A(n10079), .B(n753), .Y(n782) );
  INVX1 U6749 ( .A(n782), .Y(n7249) );
  INVX1 U6750 ( .A(n7252), .Y(n7250) );
  INVX1 U6751 ( .A(n7250), .Y(n7251) );
  AND2X1 U6752 ( .A(n10082), .B(n753), .Y(n781) );
  INVX1 U6753 ( .A(n781), .Y(n7252) );
  INVX1 U6754 ( .A(n7255), .Y(n7253) );
  INVX1 U6755 ( .A(n7253), .Y(n7254) );
  AND2X1 U6756 ( .A(n10085), .B(n753), .Y(n780) );
  INVX1 U6757 ( .A(n780), .Y(n7255) );
  INVX1 U6758 ( .A(n7258), .Y(n7256) );
  INVX1 U6759 ( .A(n7256), .Y(n7257) );
  AND2X1 U6760 ( .A(n10088), .B(n753), .Y(n779) );
  INVX1 U6761 ( .A(n779), .Y(n7258) );
  INVX1 U6762 ( .A(n7261), .Y(n7259) );
  INVX1 U6763 ( .A(n7259), .Y(n7260) );
  AND2X1 U6764 ( .A(n10091), .B(n753), .Y(n778) );
  INVX1 U6765 ( .A(n778), .Y(n7261) );
  INVX1 U6766 ( .A(n7264), .Y(n7262) );
  INVX1 U6767 ( .A(n7262), .Y(n7263) );
  AND2X1 U6768 ( .A(n10094), .B(n753), .Y(n777) );
  INVX1 U6769 ( .A(n777), .Y(n7264) );
  INVX1 U6770 ( .A(n7267), .Y(n7265) );
  INVX1 U6771 ( .A(n7265), .Y(n7266) );
  AND2X1 U6772 ( .A(n10097), .B(n753), .Y(n776) );
  INVX1 U6773 ( .A(n776), .Y(n7267) );
  INVX1 U6774 ( .A(n7270), .Y(n7268) );
  INVX1 U6775 ( .A(n7268), .Y(n7269) );
  AND2X1 U6776 ( .A(n10100), .B(n753), .Y(n775) );
  INVX1 U6777 ( .A(n775), .Y(n7270) );
  INVX1 U6778 ( .A(n7273), .Y(n7271) );
  INVX1 U6779 ( .A(n7271), .Y(n7272) );
  AND2X1 U6780 ( .A(n10103), .B(n753), .Y(n774) );
  INVX1 U6781 ( .A(n774), .Y(n7273) );
  INVX1 U6782 ( .A(n7276), .Y(n7274) );
  INVX1 U6783 ( .A(n7274), .Y(n7275) );
  AND2X1 U6784 ( .A(n10106), .B(n753), .Y(n773) );
  INVX1 U6785 ( .A(n773), .Y(n7276) );
  INVX1 U6786 ( .A(n7279), .Y(n7277) );
  INVX1 U6787 ( .A(n7277), .Y(n7278) );
  AND2X1 U6788 ( .A(n10109), .B(n753), .Y(n772) );
  INVX1 U6789 ( .A(n772), .Y(n7279) );
  INVX1 U6790 ( .A(n7282), .Y(n7280) );
  INVX1 U6791 ( .A(n7280), .Y(n7281) );
  AND2X1 U6792 ( .A(n10112), .B(n753), .Y(n771) );
  INVX1 U6793 ( .A(n771), .Y(n7282) );
  INVX1 U6794 ( .A(n7285), .Y(n7283) );
  INVX1 U6795 ( .A(n7283), .Y(n7284) );
  AND2X1 U6796 ( .A(n10115), .B(n753), .Y(n770) );
  INVX1 U6797 ( .A(n770), .Y(n7285) );
  INVX1 U6798 ( .A(n7288), .Y(n7286) );
  INVX1 U6799 ( .A(n7286), .Y(n7287) );
  AND2X1 U6800 ( .A(n10118), .B(n753), .Y(n769) );
  INVX1 U6801 ( .A(n769), .Y(n7288) );
  INVX1 U6802 ( .A(n7291), .Y(n7289) );
  INVX1 U6803 ( .A(n7289), .Y(n7290) );
  AND2X1 U6804 ( .A(n10121), .B(n753), .Y(n768) );
  INVX1 U6805 ( .A(n768), .Y(n7291) );
  INVX1 U6806 ( .A(n7294), .Y(n7292) );
  INVX1 U6807 ( .A(n7292), .Y(n7293) );
  AND2X1 U6808 ( .A(n10124), .B(n753), .Y(n767) );
  INVX1 U6809 ( .A(n767), .Y(n7294) );
  INVX1 U6810 ( .A(n7297), .Y(n7295) );
  INVX1 U6811 ( .A(n7295), .Y(n7296) );
  AND2X1 U6812 ( .A(n10127), .B(n753), .Y(n766) );
  INVX1 U6813 ( .A(n766), .Y(n7297) );
  INVX1 U6814 ( .A(n7300), .Y(n7298) );
  INVX1 U6815 ( .A(n7298), .Y(n7299) );
  AND2X1 U6816 ( .A(n10130), .B(n753), .Y(n765) );
  INVX1 U6817 ( .A(n765), .Y(n7300) );
  INVX1 U6818 ( .A(n7303), .Y(n7301) );
  INVX1 U6819 ( .A(n7301), .Y(n7302) );
  AND2X1 U6820 ( .A(n10133), .B(n753), .Y(n764) );
  INVX1 U6821 ( .A(n764), .Y(n7303) );
  INVX1 U6822 ( .A(n7306), .Y(n7304) );
  INVX1 U6823 ( .A(n7304), .Y(n7305) );
  AND2X1 U6824 ( .A(n10136), .B(n753), .Y(n763) );
  INVX1 U6825 ( .A(n763), .Y(n7306) );
  INVX1 U6826 ( .A(n7309), .Y(n7307) );
  INVX1 U6827 ( .A(n7307), .Y(n7308) );
  AND2X1 U6828 ( .A(n10139), .B(n753), .Y(n762) );
  INVX1 U6829 ( .A(n762), .Y(n7309) );
  INVX1 U6830 ( .A(n7312), .Y(n7310) );
  INVX1 U6831 ( .A(n7310), .Y(n7311) );
  AND2X1 U6832 ( .A(n10142), .B(n753), .Y(n761) );
  INVX1 U6833 ( .A(n761), .Y(n7312) );
  INVX1 U6834 ( .A(n7315), .Y(n7313) );
  INVX1 U6835 ( .A(n7313), .Y(n7314) );
  AND2X1 U6836 ( .A(n10145), .B(n753), .Y(n760) );
  INVX1 U6837 ( .A(n760), .Y(n7315) );
  INVX1 U6838 ( .A(n7318), .Y(n7316) );
  INVX1 U6839 ( .A(n7316), .Y(n7317) );
  AND2X1 U6840 ( .A(n10148), .B(n753), .Y(n759) );
  INVX1 U6841 ( .A(n759), .Y(n7318) );
  INVX1 U6842 ( .A(n7321), .Y(n7319) );
  INVX1 U6843 ( .A(n7319), .Y(n7320) );
  AND2X1 U6844 ( .A(n10151), .B(n753), .Y(n758) );
  INVX1 U6845 ( .A(n758), .Y(n7321) );
  INVX1 U6846 ( .A(n7324), .Y(n7322) );
  INVX1 U6847 ( .A(n7322), .Y(n7323) );
  AND2X1 U6848 ( .A(n10154), .B(n753), .Y(n757) );
  INVX1 U6849 ( .A(n757), .Y(n7324) );
  INVX1 U6850 ( .A(n7327), .Y(n7325) );
  INVX1 U6851 ( .A(n7325), .Y(n7326) );
  AND2X1 U6852 ( .A(n10157), .B(n753), .Y(n756) );
  INVX1 U6853 ( .A(n756), .Y(n7327) );
  INVX1 U6854 ( .A(n7330), .Y(n7328) );
  INVX1 U6855 ( .A(n7328), .Y(n7329) );
  AND2X1 U6856 ( .A(n10160), .B(n753), .Y(n755) );
  INVX1 U6857 ( .A(n755), .Y(n7330) );
  INVX1 U6858 ( .A(n7333), .Y(n7331) );
  INVX1 U6859 ( .A(n7331), .Y(n7332) );
  AND2X1 U6860 ( .A(n10163), .B(n753), .Y(n754) );
  INVX1 U6861 ( .A(n754), .Y(n7333) );
  INVX1 U6862 ( .A(n7336), .Y(n7334) );
  INVX1 U6863 ( .A(n7334), .Y(n7335) );
  AND2X1 U6864 ( .A(n12190), .B(n710), .Y(n752) );
  INVX1 U6865 ( .A(n752), .Y(n7336) );
  INVX1 U6866 ( .A(n7339), .Y(n7337) );
  INVX1 U6867 ( .A(n7337), .Y(n7338) );
  AND2X1 U6868 ( .A(n12193), .B(n710), .Y(n751) );
  INVX1 U6869 ( .A(n751), .Y(n7339) );
  INVX1 U6870 ( .A(n7342), .Y(n7340) );
  INVX1 U6871 ( .A(n7340), .Y(n7341) );
  AND2X1 U6872 ( .A(n12196), .B(n710), .Y(n750) );
  INVX1 U6873 ( .A(n750), .Y(n7342) );
  INVX1 U6874 ( .A(n7345), .Y(n7343) );
  INVX1 U6875 ( .A(n7343), .Y(n7344) );
  AND2X1 U6876 ( .A(n12199), .B(n710), .Y(n749) );
  INVX1 U6877 ( .A(n749), .Y(n7345) );
  INVX1 U6878 ( .A(n7348), .Y(n7346) );
  INVX1 U6879 ( .A(n7346), .Y(n7347) );
  AND2X1 U6880 ( .A(n12202), .B(n710), .Y(n748) );
  INVX1 U6881 ( .A(n748), .Y(n7348) );
  INVX1 U6882 ( .A(n7351), .Y(n7349) );
  INVX1 U6883 ( .A(n7349), .Y(n7350) );
  AND2X1 U6884 ( .A(n12205), .B(n710), .Y(n747) );
  INVX1 U6885 ( .A(n747), .Y(n7351) );
  INVX1 U6886 ( .A(n7354), .Y(n7352) );
  INVX1 U6887 ( .A(n7352), .Y(n7353) );
  AND2X1 U6888 ( .A(n12208), .B(n710), .Y(n746) );
  INVX1 U6889 ( .A(n746), .Y(n7354) );
  INVX1 U6890 ( .A(n7357), .Y(n7355) );
  INVX1 U6891 ( .A(n7355), .Y(n7356) );
  AND2X1 U6892 ( .A(n12211), .B(n710), .Y(n745) );
  INVX1 U6893 ( .A(n745), .Y(n7357) );
  INVX1 U6894 ( .A(n7360), .Y(n7358) );
  INVX1 U6895 ( .A(n7358), .Y(n7359) );
  AND2X1 U6896 ( .A(n12214), .B(n710), .Y(n744) );
  INVX1 U6897 ( .A(n744), .Y(n7360) );
  INVX1 U6898 ( .A(n7363), .Y(n7361) );
  INVX1 U6899 ( .A(n7361), .Y(n7362) );
  AND2X1 U6900 ( .A(n12217), .B(n710), .Y(n743) );
  INVX1 U6901 ( .A(n743), .Y(n7363) );
  INVX1 U6902 ( .A(n7366), .Y(n7364) );
  INVX1 U6903 ( .A(n7364), .Y(n7365) );
  AND2X1 U6904 ( .A(n12220), .B(n710), .Y(n742) );
  INVX1 U6905 ( .A(n742), .Y(n7366) );
  INVX1 U6906 ( .A(n7369), .Y(n7367) );
  INVX1 U6907 ( .A(n7367), .Y(n7368) );
  AND2X1 U6908 ( .A(n12223), .B(n710), .Y(n741) );
  INVX1 U6909 ( .A(n741), .Y(n7369) );
  INVX1 U6910 ( .A(n7372), .Y(n7370) );
  INVX1 U6911 ( .A(n7370), .Y(n7371) );
  AND2X1 U6912 ( .A(n12226), .B(n710), .Y(n740) );
  INVX1 U6913 ( .A(n740), .Y(n7372) );
  INVX1 U6914 ( .A(n7375), .Y(n7373) );
  INVX1 U6915 ( .A(n7373), .Y(n7374) );
  AND2X1 U6916 ( .A(n12229), .B(n710), .Y(n739) );
  INVX1 U6917 ( .A(n739), .Y(n7375) );
  INVX1 U6918 ( .A(n7378), .Y(n7376) );
  INVX1 U6919 ( .A(n7376), .Y(n7377) );
  AND2X1 U6920 ( .A(n12232), .B(n710), .Y(n738) );
  INVX1 U6921 ( .A(n738), .Y(n7378) );
  INVX1 U6922 ( .A(n7381), .Y(n7379) );
  INVX1 U6923 ( .A(n7379), .Y(n7380) );
  AND2X1 U6924 ( .A(n12235), .B(n710), .Y(n737) );
  INVX1 U6925 ( .A(n737), .Y(n7381) );
  INVX1 U6926 ( .A(n7384), .Y(n7382) );
  INVX1 U6927 ( .A(n7382), .Y(n7383) );
  AND2X1 U6928 ( .A(n12238), .B(n710), .Y(n736) );
  INVX1 U6929 ( .A(n736), .Y(n7384) );
  INVX1 U6930 ( .A(n7387), .Y(n7385) );
  INVX1 U6931 ( .A(n7385), .Y(n7386) );
  AND2X1 U6932 ( .A(n12241), .B(n710), .Y(n735) );
  INVX1 U6933 ( .A(n735), .Y(n7387) );
  INVX1 U6934 ( .A(n7390), .Y(n7388) );
  INVX1 U6935 ( .A(n7388), .Y(n7389) );
  AND2X1 U6936 ( .A(n12244), .B(n710), .Y(n734) );
  INVX1 U6937 ( .A(n734), .Y(n7390) );
  INVX1 U6938 ( .A(n7393), .Y(n7391) );
  INVX1 U6939 ( .A(n7391), .Y(n7392) );
  AND2X1 U6940 ( .A(n12247), .B(n710), .Y(n733) );
  INVX1 U6941 ( .A(n733), .Y(n7393) );
  INVX1 U6942 ( .A(n7396), .Y(n7394) );
  INVX1 U6943 ( .A(n7394), .Y(n7395) );
  AND2X1 U6944 ( .A(n12250), .B(n710), .Y(n732) );
  INVX1 U6945 ( .A(n732), .Y(n7396) );
  INVX1 U6946 ( .A(n7399), .Y(n7397) );
  INVX1 U6947 ( .A(n7397), .Y(n7398) );
  AND2X1 U6948 ( .A(n12253), .B(n710), .Y(n731) );
  INVX1 U6949 ( .A(n731), .Y(n7399) );
  INVX1 U6950 ( .A(n7402), .Y(n7400) );
  INVX1 U6951 ( .A(n7400), .Y(n7401) );
  AND2X1 U6952 ( .A(n12256), .B(n710), .Y(n730) );
  INVX1 U6953 ( .A(n730), .Y(n7402) );
  INVX1 U6954 ( .A(n7405), .Y(n7403) );
  INVX1 U6955 ( .A(n7403), .Y(n7404) );
  AND2X1 U6956 ( .A(n12259), .B(n710), .Y(n729) );
  INVX1 U6957 ( .A(n729), .Y(n7405) );
  INVX1 U6958 ( .A(n7408), .Y(n7406) );
  INVX1 U6959 ( .A(n7406), .Y(n7407) );
  AND2X1 U6960 ( .A(n12262), .B(n710), .Y(n728) );
  INVX1 U6961 ( .A(n728), .Y(n7408) );
  INVX1 U6962 ( .A(n7411), .Y(n7409) );
  INVX1 U6963 ( .A(n7409), .Y(n7410) );
  AND2X1 U6964 ( .A(n12265), .B(n710), .Y(n727) );
  INVX1 U6965 ( .A(n727), .Y(n7411) );
  INVX1 U6966 ( .A(n7414), .Y(n7412) );
  INVX1 U6967 ( .A(n7412), .Y(n7413) );
  AND2X1 U6968 ( .A(n12268), .B(n710), .Y(n726) );
  INVX1 U6969 ( .A(n726), .Y(n7414) );
  INVX1 U6970 ( .A(n7417), .Y(n7415) );
  INVX1 U6971 ( .A(n7415), .Y(n7416) );
  AND2X1 U6972 ( .A(n12271), .B(n710), .Y(n725) );
  INVX1 U6973 ( .A(n725), .Y(n7417) );
  INVX1 U6974 ( .A(n7420), .Y(n7418) );
  INVX1 U6975 ( .A(n7418), .Y(n7419) );
  AND2X1 U6976 ( .A(n12274), .B(n710), .Y(n724) );
  INVX1 U6977 ( .A(n724), .Y(n7420) );
  INVX1 U6978 ( .A(n7423), .Y(n7421) );
  INVX1 U6979 ( .A(n7421), .Y(n7422) );
  AND2X1 U6980 ( .A(n12277), .B(n710), .Y(n723) );
  INVX1 U6981 ( .A(n723), .Y(n7423) );
  INVX1 U6982 ( .A(n7426), .Y(n7424) );
  INVX1 U6983 ( .A(n7424), .Y(n7425) );
  AND2X1 U6984 ( .A(n12280), .B(n710), .Y(n722) );
  INVX1 U6985 ( .A(n722), .Y(n7426) );
  INVX1 U6986 ( .A(n7429), .Y(n7427) );
  INVX1 U6987 ( .A(n7427), .Y(n7428) );
  AND2X1 U6988 ( .A(n12283), .B(n710), .Y(n721) );
  INVX1 U6989 ( .A(n721), .Y(n7429) );
  INVX1 U6990 ( .A(n7432), .Y(n7430) );
  INVX1 U6991 ( .A(n7430), .Y(n7431) );
  AND2X1 U6992 ( .A(n12286), .B(n710), .Y(n720) );
  INVX1 U6993 ( .A(n720), .Y(n7432) );
  INVX1 U6994 ( .A(n7435), .Y(n7433) );
  INVX1 U6995 ( .A(n7433), .Y(n7434) );
  AND2X1 U6996 ( .A(n12289), .B(n710), .Y(n719) );
  INVX1 U6997 ( .A(n719), .Y(n7435) );
  INVX1 U6998 ( .A(n7438), .Y(n7436) );
  INVX1 U6999 ( .A(n7436), .Y(n7437) );
  AND2X1 U7000 ( .A(n12292), .B(n710), .Y(n718) );
  INVX1 U7001 ( .A(n718), .Y(n7438) );
  INVX1 U7002 ( .A(n7441), .Y(n7439) );
  INVX1 U7003 ( .A(n7439), .Y(n7440) );
  AND2X1 U7004 ( .A(n12295), .B(n710), .Y(n717) );
  INVX1 U7005 ( .A(n717), .Y(n7441) );
  INVX1 U7006 ( .A(n7444), .Y(n7442) );
  INVX1 U7007 ( .A(n7442), .Y(n7443) );
  AND2X1 U7008 ( .A(n12298), .B(n710), .Y(n716) );
  INVX1 U7009 ( .A(n716), .Y(n7444) );
  INVX1 U7010 ( .A(n7447), .Y(n7445) );
  INVX1 U7011 ( .A(n7445), .Y(n7446) );
  AND2X1 U7012 ( .A(n12301), .B(n710), .Y(n715) );
  INVX1 U7013 ( .A(n715), .Y(n7447) );
  INVX1 U7014 ( .A(n7450), .Y(n7448) );
  INVX1 U7015 ( .A(n7448), .Y(n7449) );
  AND2X1 U7016 ( .A(n12304), .B(n710), .Y(n714) );
  INVX1 U7017 ( .A(n714), .Y(n7450) );
  INVX1 U7018 ( .A(n7453), .Y(n7451) );
  INVX1 U7019 ( .A(n7451), .Y(n7452) );
  AND2X1 U7020 ( .A(n12307), .B(n710), .Y(n713) );
  INVX1 U7021 ( .A(n713), .Y(n7453) );
  INVX1 U7022 ( .A(n7456), .Y(n7454) );
  INVX1 U7023 ( .A(n7454), .Y(n7455) );
  AND2X1 U7024 ( .A(n12310), .B(n710), .Y(n712) );
  INVX1 U7025 ( .A(n712), .Y(n7456) );
  INVX1 U7026 ( .A(n7459), .Y(n7457) );
  INVX1 U7027 ( .A(n7457), .Y(n7458) );
  AND2X1 U7028 ( .A(n12313), .B(n710), .Y(n711) );
  INVX1 U7029 ( .A(n711), .Y(n7459) );
  INVX1 U7030 ( .A(n7462), .Y(n7460) );
  INVX1 U7031 ( .A(n7460), .Y(n7461) );
  AND2X1 U7032 ( .A(n10166), .B(n666), .Y(n708) );
  INVX1 U7033 ( .A(n708), .Y(n7462) );
  INVX1 U7034 ( .A(n7465), .Y(n7463) );
  INVX1 U7035 ( .A(n7463), .Y(n7464) );
  AND2X1 U7036 ( .A(n10169), .B(n666), .Y(n707) );
  INVX1 U7037 ( .A(n707), .Y(n7465) );
  INVX1 U7038 ( .A(n7468), .Y(n7466) );
  INVX1 U7039 ( .A(n7466), .Y(n7467) );
  AND2X1 U7040 ( .A(n10172), .B(n666), .Y(n706) );
  INVX1 U7041 ( .A(n706), .Y(n7468) );
  INVX1 U7042 ( .A(n7471), .Y(n7469) );
  INVX1 U7043 ( .A(n7469), .Y(n7470) );
  AND2X1 U7044 ( .A(n10175), .B(n666), .Y(n705) );
  INVX1 U7045 ( .A(n705), .Y(n7471) );
  INVX1 U7046 ( .A(n7474), .Y(n7472) );
  INVX1 U7047 ( .A(n7472), .Y(n7473) );
  AND2X1 U7048 ( .A(n10178), .B(n666), .Y(n704) );
  INVX1 U7049 ( .A(n704), .Y(n7474) );
  INVX1 U7050 ( .A(n7477), .Y(n7475) );
  INVX1 U7051 ( .A(n7475), .Y(n7476) );
  AND2X1 U7052 ( .A(n10181), .B(n666), .Y(n703) );
  INVX1 U7053 ( .A(n703), .Y(n7477) );
  INVX1 U7054 ( .A(n7480), .Y(n7478) );
  INVX1 U7055 ( .A(n7478), .Y(n7479) );
  AND2X1 U7056 ( .A(n10184), .B(n666), .Y(n702) );
  INVX1 U7057 ( .A(n702), .Y(n7480) );
  INVX1 U7058 ( .A(n7483), .Y(n7481) );
  INVX1 U7059 ( .A(n7481), .Y(n7482) );
  AND2X1 U7060 ( .A(n10187), .B(n666), .Y(n701) );
  INVX1 U7061 ( .A(n701), .Y(n7483) );
  INVX1 U7062 ( .A(n7486), .Y(n7484) );
  INVX1 U7063 ( .A(n7484), .Y(n7485) );
  AND2X1 U7064 ( .A(n10190), .B(n666), .Y(n700) );
  INVX1 U7065 ( .A(n700), .Y(n7486) );
  INVX1 U7066 ( .A(n7489), .Y(n7487) );
  INVX1 U7067 ( .A(n7487), .Y(n7488) );
  AND2X1 U7068 ( .A(n10193), .B(n666), .Y(n699) );
  INVX1 U7069 ( .A(n699), .Y(n7489) );
  INVX1 U7070 ( .A(n7492), .Y(n7490) );
  INVX1 U7071 ( .A(n7490), .Y(n7491) );
  AND2X1 U7072 ( .A(n10196), .B(n666), .Y(n698) );
  INVX1 U7073 ( .A(n698), .Y(n7492) );
  INVX1 U7074 ( .A(n7495), .Y(n7493) );
  INVX1 U7075 ( .A(n7493), .Y(n7494) );
  AND2X1 U7076 ( .A(n10199), .B(n666), .Y(n697) );
  INVX1 U7077 ( .A(n697), .Y(n7495) );
  INVX1 U7078 ( .A(n7498), .Y(n7496) );
  INVX1 U7079 ( .A(n7496), .Y(n7497) );
  AND2X1 U7080 ( .A(n10202), .B(n666), .Y(n696) );
  INVX1 U7081 ( .A(n696), .Y(n7498) );
  INVX1 U7082 ( .A(n7501), .Y(n7499) );
  INVX1 U7083 ( .A(n7499), .Y(n7500) );
  AND2X1 U7084 ( .A(n10205), .B(n666), .Y(n695) );
  INVX1 U7085 ( .A(n695), .Y(n7501) );
  INVX1 U7086 ( .A(n7504), .Y(n7502) );
  INVX1 U7087 ( .A(n7502), .Y(n7503) );
  AND2X1 U7088 ( .A(n10208), .B(n666), .Y(n694) );
  INVX1 U7089 ( .A(n694), .Y(n7504) );
  INVX1 U7090 ( .A(n7507), .Y(n7505) );
  INVX1 U7091 ( .A(n7505), .Y(n7506) );
  AND2X1 U7092 ( .A(n10211), .B(n666), .Y(n693) );
  INVX1 U7093 ( .A(n693), .Y(n7507) );
  INVX1 U7094 ( .A(n7510), .Y(n7508) );
  INVX1 U7095 ( .A(n7508), .Y(n7509) );
  AND2X1 U7096 ( .A(n10214), .B(n666), .Y(n692) );
  INVX1 U7097 ( .A(n692), .Y(n7510) );
  INVX1 U7098 ( .A(n7513), .Y(n7511) );
  INVX1 U7099 ( .A(n7511), .Y(n7512) );
  AND2X1 U7100 ( .A(n10217), .B(n666), .Y(n691) );
  INVX1 U7101 ( .A(n691), .Y(n7513) );
  INVX1 U7102 ( .A(n7516), .Y(n7514) );
  INVX1 U7103 ( .A(n7514), .Y(n7515) );
  AND2X1 U7104 ( .A(n10220), .B(n666), .Y(n690) );
  INVX1 U7105 ( .A(n690), .Y(n7516) );
  INVX1 U7106 ( .A(n7519), .Y(n7517) );
  INVX1 U7107 ( .A(n7517), .Y(n7518) );
  AND2X1 U7108 ( .A(n10223), .B(n666), .Y(n689) );
  INVX1 U7109 ( .A(n689), .Y(n7519) );
  INVX1 U7110 ( .A(n7522), .Y(n7520) );
  INVX1 U7111 ( .A(n7520), .Y(n7521) );
  AND2X1 U7112 ( .A(n10226), .B(n666), .Y(n688) );
  INVX1 U7113 ( .A(n688), .Y(n7522) );
  INVX1 U7114 ( .A(n7525), .Y(n7523) );
  INVX1 U7115 ( .A(n7523), .Y(n7524) );
  AND2X1 U7116 ( .A(n10229), .B(n666), .Y(n687) );
  INVX1 U7117 ( .A(n687), .Y(n7525) );
  INVX1 U7118 ( .A(n7528), .Y(n7526) );
  INVX1 U7119 ( .A(n7526), .Y(n7527) );
  AND2X1 U7120 ( .A(n10232), .B(n666), .Y(n686) );
  INVX1 U7121 ( .A(n686), .Y(n7528) );
  INVX1 U7122 ( .A(n7531), .Y(n7529) );
  INVX1 U7123 ( .A(n7529), .Y(n7530) );
  AND2X1 U7124 ( .A(n10235), .B(n666), .Y(n685) );
  INVX1 U7125 ( .A(n685), .Y(n7531) );
  INVX1 U7126 ( .A(n7534), .Y(n7532) );
  INVX1 U7127 ( .A(n7532), .Y(n7533) );
  AND2X1 U7128 ( .A(n10238), .B(n666), .Y(n684) );
  INVX1 U7129 ( .A(n684), .Y(n7534) );
  INVX1 U7130 ( .A(n7537), .Y(n7535) );
  INVX1 U7131 ( .A(n7535), .Y(n7536) );
  AND2X1 U7132 ( .A(n10241), .B(n666), .Y(n683) );
  INVX1 U7133 ( .A(n683), .Y(n7537) );
  INVX1 U7134 ( .A(n7540), .Y(n7538) );
  INVX1 U7135 ( .A(n7538), .Y(n7539) );
  AND2X1 U7136 ( .A(n10244), .B(n666), .Y(n682) );
  INVX1 U7137 ( .A(n682), .Y(n7540) );
  INVX1 U7138 ( .A(n7543), .Y(n7541) );
  INVX1 U7139 ( .A(n7541), .Y(n7542) );
  AND2X1 U7140 ( .A(n10247), .B(n666), .Y(n681) );
  INVX1 U7141 ( .A(n681), .Y(n7543) );
  INVX1 U7142 ( .A(n7546), .Y(n7544) );
  INVX1 U7143 ( .A(n7544), .Y(n7545) );
  AND2X1 U7144 ( .A(n10250), .B(n666), .Y(n680) );
  INVX1 U7145 ( .A(n680), .Y(n7546) );
  INVX1 U7146 ( .A(n7549), .Y(n7547) );
  INVX1 U7147 ( .A(n7547), .Y(n7548) );
  AND2X1 U7148 ( .A(n10253), .B(n666), .Y(n679) );
  INVX1 U7149 ( .A(n679), .Y(n7549) );
  INVX1 U7150 ( .A(n7552), .Y(n7550) );
  INVX1 U7151 ( .A(n7550), .Y(n7551) );
  AND2X1 U7152 ( .A(n10256), .B(n666), .Y(n678) );
  INVX1 U7153 ( .A(n678), .Y(n7552) );
  INVX1 U7154 ( .A(n7555), .Y(n7553) );
  INVX1 U7155 ( .A(n7553), .Y(n7554) );
  AND2X1 U7156 ( .A(n10259), .B(n666), .Y(n677) );
  INVX1 U7157 ( .A(n677), .Y(n7555) );
  INVX1 U7158 ( .A(n7558), .Y(n7556) );
  INVX1 U7159 ( .A(n7556), .Y(n7557) );
  AND2X1 U7160 ( .A(n10262), .B(n666), .Y(n676) );
  INVX1 U7161 ( .A(n676), .Y(n7558) );
  INVX1 U7162 ( .A(n7561), .Y(n7559) );
  INVX1 U7163 ( .A(n7559), .Y(n7560) );
  AND2X1 U7164 ( .A(n10265), .B(n666), .Y(n675) );
  INVX1 U7165 ( .A(n675), .Y(n7561) );
  INVX1 U7166 ( .A(n7564), .Y(n7562) );
  INVX1 U7167 ( .A(n7562), .Y(n7563) );
  AND2X1 U7168 ( .A(n10268), .B(n666), .Y(n674) );
  INVX1 U7169 ( .A(n674), .Y(n7564) );
  INVX1 U7170 ( .A(n7567), .Y(n7565) );
  INVX1 U7171 ( .A(n7565), .Y(n7566) );
  AND2X1 U7172 ( .A(n10271), .B(n666), .Y(n673) );
  INVX1 U7173 ( .A(n673), .Y(n7567) );
  INVX1 U7174 ( .A(n7570), .Y(n7568) );
  INVX1 U7175 ( .A(n7568), .Y(n7569) );
  AND2X1 U7176 ( .A(n10274), .B(n666), .Y(n672) );
  INVX1 U7177 ( .A(n672), .Y(n7570) );
  INVX1 U7178 ( .A(n7573), .Y(n7571) );
  INVX1 U7179 ( .A(n7571), .Y(n7572) );
  AND2X1 U7180 ( .A(n10277), .B(n666), .Y(n671) );
  INVX1 U7181 ( .A(n671), .Y(n7573) );
  INVX1 U7182 ( .A(n7576), .Y(n7574) );
  INVX1 U7183 ( .A(n7574), .Y(n7575) );
  AND2X1 U7184 ( .A(n10280), .B(n666), .Y(n670) );
  INVX1 U7185 ( .A(n670), .Y(n7576) );
  INVX1 U7186 ( .A(n7579), .Y(n7577) );
  INVX1 U7187 ( .A(n7577), .Y(n7578) );
  AND2X1 U7188 ( .A(n10283), .B(n666), .Y(n669) );
  INVX1 U7189 ( .A(n669), .Y(n7579) );
  INVX1 U7190 ( .A(n7582), .Y(n7580) );
  INVX1 U7191 ( .A(n7580), .Y(n7581) );
  AND2X1 U7192 ( .A(n10286), .B(n666), .Y(n668) );
  INVX1 U7193 ( .A(n668), .Y(n7582) );
  INVX1 U7194 ( .A(n7585), .Y(n7583) );
  INVX1 U7195 ( .A(n7583), .Y(n7584) );
  AND2X1 U7196 ( .A(n10289), .B(n666), .Y(n667) );
  INVX1 U7197 ( .A(n667), .Y(n7585) );
  INVX1 U7198 ( .A(n7588), .Y(n7586) );
  INVX1 U7199 ( .A(n7586), .Y(n7587) );
  AND2X1 U7200 ( .A(n12316), .B(n621), .Y(n663) );
  INVX1 U7201 ( .A(n663), .Y(n7588) );
  INVX1 U7202 ( .A(n7591), .Y(n7589) );
  INVX1 U7203 ( .A(n7589), .Y(n7590) );
  AND2X1 U7204 ( .A(n12319), .B(n621), .Y(n662) );
  INVX1 U7205 ( .A(n662), .Y(n7591) );
  INVX1 U7206 ( .A(n7594), .Y(n7592) );
  INVX1 U7207 ( .A(n7592), .Y(n7593) );
  AND2X1 U7208 ( .A(n12322), .B(n621), .Y(n661) );
  INVX1 U7209 ( .A(n661), .Y(n7594) );
  INVX1 U7210 ( .A(n7597), .Y(n7595) );
  INVX1 U7211 ( .A(n7595), .Y(n7596) );
  AND2X1 U7212 ( .A(n12325), .B(n621), .Y(n660) );
  INVX1 U7213 ( .A(n660), .Y(n7597) );
  INVX1 U7214 ( .A(n7600), .Y(n7598) );
  INVX1 U7215 ( .A(n7598), .Y(n7599) );
  AND2X1 U7216 ( .A(n12328), .B(n621), .Y(n659) );
  INVX1 U7217 ( .A(n659), .Y(n7600) );
  INVX1 U7218 ( .A(n7603), .Y(n7601) );
  INVX1 U7219 ( .A(n7601), .Y(n7602) );
  AND2X1 U7220 ( .A(n12331), .B(n621), .Y(n658) );
  INVX1 U7221 ( .A(n658), .Y(n7603) );
  INVX1 U7222 ( .A(n7606), .Y(n7604) );
  INVX1 U7223 ( .A(n7604), .Y(n7605) );
  AND2X1 U7224 ( .A(n12334), .B(n621), .Y(n657) );
  INVX1 U7225 ( .A(n657), .Y(n7606) );
  INVX1 U7226 ( .A(n7609), .Y(n7607) );
  INVX1 U7227 ( .A(n7607), .Y(n7608) );
  AND2X1 U7228 ( .A(n12337), .B(n621), .Y(n656) );
  INVX1 U7229 ( .A(n656), .Y(n7609) );
  INVX1 U7230 ( .A(n7612), .Y(n7610) );
  INVX1 U7231 ( .A(n7610), .Y(n7611) );
  AND2X1 U7232 ( .A(n12340), .B(n621), .Y(n655) );
  INVX1 U7233 ( .A(n655), .Y(n7612) );
  INVX1 U7234 ( .A(n7615), .Y(n7613) );
  INVX1 U7235 ( .A(n7613), .Y(n7614) );
  AND2X1 U7236 ( .A(n12343), .B(n621), .Y(n654) );
  INVX1 U7237 ( .A(n654), .Y(n7615) );
  INVX1 U7238 ( .A(n7618), .Y(n7616) );
  INVX1 U7239 ( .A(n7616), .Y(n7617) );
  AND2X1 U7240 ( .A(n12346), .B(n621), .Y(n653) );
  INVX1 U7241 ( .A(n653), .Y(n7618) );
  INVX1 U7242 ( .A(n7621), .Y(n7619) );
  INVX1 U7243 ( .A(n7619), .Y(n7620) );
  AND2X1 U7244 ( .A(n12349), .B(n621), .Y(n652) );
  INVX1 U7245 ( .A(n652), .Y(n7621) );
  INVX1 U7246 ( .A(n7624), .Y(n7622) );
  INVX1 U7247 ( .A(n7622), .Y(n7623) );
  AND2X1 U7248 ( .A(n12352), .B(n621), .Y(n651) );
  INVX1 U7249 ( .A(n651), .Y(n7624) );
  INVX1 U7250 ( .A(n7627), .Y(n7625) );
  INVX1 U7251 ( .A(n7625), .Y(n7626) );
  AND2X1 U7252 ( .A(n12355), .B(n621), .Y(n650) );
  INVX1 U7253 ( .A(n650), .Y(n7627) );
  INVX1 U7254 ( .A(n7630), .Y(n7628) );
  INVX1 U7255 ( .A(n7628), .Y(n7629) );
  AND2X1 U7256 ( .A(n12358), .B(n621), .Y(n649) );
  INVX1 U7257 ( .A(n649), .Y(n7630) );
  INVX1 U7258 ( .A(n7633), .Y(n7631) );
  INVX1 U7259 ( .A(n7631), .Y(n7632) );
  AND2X1 U7260 ( .A(n12361), .B(n621), .Y(n648) );
  INVX1 U7261 ( .A(n648), .Y(n7633) );
  INVX1 U7262 ( .A(n7636), .Y(n7634) );
  INVX1 U7263 ( .A(n7634), .Y(n7635) );
  AND2X1 U7264 ( .A(n12364), .B(n621), .Y(n647) );
  INVX1 U7265 ( .A(n647), .Y(n7636) );
  INVX1 U7266 ( .A(n7639), .Y(n7637) );
  INVX1 U7267 ( .A(n7637), .Y(n7638) );
  AND2X1 U7268 ( .A(n12367), .B(n621), .Y(n646) );
  INVX1 U7269 ( .A(n646), .Y(n7639) );
  INVX1 U7270 ( .A(n7642), .Y(n7640) );
  INVX1 U7271 ( .A(n7640), .Y(n7641) );
  AND2X1 U7272 ( .A(n12370), .B(n621), .Y(n645) );
  INVX1 U7273 ( .A(n645), .Y(n7642) );
  INVX1 U7274 ( .A(n7645), .Y(n7643) );
  INVX1 U7275 ( .A(n7643), .Y(n7644) );
  AND2X1 U7276 ( .A(n12373), .B(n621), .Y(n644) );
  INVX1 U7277 ( .A(n644), .Y(n7645) );
  INVX1 U7278 ( .A(n7648), .Y(n7646) );
  INVX1 U7279 ( .A(n7646), .Y(n7647) );
  AND2X1 U7280 ( .A(n12376), .B(n621), .Y(n643) );
  INVX1 U7281 ( .A(n643), .Y(n7648) );
  INVX1 U7282 ( .A(n7651), .Y(n7649) );
  INVX1 U7283 ( .A(n7649), .Y(n7650) );
  AND2X1 U7284 ( .A(n12379), .B(n621), .Y(n642) );
  INVX1 U7285 ( .A(n642), .Y(n7651) );
  INVX1 U7286 ( .A(n7654), .Y(n7652) );
  INVX1 U7287 ( .A(n7652), .Y(n7653) );
  AND2X1 U7288 ( .A(n12382), .B(n621), .Y(n641) );
  INVX1 U7289 ( .A(n641), .Y(n7654) );
  INVX1 U7290 ( .A(n7657), .Y(n7655) );
  INVX1 U7291 ( .A(n7655), .Y(n7656) );
  AND2X1 U7292 ( .A(n12385), .B(n621), .Y(n640) );
  INVX1 U7293 ( .A(n640), .Y(n7657) );
  INVX1 U7294 ( .A(n7660), .Y(n7658) );
  INVX1 U7295 ( .A(n7658), .Y(n7659) );
  AND2X1 U7296 ( .A(n12388), .B(n621), .Y(n639) );
  INVX1 U7297 ( .A(n639), .Y(n7660) );
  INVX1 U7298 ( .A(n7663), .Y(n7661) );
  INVX1 U7299 ( .A(n7661), .Y(n7662) );
  AND2X1 U7300 ( .A(n12391), .B(n621), .Y(n638) );
  INVX1 U7301 ( .A(n638), .Y(n7663) );
  INVX1 U7302 ( .A(n7666), .Y(n7664) );
  INVX1 U7303 ( .A(n7664), .Y(n7665) );
  AND2X1 U7304 ( .A(n12394), .B(n621), .Y(n637) );
  INVX1 U7305 ( .A(n637), .Y(n7666) );
  INVX1 U7306 ( .A(n7669), .Y(n7667) );
  INVX1 U7307 ( .A(n7667), .Y(n7668) );
  AND2X1 U7308 ( .A(n12397), .B(n621), .Y(n636) );
  INVX1 U7309 ( .A(n636), .Y(n7669) );
  INVX1 U7310 ( .A(n7672), .Y(n7670) );
  INVX1 U7311 ( .A(n7670), .Y(n7671) );
  AND2X1 U7312 ( .A(n12400), .B(n621), .Y(n635) );
  INVX1 U7313 ( .A(n635), .Y(n7672) );
  INVX1 U7314 ( .A(n7675), .Y(n7673) );
  INVX1 U7315 ( .A(n7673), .Y(n7674) );
  AND2X1 U7316 ( .A(n12403), .B(n621), .Y(n634) );
  INVX1 U7317 ( .A(n634), .Y(n7675) );
  INVX1 U7318 ( .A(n7678), .Y(n7676) );
  INVX1 U7319 ( .A(n7676), .Y(n7677) );
  AND2X1 U7320 ( .A(n12406), .B(n621), .Y(n633) );
  INVX1 U7321 ( .A(n633), .Y(n7678) );
  INVX1 U7322 ( .A(n7681), .Y(n7679) );
  INVX1 U7323 ( .A(n7679), .Y(n7680) );
  AND2X1 U7324 ( .A(n12409), .B(n621), .Y(n632) );
  INVX1 U7325 ( .A(n632), .Y(n7681) );
  INVX1 U7326 ( .A(n7684), .Y(n7682) );
  INVX1 U7327 ( .A(n7682), .Y(n7683) );
  AND2X1 U7328 ( .A(n12412), .B(n621), .Y(n631) );
  INVX1 U7329 ( .A(n631), .Y(n7684) );
  INVX1 U7330 ( .A(n7687), .Y(n7685) );
  INVX1 U7331 ( .A(n7685), .Y(n7686) );
  AND2X1 U7332 ( .A(n12415), .B(n621), .Y(n630) );
  INVX1 U7333 ( .A(n630), .Y(n7687) );
  INVX1 U7334 ( .A(n7690), .Y(n7688) );
  INVX1 U7335 ( .A(n7688), .Y(n7689) );
  AND2X1 U7336 ( .A(n12418), .B(n621), .Y(n629) );
  INVX1 U7337 ( .A(n629), .Y(n7690) );
  INVX1 U7338 ( .A(n7693), .Y(n7691) );
  INVX1 U7339 ( .A(n7691), .Y(n7692) );
  AND2X1 U7340 ( .A(n12421), .B(n621), .Y(n628) );
  INVX1 U7341 ( .A(n628), .Y(n7693) );
  INVX1 U7342 ( .A(n7696), .Y(n7694) );
  INVX1 U7343 ( .A(n7694), .Y(n7695) );
  AND2X1 U7344 ( .A(n12424), .B(n621), .Y(n627) );
  INVX1 U7345 ( .A(n627), .Y(n7696) );
  INVX1 U7346 ( .A(n7699), .Y(n7697) );
  INVX1 U7347 ( .A(n7697), .Y(n7698) );
  AND2X1 U7348 ( .A(n12427), .B(n621), .Y(n626) );
  INVX1 U7349 ( .A(n626), .Y(n7699) );
  INVX1 U7350 ( .A(n7702), .Y(n7700) );
  INVX1 U7351 ( .A(n7700), .Y(n7701) );
  AND2X1 U7352 ( .A(n12430), .B(n621), .Y(n625) );
  INVX1 U7353 ( .A(n625), .Y(n7702) );
  INVX1 U7354 ( .A(n7705), .Y(n7703) );
  INVX1 U7355 ( .A(n7703), .Y(n7704) );
  AND2X1 U7356 ( .A(n12433), .B(n621), .Y(n624) );
  INVX1 U7357 ( .A(n624), .Y(n7705) );
  INVX1 U7358 ( .A(n7708), .Y(n7706) );
  INVX1 U7359 ( .A(n7706), .Y(n7707) );
  AND2X1 U7360 ( .A(n12436), .B(n621), .Y(n623) );
  INVX1 U7361 ( .A(n623), .Y(n7708) );
  INVX1 U7362 ( .A(n7711), .Y(n7709) );
  INVX1 U7363 ( .A(n7709), .Y(n7710) );
  AND2X1 U7364 ( .A(n12439), .B(n621), .Y(n622) );
  INVX1 U7365 ( .A(n622), .Y(n7711) );
  INVX1 U7366 ( .A(n7714), .Y(n7712) );
  INVX1 U7367 ( .A(n7712), .Y(n7713) );
  AND2X1 U7368 ( .A(n10292), .B(n577), .Y(n619) );
  INVX1 U7369 ( .A(n619), .Y(n7714) );
  INVX1 U7370 ( .A(n7717), .Y(n7715) );
  INVX1 U7371 ( .A(n7715), .Y(n7716) );
  AND2X1 U7372 ( .A(n10295), .B(n577), .Y(n618) );
  INVX1 U7373 ( .A(n618), .Y(n7717) );
  INVX1 U7374 ( .A(n7720), .Y(n7718) );
  INVX1 U7375 ( .A(n7718), .Y(n7719) );
  AND2X1 U7376 ( .A(n10298), .B(n577), .Y(n617) );
  INVX1 U7377 ( .A(n617), .Y(n7720) );
  INVX1 U7378 ( .A(n7723), .Y(n7721) );
  INVX1 U7379 ( .A(n7721), .Y(n7722) );
  AND2X1 U7380 ( .A(n10301), .B(n577), .Y(n616) );
  INVX1 U7381 ( .A(n616), .Y(n7723) );
  INVX1 U7382 ( .A(n7726), .Y(n7724) );
  INVX1 U7383 ( .A(n7724), .Y(n7725) );
  AND2X1 U7384 ( .A(n10304), .B(n577), .Y(n615) );
  INVX1 U7385 ( .A(n615), .Y(n7726) );
  INVX1 U7386 ( .A(n7729), .Y(n7727) );
  INVX1 U7387 ( .A(n7727), .Y(n7728) );
  AND2X1 U7388 ( .A(n10307), .B(n577), .Y(n614) );
  INVX1 U7389 ( .A(n614), .Y(n7729) );
  INVX1 U7390 ( .A(n7732), .Y(n7730) );
  INVX1 U7391 ( .A(n7730), .Y(n7731) );
  AND2X1 U7392 ( .A(n10310), .B(n577), .Y(n613) );
  INVX1 U7393 ( .A(n613), .Y(n7732) );
  INVX1 U7394 ( .A(n7735), .Y(n7733) );
  INVX1 U7395 ( .A(n7733), .Y(n7734) );
  AND2X1 U7396 ( .A(n10313), .B(n577), .Y(n612) );
  INVX1 U7397 ( .A(n612), .Y(n7735) );
  INVX1 U7398 ( .A(n7738), .Y(n7736) );
  INVX1 U7399 ( .A(n7736), .Y(n7737) );
  AND2X1 U7400 ( .A(n10316), .B(n577), .Y(n611) );
  INVX1 U7401 ( .A(n611), .Y(n7738) );
  INVX1 U7402 ( .A(n7741), .Y(n7739) );
  INVX1 U7403 ( .A(n7739), .Y(n7740) );
  AND2X1 U7404 ( .A(n10319), .B(n577), .Y(n610) );
  INVX1 U7405 ( .A(n610), .Y(n7741) );
  INVX1 U7406 ( .A(n7744), .Y(n7742) );
  INVX1 U7407 ( .A(n7742), .Y(n7743) );
  AND2X1 U7408 ( .A(n10322), .B(n577), .Y(n609) );
  INVX1 U7409 ( .A(n609), .Y(n7744) );
  INVX1 U7410 ( .A(n7747), .Y(n7745) );
  INVX1 U7411 ( .A(n7745), .Y(n7746) );
  AND2X1 U7412 ( .A(n10325), .B(n577), .Y(n608) );
  INVX1 U7413 ( .A(n608), .Y(n7747) );
  INVX1 U7414 ( .A(n7750), .Y(n7748) );
  INVX1 U7415 ( .A(n7748), .Y(n7749) );
  AND2X1 U7416 ( .A(n10328), .B(n577), .Y(n607) );
  INVX1 U7417 ( .A(n607), .Y(n7750) );
  INVX1 U7418 ( .A(n7753), .Y(n7751) );
  INVX1 U7419 ( .A(n7751), .Y(n7752) );
  AND2X1 U7420 ( .A(n10331), .B(n577), .Y(n606) );
  INVX1 U7421 ( .A(n606), .Y(n7753) );
  INVX1 U7422 ( .A(n7756), .Y(n7754) );
  INVX1 U7423 ( .A(n7754), .Y(n7755) );
  AND2X1 U7424 ( .A(n10334), .B(n577), .Y(n605) );
  INVX1 U7425 ( .A(n605), .Y(n7756) );
  INVX1 U7426 ( .A(n7759), .Y(n7757) );
  INVX1 U7427 ( .A(n7757), .Y(n7758) );
  AND2X1 U7428 ( .A(n10337), .B(n577), .Y(n604) );
  INVX1 U7429 ( .A(n604), .Y(n7759) );
  INVX1 U7430 ( .A(n7762), .Y(n7760) );
  INVX1 U7431 ( .A(n7760), .Y(n7761) );
  AND2X1 U7432 ( .A(n10340), .B(n577), .Y(n603) );
  INVX1 U7433 ( .A(n603), .Y(n7762) );
  INVX1 U7434 ( .A(n7765), .Y(n7763) );
  INVX1 U7435 ( .A(n7763), .Y(n7764) );
  AND2X1 U7436 ( .A(n10343), .B(n577), .Y(n602) );
  INVX1 U7437 ( .A(n602), .Y(n7765) );
  INVX1 U7438 ( .A(n7768), .Y(n7766) );
  INVX1 U7439 ( .A(n7766), .Y(n7767) );
  AND2X1 U7440 ( .A(n10346), .B(n577), .Y(n601) );
  INVX1 U7441 ( .A(n601), .Y(n7768) );
  INVX1 U7442 ( .A(n7771), .Y(n7769) );
  INVX1 U7443 ( .A(n7769), .Y(n7770) );
  AND2X1 U7444 ( .A(n10349), .B(n577), .Y(n600) );
  INVX1 U7445 ( .A(n600), .Y(n7771) );
  INVX1 U7446 ( .A(n7774), .Y(n7772) );
  INVX1 U7447 ( .A(n7772), .Y(n7773) );
  AND2X1 U7448 ( .A(n10352), .B(n577), .Y(n599) );
  INVX1 U7449 ( .A(n599), .Y(n7774) );
  INVX1 U7450 ( .A(n7777), .Y(n7775) );
  INVX1 U7451 ( .A(n7775), .Y(n7776) );
  AND2X1 U7452 ( .A(n10355), .B(n577), .Y(n598) );
  INVX1 U7453 ( .A(n598), .Y(n7777) );
  INVX1 U7454 ( .A(n7780), .Y(n7778) );
  INVX1 U7455 ( .A(n7778), .Y(n7779) );
  AND2X1 U7456 ( .A(n10358), .B(n577), .Y(n597) );
  INVX1 U7457 ( .A(n597), .Y(n7780) );
  INVX1 U7458 ( .A(n7783), .Y(n7781) );
  INVX1 U7459 ( .A(n7781), .Y(n7782) );
  AND2X1 U7460 ( .A(n10361), .B(n577), .Y(n596) );
  INVX1 U7461 ( .A(n596), .Y(n7783) );
  INVX1 U7462 ( .A(n7786), .Y(n7784) );
  INVX1 U7463 ( .A(n7784), .Y(n7785) );
  AND2X1 U7464 ( .A(n10364), .B(n577), .Y(n595) );
  INVX1 U7465 ( .A(n595), .Y(n7786) );
  INVX1 U7466 ( .A(n7789), .Y(n7787) );
  INVX1 U7467 ( .A(n7787), .Y(n7788) );
  AND2X1 U7468 ( .A(n10367), .B(n577), .Y(n594) );
  INVX1 U7469 ( .A(n594), .Y(n7789) );
  INVX1 U7470 ( .A(n7792), .Y(n7790) );
  INVX1 U7471 ( .A(n7790), .Y(n7791) );
  AND2X1 U7472 ( .A(n10370), .B(n577), .Y(n593) );
  INVX1 U7473 ( .A(n593), .Y(n7792) );
  INVX1 U7474 ( .A(n7795), .Y(n7793) );
  INVX1 U7475 ( .A(n7793), .Y(n7794) );
  AND2X1 U7476 ( .A(n10373), .B(n577), .Y(n592) );
  INVX1 U7477 ( .A(n592), .Y(n7795) );
  INVX1 U7478 ( .A(n7798), .Y(n7796) );
  INVX1 U7479 ( .A(n7796), .Y(n7797) );
  AND2X1 U7480 ( .A(n10376), .B(n577), .Y(n591) );
  INVX1 U7481 ( .A(n591), .Y(n7798) );
  INVX1 U7482 ( .A(n7801), .Y(n7799) );
  INVX1 U7483 ( .A(n7799), .Y(n7800) );
  AND2X1 U7484 ( .A(n10379), .B(n577), .Y(n590) );
  INVX1 U7485 ( .A(n590), .Y(n7801) );
  INVX1 U7486 ( .A(n7804), .Y(n7802) );
  INVX1 U7487 ( .A(n7802), .Y(n7803) );
  AND2X1 U7488 ( .A(n10382), .B(n577), .Y(n589) );
  INVX1 U7489 ( .A(n589), .Y(n7804) );
  INVX1 U7490 ( .A(n7807), .Y(n7805) );
  INVX1 U7491 ( .A(n7805), .Y(n7806) );
  AND2X1 U7492 ( .A(n10385), .B(n577), .Y(n588) );
  INVX1 U7493 ( .A(n588), .Y(n7807) );
  INVX1 U7494 ( .A(n7810), .Y(n7808) );
  INVX1 U7495 ( .A(n7808), .Y(n7809) );
  AND2X1 U7496 ( .A(n10388), .B(n577), .Y(n587) );
  INVX1 U7497 ( .A(n587), .Y(n7810) );
  INVX1 U7498 ( .A(n7813), .Y(n7811) );
  INVX1 U7499 ( .A(n7811), .Y(n7812) );
  AND2X1 U7500 ( .A(n10391), .B(n577), .Y(n586) );
  INVX1 U7501 ( .A(n586), .Y(n7813) );
  INVX1 U7502 ( .A(n7816), .Y(n7814) );
  INVX1 U7503 ( .A(n7814), .Y(n7815) );
  AND2X1 U7504 ( .A(n10394), .B(n577), .Y(n585) );
  INVX1 U7505 ( .A(n585), .Y(n7816) );
  INVX1 U7506 ( .A(n7819), .Y(n7817) );
  INVX1 U7507 ( .A(n7817), .Y(n7818) );
  AND2X1 U7508 ( .A(n10397), .B(n577), .Y(n584) );
  INVX1 U7509 ( .A(n584), .Y(n7819) );
  INVX1 U7510 ( .A(n7822), .Y(n7820) );
  INVX1 U7511 ( .A(n7820), .Y(n7821) );
  AND2X1 U7512 ( .A(n10400), .B(n577), .Y(n583) );
  INVX1 U7513 ( .A(n583), .Y(n7822) );
  INVX1 U7514 ( .A(n7825), .Y(n7823) );
  INVX1 U7515 ( .A(n7823), .Y(n7824) );
  AND2X1 U7516 ( .A(n10403), .B(n577), .Y(n582) );
  INVX1 U7517 ( .A(n582), .Y(n7825) );
  INVX1 U7518 ( .A(n7828), .Y(n7826) );
  INVX1 U7519 ( .A(n7826), .Y(n7827) );
  AND2X1 U7520 ( .A(n10406), .B(n577), .Y(n581) );
  INVX1 U7521 ( .A(n581), .Y(n7828) );
  INVX1 U7522 ( .A(n7831), .Y(n7829) );
  INVX1 U7523 ( .A(n7829), .Y(n7830) );
  AND2X1 U7524 ( .A(n10409), .B(n577), .Y(n580) );
  INVX1 U7525 ( .A(n580), .Y(n7831) );
  INVX1 U7526 ( .A(n7834), .Y(n7832) );
  INVX1 U7527 ( .A(n7832), .Y(n7833) );
  AND2X1 U7528 ( .A(n10412), .B(n577), .Y(n579) );
  INVX1 U7529 ( .A(n579), .Y(n7834) );
  INVX1 U7530 ( .A(n7837), .Y(n7835) );
  INVX1 U7531 ( .A(n7835), .Y(n7836) );
  AND2X1 U7532 ( .A(n10415), .B(n577), .Y(n578) );
  INVX1 U7533 ( .A(n578), .Y(n7837) );
  INVX1 U7534 ( .A(n7840), .Y(n7838) );
  INVX1 U7535 ( .A(n7838), .Y(n7839) );
  AND2X1 U7536 ( .A(n12442), .B(n533), .Y(n575) );
  INVX1 U7537 ( .A(n575), .Y(n7840) );
  INVX1 U7538 ( .A(n7843), .Y(n7841) );
  INVX1 U7539 ( .A(n7841), .Y(n7842) );
  AND2X1 U7540 ( .A(n12445), .B(n533), .Y(n574) );
  INVX1 U7541 ( .A(n574), .Y(n7843) );
  INVX1 U7542 ( .A(n7846), .Y(n7844) );
  INVX1 U7543 ( .A(n7844), .Y(n7845) );
  AND2X1 U7544 ( .A(n12448), .B(n533), .Y(n573) );
  INVX1 U7545 ( .A(n573), .Y(n7846) );
  INVX1 U7546 ( .A(n7849), .Y(n7847) );
  INVX1 U7547 ( .A(n7847), .Y(n7848) );
  AND2X1 U7548 ( .A(n12451), .B(n533), .Y(n572) );
  INVX1 U7549 ( .A(n572), .Y(n7849) );
  INVX1 U7550 ( .A(n7852), .Y(n7850) );
  INVX1 U7551 ( .A(n7850), .Y(n7851) );
  AND2X1 U7552 ( .A(n12454), .B(n533), .Y(n571) );
  INVX1 U7553 ( .A(n571), .Y(n7852) );
  INVX1 U7554 ( .A(n7855), .Y(n7853) );
  INVX1 U7555 ( .A(n7853), .Y(n7854) );
  AND2X1 U7556 ( .A(n12457), .B(n533), .Y(n570) );
  INVX1 U7557 ( .A(n570), .Y(n7855) );
  INVX1 U7558 ( .A(n7858), .Y(n7856) );
  INVX1 U7559 ( .A(n7856), .Y(n7857) );
  AND2X1 U7560 ( .A(n12460), .B(n533), .Y(n569) );
  INVX1 U7561 ( .A(n569), .Y(n7858) );
  INVX1 U7562 ( .A(n7861), .Y(n7859) );
  INVX1 U7563 ( .A(n7859), .Y(n7860) );
  AND2X1 U7564 ( .A(n12463), .B(n533), .Y(n568) );
  INVX1 U7565 ( .A(n568), .Y(n7861) );
  INVX1 U7566 ( .A(n7864), .Y(n7862) );
  INVX1 U7567 ( .A(n7862), .Y(n7863) );
  AND2X1 U7568 ( .A(n12466), .B(n533), .Y(n567) );
  INVX1 U7569 ( .A(n567), .Y(n7864) );
  INVX1 U7570 ( .A(n7867), .Y(n7865) );
  INVX1 U7571 ( .A(n7865), .Y(n7866) );
  AND2X1 U7572 ( .A(n12469), .B(n533), .Y(n566) );
  INVX1 U7573 ( .A(n566), .Y(n7867) );
  INVX1 U7574 ( .A(n7870), .Y(n7868) );
  INVX1 U7575 ( .A(n7868), .Y(n7869) );
  AND2X1 U7576 ( .A(n12472), .B(n533), .Y(n565) );
  INVX1 U7577 ( .A(n565), .Y(n7870) );
  INVX1 U7578 ( .A(n7873), .Y(n7871) );
  INVX1 U7579 ( .A(n7871), .Y(n7872) );
  AND2X1 U7580 ( .A(n12475), .B(n533), .Y(n564) );
  INVX1 U7581 ( .A(n564), .Y(n7873) );
  INVX1 U7582 ( .A(n7876), .Y(n7874) );
  INVX1 U7583 ( .A(n7874), .Y(n7875) );
  AND2X1 U7584 ( .A(n12478), .B(n533), .Y(n563) );
  INVX1 U7585 ( .A(n563), .Y(n7876) );
  INVX1 U7586 ( .A(n7879), .Y(n7877) );
  INVX1 U7587 ( .A(n7877), .Y(n7878) );
  AND2X1 U7588 ( .A(n12481), .B(n533), .Y(n562) );
  INVX1 U7589 ( .A(n562), .Y(n7879) );
  INVX1 U7590 ( .A(n7882), .Y(n7880) );
  INVX1 U7591 ( .A(n7880), .Y(n7881) );
  AND2X1 U7592 ( .A(n12484), .B(n533), .Y(n561) );
  INVX1 U7593 ( .A(n561), .Y(n7882) );
  INVX1 U7594 ( .A(n7885), .Y(n7883) );
  INVX1 U7595 ( .A(n7883), .Y(n7884) );
  AND2X1 U7596 ( .A(n12487), .B(n533), .Y(n560) );
  INVX1 U7597 ( .A(n560), .Y(n7885) );
  INVX1 U7598 ( .A(n7888), .Y(n7886) );
  INVX1 U7599 ( .A(n7886), .Y(n7887) );
  AND2X1 U7600 ( .A(n12490), .B(n533), .Y(n559) );
  INVX1 U7601 ( .A(n559), .Y(n7888) );
  INVX1 U7602 ( .A(n7891), .Y(n7889) );
  INVX1 U7603 ( .A(n7889), .Y(n7890) );
  AND2X1 U7604 ( .A(n12493), .B(n533), .Y(n558) );
  INVX1 U7605 ( .A(n558), .Y(n7891) );
  INVX1 U7606 ( .A(n7894), .Y(n7892) );
  INVX1 U7607 ( .A(n7892), .Y(n7893) );
  AND2X1 U7608 ( .A(n12496), .B(n533), .Y(n557) );
  INVX1 U7609 ( .A(n557), .Y(n7894) );
  INVX1 U7610 ( .A(n7897), .Y(n7895) );
  INVX1 U7611 ( .A(n7895), .Y(n7896) );
  AND2X1 U7612 ( .A(n12499), .B(n533), .Y(n556) );
  INVX1 U7613 ( .A(n556), .Y(n7897) );
  INVX1 U7614 ( .A(n7900), .Y(n7898) );
  INVX1 U7615 ( .A(n7898), .Y(n7899) );
  AND2X1 U7616 ( .A(n12502), .B(n533), .Y(n555) );
  INVX1 U7617 ( .A(n555), .Y(n7900) );
  INVX1 U7618 ( .A(n7903), .Y(n7901) );
  INVX1 U7619 ( .A(n7901), .Y(n7902) );
  AND2X1 U7620 ( .A(n12505), .B(n533), .Y(n554) );
  INVX1 U7621 ( .A(n554), .Y(n7903) );
  INVX1 U7622 ( .A(n7906), .Y(n7904) );
  INVX1 U7623 ( .A(n7904), .Y(n7905) );
  AND2X1 U7624 ( .A(n12508), .B(n533), .Y(n553) );
  INVX1 U7625 ( .A(n553), .Y(n7906) );
  INVX1 U7626 ( .A(n7909), .Y(n7907) );
  INVX1 U7627 ( .A(n7907), .Y(n7908) );
  AND2X1 U7628 ( .A(n12511), .B(n533), .Y(n552) );
  INVX1 U7629 ( .A(n552), .Y(n7909) );
  INVX1 U7630 ( .A(n7912), .Y(n7910) );
  INVX1 U7631 ( .A(n7910), .Y(n7911) );
  AND2X1 U7632 ( .A(n12514), .B(n533), .Y(n551) );
  INVX1 U7633 ( .A(n551), .Y(n7912) );
  INVX1 U7634 ( .A(n7915), .Y(n7913) );
  INVX1 U7635 ( .A(n7913), .Y(n7914) );
  AND2X1 U7636 ( .A(n12517), .B(n533), .Y(n550) );
  INVX1 U7637 ( .A(n550), .Y(n7915) );
  INVX1 U7638 ( .A(n7918), .Y(n7916) );
  INVX1 U7639 ( .A(n7916), .Y(n7917) );
  AND2X1 U7640 ( .A(n12520), .B(n533), .Y(n549) );
  INVX1 U7641 ( .A(n549), .Y(n7918) );
  INVX1 U7642 ( .A(n7921), .Y(n7919) );
  INVX1 U7643 ( .A(n7919), .Y(n7920) );
  AND2X1 U7644 ( .A(n12523), .B(n533), .Y(n548) );
  INVX1 U7645 ( .A(n548), .Y(n7921) );
  INVX1 U7646 ( .A(n7924), .Y(n7922) );
  INVX1 U7647 ( .A(n7922), .Y(n7923) );
  AND2X1 U7648 ( .A(n12526), .B(n533), .Y(n547) );
  INVX1 U7649 ( .A(n547), .Y(n7924) );
  INVX1 U7650 ( .A(n7927), .Y(n7925) );
  INVX1 U7651 ( .A(n7925), .Y(n7926) );
  AND2X1 U7652 ( .A(n12529), .B(n533), .Y(n546) );
  INVX1 U7653 ( .A(n546), .Y(n7927) );
  INVX1 U7654 ( .A(n7930), .Y(n7928) );
  INVX1 U7655 ( .A(n7928), .Y(n7929) );
  AND2X1 U7656 ( .A(n12532), .B(n533), .Y(n545) );
  INVX1 U7657 ( .A(n545), .Y(n7930) );
  INVX1 U7658 ( .A(n7933), .Y(n7931) );
  INVX1 U7659 ( .A(n7931), .Y(n7932) );
  AND2X1 U7660 ( .A(n12535), .B(n533), .Y(n544) );
  INVX1 U7661 ( .A(n544), .Y(n7933) );
  INVX1 U7662 ( .A(n7936), .Y(n7934) );
  INVX1 U7663 ( .A(n7934), .Y(n7935) );
  AND2X1 U7664 ( .A(n12538), .B(n533), .Y(n543) );
  INVX1 U7665 ( .A(n543), .Y(n7936) );
  INVX1 U7666 ( .A(n7939), .Y(n7937) );
  INVX1 U7667 ( .A(n7937), .Y(n7938) );
  AND2X1 U7668 ( .A(n12541), .B(n533), .Y(n542) );
  INVX1 U7669 ( .A(n542), .Y(n7939) );
  INVX1 U7670 ( .A(n7942), .Y(n7940) );
  INVX1 U7671 ( .A(n7940), .Y(n7941) );
  AND2X1 U7672 ( .A(n12544), .B(n533), .Y(n541) );
  INVX1 U7673 ( .A(n541), .Y(n7942) );
  INVX1 U7674 ( .A(n7945), .Y(n7943) );
  INVX1 U7675 ( .A(n7943), .Y(n7944) );
  AND2X1 U7676 ( .A(n12547), .B(n533), .Y(n540) );
  INVX1 U7677 ( .A(n540), .Y(n7945) );
  INVX1 U7678 ( .A(n7948), .Y(n7946) );
  INVX1 U7679 ( .A(n7946), .Y(n7947) );
  AND2X1 U7680 ( .A(n12550), .B(n533), .Y(n539) );
  INVX1 U7681 ( .A(n539), .Y(n7948) );
  INVX1 U7682 ( .A(n7951), .Y(n7949) );
  INVX1 U7683 ( .A(n7949), .Y(n7950) );
  AND2X1 U7684 ( .A(n12553), .B(n533), .Y(n538) );
  INVX1 U7685 ( .A(n538), .Y(n7951) );
  INVX1 U7686 ( .A(n7954), .Y(n7952) );
  INVX1 U7687 ( .A(n7952), .Y(n7953) );
  AND2X1 U7688 ( .A(n12556), .B(n533), .Y(n537) );
  INVX1 U7689 ( .A(n537), .Y(n7954) );
  INVX1 U7690 ( .A(n7957), .Y(n7955) );
  INVX1 U7691 ( .A(n7955), .Y(n7956) );
  AND2X1 U7692 ( .A(n12559), .B(n533), .Y(n536) );
  INVX1 U7693 ( .A(n536), .Y(n7957) );
  INVX1 U7694 ( .A(n7960), .Y(n7958) );
  INVX1 U7695 ( .A(n7958), .Y(n7959) );
  AND2X1 U7696 ( .A(n12562), .B(n533), .Y(n535) );
  INVX1 U7697 ( .A(n535), .Y(n7960) );
  INVX1 U7698 ( .A(n7963), .Y(n7961) );
  INVX1 U7699 ( .A(n7961), .Y(n7962) );
  AND2X1 U7700 ( .A(n12565), .B(n533), .Y(n534) );
  INVX1 U7701 ( .A(n534), .Y(n7963) );
  INVX1 U7702 ( .A(n7966), .Y(n7964) );
  INVX1 U7703 ( .A(n7964), .Y(n7965) );
  AND2X1 U7704 ( .A(n10418), .B(n489), .Y(n531) );
  INVX1 U7705 ( .A(n531), .Y(n7966) );
  INVX1 U7706 ( .A(n7969), .Y(n7967) );
  INVX1 U7707 ( .A(n7967), .Y(n7968) );
  AND2X1 U7708 ( .A(n10421), .B(n489), .Y(n530) );
  INVX1 U7709 ( .A(n530), .Y(n7969) );
  INVX1 U7710 ( .A(n7972), .Y(n7970) );
  INVX1 U7711 ( .A(n7970), .Y(n7971) );
  AND2X1 U7712 ( .A(n10424), .B(n489), .Y(n529) );
  INVX1 U7713 ( .A(n529), .Y(n7972) );
  INVX1 U7714 ( .A(n7975), .Y(n7973) );
  INVX1 U7715 ( .A(n7973), .Y(n7974) );
  AND2X1 U7716 ( .A(n10427), .B(n489), .Y(n528) );
  INVX1 U7717 ( .A(n528), .Y(n7975) );
  INVX1 U7718 ( .A(n7978), .Y(n7976) );
  INVX1 U7719 ( .A(n7976), .Y(n7977) );
  AND2X1 U7720 ( .A(n10430), .B(n489), .Y(n527) );
  INVX1 U7721 ( .A(n527), .Y(n7978) );
  INVX1 U7722 ( .A(n7981), .Y(n7979) );
  INVX1 U7723 ( .A(n7979), .Y(n7980) );
  AND2X1 U7724 ( .A(n10433), .B(n489), .Y(n526) );
  INVX1 U7725 ( .A(n526), .Y(n7981) );
  INVX1 U7726 ( .A(n7984), .Y(n7982) );
  INVX1 U7727 ( .A(n7982), .Y(n7983) );
  AND2X1 U7728 ( .A(n10436), .B(n489), .Y(n525) );
  INVX1 U7729 ( .A(n525), .Y(n7984) );
  INVX1 U7730 ( .A(n7987), .Y(n7985) );
  INVX1 U7731 ( .A(n7985), .Y(n7986) );
  AND2X1 U7732 ( .A(n10439), .B(n489), .Y(n524) );
  INVX1 U7733 ( .A(n524), .Y(n7987) );
  INVX1 U7734 ( .A(n7990), .Y(n7988) );
  INVX1 U7735 ( .A(n7988), .Y(n7989) );
  AND2X1 U7736 ( .A(n10442), .B(n489), .Y(n523) );
  INVX1 U7737 ( .A(n523), .Y(n7990) );
  INVX1 U7738 ( .A(n7993), .Y(n7991) );
  INVX1 U7739 ( .A(n7991), .Y(n7992) );
  AND2X1 U7740 ( .A(n10445), .B(n489), .Y(n522) );
  INVX1 U7741 ( .A(n522), .Y(n7993) );
  INVX1 U7742 ( .A(n7996), .Y(n7994) );
  INVX1 U7743 ( .A(n7994), .Y(n7995) );
  AND2X1 U7744 ( .A(n10448), .B(n489), .Y(n521) );
  INVX1 U7745 ( .A(n521), .Y(n7996) );
  INVX1 U7746 ( .A(n7999), .Y(n7997) );
  INVX1 U7747 ( .A(n7997), .Y(n7998) );
  AND2X1 U7748 ( .A(n10451), .B(n489), .Y(n520) );
  INVX1 U7749 ( .A(n520), .Y(n7999) );
  INVX1 U7750 ( .A(n8002), .Y(n8000) );
  INVX1 U7751 ( .A(n8000), .Y(n8001) );
  AND2X1 U7752 ( .A(n10454), .B(n489), .Y(n519) );
  INVX1 U7753 ( .A(n519), .Y(n8002) );
  INVX1 U7754 ( .A(n8005), .Y(n8003) );
  INVX1 U7755 ( .A(n8003), .Y(n8004) );
  AND2X1 U7756 ( .A(n10457), .B(n489), .Y(n518) );
  INVX1 U7757 ( .A(n518), .Y(n8005) );
  INVX1 U7758 ( .A(n8008), .Y(n8006) );
  INVX1 U7759 ( .A(n8006), .Y(n8007) );
  AND2X1 U7760 ( .A(n10460), .B(n489), .Y(n517) );
  INVX1 U7761 ( .A(n517), .Y(n8008) );
  INVX1 U7762 ( .A(n8011), .Y(n8009) );
  INVX1 U7763 ( .A(n8009), .Y(n8010) );
  AND2X1 U7764 ( .A(n10463), .B(n489), .Y(n516) );
  INVX1 U7765 ( .A(n516), .Y(n8011) );
  INVX1 U7766 ( .A(n8014), .Y(n8012) );
  INVX1 U7767 ( .A(n8012), .Y(n8013) );
  AND2X1 U7768 ( .A(n10466), .B(n489), .Y(n515) );
  INVX1 U7769 ( .A(n515), .Y(n8014) );
  INVX1 U7770 ( .A(n8017), .Y(n8015) );
  INVX1 U7771 ( .A(n8015), .Y(n8016) );
  AND2X1 U7772 ( .A(n10469), .B(n489), .Y(n514) );
  INVX1 U7773 ( .A(n514), .Y(n8017) );
  INVX1 U7774 ( .A(n8020), .Y(n8018) );
  INVX1 U7775 ( .A(n8018), .Y(n8019) );
  AND2X1 U7776 ( .A(n10472), .B(n489), .Y(n513) );
  INVX1 U7777 ( .A(n513), .Y(n8020) );
  INVX1 U7778 ( .A(n8023), .Y(n8021) );
  INVX1 U7779 ( .A(n8021), .Y(n8022) );
  AND2X1 U7780 ( .A(n10475), .B(n489), .Y(n512) );
  INVX1 U7781 ( .A(n512), .Y(n8023) );
  INVX1 U7782 ( .A(n8026), .Y(n8024) );
  INVX1 U7783 ( .A(n8024), .Y(n8025) );
  AND2X1 U7784 ( .A(n10478), .B(n489), .Y(n511) );
  INVX1 U7785 ( .A(n511), .Y(n8026) );
  INVX1 U7786 ( .A(n8029), .Y(n8027) );
  INVX1 U7787 ( .A(n8027), .Y(n8028) );
  AND2X1 U7788 ( .A(n10481), .B(n489), .Y(n510) );
  INVX1 U7789 ( .A(n510), .Y(n8029) );
  INVX1 U7790 ( .A(n8032), .Y(n8030) );
  INVX1 U7791 ( .A(n8030), .Y(n8031) );
  AND2X1 U7792 ( .A(n10484), .B(n489), .Y(n509) );
  INVX1 U7793 ( .A(n509), .Y(n8032) );
  INVX1 U7794 ( .A(n8035), .Y(n8033) );
  INVX1 U7795 ( .A(n8033), .Y(n8034) );
  AND2X1 U7796 ( .A(n10487), .B(n489), .Y(n508) );
  INVX1 U7797 ( .A(n508), .Y(n8035) );
  INVX1 U7798 ( .A(n8038), .Y(n8036) );
  INVX1 U7799 ( .A(n8036), .Y(n8037) );
  AND2X1 U7800 ( .A(n10490), .B(n489), .Y(n507) );
  INVX1 U7801 ( .A(n507), .Y(n8038) );
  INVX1 U7802 ( .A(n8041), .Y(n8039) );
  INVX1 U7803 ( .A(n8039), .Y(n8040) );
  AND2X1 U7804 ( .A(n10493), .B(n489), .Y(n506) );
  INVX1 U7805 ( .A(n506), .Y(n8041) );
  INVX1 U7806 ( .A(n8044), .Y(n8042) );
  INVX1 U7807 ( .A(n8042), .Y(n8043) );
  AND2X1 U7808 ( .A(n10496), .B(n489), .Y(n505) );
  INVX1 U7809 ( .A(n505), .Y(n8044) );
  INVX1 U7810 ( .A(n8047), .Y(n8045) );
  INVX1 U7811 ( .A(n8045), .Y(n8046) );
  AND2X1 U7812 ( .A(n10499), .B(n489), .Y(n504) );
  INVX1 U7813 ( .A(n504), .Y(n8047) );
  INVX1 U7814 ( .A(n8050), .Y(n8048) );
  INVX1 U7815 ( .A(n8048), .Y(n8049) );
  AND2X1 U7816 ( .A(n10502), .B(n489), .Y(n503) );
  INVX1 U7817 ( .A(n503), .Y(n8050) );
  INVX1 U7818 ( .A(n8053), .Y(n8051) );
  INVX1 U7819 ( .A(n8051), .Y(n8052) );
  AND2X1 U7820 ( .A(n10505), .B(n489), .Y(n502) );
  INVX1 U7821 ( .A(n502), .Y(n8053) );
  INVX1 U7822 ( .A(n8056), .Y(n8054) );
  INVX1 U7823 ( .A(n8054), .Y(n8055) );
  AND2X1 U7824 ( .A(n10508), .B(n489), .Y(n501) );
  INVX1 U7825 ( .A(n501), .Y(n8056) );
  INVX1 U7826 ( .A(n8059), .Y(n8057) );
  INVX1 U7827 ( .A(n8057), .Y(n8058) );
  AND2X1 U7828 ( .A(n10511), .B(n489), .Y(n500) );
  INVX1 U7829 ( .A(n500), .Y(n8059) );
  INVX1 U7830 ( .A(n8062), .Y(n8060) );
  INVX1 U7831 ( .A(n8060), .Y(n8061) );
  AND2X1 U7832 ( .A(n10514), .B(n489), .Y(n499) );
  INVX1 U7833 ( .A(n499), .Y(n8062) );
  INVX1 U7834 ( .A(n8065), .Y(n8063) );
  INVX1 U7835 ( .A(n8063), .Y(n8064) );
  AND2X1 U7836 ( .A(n10517), .B(n489), .Y(n498) );
  INVX1 U7837 ( .A(n498), .Y(n8065) );
  INVX1 U7838 ( .A(n8068), .Y(n8066) );
  INVX1 U7839 ( .A(n8066), .Y(n8067) );
  AND2X1 U7840 ( .A(n10520), .B(n489), .Y(n497) );
  INVX1 U7841 ( .A(n497), .Y(n8068) );
  INVX1 U7842 ( .A(n8071), .Y(n8069) );
  INVX1 U7843 ( .A(n8069), .Y(n8070) );
  AND2X1 U7844 ( .A(n10523), .B(n489), .Y(n496) );
  INVX1 U7845 ( .A(n496), .Y(n8071) );
  INVX1 U7846 ( .A(n8074), .Y(n8072) );
  INVX1 U7847 ( .A(n8072), .Y(n8073) );
  AND2X1 U7848 ( .A(n10526), .B(n489), .Y(n495) );
  INVX1 U7849 ( .A(n495), .Y(n8074) );
  INVX1 U7850 ( .A(n8077), .Y(n8075) );
  INVX1 U7851 ( .A(n8075), .Y(n8076) );
  AND2X1 U7852 ( .A(n10529), .B(n489), .Y(n494) );
  INVX1 U7853 ( .A(n494), .Y(n8077) );
  INVX1 U7854 ( .A(n8080), .Y(n8078) );
  INVX1 U7855 ( .A(n8078), .Y(n8079) );
  AND2X1 U7856 ( .A(n10532), .B(n489), .Y(n493) );
  INVX1 U7857 ( .A(n493), .Y(n8080) );
  INVX1 U7858 ( .A(n8083), .Y(n8081) );
  INVX1 U7859 ( .A(n8081), .Y(n8082) );
  AND2X1 U7860 ( .A(n10535), .B(n489), .Y(n492) );
  INVX1 U7861 ( .A(n492), .Y(n8083) );
  INVX1 U7862 ( .A(n8086), .Y(n8084) );
  INVX1 U7863 ( .A(n8084), .Y(n8085) );
  AND2X1 U7864 ( .A(n10538), .B(n489), .Y(n491) );
  INVX1 U7865 ( .A(n491), .Y(n8086) );
  INVX1 U7866 ( .A(n8089), .Y(n8087) );
  INVX1 U7867 ( .A(n8087), .Y(n8088) );
  AND2X1 U7868 ( .A(n10541), .B(n489), .Y(n490) );
  INVX1 U7869 ( .A(n490), .Y(n8089) );
  INVX1 U7870 ( .A(n8092), .Y(n8090) );
  INVX1 U7871 ( .A(n8090), .Y(n8091) );
  AND2X1 U7872 ( .A(n12568), .B(n445), .Y(n487) );
  INVX1 U7873 ( .A(n487), .Y(n8092) );
  INVX1 U7874 ( .A(n8095), .Y(n8093) );
  INVX1 U7875 ( .A(n8093), .Y(n8094) );
  AND2X1 U7876 ( .A(n12571), .B(n445), .Y(n486) );
  INVX1 U7877 ( .A(n486), .Y(n8095) );
  INVX1 U7878 ( .A(n8098), .Y(n8096) );
  INVX1 U7879 ( .A(n8096), .Y(n8097) );
  AND2X1 U7880 ( .A(n12574), .B(n445), .Y(n485) );
  INVX1 U7881 ( .A(n485), .Y(n8098) );
  INVX1 U7882 ( .A(n8101), .Y(n8099) );
  INVX1 U7883 ( .A(n8099), .Y(n8100) );
  AND2X1 U7884 ( .A(n12577), .B(n445), .Y(n484) );
  INVX1 U7885 ( .A(n484), .Y(n8101) );
  INVX1 U7886 ( .A(n8104), .Y(n8102) );
  INVX1 U7887 ( .A(n8102), .Y(n8103) );
  AND2X1 U7888 ( .A(n12580), .B(n445), .Y(n483) );
  INVX1 U7889 ( .A(n483), .Y(n8104) );
  INVX1 U7890 ( .A(n8107), .Y(n8105) );
  INVX1 U7891 ( .A(n8105), .Y(n8106) );
  AND2X1 U7892 ( .A(n12583), .B(n445), .Y(n482) );
  INVX1 U7893 ( .A(n482), .Y(n8107) );
  INVX1 U7894 ( .A(n8110), .Y(n8108) );
  INVX1 U7895 ( .A(n8108), .Y(n8109) );
  AND2X1 U7896 ( .A(n12586), .B(n445), .Y(n481) );
  INVX1 U7897 ( .A(n481), .Y(n8110) );
  INVX1 U7898 ( .A(n8113), .Y(n8111) );
  INVX1 U7899 ( .A(n8111), .Y(n8112) );
  AND2X1 U7900 ( .A(n12589), .B(n445), .Y(n480) );
  INVX1 U7901 ( .A(n480), .Y(n8113) );
  INVX1 U7902 ( .A(n8116), .Y(n8114) );
  INVX1 U7903 ( .A(n8114), .Y(n8115) );
  AND2X1 U7904 ( .A(n12592), .B(n445), .Y(n479) );
  INVX1 U7905 ( .A(n479), .Y(n8116) );
  INVX1 U7906 ( .A(n8119), .Y(n8117) );
  INVX1 U7907 ( .A(n8117), .Y(n8118) );
  AND2X1 U7908 ( .A(n12595), .B(n445), .Y(n478) );
  INVX1 U7909 ( .A(n478), .Y(n8119) );
  INVX1 U7910 ( .A(n8122), .Y(n8120) );
  INVX1 U7911 ( .A(n8120), .Y(n8121) );
  AND2X1 U7912 ( .A(n12598), .B(n445), .Y(n477) );
  INVX1 U7913 ( .A(n477), .Y(n8122) );
  INVX1 U7914 ( .A(n8125), .Y(n8123) );
  INVX1 U7915 ( .A(n8123), .Y(n8124) );
  AND2X1 U7916 ( .A(n12601), .B(n445), .Y(n476) );
  INVX1 U7917 ( .A(n476), .Y(n8125) );
  INVX1 U7918 ( .A(n8128), .Y(n8126) );
  INVX1 U7919 ( .A(n8126), .Y(n8127) );
  AND2X1 U7920 ( .A(n12604), .B(n445), .Y(n475) );
  INVX1 U7921 ( .A(n475), .Y(n8128) );
  INVX1 U7922 ( .A(n8131), .Y(n8129) );
  INVX1 U7923 ( .A(n8129), .Y(n8130) );
  AND2X1 U7924 ( .A(n12607), .B(n445), .Y(n474) );
  INVX1 U7925 ( .A(n474), .Y(n8131) );
  INVX1 U7926 ( .A(n8134), .Y(n8132) );
  INVX1 U7927 ( .A(n8132), .Y(n8133) );
  AND2X1 U7928 ( .A(n12610), .B(n445), .Y(n473) );
  INVX1 U7929 ( .A(n473), .Y(n8134) );
  INVX1 U7930 ( .A(n8137), .Y(n8135) );
  INVX1 U7931 ( .A(n8135), .Y(n8136) );
  AND2X1 U7932 ( .A(n12613), .B(n445), .Y(n472) );
  INVX1 U7933 ( .A(n472), .Y(n8137) );
  INVX1 U7934 ( .A(n8140), .Y(n8138) );
  INVX1 U7935 ( .A(n8138), .Y(n8139) );
  AND2X1 U7936 ( .A(n12616), .B(n445), .Y(n471) );
  INVX1 U7937 ( .A(n471), .Y(n8140) );
  INVX1 U7938 ( .A(n8143), .Y(n8141) );
  INVX1 U7939 ( .A(n8141), .Y(n8142) );
  AND2X1 U7940 ( .A(n12619), .B(n445), .Y(n470) );
  INVX1 U7941 ( .A(n470), .Y(n8143) );
  INVX1 U7942 ( .A(n8146), .Y(n8144) );
  INVX1 U7943 ( .A(n8144), .Y(n8145) );
  AND2X1 U7944 ( .A(n12622), .B(n445), .Y(n469) );
  INVX1 U7945 ( .A(n469), .Y(n8146) );
  INVX1 U7946 ( .A(n8149), .Y(n8147) );
  INVX1 U7947 ( .A(n8147), .Y(n8148) );
  AND2X1 U7948 ( .A(n12625), .B(n445), .Y(n468) );
  INVX1 U7949 ( .A(n468), .Y(n8149) );
  INVX1 U7950 ( .A(n8152), .Y(n8150) );
  INVX1 U7951 ( .A(n8150), .Y(n8151) );
  AND2X1 U7952 ( .A(n12628), .B(n445), .Y(n467) );
  INVX1 U7953 ( .A(n467), .Y(n8152) );
  INVX1 U7954 ( .A(n8155), .Y(n8153) );
  INVX1 U7955 ( .A(n8153), .Y(n8154) );
  AND2X1 U7956 ( .A(n12631), .B(n445), .Y(n466) );
  INVX1 U7957 ( .A(n466), .Y(n8155) );
  INVX1 U7958 ( .A(n8158), .Y(n8156) );
  INVX1 U7959 ( .A(n8156), .Y(n8157) );
  AND2X1 U7960 ( .A(n12634), .B(n445), .Y(n465) );
  INVX1 U7961 ( .A(n465), .Y(n8158) );
  INVX1 U7962 ( .A(n8161), .Y(n8159) );
  INVX1 U7963 ( .A(n8159), .Y(n8160) );
  AND2X1 U7964 ( .A(n12637), .B(n445), .Y(n464) );
  INVX1 U7965 ( .A(n464), .Y(n8161) );
  INVX1 U7966 ( .A(n8164), .Y(n8162) );
  INVX1 U7967 ( .A(n8162), .Y(n8163) );
  AND2X1 U7968 ( .A(n12640), .B(n445), .Y(n463) );
  INVX1 U7969 ( .A(n463), .Y(n8164) );
  INVX1 U7970 ( .A(n8167), .Y(n8165) );
  INVX1 U7971 ( .A(n8165), .Y(n8166) );
  AND2X1 U7972 ( .A(n12643), .B(n445), .Y(n462) );
  INVX1 U7973 ( .A(n462), .Y(n8167) );
  INVX1 U7974 ( .A(n8170), .Y(n8168) );
  INVX1 U7975 ( .A(n8168), .Y(n8169) );
  AND2X1 U7976 ( .A(n12646), .B(n445), .Y(n461) );
  INVX1 U7977 ( .A(n461), .Y(n8170) );
  INVX1 U7978 ( .A(n8173), .Y(n8171) );
  INVX1 U7979 ( .A(n8171), .Y(n8172) );
  AND2X1 U7980 ( .A(n12649), .B(n445), .Y(n460) );
  INVX1 U7981 ( .A(n460), .Y(n8173) );
  INVX1 U7982 ( .A(n8176), .Y(n8174) );
  INVX1 U7983 ( .A(n8174), .Y(n8175) );
  AND2X1 U7984 ( .A(n12652), .B(n445), .Y(n459) );
  INVX1 U7985 ( .A(n459), .Y(n8176) );
  INVX1 U7986 ( .A(n8179), .Y(n8177) );
  INVX1 U7987 ( .A(n8177), .Y(n8178) );
  AND2X1 U7988 ( .A(n12655), .B(n445), .Y(n458) );
  INVX1 U7989 ( .A(n458), .Y(n8179) );
  INVX1 U7990 ( .A(n8182), .Y(n8180) );
  INVX1 U7991 ( .A(n8180), .Y(n8181) );
  AND2X1 U7992 ( .A(n12658), .B(n445), .Y(n457) );
  INVX1 U7993 ( .A(n457), .Y(n8182) );
  INVX1 U7994 ( .A(n8185), .Y(n8183) );
  INVX1 U7995 ( .A(n8183), .Y(n8184) );
  AND2X1 U7996 ( .A(n12661), .B(n445), .Y(n456) );
  INVX1 U7997 ( .A(n456), .Y(n8185) );
  INVX1 U7998 ( .A(n8188), .Y(n8186) );
  INVX1 U7999 ( .A(n8186), .Y(n8187) );
  AND2X1 U8000 ( .A(n12664), .B(n445), .Y(n455) );
  INVX1 U8001 ( .A(n455), .Y(n8188) );
  INVX1 U8002 ( .A(n8191), .Y(n8189) );
  INVX1 U8003 ( .A(n8189), .Y(n8190) );
  AND2X1 U8004 ( .A(n12667), .B(n445), .Y(n454) );
  INVX1 U8005 ( .A(n454), .Y(n8191) );
  INVX1 U8006 ( .A(n8194), .Y(n8192) );
  INVX1 U8007 ( .A(n8192), .Y(n8193) );
  AND2X1 U8008 ( .A(n12670), .B(n445), .Y(n453) );
  INVX1 U8009 ( .A(n453), .Y(n8194) );
  INVX1 U8010 ( .A(n8197), .Y(n8195) );
  INVX1 U8011 ( .A(n8195), .Y(n8196) );
  AND2X1 U8012 ( .A(n12673), .B(n445), .Y(n452) );
  INVX1 U8013 ( .A(n452), .Y(n8197) );
  INVX1 U8014 ( .A(n8200), .Y(n8198) );
  INVX1 U8015 ( .A(n8198), .Y(n8199) );
  AND2X1 U8016 ( .A(n12676), .B(n445), .Y(n451) );
  INVX1 U8017 ( .A(n451), .Y(n8200) );
  INVX1 U8018 ( .A(n8203), .Y(n8201) );
  INVX1 U8019 ( .A(n8201), .Y(n8202) );
  AND2X1 U8020 ( .A(n12679), .B(n445), .Y(n450) );
  INVX1 U8021 ( .A(n450), .Y(n8203) );
  INVX1 U8022 ( .A(n8206), .Y(n8204) );
  INVX1 U8023 ( .A(n8204), .Y(n8205) );
  AND2X1 U8024 ( .A(n12682), .B(n445), .Y(n449) );
  INVX1 U8025 ( .A(n449), .Y(n8206) );
  INVX1 U8026 ( .A(n8209), .Y(n8207) );
  INVX1 U8027 ( .A(n8207), .Y(n8208) );
  AND2X1 U8028 ( .A(n12685), .B(n445), .Y(n448) );
  INVX1 U8029 ( .A(n448), .Y(n8209) );
  INVX1 U8030 ( .A(n8212), .Y(n8210) );
  INVX1 U8031 ( .A(n8210), .Y(n8211) );
  AND2X1 U8032 ( .A(n12688), .B(n445), .Y(n447) );
  INVX1 U8033 ( .A(n447), .Y(n8212) );
  INVX1 U8034 ( .A(n8215), .Y(n8213) );
  INVX1 U8035 ( .A(n8213), .Y(n8214) );
  AND2X1 U8036 ( .A(n12691), .B(n445), .Y(n446) );
  INVX1 U8037 ( .A(n446), .Y(n8215) );
  INVX1 U8038 ( .A(n8218), .Y(n8216) );
  INVX1 U8039 ( .A(n8216), .Y(n8217) );
  AND2X1 U8040 ( .A(n10544), .B(n13042), .Y(n443) );
  INVX1 U8041 ( .A(n443), .Y(n8218) );
  INVX1 U8042 ( .A(n8221), .Y(n8219) );
  INVX1 U8043 ( .A(n8219), .Y(n8220) );
  AND2X1 U8044 ( .A(n10547), .B(n13043), .Y(n442) );
  INVX1 U8045 ( .A(n442), .Y(n8221) );
  INVX1 U8046 ( .A(n8224), .Y(n8222) );
  INVX1 U8047 ( .A(n8222), .Y(n8223) );
  AND2X1 U8048 ( .A(n10550), .B(n12971), .Y(n441) );
  INVX1 U8049 ( .A(n441), .Y(n8224) );
  INVX1 U8050 ( .A(n8227), .Y(n8225) );
  INVX1 U8051 ( .A(n8225), .Y(n8226) );
  AND2X1 U8052 ( .A(n10553), .B(n13042), .Y(n440) );
  INVX1 U8053 ( .A(n440), .Y(n8227) );
  INVX1 U8054 ( .A(n8230), .Y(n8228) );
  INVX1 U8055 ( .A(n8228), .Y(n8229) );
  AND2X1 U8056 ( .A(n10556), .B(n8628), .Y(n439) );
  INVX1 U8057 ( .A(n439), .Y(n8230) );
  INVX1 U8058 ( .A(n8233), .Y(n8231) );
  INVX1 U8059 ( .A(n8231), .Y(n8232) );
  AND2X1 U8060 ( .A(n10559), .B(n12960), .Y(n438) );
  INVX1 U8061 ( .A(n438), .Y(n8233) );
  INVX1 U8062 ( .A(n8236), .Y(n8234) );
  INVX1 U8063 ( .A(n8234), .Y(n8235) );
  AND2X1 U8064 ( .A(n10562), .B(n13042), .Y(n437) );
  INVX1 U8065 ( .A(n437), .Y(n8236) );
  INVX1 U8066 ( .A(n8239), .Y(n8237) );
  INVX1 U8067 ( .A(n8237), .Y(n8238) );
  AND2X1 U8068 ( .A(n10565), .B(n8664), .Y(n436) );
  INVX1 U8069 ( .A(n436), .Y(n8239) );
  INVX1 U8070 ( .A(n8242), .Y(n8240) );
  INVX1 U8071 ( .A(n8240), .Y(n8241) );
  AND2X1 U8072 ( .A(n10568), .B(n8648), .Y(n435) );
  INVX1 U8073 ( .A(n435), .Y(n8242) );
  INVX1 U8074 ( .A(n8245), .Y(n8243) );
  INVX1 U8075 ( .A(n8243), .Y(n8244) );
  AND2X1 U8076 ( .A(n10571), .B(n13042), .Y(n434) );
  INVX1 U8077 ( .A(n434), .Y(n8245) );
  INVX1 U8078 ( .A(n8248), .Y(n8246) );
  INVX1 U8079 ( .A(n8246), .Y(n8247) );
  AND2X1 U8080 ( .A(n10574), .B(n8646), .Y(n433) );
  INVX1 U8081 ( .A(n433), .Y(n8248) );
  INVX1 U8082 ( .A(n8251), .Y(n8249) );
  INVX1 U8083 ( .A(n8249), .Y(n8250) );
  AND2X1 U8084 ( .A(n10577), .B(n8764), .Y(n432) );
  INVX1 U8085 ( .A(n432), .Y(n8251) );
  INVX1 U8086 ( .A(n8254), .Y(n8252) );
  INVX1 U8087 ( .A(n8252), .Y(n8253) );
  AND2X1 U8088 ( .A(n10580), .B(n13042), .Y(n431) );
  INVX1 U8089 ( .A(n431), .Y(n8254) );
  INVX1 U8090 ( .A(n8257), .Y(n8255) );
  INVX1 U8091 ( .A(n8255), .Y(n8256) );
  AND2X1 U8092 ( .A(n10583), .B(n13024), .Y(n430) );
  INVX1 U8093 ( .A(n430), .Y(n8257) );
  INVX1 U8094 ( .A(n8260), .Y(n8258) );
  INVX1 U8095 ( .A(n8258), .Y(n8259) );
  AND2X1 U8096 ( .A(n10586), .B(n13024), .Y(n429) );
  INVX1 U8097 ( .A(n429), .Y(n8260) );
  INVX1 U8098 ( .A(n8263), .Y(n8261) );
  INVX1 U8099 ( .A(n8261), .Y(n8262) );
  AND2X1 U8100 ( .A(n10589), .B(n13042), .Y(n428) );
  INVX1 U8101 ( .A(n428), .Y(n8263) );
  INVX1 U8102 ( .A(n8266), .Y(n8264) );
  INVX1 U8103 ( .A(n8264), .Y(n8265) );
  AND2X1 U8104 ( .A(n10592), .B(n13043), .Y(n427) );
  INVX1 U8105 ( .A(n427), .Y(n8266) );
  INVX1 U8106 ( .A(n8269), .Y(n8267) );
  INVX1 U8107 ( .A(n8267), .Y(n8268) );
  AND2X1 U8108 ( .A(n10595), .B(n12971), .Y(n426) );
  INVX1 U8109 ( .A(n426), .Y(n8269) );
  INVX1 U8110 ( .A(n8272), .Y(n8270) );
  INVX1 U8111 ( .A(n8270), .Y(n8271) );
  AND2X1 U8112 ( .A(n10598), .B(n13042), .Y(n425) );
  INVX1 U8113 ( .A(n425), .Y(n8272) );
  INVX1 U8114 ( .A(n8275), .Y(n8273) );
  INVX1 U8115 ( .A(n8273), .Y(n8274) );
  AND2X1 U8116 ( .A(n10601), .B(n12960), .Y(n424) );
  INVX1 U8117 ( .A(n424), .Y(n8275) );
  INVX1 U8118 ( .A(n8278), .Y(n8276) );
  INVX1 U8119 ( .A(n8276), .Y(n8277) );
  AND2X1 U8120 ( .A(n10604), .B(n10798), .Y(n423) );
  INVX1 U8121 ( .A(n423), .Y(n8278) );
  INVX1 U8122 ( .A(n8281), .Y(n8279) );
  INVX1 U8123 ( .A(n8279), .Y(n8280) );
  AND2X1 U8124 ( .A(n10607), .B(n13042), .Y(n422) );
  INVX1 U8125 ( .A(n422), .Y(n8281) );
  INVX1 U8126 ( .A(n8284), .Y(n8282) );
  INVX1 U8127 ( .A(n8282), .Y(n8283) );
  AND2X1 U8128 ( .A(n10610), .B(n8644), .Y(n421) );
  INVX1 U8129 ( .A(n421), .Y(n8284) );
  INVX1 U8130 ( .A(n8287), .Y(n8285) );
  INVX1 U8131 ( .A(n8285), .Y(n8286) );
  AND2X1 U8132 ( .A(n10613), .B(n13024), .Y(n420) );
  INVX1 U8133 ( .A(n420), .Y(n8287) );
  INVX1 U8134 ( .A(n8290), .Y(n8288) );
  INVX1 U8135 ( .A(n8288), .Y(n8289) );
  AND2X1 U8136 ( .A(n10616), .B(n13042), .Y(n419) );
  INVX1 U8137 ( .A(n419), .Y(n8290) );
  INVX1 U8138 ( .A(n8293), .Y(n8291) );
  INVX1 U8139 ( .A(n8291), .Y(n8292) );
  AND2X1 U8140 ( .A(n10619), .B(n8660), .Y(n418) );
  INVX1 U8141 ( .A(n418), .Y(n8293) );
  INVX1 U8142 ( .A(n8296), .Y(n8294) );
  INVX1 U8143 ( .A(n8294), .Y(n8295) );
  AND2X1 U8144 ( .A(n10622), .B(n12988), .Y(n417) );
  INVX1 U8145 ( .A(n417), .Y(n8296) );
  INVX1 U8146 ( .A(n8299), .Y(n8297) );
  INVX1 U8147 ( .A(n8297), .Y(n8298) );
  AND2X1 U8148 ( .A(n10625), .B(n13042), .Y(n416) );
  INVX1 U8149 ( .A(n416), .Y(n8299) );
  INVX1 U8150 ( .A(n8302), .Y(n8300) );
  INVX1 U8151 ( .A(n8300), .Y(n8301) );
  AND2X1 U8152 ( .A(n10628), .B(n8638), .Y(n415) );
  INVX1 U8153 ( .A(n415), .Y(n8302) );
  INVX1 U8154 ( .A(n8305), .Y(n8303) );
  INVX1 U8155 ( .A(n8303), .Y(n8304) );
  AND2X1 U8156 ( .A(n10631), .B(n12988), .Y(n414) );
  INVX1 U8157 ( .A(n414), .Y(n8305) );
  INVX1 U8158 ( .A(n8308), .Y(n8306) );
  INVX1 U8159 ( .A(n8306), .Y(n8307) );
  AND2X1 U8160 ( .A(n10634), .B(n13042), .Y(n413) );
  INVX1 U8161 ( .A(n413), .Y(n8308) );
  INVX1 U8162 ( .A(n8311), .Y(n8309) );
  INVX1 U8163 ( .A(n8309), .Y(n8310) );
  AND2X1 U8164 ( .A(n10637), .B(n8650), .Y(n412) );
  INVX1 U8165 ( .A(n412), .Y(n8311) );
  INVX1 U8166 ( .A(n8314), .Y(n8312) );
  INVX1 U8167 ( .A(n8312), .Y(n8313) );
  AND2X1 U8168 ( .A(n10640), .B(n13024), .Y(n411) );
  INVX1 U8169 ( .A(n411), .Y(n8314) );
  INVX1 U8170 ( .A(n8317), .Y(n8315) );
  INVX1 U8171 ( .A(n8315), .Y(n8316) );
  AND2X1 U8172 ( .A(n10643), .B(n13042), .Y(n410) );
  INVX1 U8173 ( .A(n410), .Y(n8317) );
  INVX1 U8174 ( .A(n8320), .Y(n8318) );
  INVX1 U8175 ( .A(n8318), .Y(n8319) );
  AND2X1 U8176 ( .A(n10646), .B(n12971), .Y(n409) );
  INVX1 U8177 ( .A(n409), .Y(n8320) );
  INVX1 U8178 ( .A(n8323), .Y(n8321) );
  INVX1 U8179 ( .A(n8321), .Y(n8322) );
  AND2X1 U8180 ( .A(n10649), .B(n12971), .Y(n408) );
  INVX1 U8181 ( .A(n408), .Y(n8323) );
  INVX1 U8182 ( .A(n8326), .Y(n8324) );
  INVX1 U8183 ( .A(n8324), .Y(n8325) );
  AND2X1 U8184 ( .A(n10652), .B(n13042), .Y(n407) );
  INVX1 U8185 ( .A(n407), .Y(n8326) );
  INVX1 U8186 ( .A(n8329), .Y(n8327) );
  INVX1 U8187 ( .A(n8327), .Y(n8328) );
  AND2X1 U8188 ( .A(n10655), .B(n13024), .Y(n406) );
  INVX1 U8189 ( .A(n406), .Y(n8329) );
  INVX1 U8190 ( .A(n8332), .Y(n8330) );
  INVX1 U8191 ( .A(n8330), .Y(n8331) );
  AND2X1 U8192 ( .A(n10658), .B(n8764), .Y(n405) );
  INVX1 U8193 ( .A(n405), .Y(n8332) );
  INVX1 U8194 ( .A(n8335), .Y(n8333) );
  INVX1 U8195 ( .A(n8333), .Y(n8334) );
  AND2X1 U8196 ( .A(n10661), .B(n13042), .Y(n404) );
  INVX1 U8197 ( .A(n404), .Y(n8335) );
  INVX1 U8198 ( .A(n8338), .Y(n8336) );
  INVX1 U8199 ( .A(n8336), .Y(n8337) );
  AND2X1 U8200 ( .A(n10664), .B(n13043), .Y(n403) );
  INVX1 U8201 ( .A(n403), .Y(n8338) );
  INVX1 U8202 ( .A(n8341), .Y(n8339) );
  INVX1 U8203 ( .A(n8339), .Y(n8340) );
  AND2X1 U8204 ( .A(n10667), .B(n13024), .Y(n402) );
  INVX1 U8205 ( .A(n402), .Y(n8341) );
  INVX1 U8206 ( .A(n8344), .Y(n8342) );
  INVX1 U8207 ( .A(n8342), .Y(n8343) );
  AND2X1 U8208 ( .A(n12694), .B(n357), .Y(n399) );
  INVX1 U8209 ( .A(n399), .Y(n8344) );
  INVX1 U8210 ( .A(n8347), .Y(n8345) );
  INVX1 U8211 ( .A(n8345), .Y(n8346) );
  AND2X1 U8212 ( .A(n12697), .B(n357), .Y(n398) );
  INVX1 U8213 ( .A(n398), .Y(n8347) );
  INVX1 U8214 ( .A(n8350), .Y(n8348) );
  INVX1 U8215 ( .A(n8348), .Y(n8349) );
  AND2X1 U8216 ( .A(n12700), .B(n357), .Y(n397) );
  INVX1 U8217 ( .A(n397), .Y(n8350) );
  INVX1 U8218 ( .A(n8353), .Y(n8351) );
  INVX1 U8219 ( .A(n8351), .Y(n8352) );
  AND2X1 U8220 ( .A(n12703), .B(n357), .Y(n396) );
  INVX1 U8221 ( .A(n396), .Y(n8353) );
  INVX1 U8222 ( .A(n8356), .Y(n8354) );
  INVX1 U8223 ( .A(n8354), .Y(n8355) );
  AND2X1 U8224 ( .A(n12706), .B(n357), .Y(n395) );
  INVX1 U8225 ( .A(n395), .Y(n8356) );
  INVX1 U8226 ( .A(n8359), .Y(n8357) );
  INVX1 U8227 ( .A(n8357), .Y(n8358) );
  AND2X1 U8228 ( .A(n12709), .B(n357), .Y(n394) );
  INVX1 U8229 ( .A(n394), .Y(n8359) );
  INVX1 U8230 ( .A(n8362), .Y(n8360) );
  INVX1 U8231 ( .A(n8360), .Y(n8361) );
  AND2X1 U8232 ( .A(n12712), .B(n357), .Y(n393) );
  INVX1 U8233 ( .A(n393), .Y(n8362) );
  INVX1 U8234 ( .A(n8365), .Y(n8363) );
  INVX1 U8235 ( .A(n8363), .Y(n8364) );
  AND2X1 U8236 ( .A(n12715), .B(n357), .Y(n392) );
  INVX1 U8237 ( .A(n392), .Y(n8365) );
  INVX1 U8238 ( .A(n8368), .Y(n8366) );
  INVX1 U8239 ( .A(n8366), .Y(n8367) );
  AND2X1 U8240 ( .A(n12718), .B(n357), .Y(n391) );
  INVX1 U8241 ( .A(n391), .Y(n8368) );
  INVX1 U8242 ( .A(n8371), .Y(n8369) );
  INVX1 U8243 ( .A(n8369), .Y(n8370) );
  AND2X1 U8244 ( .A(n12721), .B(n357), .Y(n390) );
  INVX1 U8245 ( .A(n390), .Y(n8371) );
  INVX1 U8246 ( .A(n8374), .Y(n8372) );
  INVX1 U8247 ( .A(n8372), .Y(n8373) );
  AND2X1 U8248 ( .A(n12724), .B(n357), .Y(n389) );
  INVX1 U8249 ( .A(n389), .Y(n8374) );
  INVX1 U8250 ( .A(n8377), .Y(n8375) );
  INVX1 U8251 ( .A(n8375), .Y(n8376) );
  AND2X1 U8252 ( .A(n12727), .B(n357), .Y(n388) );
  INVX1 U8253 ( .A(n388), .Y(n8377) );
  INVX1 U8254 ( .A(n8380), .Y(n8378) );
  INVX1 U8255 ( .A(n8378), .Y(n8379) );
  AND2X1 U8256 ( .A(n12730), .B(n357), .Y(n387) );
  INVX1 U8257 ( .A(n387), .Y(n8380) );
  INVX1 U8258 ( .A(n8383), .Y(n8381) );
  INVX1 U8259 ( .A(n8381), .Y(n8382) );
  AND2X1 U8260 ( .A(n12733), .B(n357), .Y(n386) );
  INVX1 U8261 ( .A(n386), .Y(n8383) );
  INVX1 U8262 ( .A(n8386), .Y(n8384) );
  INVX1 U8263 ( .A(n8384), .Y(n8385) );
  AND2X1 U8264 ( .A(n12736), .B(n357), .Y(n385) );
  INVX1 U8265 ( .A(n385), .Y(n8386) );
  INVX1 U8266 ( .A(n8389), .Y(n8387) );
  INVX1 U8267 ( .A(n8387), .Y(n8388) );
  AND2X1 U8268 ( .A(n12739), .B(n357), .Y(n384) );
  INVX1 U8269 ( .A(n384), .Y(n8389) );
  INVX1 U8270 ( .A(n8392), .Y(n8390) );
  INVX1 U8271 ( .A(n8390), .Y(n8391) );
  AND2X1 U8272 ( .A(n12742), .B(n357), .Y(n383) );
  INVX1 U8273 ( .A(n383), .Y(n8392) );
  INVX1 U8274 ( .A(n8395), .Y(n8393) );
  INVX1 U8275 ( .A(n8393), .Y(n8394) );
  AND2X1 U8276 ( .A(n12745), .B(n357), .Y(n382) );
  INVX1 U8277 ( .A(n382), .Y(n8395) );
  INVX1 U8278 ( .A(n8398), .Y(n8396) );
  INVX1 U8279 ( .A(n8396), .Y(n8397) );
  AND2X1 U8280 ( .A(n12748), .B(n357), .Y(n381) );
  INVX1 U8281 ( .A(n381), .Y(n8398) );
  INVX1 U8282 ( .A(n8401), .Y(n8399) );
  INVX1 U8283 ( .A(n8399), .Y(n8400) );
  AND2X1 U8284 ( .A(n12751), .B(n357), .Y(n380) );
  INVX1 U8285 ( .A(n380), .Y(n8401) );
  INVX1 U8286 ( .A(n8404), .Y(n8402) );
  INVX1 U8287 ( .A(n8402), .Y(n8403) );
  AND2X1 U8288 ( .A(n12754), .B(n357), .Y(n379) );
  INVX1 U8289 ( .A(n379), .Y(n8404) );
  INVX1 U8290 ( .A(n8407), .Y(n8405) );
  INVX1 U8291 ( .A(n8405), .Y(n8406) );
  AND2X1 U8292 ( .A(n12757), .B(n357), .Y(n378) );
  INVX1 U8293 ( .A(n378), .Y(n8407) );
  INVX1 U8294 ( .A(n8410), .Y(n8408) );
  INVX1 U8295 ( .A(n8408), .Y(n8409) );
  AND2X1 U8296 ( .A(n12760), .B(n357), .Y(n377) );
  INVX1 U8297 ( .A(n377), .Y(n8410) );
  INVX1 U8298 ( .A(n8413), .Y(n8411) );
  INVX1 U8299 ( .A(n8411), .Y(n8412) );
  AND2X1 U8300 ( .A(n12763), .B(n357), .Y(n376) );
  INVX1 U8301 ( .A(n376), .Y(n8413) );
  INVX1 U8302 ( .A(n8416), .Y(n8414) );
  INVX1 U8303 ( .A(n8414), .Y(n8415) );
  AND2X1 U8304 ( .A(n12766), .B(n357), .Y(n375) );
  INVX1 U8305 ( .A(n375), .Y(n8416) );
  INVX1 U8306 ( .A(n8419), .Y(n8417) );
  INVX1 U8307 ( .A(n8417), .Y(n8418) );
  AND2X1 U8308 ( .A(n12769), .B(n357), .Y(n374) );
  INVX1 U8309 ( .A(n374), .Y(n8419) );
  INVX1 U8310 ( .A(n8422), .Y(n8420) );
  INVX1 U8311 ( .A(n8420), .Y(n8421) );
  AND2X1 U8312 ( .A(n12772), .B(n357), .Y(n373) );
  INVX1 U8313 ( .A(n373), .Y(n8422) );
  INVX1 U8314 ( .A(n8425), .Y(n8423) );
  INVX1 U8315 ( .A(n8423), .Y(n8424) );
  AND2X1 U8316 ( .A(n12775), .B(n357), .Y(n372) );
  INVX1 U8317 ( .A(n372), .Y(n8425) );
  INVX1 U8318 ( .A(n8428), .Y(n8426) );
  INVX1 U8319 ( .A(n8426), .Y(n8427) );
  AND2X1 U8320 ( .A(n12778), .B(n357), .Y(n371) );
  INVX1 U8321 ( .A(n371), .Y(n8428) );
  INVX1 U8322 ( .A(n8431), .Y(n8429) );
  INVX1 U8323 ( .A(n8429), .Y(n8430) );
  AND2X1 U8324 ( .A(n12781), .B(n357), .Y(n370) );
  INVX1 U8325 ( .A(n370), .Y(n8431) );
  INVX1 U8326 ( .A(n8434), .Y(n8432) );
  INVX1 U8327 ( .A(n8432), .Y(n8433) );
  AND2X1 U8328 ( .A(n12784), .B(n357), .Y(n369) );
  INVX1 U8329 ( .A(n369), .Y(n8434) );
  INVX1 U8330 ( .A(n8437), .Y(n8435) );
  INVX1 U8331 ( .A(n8435), .Y(n8436) );
  AND2X1 U8332 ( .A(n12787), .B(n357), .Y(n368) );
  INVX1 U8333 ( .A(n368), .Y(n8437) );
  INVX1 U8334 ( .A(n8440), .Y(n8438) );
  INVX1 U8335 ( .A(n8438), .Y(n8439) );
  AND2X1 U8336 ( .A(n12790), .B(n357), .Y(n367) );
  INVX1 U8337 ( .A(n367), .Y(n8440) );
  INVX1 U8338 ( .A(n8443), .Y(n8441) );
  INVX1 U8339 ( .A(n8441), .Y(n8442) );
  AND2X1 U8340 ( .A(n12793), .B(n357), .Y(n366) );
  INVX1 U8341 ( .A(n366), .Y(n8443) );
  INVX1 U8342 ( .A(n8446), .Y(n8444) );
  INVX1 U8343 ( .A(n8444), .Y(n8445) );
  AND2X1 U8344 ( .A(n12796), .B(n357), .Y(n365) );
  INVX1 U8345 ( .A(n365), .Y(n8446) );
  INVX1 U8346 ( .A(n8449), .Y(n8447) );
  INVX1 U8347 ( .A(n8447), .Y(n8448) );
  AND2X1 U8348 ( .A(n12799), .B(n357), .Y(n364) );
  INVX1 U8349 ( .A(n364), .Y(n8449) );
  INVX1 U8350 ( .A(n8452), .Y(n8450) );
  INVX1 U8351 ( .A(n8450), .Y(n8451) );
  AND2X1 U8352 ( .A(n12802), .B(n357), .Y(n363) );
  INVX1 U8353 ( .A(n363), .Y(n8452) );
  INVX1 U8354 ( .A(n8455), .Y(n8453) );
  INVX1 U8355 ( .A(n8453), .Y(n8454) );
  AND2X1 U8356 ( .A(n12805), .B(n357), .Y(n362) );
  INVX1 U8357 ( .A(n362), .Y(n8455) );
  INVX1 U8358 ( .A(n8458), .Y(n8456) );
  INVX1 U8359 ( .A(n8456), .Y(n8457) );
  AND2X1 U8360 ( .A(n12808), .B(n357), .Y(n361) );
  INVX1 U8361 ( .A(n361), .Y(n8458) );
  INVX1 U8362 ( .A(n8461), .Y(n8459) );
  INVX1 U8363 ( .A(n8459), .Y(n8460) );
  AND2X1 U8364 ( .A(n12811), .B(n357), .Y(n360) );
  INVX1 U8365 ( .A(n360), .Y(n8461) );
  INVX1 U8366 ( .A(n8464), .Y(n8462) );
  INVX1 U8367 ( .A(n8462), .Y(n8463) );
  AND2X1 U8368 ( .A(n12814), .B(n357), .Y(n359) );
  INVX1 U8369 ( .A(n359), .Y(n8464) );
  INVX1 U8370 ( .A(n8467), .Y(n8465) );
  INVX1 U8371 ( .A(n8465), .Y(n8466) );
  AND2X1 U8372 ( .A(n12817), .B(n357), .Y(n358) );
  INVX1 U8373 ( .A(n358), .Y(n8467) );
  INVX1 U8374 ( .A(n8470), .Y(n8468) );
  INVX1 U8375 ( .A(n8468), .Y(n8469) );
  AND2X1 U8376 ( .A(n10670), .B(n270), .Y(n354) );
  INVX1 U8377 ( .A(n354), .Y(n8470) );
  INVX1 U8378 ( .A(n8473), .Y(n8471) );
  INVX1 U8379 ( .A(n8471), .Y(n8472) );
  AND2X1 U8380 ( .A(n10673), .B(n270), .Y(n352) );
  INVX1 U8381 ( .A(n352), .Y(n8473) );
  INVX1 U8382 ( .A(n8476), .Y(n8474) );
  INVX1 U8383 ( .A(n8474), .Y(n8475) );
  AND2X1 U8384 ( .A(n10676), .B(n270), .Y(n350) );
  INVX1 U8385 ( .A(n350), .Y(n8476) );
  INVX1 U8386 ( .A(n8479), .Y(n8477) );
  INVX1 U8387 ( .A(n8477), .Y(n8478) );
  AND2X1 U8388 ( .A(n10679), .B(n270), .Y(n348) );
  INVX1 U8389 ( .A(n348), .Y(n8479) );
  INVX1 U8390 ( .A(n8482), .Y(n8480) );
  INVX1 U8391 ( .A(n8480), .Y(n8481) );
  AND2X1 U8392 ( .A(n10682), .B(n270), .Y(n346) );
  INVX1 U8393 ( .A(n346), .Y(n8482) );
  INVX1 U8394 ( .A(n8485), .Y(n8483) );
  INVX1 U8395 ( .A(n8483), .Y(n8484) );
  AND2X1 U8396 ( .A(n10685), .B(n270), .Y(n344) );
  INVX1 U8397 ( .A(n344), .Y(n8485) );
  INVX1 U8398 ( .A(n8488), .Y(n8486) );
  INVX1 U8399 ( .A(n8486), .Y(n8487) );
  AND2X1 U8400 ( .A(n10688), .B(n270), .Y(n342) );
  INVX1 U8401 ( .A(n342), .Y(n8488) );
  INVX1 U8402 ( .A(n8491), .Y(n8489) );
  INVX1 U8403 ( .A(n8489), .Y(n8490) );
  AND2X1 U8404 ( .A(n10691), .B(n270), .Y(n340) );
  INVX1 U8405 ( .A(n340), .Y(n8491) );
  INVX1 U8406 ( .A(n8494), .Y(n8492) );
  INVX1 U8407 ( .A(n8492), .Y(n8493) );
  AND2X1 U8408 ( .A(n10694), .B(n270), .Y(n338) );
  INVX1 U8409 ( .A(n338), .Y(n8494) );
  INVX1 U8410 ( .A(n8497), .Y(n8495) );
  INVX1 U8411 ( .A(n8495), .Y(n8496) );
  AND2X1 U8412 ( .A(n10697), .B(n270), .Y(n336) );
  INVX1 U8413 ( .A(n336), .Y(n8497) );
  INVX1 U8414 ( .A(n8500), .Y(n8498) );
  INVX1 U8415 ( .A(n8498), .Y(n8499) );
  AND2X1 U8416 ( .A(n10700), .B(n270), .Y(n334) );
  INVX1 U8417 ( .A(n334), .Y(n8500) );
  INVX1 U8418 ( .A(n8503), .Y(n8501) );
  INVX1 U8419 ( .A(n8501), .Y(n8502) );
  AND2X1 U8420 ( .A(n10703), .B(n270), .Y(n332) );
  INVX1 U8421 ( .A(n332), .Y(n8503) );
  INVX1 U8422 ( .A(n8506), .Y(n8504) );
  INVX1 U8423 ( .A(n8504), .Y(n8505) );
  AND2X1 U8424 ( .A(n10706), .B(n270), .Y(n330) );
  INVX1 U8425 ( .A(n330), .Y(n8506) );
  INVX1 U8426 ( .A(n8509), .Y(n8507) );
  INVX1 U8427 ( .A(n8507), .Y(n8508) );
  AND2X1 U8428 ( .A(n10709), .B(n270), .Y(n328) );
  INVX1 U8429 ( .A(n328), .Y(n8509) );
  INVX1 U8430 ( .A(n8512), .Y(n8510) );
  INVX1 U8431 ( .A(n8510), .Y(n8511) );
  AND2X1 U8432 ( .A(n10712), .B(n270), .Y(n326) );
  INVX1 U8433 ( .A(n326), .Y(n8512) );
  INVX1 U8434 ( .A(n8515), .Y(n8513) );
  INVX1 U8435 ( .A(n8513), .Y(n8514) );
  AND2X1 U8436 ( .A(n10715), .B(n270), .Y(n324) );
  INVX1 U8437 ( .A(n324), .Y(n8515) );
  INVX1 U8438 ( .A(n8518), .Y(n8516) );
  INVX1 U8439 ( .A(n8516), .Y(n8517) );
  AND2X1 U8440 ( .A(n10718), .B(n270), .Y(n322) );
  INVX1 U8441 ( .A(n322), .Y(n8518) );
  INVX1 U8442 ( .A(n8521), .Y(n8519) );
  INVX1 U8443 ( .A(n8519), .Y(n8520) );
  AND2X1 U8444 ( .A(n10721), .B(n270), .Y(n320) );
  INVX1 U8445 ( .A(n320), .Y(n8521) );
  INVX1 U8446 ( .A(n8524), .Y(n8522) );
  INVX1 U8447 ( .A(n8522), .Y(n8523) );
  AND2X1 U8448 ( .A(n10724), .B(n270), .Y(n318) );
  INVX1 U8449 ( .A(n318), .Y(n8524) );
  INVX1 U8450 ( .A(n8527), .Y(n8525) );
  INVX1 U8451 ( .A(n8525), .Y(n8526) );
  AND2X1 U8452 ( .A(n10727), .B(n270), .Y(n316) );
  INVX1 U8453 ( .A(n316), .Y(n8527) );
  INVX1 U8454 ( .A(n8530), .Y(n8528) );
  INVX1 U8455 ( .A(n8528), .Y(n8529) );
  AND2X1 U8456 ( .A(n10730), .B(n270), .Y(n314) );
  INVX1 U8457 ( .A(n314), .Y(n8530) );
  INVX1 U8458 ( .A(n8533), .Y(n8531) );
  INVX1 U8459 ( .A(n8531), .Y(n8532) );
  AND2X1 U8460 ( .A(n10733), .B(n270), .Y(n312) );
  INVX1 U8461 ( .A(n312), .Y(n8533) );
  INVX1 U8462 ( .A(n8536), .Y(n8534) );
  INVX1 U8463 ( .A(n8534), .Y(n8535) );
  AND2X1 U8464 ( .A(n10736), .B(n270), .Y(n310) );
  INVX1 U8465 ( .A(n310), .Y(n8536) );
  INVX1 U8466 ( .A(n8539), .Y(n8537) );
  INVX1 U8467 ( .A(n8537), .Y(n8538) );
  AND2X1 U8468 ( .A(n10739), .B(n270), .Y(n308) );
  INVX1 U8469 ( .A(n308), .Y(n8539) );
  INVX1 U8470 ( .A(n8542), .Y(n8540) );
  INVX1 U8471 ( .A(n8540), .Y(n8541) );
  AND2X1 U8472 ( .A(n10742), .B(n270), .Y(n306) );
  INVX1 U8473 ( .A(n306), .Y(n8542) );
  INVX1 U8474 ( .A(n8545), .Y(n8543) );
  INVX1 U8475 ( .A(n8543), .Y(n8544) );
  AND2X1 U8476 ( .A(n10745), .B(n270), .Y(n304) );
  INVX1 U8477 ( .A(n304), .Y(n8545) );
  INVX1 U8478 ( .A(n8548), .Y(n8546) );
  INVX1 U8479 ( .A(n8546), .Y(n8547) );
  AND2X1 U8480 ( .A(n10748), .B(n270), .Y(n302) );
  INVX1 U8481 ( .A(n302), .Y(n8548) );
  INVX1 U8482 ( .A(n8551), .Y(n8549) );
  INVX1 U8483 ( .A(n8549), .Y(n8550) );
  AND2X1 U8484 ( .A(n10751), .B(n270), .Y(n300) );
  INVX1 U8485 ( .A(n300), .Y(n8551) );
  INVX1 U8486 ( .A(n8554), .Y(n8552) );
  INVX1 U8487 ( .A(n8552), .Y(n8553) );
  AND2X1 U8488 ( .A(n10754), .B(n270), .Y(n298) );
  INVX1 U8489 ( .A(n298), .Y(n8554) );
  INVX1 U8490 ( .A(n8557), .Y(n8555) );
  INVX1 U8491 ( .A(n8555), .Y(n8556) );
  AND2X1 U8492 ( .A(n10757), .B(n270), .Y(n296) );
  INVX1 U8493 ( .A(n296), .Y(n8557) );
  INVX1 U8494 ( .A(n8560), .Y(n8558) );
  INVX1 U8495 ( .A(n8558), .Y(n8559) );
  AND2X1 U8496 ( .A(n10760), .B(n270), .Y(n294) );
  INVX1 U8497 ( .A(n294), .Y(n8560) );
  INVX1 U8498 ( .A(n8563), .Y(n8561) );
  INVX1 U8499 ( .A(n8561), .Y(n8562) );
  AND2X1 U8500 ( .A(n10763), .B(n270), .Y(n292) );
  INVX1 U8501 ( .A(n292), .Y(n8563) );
  INVX1 U8502 ( .A(n8566), .Y(n8564) );
  INVX1 U8503 ( .A(n8564), .Y(n8565) );
  AND2X1 U8504 ( .A(n10766), .B(n270), .Y(n290) );
  INVX1 U8505 ( .A(n290), .Y(n8566) );
  INVX1 U8506 ( .A(n8569), .Y(n8567) );
  INVX1 U8507 ( .A(n8567), .Y(n8568) );
  AND2X1 U8508 ( .A(n10769), .B(n270), .Y(n288) );
  INVX1 U8509 ( .A(n288), .Y(n8569) );
  INVX1 U8510 ( .A(n8572), .Y(n8570) );
  INVX1 U8511 ( .A(n8570), .Y(n8571) );
  AND2X1 U8512 ( .A(n10772), .B(n270), .Y(n286) );
  INVX1 U8513 ( .A(n286), .Y(n8572) );
  INVX1 U8514 ( .A(n8575), .Y(n8573) );
  INVX1 U8515 ( .A(n8573), .Y(n8574) );
  AND2X1 U8516 ( .A(n10775), .B(n270), .Y(n284) );
  INVX1 U8517 ( .A(n284), .Y(n8575) );
  INVX1 U8518 ( .A(n8578), .Y(n8576) );
  INVX1 U8519 ( .A(n8576), .Y(n8577) );
  AND2X1 U8520 ( .A(n10778), .B(n270), .Y(n282) );
  INVX1 U8521 ( .A(n282), .Y(n8578) );
  INVX1 U8522 ( .A(n8581), .Y(n8579) );
  INVX1 U8523 ( .A(n8579), .Y(n8580) );
  AND2X1 U8524 ( .A(n10781), .B(n270), .Y(n280) );
  INVX1 U8525 ( .A(n280), .Y(n8581) );
  INVX1 U8526 ( .A(n8584), .Y(n8582) );
  INVX1 U8527 ( .A(n8582), .Y(n8583) );
  AND2X1 U8528 ( .A(n10784), .B(n270), .Y(n278) );
  INVX1 U8529 ( .A(n278), .Y(n8584) );
  INVX1 U8530 ( .A(n8587), .Y(n8585) );
  INVX1 U8531 ( .A(n8585), .Y(n8586) );
  AND2X1 U8532 ( .A(n10787), .B(n270), .Y(n276) );
  INVX1 U8533 ( .A(n276), .Y(n8587) );
  INVX1 U8534 ( .A(n8590), .Y(n8588) );
  INVX1 U8535 ( .A(n8588), .Y(n8589) );
  AND2X1 U8536 ( .A(n10790), .B(n270), .Y(n274) );
  INVX1 U8537 ( .A(n274), .Y(n8590) );
  INVX1 U8538 ( .A(n8593), .Y(n8591) );
  INVX1 U8539 ( .A(n8591), .Y(n8592) );
  AND2X1 U8540 ( .A(n10793), .B(n270), .Y(n272) );
  INVX1 U8541 ( .A(n272), .Y(n8593) );
  INVX1 U8542 ( .A(n8596), .Y(n8594) );
  INVX1 U8543 ( .A(n8594), .Y(n8595) );
  AND2X1 U8544 ( .A(n13357), .B(n201), .Y(n269) );
  INVX1 U8545 ( .A(n269), .Y(n8596) );
  INVX1 U8546 ( .A(n8599), .Y(n8597) );
  INVX1 U8547 ( .A(n8597), .Y(n8598) );
  AND2X1 U8548 ( .A(n118), .B(n201), .Y(n267) );
  INVX1 U8549 ( .A(n267), .Y(n8599) );
  INVX1 U8550 ( .A(n8602), .Y(n8600) );
  INVX1 U8551 ( .A(n8600), .Y(n8601) );
  AND2X1 U8552 ( .A(n38), .B(n253), .Y(n265) );
  INVX1 U8553 ( .A(n265), .Y(n8602) );
  INVX1 U8554 ( .A(n8605), .Y(n8603) );
  INVX1 U8555 ( .A(n8603), .Y(n8604) );
  AND2X1 U8556 ( .A(n34), .B(n253), .Y(n261) );
  INVX1 U8557 ( .A(n261), .Y(n8605) );
  INVX1 U8558 ( .A(n8608), .Y(n8606) );
  INVX1 U8559 ( .A(n8606), .Y(n8607) );
  AND2X1 U8560 ( .A(n35), .B(n253), .Y(n259) );
  INVX1 U8561 ( .A(n259), .Y(n8608) );
  INVX1 U8562 ( .A(n8611), .Y(n8609) );
  INVX1 U8563 ( .A(n8609), .Y(n8610) );
  AND2X1 U8564 ( .A(n36), .B(n253), .Y(n257) );
  INVX1 U8565 ( .A(n257), .Y(n8611) );
  INVX1 U8566 ( .A(n8614), .Y(n8612) );
  INVX1 U8567 ( .A(n8612), .Y(n8613) );
  AND2X1 U8568 ( .A(n37), .B(n253), .Y(n255) );
  INVX1 U8569 ( .A(n255), .Y(n8614) );
  INVX1 U8570 ( .A(n8617), .Y(n8615) );
  INVX1 U8571 ( .A(n8615), .Y(n8616) );
  AND2X1 U8572 ( .A(n114), .B(n201), .Y(n209) );
  INVX1 U8573 ( .A(n209), .Y(n8617) );
  INVX1 U8574 ( .A(n8620), .Y(n8618) );
  INVX1 U8575 ( .A(n8618), .Y(n8619) );
  AND2X1 U8576 ( .A(n115), .B(n201), .Y(n207) );
  INVX1 U8577 ( .A(n207), .Y(n8620) );
  INVX1 U8578 ( .A(n8623), .Y(n8621) );
  INVX1 U8579 ( .A(n8621), .Y(n8622) );
  AND2X1 U8580 ( .A(n116), .B(n201), .Y(n205) );
  INVX1 U8581 ( .A(n205), .Y(n8623) );
  INVX1 U8582 ( .A(n8626), .Y(n8624) );
  INVX1 U8583 ( .A(n8624), .Y(n8625) );
  AND2X1 U8584 ( .A(n117), .B(n201), .Y(n203) );
  INVX1 U8585 ( .A(n203), .Y(n8626) );
  INVX1 U8586 ( .A(n13043), .Y(n8627) );
  INVX1 U8587 ( .A(n8627), .Y(n8628) );
  INVX1 U8588 ( .A(n10802), .Y(n8629) );
  INVX1 U8589 ( .A(n8629), .Y(n8630) );
  INVX1 U8590 ( .A(n10800), .Y(n8631) );
  INVX1 U8591 ( .A(n8631), .Y(n8632) );
  INVX1 U8592 ( .A(n13039), .Y(n8633) );
  INVX1 U8593 ( .A(n8633), .Y(n8634) );
  INVX1 U8594 ( .A(n13035), .Y(n8635) );
  INVX1 U8595 ( .A(n8635), .Y(n8636) );
  INVX1 U8596 ( .A(n8770), .Y(n8637) );
  INVX1 U8597 ( .A(n8637), .Y(n8638) );
  INVX1 U8598 ( .A(n13039), .Y(n8639) );
  INVX1 U8599 ( .A(n8639), .Y(n8640) );
  INVX1 U8600 ( .A(n13035), .Y(n8641) );
  INVX1 U8601 ( .A(n8641), .Y(n8642) );
  INVX1 U8602 ( .A(n13043), .Y(n8643) );
  INVX1 U8603 ( .A(n8643), .Y(n8644) );
  INVX1 U8604 ( .A(n12960), .Y(n8645) );
  INVX1 U8605 ( .A(n8645), .Y(n8646) );
  INVX1 U8606 ( .A(n8770), .Y(n8647) );
  INVX1 U8607 ( .A(n8647), .Y(n8648) );
  INVX1 U8608 ( .A(n8770), .Y(n8649) );
  INVX1 U8609 ( .A(n8649), .Y(n8650) );
  INVX1 U8610 ( .A(n10800), .Y(n8651) );
  INVX1 U8611 ( .A(n8651), .Y(n8652) );
  INVX1 U8612 ( .A(n10802), .Y(n8653) );
  INVX1 U8613 ( .A(n8653), .Y(n8654) );
  INVX1 U8614 ( .A(n13035), .Y(n8655) );
  INVX1 U8615 ( .A(n8655), .Y(n8656) );
  INVX1 U8616 ( .A(n13039), .Y(n8657) );
  INVX1 U8617 ( .A(n8657), .Y(n8658) );
  INVX1 U8618 ( .A(n13043), .Y(n8659) );
  INVX1 U8619 ( .A(n8659), .Y(n8660) );
  INVX1 U8620 ( .A(n10796), .Y(n8661) );
  INVX1 U8621 ( .A(n8661), .Y(n8662) );
  INVX1 U8622 ( .A(n8770), .Y(n8663) );
  INVX1 U8623 ( .A(n8663), .Y(n8664) );
  INVX1 U8624 ( .A(n10800), .Y(n8665) );
  INVX1 U8625 ( .A(n8665), .Y(n8666) );
  INVX1 U8626 ( .A(n10802), .Y(n8667) );
  INVX1 U8627 ( .A(n8667), .Y(n8668) );
  INVX1 U8628 ( .A(n1705), .Y(n1401) );
  AND2X1 U8629 ( .A(n1401), .B(n13007), .Y(n13080) );
  AND2X1 U8630 ( .A(n1401), .B(n13004), .Y(n13081) );
  AND2X1 U8631 ( .A(n1401), .B(n13001), .Y(n13082) );
  AND2X1 U8632 ( .A(n1401), .B(n620), .Y(n13078) );
  INVX1 U8633 ( .A(n39), .Y(n8670) );
  INVX1 U8634 ( .A(n10802), .Y(n8671) );
  INVX1 U8635 ( .A(n8671), .Y(n8672) );
  INVX1 U8636 ( .A(n10800), .Y(n8673) );
  INVX1 U8637 ( .A(n8673), .Y(n8674) );
  INVX1 U8638 ( .A(n8708), .Y(n8675) );
  INVX1 U8639 ( .A(n8675), .Y(n8676) );
  INVX1 U8640 ( .A(n8684), .Y(n8677) );
  INVX1 U8641 ( .A(n8677), .Y(n8678) );
  INVX1 U8642 ( .A(n10800), .Y(n8679) );
  INVX1 U8643 ( .A(n8679), .Y(n8680) );
  INVX1 U8644 ( .A(n10802), .Y(n8681) );
  INVX1 U8645 ( .A(n8681), .Y(n8682) );
  INVX1 U8646 ( .A(n13043), .Y(n8683) );
  INVX1 U8647 ( .A(n8683), .Y(n8684) );
  INVX1 U8648 ( .A(n8714), .Y(n8685) );
  INVX1 U8649 ( .A(n8685), .Y(n8686) );
  INVX1 U8650 ( .A(n12960), .Y(n8687) );
  INVX1 U8651 ( .A(n8687), .Y(n8688) );
  INVX1 U8652 ( .A(n8708), .Y(n8689) );
  INVX1 U8653 ( .A(n8689), .Y(n8690) );
  INVX1 U8654 ( .A(n10800), .Y(n8691) );
  INVX1 U8655 ( .A(n8691), .Y(n8692) );
  INVX1 U8656 ( .A(n10802), .Y(n8693) );
  INVX1 U8657 ( .A(n8693), .Y(n8694) );
  INVX1 U8658 ( .A(n8720), .Y(n8695) );
  INVX1 U8659 ( .A(n8695), .Y(n8696) );
  INVX1 U8660 ( .A(n10800), .Y(n8697) );
  INVX1 U8661 ( .A(n8697), .Y(n8698) );
  INVX1 U8662 ( .A(n10800), .Y(n8699) );
  INVX1 U8663 ( .A(n8699), .Y(n8700) );
  INVX1 U8664 ( .A(n10802), .Y(n8701) );
  INVX1 U8665 ( .A(n8701), .Y(n8702) );
  INVX1 U8666 ( .A(n10802), .Y(n8703) );
  INVX1 U8667 ( .A(n8703), .Y(n8704) );
  INVX1 U8668 ( .A(n8714), .Y(n8705) );
  INVX1 U8669 ( .A(n8705), .Y(n8706) );
  INVX1 U8670 ( .A(n13043), .Y(n8707) );
  INVX1 U8671 ( .A(n8707), .Y(n8708) );
  INVX1 U8672 ( .A(n10802), .Y(n8709) );
  INVX1 U8673 ( .A(n8709), .Y(n8710) );
  INVX1 U8674 ( .A(n10800), .Y(n8711) );
  INVX1 U8675 ( .A(n8711), .Y(n8712) );
  INVX1 U8676 ( .A(n10796), .Y(n8713) );
  INVX1 U8677 ( .A(n8713), .Y(n8714) );
  INVX1 U8678 ( .A(n10802), .Y(n8715) );
  INVX1 U8679 ( .A(n8715), .Y(n8716) );
  INVX1 U8680 ( .A(n10800), .Y(n8717) );
  INVX1 U8681 ( .A(n8717), .Y(n8718) );
  INVX1 U8682 ( .A(n13043), .Y(n8719) );
  INVX1 U8683 ( .A(n8719), .Y(n8720) );
  INVX1 U8684 ( .A(n10800), .Y(n8721) );
  INVX1 U8685 ( .A(n8721), .Y(n8722) );
  INVX1 U8686 ( .A(n10802), .Y(n8723) );
  INVX1 U8687 ( .A(n8723), .Y(n8724) );
  INVX1 U8688 ( .A(n8727), .Y(n8725) );
  INVX1 U8689 ( .A(n8725), .Y(n8726) );
  BUFX2 U8690 ( .A(n1718), .Y(n8727) );
  INVX1 U8691 ( .A(n13061), .Y(n8728) );
  INVX1 U8692 ( .A(n8728), .Y(n8729) );
  INVX1 U8693 ( .A(n8732), .Y(n8730) );
  INVX1 U8694 ( .A(n8730), .Y(n8731) );
  OR2X1 U8695 ( .A(n1711), .B(n1712), .Y(n1710) );
  INVX1 U8696 ( .A(n1710), .Y(n8732) );
  INVX1 U8697 ( .A(n8735), .Y(n8733) );
  INVX1 U8698 ( .A(n8733), .Y(n8734) );
  BUFX2 U8699 ( .A(wr_ptr_gray_ss[2]), .Y(n8735) );
  INVX1 U8700 ( .A(n8738), .Y(n8736) );
  INVX1 U8701 ( .A(n8736), .Y(n8737) );
  BUFX2 U8702 ( .A(wr_ptr_gray_ss[4]), .Y(n8738) );
  INVX1 U8703 ( .A(n8741), .Y(n8739) );
  INVX1 U8704 ( .A(n8739), .Y(n8740) );
  BUFX2 U8705 ( .A(wr_ptr_gray_ss[3]), .Y(n8741) );
  INVX1 U8706 ( .A(n8744), .Y(n8742) );
  INVX1 U8707 ( .A(n8742), .Y(n8743) );
  BUFX2 U8708 ( .A(wr_ptr_gray_ss[0]), .Y(n8744) );
  INVX1 U8709 ( .A(n8756), .Y(n8745) );
  INVX1 U8710 ( .A(n8745), .Y(n8746) );
  INVX1 U8711 ( .A(n8754), .Y(n8747) );
  INVX1 U8712 ( .A(n8747), .Y(n8748) );
  INVX1 U8713 ( .A(n13024), .Y(n8749) );
  INVX1 U8714 ( .A(n8749), .Y(n8750) );
  INVX1 U8715 ( .A(n8764), .Y(n8751) );
  INVX1 U8716 ( .A(n8751), .Y(n8752) );
  INVX1 U8717 ( .A(n268), .Y(n8753) );
  INVX1 U8718 ( .A(n8753), .Y(n8754) );
  INVX1 U8719 ( .A(n796), .Y(n8755) );
  INVX1 U8720 ( .A(n8755), .Y(n8756) );
  INVX1 U8721 ( .A(n8766), .Y(n8757) );
  INVX1 U8722 ( .A(n8757), .Y(n8758) );
  INVX1 U8723 ( .A(n8768), .Y(n8759) );
  INVX1 U8724 ( .A(n8759), .Y(n8760) );
  INVX1 U8725 ( .A(n13045), .Y(n8761) );
  INVX1 U8726 ( .A(n8761), .Y(n8762) );
  INVX8 U8727 ( .A(n13044), .Y(n13045) );
  INVX1 U8728 ( .A(n8750), .Y(n8763) );
  INVX1 U8729 ( .A(n8763), .Y(n8764) );
  INVX1 U8730 ( .A(n8746), .Y(n8765) );
  INVX1 U8731 ( .A(n8765), .Y(n8766) );
  INVX1 U8732 ( .A(n8748), .Y(n8767) );
  INVX1 U8733 ( .A(n8767), .Y(n8768) );
  INVX1 U8734 ( .A(n8752), .Y(n8769) );
  INVX1 U8735 ( .A(n8769), .Y(n8770) );
  INVX1 U8736 ( .A(n8760), .Y(n8771) );
  INVX1 U8737 ( .A(n8771), .Y(n8772) );
  INVX1 U8738 ( .A(n8758), .Y(n8774) );
  INVX1 U8739 ( .A(n8774), .Y(n8775) );
  INVX1 U8740 ( .A(n13062), .Y(n8777) );
  INVX1 U8741 ( .A(n40), .Y(n13062) );
  INVX1 U8742 ( .A(n12976), .Y(n8778) );
  INVX1 U8743 ( .A(n8781), .Y(n8779) );
  INVX1 U8744 ( .A(n8779), .Y(n8780) );
  BUFX2 U8745 ( .A(fifo[42]), .Y(n8781) );
  INVX1 U8746 ( .A(n8784), .Y(n8782) );
  INVX1 U8747 ( .A(n8782), .Y(n8783) );
  BUFX2 U8748 ( .A(fifo[43]), .Y(n8784) );
  INVX1 U8749 ( .A(n8787), .Y(n8785) );
  INVX1 U8750 ( .A(n8785), .Y(n8786) );
  BUFX2 U8751 ( .A(fifo[44]), .Y(n8787) );
  INVX1 U8752 ( .A(n8790), .Y(n8788) );
  INVX1 U8753 ( .A(n8788), .Y(n8789) );
  BUFX2 U8754 ( .A(fifo[45]), .Y(n8790) );
  INVX1 U8755 ( .A(n8793), .Y(n8791) );
  INVX1 U8756 ( .A(n8791), .Y(n8792) );
  BUFX2 U8757 ( .A(fifo[46]), .Y(n8793) );
  INVX1 U8758 ( .A(n8796), .Y(n8794) );
  INVX1 U8759 ( .A(n8794), .Y(n8795) );
  BUFX2 U8760 ( .A(fifo[47]), .Y(n8796) );
  INVX1 U8761 ( .A(n8799), .Y(n8797) );
  INVX1 U8762 ( .A(n8797), .Y(n8798) );
  BUFX2 U8763 ( .A(fifo[48]), .Y(n8799) );
  INVX1 U8764 ( .A(n8802), .Y(n8800) );
  INVX1 U8765 ( .A(n8800), .Y(n8801) );
  BUFX2 U8766 ( .A(fifo[49]), .Y(n8802) );
  INVX1 U8767 ( .A(n8805), .Y(n8803) );
  INVX1 U8768 ( .A(n8803), .Y(n8804) );
  BUFX2 U8769 ( .A(fifo[50]), .Y(n8805) );
  INVX1 U8770 ( .A(n8808), .Y(n8806) );
  INVX1 U8771 ( .A(n8806), .Y(n8807) );
  BUFX2 U8772 ( .A(fifo[51]), .Y(n8808) );
  INVX1 U8773 ( .A(n8811), .Y(n8809) );
  INVX1 U8774 ( .A(n8809), .Y(n8810) );
  BUFX2 U8775 ( .A(fifo[52]), .Y(n8811) );
  INVX1 U8776 ( .A(n8814), .Y(n8812) );
  INVX1 U8777 ( .A(n8812), .Y(n8813) );
  BUFX2 U8778 ( .A(fifo[53]), .Y(n8814) );
  INVX1 U8779 ( .A(n8817), .Y(n8815) );
  INVX1 U8780 ( .A(n8815), .Y(n8816) );
  BUFX2 U8781 ( .A(fifo[54]), .Y(n8817) );
  INVX1 U8782 ( .A(n8820), .Y(n8818) );
  INVX1 U8783 ( .A(n8818), .Y(n8819) );
  BUFX2 U8784 ( .A(fifo[55]), .Y(n8820) );
  INVX1 U8785 ( .A(n8823), .Y(n8821) );
  INVX1 U8786 ( .A(n8821), .Y(n8822) );
  BUFX2 U8787 ( .A(fifo[56]), .Y(n8823) );
  INVX1 U8788 ( .A(n8826), .Y(n8824) );
  INVX1 U8789 ( .A(n8824), .Y(n8825) );
  BUFX2 U8790 ( .A(fifo[57]), .Y(n8826) );
  INVX1 U8791 ( .A(n8829), .Y(n8827) );
  INVX1 U8792 ( .A(n8827), .Y(n8828) );
  BUFX2 U8793 ( .A(fifo[58]), .Y(n8829) );
  INVX1 U8794 ( .A(n8832), .Y(n8830) );
  INVX1 U8795 ( .A(n8830), .Y(n8831) );
  BUFX2 U8796 ( .A(fifo[59]), .Y(n8832) );
  INVX1 U8797 ( .A(n8835), .Y(n8833) );
  INVX1 U8798 ( .A(n8833), .Y(n8834) );
  BUFX2 U8799 ( .A(fifo[60]), .Y(n8835) );
  INVX1 U8800 ( .A(n8838), .Y(n8836) );
  INVX1 U8801 ( .A(n8836), .Y(n8837) );
  BUFX2 U8802 ( .A(fifo[61]), .Y(n8838) );
  INVX1 U8803 ( .A(n8841), .Y(n8839) );
  INVX1 U8804 ( .A(n8839), .Y(n8840) );
  BUFX2 U8805 ( .A(fifo[62]), .Y(n8841) );
  INVX1 U8806 ( .A(n8844), .Y(n8842) );
  INVX1 U8807 ( .A(n8842), .Y(n8843) );
  BUFX2 U8808 ( .A(fifo[63]), .Y(n8844) );
  INVX1 U8809 ( .A(n8847), .Y(n8845) );
  INVX1 U8810 ( .A(n8845), .Y(n8846) );
  BUFX2 U8811 ( .A(fifo[64]), .Y(n8847) );
  INVX1 U8812 ( .A(n8850), .Y(n8848) );
  INVX1 U8813 ( .A(n8848), .Y(n8849) );
  BUFX2 U8814 ( .A(fifo[65]), .Y(n8850) );
  INVX1 U8815 ( .A(n8853), .Y(n8851) );
  INVX1 U8816 ( .A(n8851), .Y(n8852) );
  BUFX2 U8817 ( .A(fifo[66]), .Y(n8853) );
  INVX1 U8818 ( .A(n8856), .Y(n8854) );
  INVX1 U8819 ( .A(n8854), .Y(n8855) );
  BUFX2 U8820 ( .A(fifo[67]), .Y(n8856) );
  INVX1 U8821 ( .A(n8859), .Y(n8857) );
  INVX1 U8822 ( .A(n8857), .Y(n8858) );
  BUFX2 U8823 ( .A(fifo[68]), .Y(n8859) );
  INVX1 U8824 ( .A(n8862), .Y(n8860) );
  INVX1 U8825 ( .A(n8860), .Y(n8861) );
  BUFX2 U8826 ( .A(fifo[69]), .Y(n8862) );
  INVX1 U8827 ( .A(n8865), .Y(n8863) );
  INVX1 U8828 ( .A(n8863), .Y(n8864) );
  BUFX2 U8829 ( .A(fifo[70]), .Y(n8865) );
  INVX1 U8830 ( .A(n8868), .Y(n8866) );
  INVX1 U8831 ( .A(n8866), .Y(n8867) );
  BUFX2 U8832 ( .A(fifo[71]), .Y(n8868) );
  INVX1 U8833 ( .A(n8871), .Y(n8869) );
  INVX1 U8834 ( .A(n8869), .Y(n8870) );
  BUFX2 U8835 ( .A(fifo[72]), .Y(n8871) );
  INVX1 U8836 ( .A(n8874), .Y(n8872) );
  INVX1 U8837 ( .A(n8872), .Y(n8873) );
  BUFX2 U8838 ( .A(fifo[73]), .Y(n8874) );
  INVX1 U8839 ( .A(n8877), .Y(n8875) );
  INVX1 U8840 ( .A(n8875), .Y(n8876) );
  BUFX2 U8841 ( .A(fifo[74]), .Y(n8877) );
  INVX1 U8842 ( .A(n8880), .Y(n8878) );
  INVX1 U8843 ( .A(n8878), .Y(n8879) );
  BUFX2 U8844 ( .A(fifo[75]), .Y(n8880) );
  INVX1 U8845 ( .A(n8883), .Y(n8881) );
  INVX1 U8846 ( .A(n8881), .Y(n8882) );
  BUFX2 U8847 ( .A(fifo[76]), .Y(n8883) );
  INVX1 U8848 ( .A(n8886), .Y(n8884) );
  INVX1 U8849 ( .A(n8884), .Y(n8885) );
  BUFX2 U8850 ( .A(fifo[77]), .Y(n8886) );
  INVX1 U8851 ( .A(n8889), .Y(n8887) );
  INVX1 U8852 ( .A(n8887), .Y(n8888) );
  BUFX2 U8853 ( .A(fifo[78]), .Y(n8889) );
  INVX1 U8854 ( .A(n8892), .Y(n8890) );
  INVX1 U8855 ( .A(n8890), .Y(n8891) );
  BUFX2 U8856 ( .A(fifo[79]), .Y(n8892) );
  INVX1 U8857 ( .A(n8895), .Y(n8893) );
  INVX1 U8858 ( .A(n8893), .Y(n8894) );
  BUFX2 U8859 ( .A(fifo[80]), .Y(n8895) );
  INVX1 U8860 ( .A(n8898), .Y(n8896) );
  INVX1 U8861 ( .A(n8896), .Y(n8897) );
  BUFX2 U8862 ( .A(fifo[81]), .Y(n8898) );
  INVX1 U8863 ( .A(n8901), .Y(n8899) );
  INVX1 U8864 ( .A(n8899), .Y(n8900) );
  BUFX2 U8865 ( .A(fifo[82]), .Y(n8901) );
  INVX1 U8866 ( .A(n8904), .Y(n8902) );
  INVX1 U8867 ( .A(n8902), .Y(n8903) );
  BUFX2 U8868 ( .A(fifo[83]), .Y(n8904) );
  INVX1 U8869 ( .A(n8907), .Y(n8905) );
  INVX1 U8870 ( .A(n8905), .Y(n8906) );
  BUFX2 U8871 ( .A(fifo[126]), .Y(n8907) );
  INVX1 U8872 ( .A(n8910), .Y(n8908) );
  INVX1 U8873 ( .A(n8908), .Y(n8909) );
  BUFX2 U8874 ( .A(fifo[127]), .Y(n8910) );
  INVX1 U8875 ( .A(n8913), .Y(n8911) );
  INVX1 U8876 ( .A(n8911), .Y(n8912) );
  BUFX2 U8877 ( .A(fifo[128]), .Y(n8913) );
  INVX1 U8878 ( .A(n8916), .Y(n8914) );
  INVX1 U8879 ( .A(n8914), .Y(n8915) );
  BUFX2 U8880 ( .A(fifo[129]), .Y(n8916) );
  INVX1 U8881 ( .A(n8919), .Y(n8917) );
  INVX1 U8882 ( .A(n8917), .Y(n8918) );
  BUFX2 U8883 ( .A(fifo[130]), .Y(n8919) );
  INVX1 U8884 ( .A(n8922), .Y(n8920) );
  INVX1 U8885 ( .A(n8920), .Y(n8921) );
  BUFX2 U8886 ( .A(fifo[131]), .Y(n8922) );
  INVX1 U8887 ( .A(n8925), .Y(n8923) );
  INVX1 U8888 ( .A(n8923), .Y(n8924) );
  BUFX2 U8889 ( .A(fifo[132]), .Y(n8925) );
  INVX1 U8890 ( .A(n8928), .Y(n8926) );
  INVX1 U8891 ( .A(n8926), .Y(n8927) );
  BUFX2 U8892 ( .A(fifo[133]), .Y(n8928) );
  INVX1 U8893 ( .A(n8931), .Y(n8929) );
  INVX1 U8894 ( .A(n8929), .Y(n8930) );
  BUFX2 U8895 ( .A(fifo[134]), .Y(n8931) );
  INVX1 U8896 ( .A(n8934), .Y(n8932) );
  INVX1 U8897 ( .A(n8932), .Y(n8933) );
  BUFX2 U8898 ( .A(fifo[135]), .Y(n8934) );
  INVX1 U8899 ( .A(n8937), .Y(n8935) );
  INVX1 U8900 ( .A(n8935), .Y(n8936) );
  BUFX2 U8901 ( .A(fifo[136]), .Y(n8937) );
  INVX1 U8902 ( .A(n8940), .Y(n8938) );
  INVX1 U8903 ( .A(n8938), .Y(n8939) );
  BUFX2 U8904 ( .A(fifo[137]), .Y(n8940) );
  INVX1 U8905 ( .A(n8943), .Y(n8941) );
  INVX1 U8906 ( .A(n8941), .Y(n8942) );
  BUFX2 U8907 ( .A(fifo[138]), .Y(n8943) );
  INVX1 U8908 ( .A(n8946), .Y(n8944) );
  INVX1 U8909 ( .A(n8944), .Y(n8945) );
  BUFX2 U8910 ( .A(fifo[139]), .Y(n8946) );
  INVX1 U8911 ( .A(n8949), .Y(n8947) );
  INVX1 U8912 ( .A(n8947), .Y(n8948) );
  BUFX2 U8913 ( .A(fifo[140]), .Y(n8949) );
  INVX1 U8914 ( .A(n8952), .Y(n8950) );
  INVX1 U8915 ( .A(n8950), .Y(n8951) );
  BUFX2 U8916 ( .A(fifo[141]), .Y(n8952) );
  INVX1 U8917 ( .A(n8955), .Y(n8953) );
  INVX1 U8918 ( .A(n8953), .Y(n8954) );
  BUFX2 U8919 ( .A(fifo[142]), .Y(n8955) );
  INVX1 U8920 ( .A(n8958), .Y(n8956) );
  INVX1 U8921 ( .A(n8956), .Y(n8957) );
  BUFX2 U8922 ( .A(fifo[143]), .Y(n8958) );
  INVX1 U8923 ( .A(n8961), .Y(n8959) );
  INVX1 U8924 ( .A(n8959), .Y(n8960) );
  BUFX2 U8925 ( .A(fifo[144]), .Y(n8961) );
  INVX1 U8926 ( .A(n8964), .Y(n8962) );
  INVX1 U8927 ( .A(n8962), .Y(n8963) );
  BUFX2 U8928 ( .A(fifo[145]), .Y(n8964) );
  INVX1 U8929 ( .A(n8967), .Y(n8965) );
  INVX1 U8930 ( .A(n8965), .Y(n8966) );
  BUFX2 U8931 ( .A(fifo[146]), .Y(n8967) );
  INVX1 U8932 ( .A(n8970), .Y(n8968) );
  INVX1 U8933 ( .A(n8968), .Y(n8969) );
  BUFX2 U8934 ( .A(fifo[147]), .Y(n8970) );
  INVX1 U8935 ( .A(n8973), .Y(n8971) );
  INVX1 U8936 ( .A(n8971), .Y(n8972) );
  BUFX2 U8937 ( .A(fifo[148]), .Y(n8973) );
  INVX1 U8938 ( .A(n8976), .Y(n8974) );
  INVX1 U8939 ( .A(n8974), .Y(n8975) );
  BUFX2 U8940 ( .A(fifo[149]), .Y(n8976) );
  INVX1 U8941 ( .A(n8979), .Y(n8977) );
  INVX1 U8942 ( .A(n8977), .Y(n8978) );
  BUFX2 U8943 ( .A(fifo[150]), .Y(n8979) );
  INVX1 U8944 ( .A(n8982), .Y(n8980) );
  INVX1 U8945 ( .A(n8980), .Y(n8981) );
  BUFX2 U8946 ( .A(fifo[151]), .Y(n8982) );
  INVX1 U8947 ( .A(n8985), .Y(n8983) );
  INVX1 U8948 ( .A(n8983), .Y(n8984) );
  BUFX2 U8949 ( .A(fifo[152]), .Y(n8985) );
  INVX1 U8950 ( .A(n8988), .Y(n8986) );
  INVX1 U8951 ( .A(n8986), .Y(n8987) );
  BUFX2 U8952 ( .A(fifo[153]), .Y(n8988) );
  INVX1 U8953 ( .A(n8991), .Y(n8989) );
  INVX1 U8954 ( .A(n8989), .Y(n8990) );
  BUFX2 U8955 ( .A(fifo[154]), .Y(n8991) );
  INVX1 U8956 ( .A(n8994), .Y(n8992) );
  INVX1 U8957 ( .A(n8992), .Y(n8993) );
  BUFX2 U8958 ( .A(fifo[155]), .Y(n8994) );
  INVX1 U8959 ( .A(n8997), .Y(n8995) );
  INVX1 U8960 ( .A(n8995), .Y(n8996) );
  BUFX2 U8961 ( .A(fifo[156]), .Y(n8997) );
  INVX1 U8962 ( .A(n9000), .Y(n8998) );
  INVX1 U8963 ( .A(n8998), .Y(n8999) );
  BUFX2 U8964 ( .A(fifo[157]), .Y(n9000) );
  INVX1 U8965 ( .A(n9003), .Y(n9001) );
  INVX1 U8966 ( .A(n9001), .Y(n9002) );
  BUFX2 U8967 ( .A(fifo[158]), .Y(n9003) );
  INVX1 U8968 ( .A(n9006), .Y(n9004) );
  INVX1 U8969 ( .A(n9004), .Y(n9005) );
  BUFX2 U8970 ( .A(fifo[159]), .Y(n9006) );
  INVX1 U8971 ( .A(n9009), .Y(n9007) );
  INVX1 U8972 ( .A(n9007), .Y(n9008) );
  BUFX2 U8973 ( .A(fifo[160]), .Y(n9009) );
  INVX1 U8974 ( .A(n9012), .Y(n9010) );
  INVX1 U8975 ( .A(n9010), .Y(n9011) );
  BUFX2 U8976 ( .A(fifo[161]), .Y(n9012) );
  INVX1 U8977 ( .A(n9015), .Y(n9013) );
  INVX1 U8978 ( .A(n9013), .Y(n9014) );
  BUFX2 U8979 ( .A(fifo[162]), .Y(n9015) );
  INVX1 U8980 ( .A(n9018), .Y(n9016) );
  INVX1 U8981 ( .A(n9016), .Y(n9017) );
  BUFX2 U8982 ( .A(fifo[163]), .Y(n9018) );
  INVX1 U8983 ( .A(n9021), .Y(n9019) );
  INVX1 U8984 ( .A(n9019), .Y(n9020) );
  BUFX2 U8985 ( .A(fifo[164]), .Y(n9021) );
  INVX1 U8986 ( .A(n9024), .Y(n9022) );
  INVX1 U8987 ( .A(n9022), .Y(n9023) );
  BUFX2 U8988 ( .A(fifo[165]), .Y(n9024) );
  INVX1 U8989 ( .A(n9027), .Y(n9025) );
  INVX1 U8990 ( .A(n9025), .Y(n9026) );
  BUFX2 U8991 ( .A(fifo[166]), .Y(n9027) );
  INVX1 U8992 ( .A(n9030), .Y(n9028) );
  INVX1 U8993 ( .A(n9028), .Y(n9029) );
  BUFX2 U8994 ( .A(fifo[167]), .Y(n9030) );
  INVX1 U8995 ( .A(n9033), .Y(n9031) );
  INVX1 U8996 ( .A(n9031), .Y(n9032) );
  BUFX2 U8997 ( .A(fifo[210]), .Y(n9033) );
  INVX1 U8998 ( .A(n9036), .Y(n9034) );
  INVX1 U8999 ( .A(n9034), .Y(n9035) );
  BUFX2 U9000 ( .A(fifo[211]), .Y(n9036) );
  INVX1 U9001 ( .A(n9039), .Y(n9037) );
  INVX1 U9002 ( .A(n9037), .Y(n9038) );
  BUFX2 U9003 ( .A(fifo[212]), .Y(n9039) );
  INVX1 U9004 ( .A(n9042), .Y(n9040) );
  INVX1 U9005 ( .A(n9040), .Y(n9041) );
  BUFX2 U9006 ( .A(fifo[213]), .Y(n9042) );
  INVX1 U9007 ( .A(n9045), .Y(n9043) );
  INVX1 U9008 ( .A(n9043), .Y(n9044) );
  BUFX2 U9009 ( .A(fifo[214]), .Y(n9045) );
  INVX1 U9010 ( .A(n9048), .Y(n9046) );
  INVX1 U9011 ( .A(n9046), .Y(n9047) );
  BUFX2 U9012 ( .A(fifo[215]), .Y(n9048) );
  INVX1 U9013 ( .A(n9051), .Y(n9049) );
  INVX1 U9014 ( .A(n9049), .Y(n9050) );
  BUFX2 U9015 ( .A(fifo[216]), .Y(n9051) );
  INVX1 U9016 ( .A(n9054), .Y(n9052) );
  INVX1 U9017 ( .A(n9052), .Y(n9053) );
  BUFX2 U9018 ( .A(fifo[217]), .Y(n9054) );
  INVX1 U9019 ( .A(n9057), .Y(n9055) );
  INVX1 U9020 ( .A(n9055), .Y(n9056) );
  BUFX2 U9021 ( .A(fifo[218]), .Y(n9057) );
  INVX1 U9022 ( .A(n9060), .Y(n9058) );
  INVX1 U9023 ( .A(n9058), .Y(n9059) );
  BUFX2 U9024 ( .A(fifo[219]), .Y(n9060) );
  INVX1 U9025 ( .A(n9063), .Y(n9061) );
  INVX1 U9026 ( .A(n9061), .Y(n9062) );
  BUFX2 U9027 ( .A(fifo[220]), .Y(n9063) );
  INVX1 U9028 ( .A(n9066), .Y(n9064) );
  INVX1 U9029 ( .A(n9064), .Y(n9065) );
  BUFX2 U9030 ( .A(fifo[221]), .Y(n9066) );
  INVX1 U9031 ( .A(n9069), .Y(n9067) );
  INVX1 U9032 ( .A(n9067), .Y(n9068) );
  BUFX2 U9033 ( .A(fifo[222]), .Y(n9069) );
  INVX1 U9034 ( .A(n9072), .Y(n9070) );
  INVX1 U9035 ( .A(n9070), .Y(n9071) );
  BUFX2 U9036 ( .A(fifo[223]), .Y(n9072) );
  INVX1 U9037 ( .A(n9075), .Y(n9073) );
  INVX1 U9038 ( .A(n9073), .Y(n9074) );
  BUFX2 U9039 ( .A(fifo[224]), .Y(n9075) );
  INVX1 U9040 ( .A(n9078), .Y(n9076) );
  INVX1 U9041 ( .A(n9076), .Y(n9077) );
  BUFX2 U9042 ( .A(fifo[225]), .Y(n9078) );
  INVX1 U9043 ( .A(n9081), .Y(n9079) );
  INVX1 U9044 ( .A(n9079), .Y(n9080) );
  BUFX2 U9045 ( .A(fifo[226]), .Y(n9081) );
  INVX1 U9046 ( .A(n9084), .Y(n9082) );
  INVX1 U9047 ( .A(n9082), .Y(n9083) );
  BUFX2 U9048 ( .A(fifo[227]), .Y(n9084) );
  INVX1 U9049 ( .A(n9087), .Y(n9085) );
  INVX1 U9050 ( .A(n9085), .Y(n9086) );
  BUFX2 U9051 ( .A(fifo[228]), .Y(n9087) );
  INVX1 U9052 ( .A(n9090), .Y(n9088) );
  INVX1 U9053 ( .A(n9088), .Y(n9089) );
  BUFX2 U9054 ( .A(fifo[229]), .Y(n9090) );
  INVX1 U9055 ( .A(n9093), .Y(n9091) );
  INVX1 U9056 ( .A(n9091), .Y(n9092) );
  BUFX2 U9057 ( .A(fifo[230]), .Y(n9093) );
  INVX1 U9058 ( .A(n9096), .Y(n9094) );
  INVX1 U9059 ( .A(n9094), .Y(n9095) );
  BUFX2 U9060 ( .A(fifo[231]), .Y(n9096) );
  INVX1 U9061 ( .A(n9099), .Y(n9097) );
  INVX1 U9062 ( .A(n9097), .Y(n9098) );
  BUFX2 U9063 ( .A(fifo[232]), .Y(n9099) );
  INVX1 U9064 ( .A(n9102), .Y(n9100) );
  INVX1 U9065 ( .A(n9100), .Y(n9101) );
  BUFX2 U9066 ( .A(fifo[233]), .Y(n9102) );
  INVX1 U9067 ( .A(n9105), .Y(n9103) );
  INVX1 U9068 ( .A(n9103), .Y(n9104) );
  BUFX2 U9069 ( .A(fifo[234]), .Y(n9105) );
  INVX1 U9070 ( .A(n9108), .Y(n9106) );
  INVX1 U9071 ( .A(n9106), .Y(n9107) );
  BUFX2 U9072 ( .A(fifo[235]), .Y(n9108) );
  INVX1 U9073 ( .A(n9111), .Y(n9109) );
  INVX1 U9074 ( .A(n9109), .Y(n9110) );
  BUFX2 U9075 ( .A(fifo[236]), .Y(n9111) );
  INVX1 U9076 ( .A(n9114), .Y(n9112) );
  INVX1 U9077 ( .A(n9112), .Y(n9113) );
  BUFX2 U9078 ( .A(fifo[237]), .Y(n9114) );
  INVX1 U9079 ( .A(n9117), .Y(n9115) );
  INVX1 U9080 ( .A(n9115), .Y(n9116) );
  BUFX2 U9081 ( .A(fifo[238]), .Y(n9117) );
  INVX1 U9082 ( .A(n9120), .Y(n9118) );
  INVX1 U9083 ( .A(n9118), .Y(n9119) );
  BUFX2 U9084 ( .A(fifo[239]), .Y(n9120) );
  INVX1 U9085 ( .A(n9123), .Y(n9121) );
  INVX1 U9086 ( .A(n9121), .Y(n9122) );
  BUFX2 U9087 ( .A(fifo[240]), .Y(n9123) );
  INVX1 U9088 ( .A(n9126), .Y(n9124) );
  INVX1 U9089 ( .A(n9124), .Y(n9125) );
  BUFX2 U9090 ( .A(fifo[241]), .Y(n9126) );
  INVX1 U9091 ( .A(n9129), .Y(n9127) );
  INVX1 U9092 ( .A(n9127), .Y(n9128) );
  BUFX2 U9093 ( .A(fifo[242]), .Y(n9129) );
  INVX1 U9094 ( .A(n9132), .Y(n9130) );
  INVX1 U9095 ( .A(n9130), .Y(n9131) );
  BUFX2 U9096 ( .A(fifo[243]), .Y(n9132) );
  INVX1 U9097 ( .A(n9135), .Y(n9133) );
  INVX1 U9098 ( .A(n9133), .Y(n9134) );
  BUFX2 U9099 ( .A(fifo[244]), .Y(n9135) );
  INVX1 U9100 ( .A(n9138), .Y(n9136) );
  INVX1 U9101 ( .A(n9136), .Y(n9137) );
  BUFX2 U9102 ( .A(fifo[245]), .Y(n9138) );
  INVX1 U9103 ( .A(n9141), .Y(n9139) );
  INVX1 U9104 ( .A(n9139), .Y(n9140) );
  BUFX2 U9105 ( .A(fifo[246]), .Y(n9141) );
  INVX1 U9106 ( .A(n9144), .Y(n9142) );
  INVX1 U9107 ( .A(n9142), .Y(n9143) );
  BUFX2 U9108 ( .A(fifo[247]), .Y(n9144) );
  INVX1 U9109 ( .A(n9147), .Y(n9145) );
  INVX1 U9110 ( .A(n9145), .Y(n9146) );
  BUFX2 U9111 ( .A(fifo[248]), .Y(n9147) );
  INVX1 U9112 ( .A(n9150), .Y(n9148) );
  INVX1 U9113 ( .A(n9148), .Y(n9149) );
  BUFX2 U9114 ( .A(fifo[249]), .Y(n9150) );
  INVX1 U9115 ( .A(n9153), .Y(n9151) );
  INVX1 U9116 ( .A(n9151), .Y(n9152) );
  BUFX2 U9117 ( .A(fifo[250]), .Y(n9153) );
  INVX1 U9118 ( .A(n9156), .Y(n9154) );
  INVX1 U9119 ( .A(n9154), .Y(n9155) );
  BUFX2 U9120 ( .A(fifo[251]), .Y(n9156) );
  INVX1 U9121 ( .A(n9159), .Y(n9157) );
  INVX1 U9122 ( .A(n9157), .Y(n9158) );
  BUFX2 U9123 ( .A(fifo[294]), .Y(n9159) );
  INVX1 U9124 ( .A(n9162), .Y(n9160) );
  INVX1 U9125 ( .A(n9160), .Y(n9161) );
  BUFX2 U9126 ( .A(fifo[295]), .Y(n9162) );
  INVX1 U9127 ( .A(n9165), .Y(n9163) );
  INVX1 U9128 ( .A(n9163), .Y(n9164) );
  BUFX2 U9129 ( .A(fifo[296]), .Y(n9165) );
  INVX1 U9130 ( .A(n9168), .Y(n9166) );
  INVX1 U9131 ( .A(n9166), .Y(n9167) );
  BUFX2 U9132 ( .A(fifo[297]), .Y(n9168) );
  INVX1 U9133 ( .A(n9171), .Y(n9169) );
  INVX1 U9134 ( .A(n9169), .Y(n9170) );
  BUFX2 U9135 ( .A(fifo[298]), .Y(n9171) );
  INVX1 U9136 ( .A(n9174), .Y(n9172) );
  INVX1 U9137 ( .A(n9172), .Y(n9173) );
  BUFX2 U9138 ( .A(fifo[299]), .Y(n9174) );
  INVX1 U9139 ( .A(n9177), .Y(n9175) );
  INVX1 U9140 ( .A(n9175), .Y(n9176) );
  BUFX2 U9141 ( .A(fifo[300]), .Y(n9177) );
  INVX1 U9142 ( .A(n9180), .Y(n9178) );
  INVX1 U9143 ( .A(n9178), .Y(n9179) );
  BUFX2 U9144 ( .A(fifo[301]), .Y(n9180) );
  INVX1 U9145 ( .A(n9183), .Y(n9181) );
  INVX1 U9146 ( .A(n9181), .Y(n9182) );
  BUFX2 U9147 ( .A(fifo[302]), .Y(n9183) );
  INVX1 U9148 ( .A(n9186), .Y(n9184) );
  INVX1 U9149 ( .A(n9184), .Y(n9185) );
  BUFX2 U9150 ( .A(fifo[303]), .Y(n9186) );
  INVX1 U9151 ( .A(n9189), .Y(n9187) );
  INVX1 U9152 ( .A(n9187), .Y(n9188) );
  BUFX2 U9153 ( .A(fifo[304]), .Y(n9189) );
  INVX1 U9154 ( .A(n9192), .Y(n9190) );
  INVX1 U9155 ( .A(n9190), .Y(n9191) );
  BUFX2 U9156 ( .A(fifo[305]), .Y(n9192) );
  INVX1 U9157 ( .A(n9195), .Y(n9193) );
  INVX1 U9158 ( .A(n9193), .Y(n9194) );
  BUFX2 U9159 ( .A(fifo[306]), .Y(n9195) );
  INVX1 U9160 ( .A(n9198), .Y(n9196) );
  INVX1 U9161 ( .A(n9196), .Y(n9197) );
  BUFX2 U9162 ( .A(fifo[307]), .Y(n9198) );
  INVX1 U9163 ( .A(n9201), .Y(n9199) );
  INVX1 U9164 ( .A(n9199), .Y(n9200) );
  BUFX2 U9165 ( .A(fifo[308]), .Y(n9201) );
  INVX1 U9166 ( .A(n9204), .Y(n9202) );
  INVX1 U9167 ( .A(n9202), .Y(n9203) );
  BUFX2 U9168 ( .A(fifo[309]), .Y(n9204) );
  INVX1 U9169 ( .A(n9207), .Y(n9205) );
  INVX1 U9170 ( .A(n9205), .Y(n9206) );
  BUFX2 U9171 ( .A(fifo[310]), .Y(n9207) );
  INVX1 U9172 ( .A(n9210), .Y(n9208) );
  INVX1 U9173 ( .A(n9208), .Y(n9209) );
  BUFX2 U9174 ( .A(fifo[311]), .Y(n9210) );
  INVX1 U9175 ( .A(n9213), .Y(n9211) );
  INVX1 U9176 ( .A(n9211), .Y(n9212) );
  BUFX2 U9177 ( .A(fifo[312]), .Y(n9213) );
  INVX1 U9178 ( .A(n9216), .Y(n9214) );
  INVX1 U9179 ( .A(n9214), .Y(n9215) );
  BUFX2 U9180 ( .A(fifo[313]), .Y(n9216) );
  INVX1 U9181 ( .A(n9219), .Y(n9217) );
  INVX1 U9182 ( .A(n9217), .Y(n9218) );
  BUFX2 U9183 ( .A(fifo[314]), .Y(n9219) );
  INVX1 U9184 ( .A(n9222), .Y(n9220) );
  INVX1 U9185 ( .A(n9220), .Y(n9221) );
  BUFX2 U9186 ( .A(fifo[315]), .Y(n9222) );
  INVX1 U9187 ( .A(n9225), .Y(n9223) );
  INVX1 U9188 ( .A(n9223), .Y(n9224) );
  BUFX2 U9189 ( .A(fifo[316]), .Y(n9225) );
  INVX1 U9190 ( .A(n9228), .Y(n9226) );
  INVX1 U9191 ( .A(n9226), .Y(n9227) );
  BUFX2 U9192 ( .A(fifo[317]), .Y(n9228) );
  INVX1 U9193 ( .A(n9231), .Y(n9229) );
  INVX1 U9194 ( .A(n9229), .Y(n9230) );
  BUFX2 U9195 ( .A(fifo[318]), .Y(n9231) );
  INVX1 U9196 ( .A(n9234), .Y(n9232) );
  INVX1 U9197 ( .A(n9232), .Y(n9233) );
  BUFX2 U9198 ( .A(fifo[319]), .Y(n9234) );
  INVX1 U9199 ( .A(n9237), .Y(n9235) );
  INVX1 U9200 ( .A(n9235), .Y(n9236) );
  BUFX2 U9201 ( .A(fifo[320]), .Y(n9237) );
  INVX1 U9202 ( .A(n9240), .Y(n9238) );
  INVX1 U9203 ( .A(n9238), .Y(n9239) );
  BUFX2 U9204 ( .A(fifo[321]), .Y(n9240) );
  INVX1 U9205 ( .A(n9243), .Y(n9241) );
  INVX1 U9206 ( .A(n9241), .Y(n9242) );
  BUFX2 U9207 ( .A(fifo[322]), .Y(n9243) );
  INVX1 U9208 ( .A(n9246), .Y(n9244) );
  INVX1 U9209 ( .A(n9244), .Y(n9245) );
  BUFX2 U9210 ( .A(fifo[323]), .Y(n9246) );
  INVX1 U9211 ( .A(n9249), .Y(n9247) );
  INVX1 U9212 ( .A(n9247), .Y(n9248) );
  BUFX2 U9213 ( .A(fifo[324]), .Y(n9249) );
  INVX1 U9214 ( .A(n9252), .Y(n9250) );
  INVX1 U9215 ( .A(n9250), .Y(n9251) );
  BUFX2 U9216 ( .A(fifo[325]), .Y(n9252) );
  INVX1 U9217 ( .A(n9255), .Y(n9253) );
  INVX1 U9218 ( .A(n9253), .Y(n9254) );
  BUFX2 U9219 ( .A(fifo[326]), .Y(n9255) );
  INVX1 U9220 ( .A(n9258), .Y(n9256) );
  INVX1 U9221 ( .A(n9256), .Y(n9257) );
  BUFX2 U9222 ( .A(fifo[327]), .Y(n9258) );
  INVX1 U9223 ( .A(n9261), .Y(n9259) );
  INVX1 U9224 ( .A(n9259), .Y(n9260) );
  BUFX2 U9225 ( .A(fifo[328]), .Y(n9261) );
  INVX1 U9226 ( .A(n9264), .Y(n9262) );
  INVX1 U9227 ( .A(n9262), .Y(n9263) );
  BUFX2 U9228 ( .A(fifo[329]), .Y(n9264) );
  INVX1 U9229 ( .A(n9267), .Y(n9265) );
  INVX1 U9230 ( .A(n9265), .Y(n9266) );
  BUFX2 U9231 ( .A(fifo[330]), .Y(n9267) );
  INVX1 U9232 ( .A(n9270), .Y(n9268) );
  INVX1 U9233 ( .A(n9268), .Y(n9269) );
  BUFX2 U9234 ( .A(fifo[331]), .Y(n9270) );
  INVX1 U9235 ( .A(n9273), .Y(n9271) );
  INVX1 U9236 ( .A(n9271), .Y(n9272) );
  BUFX2 U9237 ( .A(fifo[332]), .Y(n9273) );
  INVX1 U9238 ( .A(n9276), .Y(n9274) );
  INVX1 U9239 ( .A(n9274), .Y(n9275) );
  BUFX2 U9240 ( .A(fifo[333]), .Y(n9276) );
  INVX1 U9241 ( .A(n9279), .Y(n9277) );
  INVX1 U9242 ( .A(n9277), .Y(n9278) );
  BUFX2 U9243 ( .A(fifo[334]), .Y(n9279) );
  INVX1 U9244 ( .A(n9282), .Y(n9280) );
  INVX1 U9245 ( .A(n9280), .Y(n9281) );
  BUFX2 U9246 ( .A(fifo[335]), .Y(n9282) );
  INVX1 U9247 ( .A(n9285), .Y(n9283) );
  INVX1 U9248 ( .A(n9283), .Y(n9284) );
  BUFX2 U9249 ( .A(fifo[378]), .Y(n9285) );
  INVX1 U9250 ( .A(n9288), .Y(n9286) );
  INVX1 U9251 ( .A(n9286), .Y(n9287) );
  BUFX2 U9252 ( .A(fifo[379]), .Y(n9288) );
  INVX1 U9253 ( .A(n9291), .Y(n9289) );
  INVX1 U9254 ( .A(n9289), .Y(n9290) );
  BUFX2 U9255 ( .A(fifo[380]), .Y(n9291) );
  INVX1 U9256 ( .A(n9294), .Y(n9292) );
  INVX1 U9257 ( .A(n9292), .Y(n9293) );
  BUFX2 U9258 ( .A(fifo[381]), .Y(n9294) );
  INVX1 U9259 ( .A(n9297), .Y(n9295) );
  INVX1 U9260 ( .A(n9295), .Y(n9296) );
  BUFX2 U9261 ( .A(fifo[382]), .Y(n9297) );
  INVX1 U9262 ( .A(n9300), .Y(n9298) );
  INVX1 U9263 ( .A(n9298), .Y(n9299) );
  BUFX2 U9264 ( .A(fifo[383]), .Y(n9300) );
  INVX1 U9265 ( .A(n9303), .Y(n9301) );
  INVX1 U9266 ( .A(n9301), .Y(n9302) );
  BUFX2 U9267 ( .A(fifo[384]), .Y(n9303) );
  INVX1 U9268 ( .A(n9306), .Y(n9304) );
  INVX1 U9269 ( .A(n9304), .Y(n9305) );
  BUFX2 U9270 ( .A(fifo[385]), .Y(n9306) );
  INVX1 U9271 ( .A(n9309), .Y(n9307) );
  INVX1 U9272 ( .A(n9307), .Y(n9308) );
  BUFX2 U9273 ( .A(fifo[386]), .Y(n9309) );
  INVX1 U9274 ( .A(n9312), .Y(n9310) );
  INVX1 U9275 ( .A(n9310), .Y(n9311) );
  BUFX2 U9276 ( .A(fifo[387]), .Y(n9312) );
  INVX1 U9277 ( .A(n9315), .Y(n9313) );
  INVX1 U9278 ( .A(n9313), .Y(n9314) );
  BUFX2 U9279 ( .A(fifo[388]), .Y(n9315) );
  INVX1 U9280 ( .A(n9318), .Y(n9316) );
  INVX1 U9281 ( .A(n9316), .Y(n9317) );
  BUFX2 U9282 ( .A(fifo[389]), .Y(n9318) );
  INVX1 U9283 ( .A(n9321), .Y(n9319) );
  INVX1 U9284 ( .A(n9319), .Y(n9320) );
  BUFX2 U9285 ( .A(fifo[390]), .Y(n9321) );
  INVX1 U9286 ( .A(n9324), .Y(n9322) );
  INVX1 U9287 ( .A(n9322), .Y(n9323) );
  BUFX2 U9288 ( .A(fifo[391]), .Y(n9324) );
  INVX1 U9289 ( .A(n9327), .Y(n9325) );
  INVX1 U9290 ( .A(n9325), .Y(n9326) );
  BUFX2 U9291 ( .A(fifo[392]), .Y(n9327) );
  INVX1 U9292 ( .A(n9330), .Y(n9328) );
  INVX1 U9293 ( .A(n9328), .Y(n9329) );
  BUFX2 U9294 ( .A(fifo[393]), .Y(n9330) );
  INVX1 U9295 ( .A(n9333), .Y(n9331) );
  INVX1 U9296 ( .A(n9331), .Y(n9332) );
  BUFX2 U9297 ( .A(fifo[394]), .Y(n9333) );
  INVX1 U9298 ( .A(n9336), .Y(n9334) );
  INVX1 U9299 ( .A(n9334), .Y(n9335) );
  BUFX2 U9300 ( .A(fifo[395]), .Y(n9336) );
  INVX1 U9301 ( .A(n9339), .Y(n9337) );
  INVX1 U9302 ( .A(n9337), .Y(n9338) );
  BUFX2 U9303 ( .A(fifo[396]), .Y(n9339) );
  INVX1 U9304 ( .A(n9342), .Y(n9340) );
  INVX1 U9305 ( .A(n9340), .Y(n9341) );
  BUFX2 U9306 ( .A(fifo[397]), .Y(n9342) );
  INVX1 U9307 ( .A(n9345), .Y(n9343) );
  INVX1 U9308 ( .A(n9343), .Y(n9344) );
  BUFX2 U9309 ( .A(fifo[398]), .Y(n9345) );
  INVX1 U9310 ( .A(n9348), .Y(n9346) );
  INVX1 U9311 ( .A(n9346), .Y(n9347) );
  BUFX2 U9312 ( .A(fifo[399]), .Y(n9348) );
  INVX1 U9313 ( .A(n9351), .Y(n9349) );
  INVX1 U9314 ( .A(n9349), .Y(n9350) );
  BUFX2 U9315 ( .A(fifo[400]), .Y(n9351) );
  INVX1 U9316 ( .A(n9354), .Y(n9352) );
  INVX1 U9317 ( .A(n9352), .Y(n9353) );
  BUFX2 U9318 ( .A(fifo[401]), .Y(n9354) );
  INVX1 U9319 ( .A(n9357), .Y(n9355) );
  INVX1 U9320 ( .A(n9355), .Y(n9356) );
  BUFX2 U9321 ( .A(fifo[402]), .Y(n9357) );
  INVX1 U9322 ( .A(n9360), .Y(n9358) );
  INVX1 U9323 ( .A(n9358), .Y(n9359) );
  BUFX2 U9324 ( .A(fifo[403]), .Y(n9360) );
  INVX1 U9325 ( .A(n9363), .Y(n9361) );
  INVX1 U9326 ( .A(n9361), .Y(n9362) );
  BUFX2 U9327 ( .A(fifo[404]), .Y(n9363) );
  INVX1 U9328 ( .A(n9366), .Y(n9364) );
  INVX1 U9329 ( .A(n9364), .Y(n9365) );
  BUFX2 U9330 ( .A(fifo[405]), .Y(n9366) );
  INVX1 U9331 ( .A(n9369), .Y(n9367) );
  INVX1 U9332 ( .A(n9367), .Y(n9368) );
  BUFX2 U9333 ( .A(fifo[406]), .Y(n9369) );
  INVX1 U9334 ( .A(n9372), .Y(n9370) );
  INVX1 U9335 ( .A(n9370), .Y(n9371) );
  BUFX2 U9336 ( .A(fifo[407]), .Y(n9372) );
  INVX1 U9337 ( .A(n9375), .Y(n9373) );
  INVX1 U9338 ( .A(n9373), .Y(n9374) );
  BUFX2 U9339 ( .A(fifo[408]), .Y(n9375) );
  INVX1 U9340 ( .A(n9378), .Y(n9376) );
  INVX1 U9341 ( .A(n9376), .Y(n9377) );
  BUFX2 U9342 ( .A(fifo[409]), .Y(n9378) );
  INVX1 U9343 ( .A(n9381), .Y(n9379) );
  INVX1 U9344 ( .A(n9379), .Y(n9380) );
  BUFX2 U9345 ( .A(fifo[410]), .Y(n9381) );
  INVX1 U9346 ( .A(n9384), .Y(n9382) );
  INVX1 U9347 ( .A(n9382), .Y(n9383) );
  BUFX2 U9348 ( .A(fifo[411]), .Y(n9384) );
  INVX1 U9349 ( .A(n9387), .Y(n9385) );
  INVX1 U9350 ( .A(n9385), .Y(n9386) );
  BUFX2 U9351 ( .A(fifo[412]), .Y(n9387) );
  INVX1 U9352 ( .A(n9390), .Y(n9388) );
  INVX1 U9353 ( .A(n9388), .Y(n9389) );
  BUFX2 U9354 ( .A(fifo[413]), .Y(n9390) );
  INVX1 U9355 ( .A(n9393), .Y(n9391) );
  INVX1 U9356 ( .A(n9391), .Y(n9392) );
  BUFX2 U9357 ( .A(fifo[414]), .Y(n9393) );
  INVX1 U9358 ( .A(n9396), .Y(n9394) );
  INVX1 U9359 ( .A(n9394), .Y(n9395) );
  BUFX2 U9360 ( .A(fifo[415]), .Y(n9396) );
  INVX1 U9361 ( .A(n9399), .Y(n9397) );
  INVX1 U9362 ( .A(n9397), .Y(n9398) );
  BUFX2 U9363 ( .A(fifo[416]), .Y(n9399) );
  INVX1 U9364 ( .A(n9402), .Y(n9400) );
  INVX1 U9365 ( .A(n9400), .Y(n9401) );
  BUFX2 U9366 ( .A(fifo[417]), .Y(n9402) );
  INVX1 U9367 ( .A(n9405), .Y(n9403) );
  INVX1 U9368 ( .A(n9403), .Y(n9404) );
  BUFX2 U9369 ( .A(fifo[418]), .Y(n9405) );
  INVX1 U9370 ( .A(n9408), .Y(n9406) );
  INVX1 U9371 ( .A(n9406), .Y(n9407) );
  BUFX2 U9372 ( .A(fifo[419]), .Y(n9408) );
  INVX1 U9373 ( .A(n9411), .Y(n9409) );
  INVX1 U9374 ( .A(n9409), .Y(n9410) );
  BUFX2 U9375 ( .A(fifo[462]), .Y(n9411) );
  INVX1 U9376 ( .A(n9414), .Y(n9412) );
  INVX1 U9377 ( .A(n9412), .Y(n9413) );
  BUFX2 U9378 ( .A(fifo[463]), .Y(n9414) );
  INVX1 U9379 ( .A(n9417), .Y(n9415) );
  INVX1 U9380 ( .A(n9415), .Y(n9416) );
  BUFX2 U9381 ( .A(fifo[464]), .Y(n9417) );
  INVX1 U9382 ( .A(n9420), .Y(n9418) );
  INVX1 U9383 ( .A(n9418), .Y(n9419) );
  BUFX2 U9384 ( .A(fifo[465]), .Y(n9420) );
  INVX1 U9385 ( .A(n9423), .Y(n9421) );
  INVX1 U9386 ( .A(n9421), .Y(n9422) );
  BUFX2 U9387 ( .A(fifo[466]), .Y(n9423) );
  INVX1 U9388 ( .A(n9426), .Y(n9424) );
  INVX1 U9389 ( .A(n9424), .Y(n9425) );
  BUFX2 U9390 ( .A(fifo[467]), .Y(n9426) );
  INVX1 U9391 ( .A(n9429), .Y(n9427) );
  INVX1 U9392 ( .A(n9427), .Y(n9428) );
  BUFX2 U9393 ( .A(fifo[468]), .Y(n9429) );
  INVX1 U9394 ( .A(n9432), .Y(n9430) );
  INVX1 U9395 ( .A(n9430), .Y(n9431) );
  BUFX2 U9396 ( .A(fifo[469]), .Y(n9432) );
  INVX1 U9397 ( .A(n9435), .Y(n9433) );
  INVX1 U9398 ( .A(n9433), .Y(n9434) );
  BUFX2 U9399 ( .A(fifo[470]), .Y(n9435) );
  INVX1 U9400 ( .A(n9438), .Y(n9436) );
  INVX1 U9401 ( .A(n9436), .Y(n9437) );
  BUFX2 U9402 ( .A(fifo[471]), .Y(n9438) );
  INVX1 U9403 ( .A(n9441), .Y(n9439) );
  INVX1 U9404 ( .A(n9439), .Y(n9440) );
  BUFX2 U9405 ( .A(fifo[472]), .Y(n9441) );
  INVX1 U9406 ( .A(n9444), .Y(n9442) );
  INVX1 U9407 ( .A(n9442), .Y(n9443) );
  BUFX2 U9408 ( .A(fifo[473]), .Y(n9444) );
  INVX1 U9409 ( .A(n9447), .Y(n9445) );
  INVX1 U9410 ( .A(n9445), .Y(n9446) );
  BUFX2 U9411 ( .A(fifo[474]), .Y(n9447) );
  INVX1 U9412 ( .A(n9450), .Y(n9448) );
  INVX1 U9413 ( .A(n9448), .Y(n9449) );
  BUFX2 U9414 ( .A(fifo[475]), .Y(n9450) );
  INVX1 U9415 ( .A(n9453), .Y(n9451) );
  INVX1 U9416 ( .A(n9451), .Y(n9452) );
  BUFX2 U9417 ( .A(fifo[476]), .Y(n9453) );
  INVX1 U9418 ( .A(n9456), .Y(n9454) );
  INVX1 U9419 ( .A(n9454), .Y(n9455) );
  BUFX2 U9420 ( .A(fifo[477]), .Y(n9456) );
  INVX1 U9421 ( .A(n9459), .Y(n9457) );
  INVX1 U9422 ( .A(n9457), .Y(n9458) );
  BUFX2 U9423 ( .A(fifo[478]), .Y(n9459) );
  INVX1 U9424 ( .A(n9462), .Y(n9460) );
  INVX1 U9425 ( .A(n9460), .Y(n9461) );
  BUFX2 U9426 ( .A(fifo[479]), .Y(n9462) );
  INVX1 U9427 ( .A(n9465), .Y(n9463) );
  INVX1 U9428 ( .A(n9463), .Y(n9464) );
  BUFX2 U9429 ( .A(fifo[480]), .Y(n9465) );
  INVX1 U9430 ( .A(n9468), .Y(n9466) );
  INVX1 U9431 ( .A(n9466), .Y(n9467) );
  BUFX2 U9432 ( .A(fifo[481]), .Y(n9468) );
  INVX1 U9433 ( .A(n9471), .Y(n9469) );
  INVX1 U9434 ( .A(n9469), .Y(n9470) );
  BUFX2 U9435 ( .A(fifo[482]), .Y(n9471) );
  INVX1 U9436 ( .A(n9474), .Y(n9472) );
  INVX1 U9437 ( .A(n9472), .Y(n9473) );
  BUFX2 U9438 ( .A(fifo[483]), .Y(n9474) );
  INVX1 U9439 ( .A(n9477), .Y(n9475) );
  INVX1 U9440 ( .A(n9475), .Y(n9476) );
  BUFX2 U9441 ( .A(fifo[484]), .Y(n9477) );
  INVX1 U9442 ( .A(n9480), .Y(n9478) );
  INVX1 U9443 ( .A(n9478), .Y(n9479) );
  BUFX2 U9444 ( .A(fifo[485]), .Y(n9480) );
  INVX1 U9445 ( .A(n9483), .Y(n9481) );
  INVX1 U9446 ( .A(n9481), .Y(n9482) );
  BUFX2 U9447 ( .A(fifo[486]), .Y(n9483) );
  INVX1 U9448 ( .A(n9486), .Y(n9484) );
  INVX1 U9449 ( .A(n9484), .Y(n9485) );
  BUFX2 U9450 ( .A(fifo[487]), .Y(n9486) );
  INVX1 U9451 ( .A(n9489), .Y(n9487) );
  INVX1 U9452 ( .A(n9487), .Y(n9488) );
  BUFX2 U9453 ( .A(fifo[488]), .Y(n9489) );
  INVX1 U9454 ( .A(n9492), .Y(n9490) );
  INVX1 U9455 ( .A(n9490), .Y(n9491) );
  BUFX2 U9456 ( .A(fifo[489]), .Y(n9492) );
  INVX1 U9457 ( .A(n9495), .Y(n9493) );
  INVX1 U9458 ( .A(n9493), .Y(n9494) );
  BUFX2 U9459 ( .A(fifo[490]), .Y(n9495) );
  INVX1 U9460 ( .A(n9498), .Y(n9496) );
  INVX1 U9461 ( .A(n9496), .Y(n9497) );
  BUFX2 U9462 ( .A(fifo[491]), .Y(n9498) );
  INVX1 U9463 ( .A(n9501), .Y(n9499) );
  INVX1 U9464 ( .A(n9499), .Y(n9500) );
  BUFX2 U9465 ( .A(fifo[492]), .Y(n9501) );
  INVX1 U9466 ( .A(n9504), .Y(n9502) );
  INVX1 U9467 ( .A(n9502), .Y(n9503) );
  BUFX2 U9468 ( .A(fifo[493]), .Y(n9504) );
  INVX1 U9469 ( .A(n9507), .Y(n9505) );
  INVX1 U9470 ( .A(n9505), .Y(n9506) );
  BUFX2 U9471 ( .A(fifo[494]), .Y(n9507) );
  INVX1 U9472 ( .A(n9510), .Y(n9508) );
  INVX1 U9473 ( .A(n9508), .Y(n9509) );
  BUFX2 U9474 ( .A(fifo[495]), .Y(n9510) );
  INVX1 U9475 ( .A(n9513), .Y(n9511) );
  INVX1 U9476 ( .A(n9511), .Y(n9512) );
  BUFX2 U9477 ( .A(fifo[496]), .Y(n9513) );
  INVX1 U9478 ( .A(n9516), .Y(n9514) );
  INVX1 U9479 ( .A(n9514), .Y(n9515) );
  BUFX2 U9480 ( .A(fifo[497]), .Y(n9516) );
  INVX1 U9481 ( .A(n9519), .Y(n9517) );
  INVX1 U9482 ( .A(n9517), .Y(n9518) );
  BUFX2 U9483 ( .A(fifo[498]), .Y(n9519) );
  INVX1 U9484 ( .A(n9522), .Y(n9520) );
  INVX1 U9485 ( .A(n9520), .Y(n9521) );
  BUFX2 U9486 ( .A(fifo[499]), .Y(n9522) );
  INVX1 U9487 ( .A(n9525), .Y(n9523) );
  INVX1 U9488 ( .A(n9523), .Y(n9524) );
  BUFX2 U9489 ( .A(fifo[500]), .Y(n9525) );
  INVX1 U9490 ( .A(n9528), .Y(n9526) );
  INVX1 U9491 ( .A(n9526), .Y(n9527) );
  BUFX2 U9492 ( .A(fifo[501]), .Y(n9528) );
  INVX1 U9493 ( .A(n9531), .Y(n9529) );
  INVX1 U9494 ( .A(n9529), .Y(n9530) );
  BUFX2 U9495 ( .A(fifo[502]), .Y(n9531) );
  INVX1 U9496 ( .A(n9534), .Y(n9532) );
  INVX1 U9497 ( .A(n9532), .Y(n9533) );
  BUFX2 U9498 ( .A(fifo[503]), .Y(n9534) );
  INVX1 U9499 ( .A(n9537), .Y(n9535) );
  INVX1 U9500 ( .A(n9535), .Y(n9536) );
  BUFX2 U9501 ( .A(fifo[546]), .Y(n9537) );
  INVX1 U9502 ( .A(n9540), .Y(n9538) );
  INVX1 U9503 ( .A(n9538), .Y(n9539) );
  BUFX2 U9504 ( .A(fifo[547]), .Y(n9540) );
  INVX1 U9505 ( .A(n9543), .Y(n9541) );
  INVX1 U9506 ( .A(n9541), .Y(n9542) );
  BUFX2 U9507 ( .A(fifo[548]), .Y(n9543) );
  INVX1 U9508 ( .A(n9546), .Y(n9544) );
  INVX1 U9509 ( .A(n9544), .Y(n9545) );
  BUFX2 U9510 ( .A(fifo[549]), .Y(n9546) );
  INVX1 U9511 ( .A(n9549), .Y(n9547) );
  INVX1 U9512 ( .A(n9547), .Y(n9548) );
  BUFX2 U9513 ( .A(fifo[550]), .Y(n9549) );
  INVX1 U9514 ( .A(n9552), .Y(n9550) );
  INVX1 U9515 ( .A(n9550), .Y(n9551) );
  BUFX2 U9516 ( .A(fifo[551]), .Y(n9552) );
  INVX1 U9517 ( .A(n9555), .Y(n9553) );
  INVX1 U9518 ( .A(n9553), .Y(n9554) );
  BUFX2 U9519 ( .A(fifo[552]), .Y(n9555) );
  INVX1 U9520 ( .A(n9558), .Y(n9556) );
  INVX1 U9521 ( .A(n9556), .Y(n9557) );
  BUFX2 U9522 ( .A(fifo[553]), .Y(n9558) );
  INVX1 U9523 ( .A(n9561), .Y(n9559) );
  INVX1 U9524 ( .A(n9559), .Y(n9560) );
  BUFX2 U9525 ( .A(fifo[554]), .Y(n9561) );
  INVX1 U9526 ( .A(n9564), .Y(n9562) );
  INVX1 U9527 ( .A(n9562), .Y(n9563) );
  BUFX2 U9528 ( .A(fifo[555]), .Y(n9564) );
  INVX1 U9529 ( .A(n9567), .Y(n9565) );
  INVX1 U9530 ( .A(n9565), .Y(n9566) );
  BUFX2 U9531 ( .A(fifo[556]), .Y(n9567) );
  INVX1 U9532 ( .A(n9570), .Y(n9568) );
  INVX1 U9533 ( .A(n9568), .Y(n9569) );
  BUFX2 U9534 ( .A(fifo[557]), .Y(n9570) );
  INVX1 U9535 ( .A(n9573), .Y(n9571) );
  INVX1 U9536 ( .A(n9571), .Y(n9572) );
  BUFX2 U9537 ( .A(fifo[558]), .Y(n9573) );
  INVX1 U9538 ( .A(n9576), .Y(n9574) );
  INVX1 U9539 ( .A(n9574), .Y(n9575) );
  BUFX2 U9540 ( .A(fifo[559]), .Y(n9576) );
  INVX1 U9541 ( .A(n9579), .Y(n9577) );
  INVX1 U9542 ( .A(n9577), .Y(n9578) );
  BUFX2 U9543 ( .A(fifo[560]), .Y(n9579) );
  INVX1 U9544 ( .A(n9582), .Y(n9580) );
  INVX1 U9545 ( .A(n9580), .Y(n9581) );
  BUFX2 U9546 ( .A(fifo[561]), .Y(n9582) );
  INVX1 U9547 ( .A(n9585), .Y(n9583) );
  INVX1 U9548 ( .A(n9583), .Y(n9584) );
  BUFX2 U9549 ( .A(fifo[562]), .Y(n9585) );
  INVX1 U9550 ( .A(n9588), .Y(n9586) );
  INVX1 U9551 ( .A(n9586), .Y(n9587) );
  BUFX2 U9552 ( .A(fifo[563]), .Y(n9588) );
  INVX1 U9553 ( .A(n9591), .Y(n9589) );
  INVX1 U9554 ( .A(n9589), .Y(n9590) );
  BUFX2 U9555 ( .A(fifo[564]), .Y(n9591) );
  INVX1 U9556 ( .A(n9594), .Y(n9592) );
  INVX1 U9557 ( .A(n9592), .Y(n9593) );
  BUFX2 U9558 ( .A(fifo[565]), .Y(n9594) );
  INVX1 U9559 ( .A(n9597), .Y(n9595) );
  INVX1 U9560 ( .A(n9595), .Y(n9596) );
  BUFX2 U9561 ( .A(fifo[566]), .Y(n9597) );
  INVX1 U9562 ( .A(n9600), .Y(n9598) );
  INVX1 U9563 ( .A(n9598), .Y(n9599) );
  BUFX2 U9564 ( .A(fifo[567]), .Y(n9600) );
  INVX1 U9565 ( .A(n9603), .Y(n9601) );
  INVX1 U9566 ( .A(n9601), .Y(n9602) );
  BUFX2 U9567 ( .A(fifo[568]), .Y(n9603) );
  INVX1 U9568 ( .A(n9606), .Y(n9604) );
  INVX1 U9569 ( .A(n9604), .Y(n9605) );
  BUFX2 U9570 ( .A(fifo[569]), .Y(n9606) );
  INVX1 U9571 ( .A(n9609), .Y(n9607) );
  INVX1 U9572 ( .A(n9607), .Y(n9608) );
  BUFX2 U9573 ( .A(fifo[570]), .Y(n9609) );
  INVX1 U9574 ( .A(n9612), .Y(n9610) );
  INVX1 U9575 ( .A(n9610), .Y(n9611) );
  BUFX2 U9576 ( .A(fifo[571]), .Y(n9612) );
  INVX1 U9577 ( .A(n9615), .Y(n9613) );
  INVX1 U9578 ( .A(n9613), .Y(n9614) );
  BUFX2 U9579 ( .A(fifo[572]), .Y(n9615) );
  INVX1 U9580 ( .A(n9618), .Y(n9616) );
  INVX1 U9581 ( .A(n9616), .Y(n9617) );
  BUFX2 U9582 ( .A(fifo[573]), .Y(n9618) );
  INVX1 U9583 ( .A(n9621), .Y(n9619) );
  INVX1 U9584 ( .A(n9619), .Y(n9620) );
  BUFX2 U9585 ( .A(fifo[574]), .Y(n9621) );
  INVX1 U9586 ( .A(n9624), .Y(n9622) );
  INVX1 U9587 ( .A(n9622), .Y(n9623) );
  BUFX2 U9588 ( .A(fifo[575]), .Y(n9624) );
  INVX1 U9589 ( .A(n9627), .Y(n9625) );
  INVX1 U9590 ( .A(n9625), .Y(n9626) );
  BUFX2 U9591 ( .A(fifo[576]), .Y(n9627) );
  INVX1 U9592 ( .A(n9630), .Y(n9628) );
  INVX1 U9593 ( .A(n9628), .Y(n9629) );
  BUFX2 U9594 ( .A(fifo[577]), .Y(n9630) );
  INVX1 U9595 ( .A(n9633), .Y(n9631) );
  INVX1 U9596 ( .A(n9631), .Y(n9632) );
  BUFX2 U9597 ( .A(fifo[578]), .Y(n9633) );
  INVX1 U9598 ( .A(n9636), .Y(n9634) );
  INVX1 U9599 ( .A(n9634), .Y(n9635) );
  BUFX2 U9600 ( .A(fifo[579]), .Y(n9636) );
  INVX1 U9601 ( .A(n9639), .Y(n9637) );
  INVX1 U9602 ( .A(n9637), .Y(n9638) );
  BUFX2 U9603 ( .A(fifo[580]), .Y(n9639) );
  INVX1 U9604 ( .A(n9642), .Y(n9640) );
  INVX1 U9605 ( .A(n9640), .Y(n9641) );
  BUFX2 U9606 ( .A(fifo[581]), .Y(n9642) );
  INVX1 U9607 ( .A(n9645), .Y(n9643) );
  INVX1 U9608 ( .A(n9643), .Y(n9644) );
  BUFX2 U9609 ( .A(fifo[582]), .Y(n9645) );
  INVX1 U9610 ( .A(n9648), .Y(n9646) );
  INVX1 U9611 ( .A(n9646), .Y(n9647) );
  BUFX2 U9612 ( .A(fifo[583]), .Y(n9648) );
  INVX1 U9613 ( .A(n9651), .Y(n9649) );
  INVX1 U9614 ( .A(n9649), .Y(n9650) );
  BUFX2 U9615 ( .A(fifo[584]), .Y(n9651) );
  INVX1 U9616 ( .A(n9654), .Y(n9652) );
  INVX1 U9617 ( .A(n9652), .Y(n9653) );
  BUFX2 U9618 ( .A(fifo[585]), .Y(n9654) );
  INVX1 U9619 ( .A(n9657), .Y(n9655) );
  INVX1 U9620 ( .A(n9655), .Y(n9656) );
  BUFX2 U9621 ( .A(fifo[586]), .Y(n9657) );
  INVX1 U9622 ( .A(n9660), .Y(n9658) );
  INVX1 U9623 ( .A(n9658), .Y(n9659) );
  BUFX2 U9624 ( .A(fifo[587]), .Y(n9660) );
  INVX1 U9625 ( .A(n9663), .Y(n9661) );
  INVX1 U9626 ( .A(n9661), .Y(n9662) );
  BUFX2 U9627 ( .A(fifo[630]), .Y(n9663) );
  INVX1 U9628 ( .A(n9666), .Y(n9664) );
  INVX1 U9629 ( .A(n9664), .Y(n9665) );
  BUFX2 U9630 ( .A(fifo[631]), .Y(n9666) );
  INVX1 U9631 ( .A(n9669), .Y(n9667) );
  INVX1 U9632 ( .A(n9667), .Y(n9668) );
  BUFX2 U9633 ( .A(fifo[632]), .Y(n9669) );
  INVX1 U9634 ( .A(n9672), .Y(n9670) );
  INVX1 U9635 ( .A(n9670), .Y(n9671) );
  BUFX2 U9636 ( .A(fifo[633]), .Y(n9672) );
  INVX1 U9637 ( .A(n9675), .Y(n9673) );
  INVX1 U9638 ( .A(n9673), .Y(n9674) );
  BUFX2 U9639 ( .A(fifo[634]), .Y(n9675) );
  INVX1 U9640 ( .A(n9678), .Y(n9676) );
  INVX1 U9641 ( .A(n9676), .Y(n9677) );
  BUFX2 U9642 ( .A(fifo[635]), .Y(n9678) );
  INVX1 U9643 ( .A(n9681), .Y(n9679) );
  INVX1 U9644 ( .A(n9679), .Y(n9680) );
  BUFX2 U9645 ( .A(fifo[636]), .Y(n9681) );
  INVX1 U9646 ( .A(n9684), .Y(n9682) );
  INVX1 U9647 ( .A(n9682), .Y(n9683) );
  BUFX2 U9648 ( .A(fifo[637]), .Y(n9684) );
  INVX1 U9649 ( .A(n9687), .Y(n9685) );
  INVX1 U9650 ( .A(n9685), .Y(n9686) );
  BUFX2 U9651 ( .A(fifo[638]), .Y(n9687) );
  INVX1 U9652 ( .A(n9690), .Y(n9688) );
  INVX1 U9653 ( .A(n9688), .Y(n9689) );
  BUFX2 U9654 ( .A(fifo[639]), .Y(n9690) );
  INVX1 U9655 ( .A(n9693), .Y(n9691) );
  INVX1 U9656 ( .A(n9691), .Y(n9692) );
  BUFX2 U9657 ( .A(fifo[640]), .Y(n9693) );
  INVX1 U9658 ( .A(n9696), .Y(n9694) );
  INVX1 U9659 ( .A(n9694), .Y(n9695) );
  BUFX2 U9660 ( .A(fifo[641]), .Y(n9696) );
  INVX1 U9661 ( .A(n9699), .Y(n9697) );
  INVX1 U9662 ( .A(n9697), .Y(n9698) );
  BUFX2 U9663 ( .A(fifo[642]), .Y(n9699) );
  INVX1 U9664 ( .A(n9702), .Y(n9700) );
  INVX1 U9665 ( .A(n9700), .Y(n9701) );
  BUFX2 U9666 ( .A(fifo[643]), .Y(n9702) );
  INVX1 U9667 ( .A(n9705), .Y(n9703) );
  INVX1 U9668 ( .A(n9703), .Y(n9704) );
  BUFX2 U9669 ( .A(fifo[644]), .Y(n9705) );
  INVX1 U9670 ( .A(n9708), .Y(n9706) );
  INVX1 U9671 ( .A(n9706), .Y(n9707) );
  BUFX2 U9672 ( .A(fifo[645]), .Y(n9708) );
  INVX1 U9673 ( .A(n9711), .Y(n9709) );
  INVX1 U9674 ( .A(n9709), .Y(n9710) );
  BUFX2 U9675 ( .A(fifo[646]), .Y(n9711) );
  INVX1 U9676 ( .A(n9714), .Y(n9712) );
  INVX1 U9677 ( .A(n9712), .Y(n9713) );
  BUFX2 U9678 ( .A(fifo[647]), .Y(n9714) );
  INVX1 U9679 ( .A(n9717), .Y(n9715) );
  INVX1 U9680 ( .A(n9715), .Y(n9716) );
  BUFX2 U9681 ( .A(fifo[648]), .Y(n9717) );
  INVX1 U9682 ( .A(n9720), .Y(n9718) );
  INVX1 U9683 ( .A(n9718), .Y(n9719) );
  BUFX2 U9684 ( .A(fifo[649]), .Y(n9720) );
  INVX1 U9685 ( .A(n9723), .Y(n9721) );
  INVX1 U9686 ( .A(n9721), .Y(n9722) );
  BUFX2 U9687 ( .A(fifo[650]), .Y(n9723) );
  INVX1 U9688 ( .A(n9726), .Y(n9724) );
  INVX1 U9689 ( .A(n9724), .Y(n9725) );
  BUFX2 U9690 ( .A(fifo[651]), .Y(n9726) );
  INVX1 U9691 ( .A(n9729), .Y(n9727) );
  INVX1 U9692 ( .A(n9727), .Y(n9728) );
  BUFX2 U9693 ( .A(fifo[652]), .Y(n9729) );
  INVX1 U9694 ( .A(n9732), .Y(n9730) );
  INVX1 U9695 ( .A(n9730), .Y(n9731) );
  BUFX2 U9696 ( .A(fifo[653]), .Y(n9732) );
  INVX1 U9697 ( .A(n9735), .Y(n9733) );
  INVX1 U9698 ( .A(n9733), .Y(n9734) );
  BUFX2 U9699 ( .A(fifo[654]), .Y(n9735) );
  INVX1 U9700 ( .A(n9738), .Y(n9736) );
  INVX1 U9701 ( .A(n9736), .Y(n9737) );
  BUFX2 U9702 ( .A(fifo[655]), .Y(n9738) );
  INVX1 U9703 ( .A(n9741), .Y(n9739) );
  INVX1 U9704 ( .A(n9739), .Y(n9740) );
  BUFX2 U9705 ( .A(fifo[656]), .Y(n9741) );
  INVX1 U9706 ( .A(n9744), .Y(n9742) );
  INVX1 U9707 ( .A(n9742), .Y(n9743) );
  BUFX2 U9708 ( .A(fifo[657]), .Y(n9744) );
  INVX1 U9709 ( .A(n9747), .Y(n9745) );
  INVX1 U9710 ( .A(n9745), .Y(n9746) );
  BUFX2 U9711 ( .A(fifo[658]), .Y(n9747) );
  INVX1 U9712 ( .A(n9750), .Y(n9748) );
  INVX1 U9713 ( .A(n9748), .Y(n9749) );
  BUFX2 U9714 ( .A(fifo[659]), .Y(n9750) );
  INVX1 U9715 ( .A(n9753), .Y(n9751) );
  INVX1 U9716 ( .A(n9751), .Y(n9752) );
  BUFX2 U9717 ( .A(fifo[660]), .Y(n9753) );
  INVX1 U9718 ( .A(n9756), .Y(n9754) );
  INVX1 U9719 ( .A(n9754), .Y(n9755) );
  BUFX2 U9720 ( .A(fifo[661]), .Y(n9756) );
  INVX1 U9721 ( .A(n9759), .Y(n9757) );
  INVX1 U9722 ( .A(n9757), .Y(n9758) );
  BUFX2 U9723 ( .A(fifo[662]), .Y(n9759) );
  INVX1 U9724 ( .A(n9762), .Y(n9760) );
  INVX1 U9725 ( .A(n9760), .Y(n9761) );
  BUFX2 U9726 ( .A(fifo[663]), .Y(n9762) );
  INVX1 U9727 ( .A(n9765), .Y(n9763) );
  INVX1 U9728 ( .A(n9763), .Y(n9764) );
  BUFX2 U9729 ( .A(fifo[664]), .Y(n9765) );
  INVX1 U9730 ( .A(n9768), .Y(n9766) );
  INVX1 U9731 ( .A(n9766), .Y(n9767) );
  BUFX2 U9732 ( .A(fifo[665]), .Y(n9768) );
  INVX1 U9733 ( .A(n9771), .Y(n9769) );
  INVX1 U9734 ( .A(n9769), .Y(n9770) );
  BUFX2 U9735 ( .A(fifo[666]), .Y(n9771) );
  INVX1 U9736 ( .A(n9774), .Y(n9772) );
  INVX1 U9737 ( .A(n9772), .Y(n9773) );
  BUFX2 U9738 ( .A(fifo[667]), .Y(n9774) );
  INVX1 U9739 ( .A(n9777), .Y(n9775) );
  INVX1 U9740 ( .A(n9775), .Y(n9776) );
  BUFX2 U9741 ( .A(fifo[668]), .Y(n9777) );
  INVX1 U9742 ( .A(n9780), .Y(n9778) );
  INVX1 U9743 ( .A(n9778), .Y(n9779) );
  BUFX2 U9744 ( .A(fifo[669]), .Y(n9780) );
  INVX1 U9745 ( .A(n9783), .Y(n9781) );
  INVX1 U9746 ( .A(n9781), .Y(n9782) );
  BUFX2 U9747 ( .A(fifo[670]), .Y(n9783) );
  INVX1 U9748 ( .A(n9786), .Y(n9784) );
  INVX1 U9749 ( .A(n9784), .Y(n9785) );
  BUFX2 U9750 ( .A(fifo[671]), .Y(n9786) );
  INVX1 U9751 ( .A(n9789), .Y(n9787) );
  INVX1 U9752 ( .A(n9787), .Y(n9788) );
  BUFX2 U9753 ( .A(fifo[714]), .Y(n9789) );
  INVX1 U9754 ( .A(n9792), .Y(n9790) );
  INVX1 U9755 ( .A(n9790), .Y(n9791) );
  BUFX2 U9756 ( .A(fifo[715]), .Y(n9792) );
  INVX1 U9757 ( .A(n9795), .Y(n9793) );
  INVX1 U9758 ( .A(n9793), .Y(n9794) );
  BUFX2 U9759 ( .A(fifo[716]), .Y(n9795) );
  INVX1 U9760 ( .A(n9798), .Y(n9796) );
  INVX1 U9761 ( .A(n9796), .Y(n9797) );
  BUFX2 U9762 ( .A(fifo[717]), .Y(n9798) );
  INVX1 U9763 ( .A(n9801), .Y(n9799) );
  INVX1 U9764 ( .A(n9799), .Y(n9800) );
  BUFX2 U9765 ( .A(fifo[718]), .Y(n9801) );
  INVX1 U9766 ( .A(n9804), .Y(n9802) );
  INVX1 U9767 ( .A(n9802), .Y(n9803) );
  BUFX2 U9768 ( .A(fifo[719]), .Y(n9804) );
  INVX1 U9769 ( .A(n9807), .Y(n9805) );
  INVX1 U9770 ( .A(n9805), .Y(n9806) );
  BUFX2 U9771 ( .A(fifo[720]), .Y(n9807) );
  INVX1 U9772 ( .A(n9810), .Y(n9808) );
  INVX1 U9773 ( .A(n9808), .Y(n9809) );
  BUFX2 U9774 ( .A(fifo[721]), .Y(n9810) );
  INVX1 U9775 ( .A(n9813), .Y(n9811) );
  INVX1 U9776 ( .A(n9811), .Y(n9812) );
  BUFX2 U9777 ( .A(fifo[722]), .Y(n9813) );
  INVX1 U9778 ( .A(n9816), .Y(n9814) );
  INVX1 U9779 ( .A(n9814), .Y(n9815) );
  BUFX2 U9780 ( .A(fifo[723]), .Y(n9816) );
  INVX1 U9781 ( .A(n9819), .Y(n9817) );
  INVX1 U9782 ( .A(n9817), .Y(n9818) );
  BUFX2 U9783 ( .A(fifo[724]), .Y(n9819) );
  INVX1 U9784 ( .A(n9822), .Y(n9820) );
  INVX1 U9785 ( .A(n9820), .Y(n9821) );
  BUFX2 U9786 ( .A(fifo[725]), .Y(n9822) );
  INVX1 U9787 ( .A(n9825), .Y(n9823) );
  INVX1 U9788 ( .A(n9823), .Y(n9824) );
  BUFX2 U9789 ( .A(fifo[726]), .Y(n9825) );
  INVX1 U9790 ( .A(n9828), .Y(n9826) );
  INVX1 U9791 ( .A(n9826), .Y(n9827) );
  BUFX2 U9792 ( .A(fifo[727]), .Y(n9828) );
  INVX1 U9793 ( .A(n9831), .Y(n9829) );
  INVX1 U9794 ( .A(n9829), .Y(n9830) );
  BUFX2 U9795 ( .A(fifo[728]), .Y(n9831) );
  INVX1 U9796 ( .A(n9834), .Y(n9832) );
  INVX1 U9797 ( .A(n9832), .Y(n9833) );
  BUFX2 U9798 ( .A(fifo[729]), .Y(n9834) );
  INVX1 U9799 ( .A(n9837), .Y(n9835) );
  INVX1 U9800 ( .A(n9835), .Y(n9836) );
  BUFX2 U9801 ( .A(fifo[730]), .Y(n9837) );
  INVX1 U9802 ( .A(n9840), .Y(n9838) );
  INVX1 U9803 ( .A(n9838), .Y(n9839) );
  BUFX2 U9804 ( .A(fifo[731]), .Y(n9840) );
  INVX1 U9805 ( .A(n9843), .Y(n9841) );
  INVX1 U9806 ( .A(n9841), .Y(n9842) );
  BUFX2 U9807 ( .A(fifo[732]), .Y(n9843) );
  INVX1 U9808 ( .A(n9846), .Y(n9844) );
  INVX1 U9809 ( .A(n9844), .Y(n9845) );
  BUFX2 U9810 ( .A(fifo[733]), .Y(n9846) );
  INVX1 U9811 ( .A(n9849), .Y(n9847) );
  INVX1 U9812 ( .A(n9847), .Y(n9848) );
  BUFX2 U9813 ( .A(fifo[734]), .Y(n9849) );
  INVX1 U9814 ( .A(n9852), .Y(n9850) );
  INVX1 U9815 ( .A(n9850), .Y(n9851) );
  BUFX2 U9816 ( .A(fifo[735]), .Y(n9852) );
  INVX1 U9817 ( .A(n9855), .Y(n9853) );
  INVX1 U9818 ( .A(n9853), .Y(n9854) );
  BUFX2 U9819 ( .A(fifo[736]), .Y(n9855) );
  INVX1 U9820 ( .A(n9858), .Y(n9856) );
  INVX1 U9821 ( .A(n9856), .Y(n9857) );
  BUFX2 U9822 ( .A(fifo[737]), .Y(n9858) );
  INVX1 U9823 ( .A(n9861), .Y(n9859) );
  INVX1 U9824 ( .A(n9859), .Y(n9860) );
  BUFX2 U9825 ( .A(fifo[738]), .Y(n9861) );
  INVX1 U9826 ( .A(n9864), .Y(n9862) );
  INVX1 U9827 ( .A(n9862), .Y(n9863) );
  BUFX2 U9828 ( .A(fifo[739]), .Y(n9864) );
  INVX1 U9829 ( .A(n9867), .Y(n9865) );
  INVX1 U9830 ( .A(n9865), .Y(n9866) );
  BUFX2 U9831 ( .A(fifo[740]), .Y(n9867) );
  INVX1 U9832 ( .A(n9870), .Y(n9868) );
  INVX1 U9833 ( .A(n9868), .Y(n9869) );
  BUFX2 U9834 ( .A(fifo[741]), .Y(n9870) );
  INVX1 U9835 ( .A(n9873), .Y(n9871) );
  INVX1 U9836 ( .A(n9871), .Y(n9872) );
  BUFX2 U9837 ( .A(fifo[742]), .Y(n9873) );
  INVX1 U9838 ( .A(n9876), .Y(n9874) );
  INVX1 U9839 ( .A(n9874), .Y(n9875) );
  BUFX2 U9840 ( .A(fifo[743]), .Y(n9876) );
  INVX1 U9841 ( .A(n9879), .Y(n9877) );
  INVX1 U9842 ( .A(n9877), .Y(n9878) );
  BUFX2 U9843 ( .A(fifo[744]), .Y(n9879) );
  INVX1 U9844 ( .A(n9882), .Y(n9880) );
  INVX1 U9845 ( .A(n9880), .Y(n9881) );
  BUFX2 U9846 ( .A(fifo[745]), .Y(n9882) );
  INVX1 U9847 ( .A(n9885), .Y(n9883) );
  INVX1 U9848 ( .A(n9883), .Y(n9884) );
  BUFX2 U9849 ( .A(fifo[746]), .Y(n9885) );
  INVX1 U9850 ( .A(n9888), .Y(n9886) );
  INVX1 U9851 ( .A(n9886), .Y(n9887) );
  BUFX2 U9852 ( .A(fifo[747]), .Y(n9888) );
  INVX1 U9853 ( .A(n9891), .Y(n9889) );
  INVX1 U9854 ( .A(n9889), .Y(n9890) );
  BUFX2 U9855 ( .A(fifo[748]), .Y(n9891) );
  INVX1 U9856 ( .A(n9894), .Y(n9892) );
  INVX1 U9857 ( .A(n9892), .Y(n9893) );
  BUFX2 U9858 ( .A(fifo[749]), .Y(n9894) );
  INVX1 U9859 ( .A(n9897), .Y(n9895) );
  INVX1 U9860 ( .A(n9895), .Y(n9896) );
  BUFX2 U9861 ( .A(fifo[750]), .Y(n9897) );
  INVX1 U9862 ( .A(n9900), .Y(n9898) );
  INVX1 U9863 ( .A(n9898), .Y(n9899) );
  BUFX2 U9864 ( .A(fifo[751]), .Y(n9900) );
  INVX1 U9865 ( .A(n9903), .Y(n9901) );
  INVX1 U9866 ( .A(n9901), .Y(n9902) );
  BUFX2 U9867 ( .A(fifo[752]), .Y(n9903) );
  INVX1 U9868 ( .A(n9906), .Y(n9904) );
  INVX1 U9869 ( .A(n9904), .Y(n9905) );
  BUFX2 U9870 ( .A(fifo[753]), .Y(n9906) );
  INVX1 U9871 ( .A(n9909), .Y(n9907) );
  INVX1 U9872 ( .A(n9907), .Y(n9908) );
  BUFX2 U9873 ( .A(fifo[754]), .Y(n9909) );
  INVX1 U9874 ( .A(n9912), .Y(n9910) );
  INVX1 U9875 ( .A(n9910), .Y(n9911) );
  BUFX2 U9876 ( .A(fifo[755]), .Y(n9912) );
  INVX1 U9877 ( .A(n9915), .Y(n9913) );
  INVX1 U9878 ( .A(n9913), .Y(n9914) );
  BUFX2 U9879 ( .A(fifo[798]), .Y(n9915) );
  INVX1 U9880 ( .A(n9918), .Y(n9916) );
  INVX1 U9881 ( .A(n9916), .Y(n9917) );
  BUFX2 U9882 ( .A(fifo[799]), .Y(n9918) );
  INVX1 U9883 ( .A(n9921), .Y(n9919) );
  INVX1 U9884 ( .A(n9919), .Y(n9920) );
  BUFX2 U9885 ( .A(fifo[800]), .Y(n9921) );
  INVX1 U9886 ( .A(n9924), .Y(n9922) );
  INVX1 U9887 ( .A(n9922), .Y(n9923) );
  BUFX2 U9888 ( .A(fifo[801]), .Y(n9924) );
  INVX1 U9889 ( .A(n9927), .Y(n9925) );
  INVX1 U9890 ( .A(n9925), .Y(n9926) );
  BUFX2 U9891 ( .A(fifo[802]), .Y(n9927) );
  INVX1 U9892 ( .A(n9930), .Y(n9928) );
  INVX1 U9893 ( .A(n9928), .Y(n9929) );
  BUFX2 U9894 ( .A(fifo[803]), .Y(n9930) );
  INVX1 U9895 ( .A(n9933), .Y(n9931) );
  INVX1 U9896 ( .A(n9931), .Y(n9932) );
  BUFX2 U9897 ( .A(fifo[804]), .Y(n9933) );
  INVX1 U9898 ( .A(n9936), .Y(n9934) );
  INVX1 U9899 ( .A(n9934), .Y(n9935) );
  BUFX2 U9900 ( .A(fifo[805]), .Y(n9936) );
  INVX1 U9901 ( .A(n9939), .Y(n9937) );
  INVX1 U9902 ( .A(n9937), .Y(n9938) );
  BUFX2 U9903 ( .A(fifo[806]), .Y(n9939) );
  INVX1 U9904 ( .A(n9942), .Y(n9940) );
  INVX1 U9905 ( .A(n9940), .Y(n9941) );
  BUFX2 U9906 ( .A(fifo[807]), .Y(n9942) );
  INVX1 U9907 ( .A(n9945), .Y(n9943) );
  INVX1 U9908 ( .A(n9943), .Y(n9944) );
  BUFX2 U9909 ( .A(fifo[808]), .Y(n9945) );
  INVX1 U9910 ( .A(n9948), .Y(n9946) );
  INVX1 U9911 ( .A(n9946), .Y(n9947) );
  BUFX2 U9912 ( .A(fifo[809]), .Y(n9948) );
  INVX1 U9913 ( .A(n9951), .Y(n9949) );
  INVX1 U9914 ( .A(n9949), .Y(n9950) );
  BUFX2 U9915 ( .A(fifo[810]), .Y(n9951) );
  INVX1 U9916 ( .A(n9954), .Y(n9952) );
  INVX1 U9917 ( .A(n9952), .Y(n9953) );
  BUFX2 U9918 ( .A(fifo[811]), .Y(n9954) );
  INVX1 U9919 ( .A(n9957), .Y(n9955) );
  INVX1 U9920 ( .A(n9955), .Y(n9956) );
  BUFX2 U9921 ( .A(fifo[812]), .Y(n9957) );
  INVX1 U9922 ( .A(n9960), .Y(n9958) );
  INVX1 U9923 ( .A(n9958), .Y(n9959) );
  BUFX2 U9924 ( .A(fifo[813]), .Y(n9960) );
  INVX1 U9925 ( .A(n9963), .Y(n9961) );
  INVX1 U9926 ( .A(n9961), .Y(n9962) );
  BUFX2 U9927 ( .A(fifo[814]), .Y(n9963) );
  INVX1 U9928 ( .A(n9966), .Y(n9964) );
  INVX1 U9929 ( .A(n9964), .Y(n9965) );
  BUFX2 U9930 ( .A(fifo[815]), .Y(n9966) );
  INVX1 U9931 ( .A(n9969), .Y(n9967) );
  INVX1 U9932 ( .A(n9967), .Y(n9968) );
  BUFX2 U9933 ( .A(fifo[816]), .Y(n9969) );
  INVX1 U9934 ( .A(n9972), .Y(n9970) );
  INVX1 U9935 ( .A(n9970), .Y(n9971) );
  BUFX2 U9936 ( .A(fifo[817]), .Y(n9972) );
  INVX1 U9937 ( .A(n9975), .Y(n9973) );
  INVX1 U9938 ( .A(n9973), .Y(n9974) );
  BUFX2 U9939 ( .A(fifo[818]), .Y(n9975) );
  INVX1 U9940 ( .A(n9978), .Y(n9976) );
  INVX1 U9941 ( .A(n9976), .Y(n9977) );
  BUFX2 U9942 ( .A(fifo[819]), .Y(n9978) );
  INVX1 U9943 ( .A(n9981), .Y(n9979) );
  INVX1 U9944 ( .A(n9979), .Y(n9980) );
  BUFX2 U9945 ( .A(fifo[820]), .Y(n9981) );
  INVX1 U9946 ( .A(n9984), .Y(n9982) );
  INVX1 U9947 ( .A(n9982), .Y(n9983) );
  BUFX2 U9948 ( .A(fifo[821]), .Y(n9984) );
  INVX1 U9949 ( .A(n9987), .Y(n9985) );
  INVX1 U9950 ( .A(n9985), .Y(n9986) );
  BUFX2 U9951 ( .A(fifo[822]), .Y(n9987) );
  INVX1 U9952 ( .A(n9990), .Y(n9988) );
  INVX1 U9953 ( .A(n9988), .Y(n9989) );
  BUFX2 U9954 ( .A(fifo[823]), .Y(n9990) );
  INVX1 U9955 ( .A(n9993), .Y(n9991) );
  INVX1 U9956 ( .A(n9991), .Y(n9992) );
  BUFX2 U9957 ( .A(fifo[824]), .Y(n9993) );
  INVX1 U9958 ( .A(n9996), .Y(n9994) );
  INVX1 U9959 ( .A(n9994), .Y(n9995) );
  BUFX2 U9960 ( .A(fifo[825]), .Y(n9996) );
  INVX1 U9961 ( .A(n9999), .Y(n9997) );
  INVX1 U9962 ( .A(n9997), .Y(n9998) );
  BUFX2 U9963 ( .A(fifo[826]), .Y(n9999) );
  INVX1 U9964 ( .A(n10002), .Y(n10000) );
  INVX1 U9965 ( .A(n10000), .Y(n10001) );
  BUFX2 U9966 ( .A(fifo[827]), .Y(n10002) );
  INVX1 U9967 ( .A(n10005), .Y(n10003) );
  INVX1 U9968 ( .A(n10003), .Y(n10004) );
  BUFX2 U9969 ( .A(fifo[828]), .Y(n10005) );
  INVX1 U9970 ( .A(n10008), .Y(n10006) );
  INVX1 U9971 ( .A(n10006), .Y(n10007) );
  BUFX2 U9972 ( .A(fifo[829]), .Y(n10008) );
  INVX1 U9973 ( .A(n10011), .Y(n10009) );
  INVX1 U9974 ( .A(n10009), .Y(n10010) );
  BUFX2 U9975 ( .A(fifo[830]), .Y(n10011) );
  INVX1 U9976 ( .A(n10014), .Y(n10012) );
  INVX1 U9977 ( .A(n10012), .Y(n10013) );
  BUFX2 U9978 ( .A(fifo[831]), .Y(n10014) );
  INVX1 U9979 ( .A(n10017), .Y(n10015) );
  INVX1 U9980 ( .A(n10015), .Y(n10016) );
  BUFX2 U9981 ( .A(fifo[832]), .Y(n10017) );
  INVX1 U9982 ( .A(n10020), .Y(n10018) );
  INVX1 U9983 ( .A(n10018), .Y(n10019) );
  BUFX2 U9984 ( .A(fifo[833]), .Y(n10020) );
  INVX1 U9985 ( .A(n10023), .Y(n10021) );
  INVX1 U9986 ( .A(n10021), .Y(n10022) );
  BUFX2 U9987 ( .A(fifo[834]), .Y(n10023) );
  INVX1 U9988 ( .A(n10026), .Y(n10024) );
  INVX1 U9989 ( .A(n10024), .Y(n10025) );
  BUFX2 U9990 ( .A(fifo[835]), .Y(n10026) );
  INVX1 U9991 ( .A(n10029), .Y(n10027) );
  INVX1 U9992 ( .A(n10027), .Y(n10028) );
  BUFX2 U9993 ( .A(fifo[836]), .Y(n10029) );
  INVX1 U9994 ( .A(n10032), .Y(n10030) );
  INVX1 U9995 ( .A(n10030), .Y(n10031) );
  BUFX2 U9996 ( .A(fifo[837]), .Y(n10032) );
  INVX1 U9997 ( .A(n10035), .Y(n10033) );
  INVX1 U9998 ( .A(n10033), .Y(n10034) );
  BUFX2 U9999 ( .A(fifo[838]), .Y(n10035) );
  INVX1 U10000 ( .A(n10038), .Y(n10036) );
  INVX1 U10001 ( .A(n10036), .Y(n10037) );
  BUFX2 U10002 ( .A(fifo[839]), .Y(n10038) );
  INVX1 U10003 ( .A(n10041), .Y(n10039) );
  INVX1 U10004 ( .A(n10039), .Y(n10040) );
  BUFX2 U10005 ( .A(fifo[882]), .Y(n10041) );
  INVX1 U10006 ( .A(n10044), .Y(n10042) );
  INVX1 U10007 ( .A(n10042), .Y(n10043) );
  BUFX2 U10008 ( .A(fifo[883]), .Y(n10044) );
  INVX1 U10009 ( .A(n10047), .Y(n10045) );
  INVX1 U10010 ( .A(n10045), .Y(n10046) );
  BUFX2 U10011 ( .A(fifo[884]), .Y(n10047) );
  INVX1 U10012 ( .A(n10050), .Y(n10048) );
  INVX1 U10013 ( .A(n10048), .Y(n10049) );
  BUFX2 U10014 ( .A(fifo[885]), .Y(n10050) );
  INVX1 U10015 ( .A(n10053), .Y(n10051) );
  INVX1 U10016 ( .A(n10051), .Y(n10052) );
  BUFX2 U10017 ( .A(fifo[886]), .Y(n10053) );
  INVX1 U10018 ( .A(n10056), .Y(n10054) );
  INVX1 U10019 ( .A(n10054), .Y(n10055) );
  BUFX2 U10020 ( .A(fifo[887]), .Y(n10056) );
  INVX1 U10021 ( .A(n10059), .Y(n10057) );
  INVX1 U10022 ( .A(n10057), .Y(n10058) );
  BUFX2 U10023 ( .A(fifo[888]), .Y(n10059) );
  INVX1 U10024 ( .A(n10062), .Y(n10060) );
  INVX1 U10025 ( .A(n10060), .Y(n10061) );
  BUFX2 U10026 ( .A(fifo[889]), .Y(n10062) );
  INVX1 U10027 ( .A(n10065), .Y(n10063) );
  INVX1 U10028 ( .A(n10063), .Y(n10064) );
  BUFX2 U10029 ( .A(fifo[890]), .Y(n10065) );
  INVX1 U10030 ( .A(n10068), .Y(n10066) );
  INVX1 U10031 ( .A(n10066), .Y(n10067) );
  BUFX2 U10032 ( .A(fifo[891]), .Y(n10068) );
  INVX1 U10033 ( .A(n10071), .Y(n10069) );
  INVX1 U10034 ( .A(n10069), .Y(n10070) );
  BUFX2 U10035 ( .A(fifo[892]), .Y(n10071) );
  INVX1 U10036 ( .A(n10074), .Y(n10072) );
  INVX1 U10037 ( .A(n10072), .Y(n10073) );
  BUFX2 U10038 ( .A(fifo[893]), .Y(n10074) );
  INVX1 U10039 ( .A(n10077), .Y(n10075) );
  INVX1 U10040 ( .A(n10075), .Y(n10076) );
  BUFX2 U10041 ( .A(fifo[894]), .Y(n10077) );
  INVX1 U10042 ( .A(n10080), .Y(n10078) );
  INVX1 U10043 ( .A(n10078), .Y(n10079) );
  BUFX2 U10044 ( .A(fifo[895]), .Y(n10080) );
  INVX1 U10045 ( .A(n10083), .Y(n10081) );
  INVX1 U10046 ( .A(n10081), .Y(n10082) );
  BUFX2 U10047 ( .A(fifo[896]), .Y(n10083) );
  INVX1 U10048 ( .A(n10086), .Y(n10084) );
  INVX1 U10049 ( .A(n10084), .Y(n10085) );
  BUFX2 U10050 ( .A(fifo[897]), .Y(n10086) );
  INVX1 U10051 ( .A(n10089), .Y(n10087) );
  INVX1 U10052 ( .A(n10087), .Y(n10088) );
  BUFX2 U10053 ( .A(fifo[898]), .Y(n10089) );
  INVX1 U10054 ( .A(n10092), .Y(n10090) );
  INVX1 U10055 ( .A(n10090), .Y(n10091) );
  BUFX2 U10056 ( .A(fifo[899]), .Y(n10092) );
  INVX1 U10057 ( .A(n10095), .Y(n10093) );
  INVX1 U10058 ( .A(n10093), .Y(n10094) );
  BUFX2 U10059 ( .A(fifo[900]), .Y(n10095) );
  INVX1 U10060 ( .A(n10098), .Y(n10096) );
  INVX1 U10061 ( .A(n10096), .Y(n10097) );
  BUFX2 U10062 ( .A(fifo[901]), .Y(n10098) );
  INVX1 U10063 ( .A(n10101), .Y(n10099) );
  INVX1 U10064 ( .A(n10099), .Y(n10100) );
  BUFX2 U10065 ( .A(fifo[902]), .Y(n10101) );
  INVX1 U10066 ( .A(n10104), .Y(n10102) );
  INVX1 U10067 ( .A(n10102), .Y(n10103) );
  BUFX2 U10068 ( .A(fifo[903]), .Y(n10104) );
  INVX1 U10069 ( .A(n10107), .Y(n10105) );
  INVX1 U10070 ( .A(n10105), .Y(n10106) );
  BUFX2 U10071 ( .A(fifo[904]), .Y(n10107) );
  INVX1 U10072 ( .A(n10110), .Y(n10108) );
  INVX1 U10073 ( .A(n10108), .Y(n10109) );
  BUFX2 U10074 ( .A(fifo[905]), .Y(n10110) );
  INVX1 U10075 ( .A(n10113), .Y(n10111) );
  INVX1 U10076 ( .A(n10111), .Y(n10112) );
  BUFX2 U10077 ( .A(fifo[906]), .Y(n10113) );
  INVX1 U10078 ( .A(n10116), .Y(n10114) );
  INVX1 U10079 ( .A(n10114), .Y(n10115) );
  BUFX2 U10080 ( .A(fifo[907]), .Y(n10116) );
  INVX1 U10081 ( .A(n10119), .Y(n10117) );
  INVX1 U10082 ( .A(n10117), .Y(n10118) );
  BUFX2 U10083 ( .A(fifo[908]), .Y(n10119) );
  INVX1 U10084 ( .A(n10122), .Y(n10120) );
  INVX1 U10085 ( .A(n10120), .Y(n10121) );
  BUFX2 U10086 ( .A(fifo[909]), .Y(n10122) );
  INVX1 U10087 ( .A(n10125), .Y(n10123) );
  INVX1 U10088 ( .A(n10123), .Y(n10124) );
  BUFX2 U10089 ( .A(fifo[910]), .Y(n10125) );
  INVX1 U10090 ( .A(n10128), .Y(n10126) );
  INVX1 U10091 ( .A(n10126), .Y(n10127) );
  BUFX2 U10092 ( .A(fifo[911]), .Y(n10128) );
  INVX1 U10093 ( .A(n10131), .Y(n10129) );
  INVX1 U10094 ( .A(n10129), .Y(n10130) );
  BUFX2 U10095 ( .A(fifo[912]), .Y(n10131) );
  INVX1 U10096 ( .A(n10134), .Y(n10132) );
  INVX1 U10097 ( .A(n10132), .Y(n10133) );
  BUFX2 U10098 ( .A(fifo[913]), .Y(n10134) );
  INVX1 U10099 ( .A(n10137), .Y(n10135) );
  INVX1 U10100 ( .A(n10135), .Y(n10136) );
  BUFX2 U10101 ( .A(fifo[914]), .Y(n10137) );
  INVX1 U10102 ( .A(n10140), .Y(n10138) );
  INVX1 U10103 ( .A(n10138), .Y(n10139) );
  BUFX2 U10104 ( .A(fifo[915]), .Y(n10140) );
  INVX1 U10105 ( .A(n10143), .Y(n10141) );
  INVX1 U10106 ( .A(n10141), .Y(n10142) );
  BUFX2 U10107 ( .A(fifo[916]), .Y(n10143) );
  INVX1 U10108 ( .A(n10146), .Y(n10144) );
  INVX1 U10109 ( .A(n10144), .Y(n10145) );
  BUFX2 U10110 ( .A(fifo[917]), .Y(n10146) );
  INVX1 U10111 ( .A(n10149), .Y(n10147) );
  INVX1 U10112 ( .A(n10147), .Y(n10148) );
  BUFX2 U10113 ( .A(fifo[918]), .Y(n10149) );
  INVX1 U10114 ( .A(n10152), .Y(n10150) );
  INVX1 U10115 ( .A(n10150), .Y(n10151) );
  BUFX2 U10116 ( .A(fifo[919]), .Y(n10152) );
  INVX1 U10117 ( .A(n10155), .Y(n10153) );
  INVX1 U10118 ( .A(n10153), .Y(n10154) );
  BUFX2 U10119 ( .A(fifo[920]), .Y(n10155) );
  INVX1 U10120 ( .A(n10158), .Y(n10156) );
  INVX1 U10121 ( .A(n10156), .Y(n10157) );
  BUFX2 U10122 ( .A(fifo[921]), .Y(n10158) );
  INVX1 U10123 ( .A(n10161), .Y(n10159) );
  INVX1 U10124 ( .A(n10159), .Y(n10160) );
  BUFX2 U10125 ( .A(fifo[922]), .Y(n10161) );
  INVX1 U10126 ( .A(n10164), .Y(n10162) );
  INVX1 U10127 ( .A(n10162), .Y(n10163) );
  BUFX2 U10128 ( .A(fifo[923]), .Y(n10164) );
  INVX1 U10129 ( .A(n10167), .Y(n10165) );
  INVX1 U10130 ( .A(n10165), .Y(n10166) );
  BUFX2 U10131 ( .A(fifo[966]), .Y(n10167) );
  INVX1 U10132 ( .A(n10170), .Y(n10168) );
  INVX1 U10133 ( .A(n10168), .Y(n10169) );
  BUFX2 U10134 ( .A(fifo[967]), .Y(n10170) );
  INVX1 U10135 ( .A(n10173), .Y(n10171) );
  INVX1 U10136 ( .A(n10171), .Y(n10172) );
  BUFX2 U10137 ( .A(fifo[968]), .Y(n10173) );
  INVX1 U10138 ( .A(n10176), .Y(n10174) );
  INVX1 U10139 ( .A(n10174), .Y(n10175) );
  BUFX2 U10140 ( .A(fifo[969]), .Y(n10176) );
  INVX1 U10141 ( .A(n10179), .Y(n10177) );
  INVX1 U10142 ( .A(n10177), .Y(n10178) );
  BUFX2 U10143 ( .A(fifo[970]), .Y(n10179) );
  INVX1 U10144 ( .A(n10182), .Y(n10180) );
  INVX1 U10145 ( .A(n10180), .Y(n10181) );
  BUFX2 U10146 ( .A(fifo[971]), .Y(n10182) );
  INVX1 U10147 ( .A(n10185), .Y(n10183) );
  INVX1 U10148 ( .A(n10183), .Y(n10184) );
  BUFX2 U10149 ( .A(fifo[972]), .Y(n10185) );
  INVX1 U10150 ( .A(n10188), .Y(n10186) );
  INVX1 U10151 ( .A(n10186), .Y(n10187) );
  BUFX2 U10152 ( .A(fifo[973]), .Y(n10188) );
  INVX1 U10153 ( .A(n10191), .Y(n10189) );
  INVX1 U10154 ( .A(n10189), .Y(n10190) );
  BUFX2 U10155 ( .A(fifo[974]), .Y(n10191) );
  INVX1 U10156 ( .A(n10194), .Y(n10192) );
  INVX1 U10157 ( .A(n10192), .Y(n10193) );
  BUFX2 U10158 ( .A(fifo[975]), .Y(n10194) );
  INVX1 U10159 ( .A(n10197), .Y(n10195) );
  INVX1 U10160 ( .A(n10195), .Y(n10196) );
  BUFX2 U10161 ( .A(fifo[976]), .Y(n10197) );
  INVX1 U10162 ( .A(n10200), .Y(n10198) );
  INVX1 U10163 ( .A(n10198), .Y(n10199) );
  BUFX2 U10164 ( .A(fifo[977]), .Y(n10200) );
  INVX1 U10165 ( .A(n10203), .Y(n10201) );
  INVX1 U10166 ( .A(n10201), .Y(n10202) );
  BUFX2 U10167 ( .A(fifo[978]), .Y(n10203) );
  INVX1 U10168 ( .A(n10206), .Y(n10204) );
  INVX1 U10169 ( .A(n10204), .Y(n10205) );
  BUFX2 U10170 ( .A(fifo[979]), .Y(n10206) );
  INVX1 U10171 ( .A(n10209), .Y(n10207) );
  INVX1 U10172 ( .A(n10207), .Y(n10208) );
  BUFX2 U10173 ( .A(fifo[980]), .Y(n10209) );
  INVX1 U10174 ( .A(n10212), .Y(n10210) );
  INVX1 U10175 ( .A(n10210), .Y(n10211) );
  BUFX2 U10176 ( .A(fifo[981]), .Y(n10212) );
  INVX1 U10177 ( .A(n10215), .Y(n10213) );
  INVX1 U10178 ( .A(n10213), .Y(n10214) );
  BUFX2 U10179 ( .A(fifo[982]), .Y(n10215) );
  INVX1 U10180 ( .A(n10218), .Y(n10216) );
  INVX1 U10181 ( .A(n10216), .Y(n10217) );
  BUFX2 U10182 ( .A(fifo[983]), .Y(n10218) );
  INVX1 U10183 ( .A(n10221), .Y(n10219) );
  INVX1 U10184 ( .A(n10219), .Y(n10220) );
  BUFX2 U10185 ( .A(fifo[984]), .Y(n10221) );
  INVX1 U10186 ( .A(n10224), .Y(n10222) );
  INVX1 U10187 ( .A(n10222), .Y(n10223) );
  BUFX2 U10188 ( .A(fifo[985]), .Y(n10224) );
  INVX1 U10189 ( .A(n10227), .Y(n10225) );
  INVX1 U10190 ( .A(n10225), .Y(n10226) );
  BUFX2 U10191 ( .A(fifo[986]), .Y(n10227) );
  INVX1 U10192 ( .A(n10230), .Y(n10228) );
  INVX1 U10193 ( .A(n10228), .Y(n10229) );
  BUFX2 U10194 ( .A(fifo[987]), .Y(n10230) );
  INVX1 U10195 ( .A(n10233), .Y(n10231) );
  INVX1 U10196 ( .A(n10231), .Y(n10232) );
  BUFX2 U10197 ( .A(fifo[988]), .Y(n10233) );
  INVX1 U10198 ( .A(n10236), .Y(n10234) );
  INVX1 U10199 ( .A(n10234), .Y(n10235) );
  BUFX2 U10200 ( .A(fifo[989]), .Y(n10236) );
  INVX1 U10201 ( .A(n10239), .Y(n10237) );
  INVX1 U10202 ( .A(n10237), .Y(n10238) );
  BUFX2 U10203 ( .A(fifo[990]), .Y(n10239) );
  INVX1 U10204 ( .A(n10242), .Y(n10240) );
  INVX1 U10205 ( .A(n10240), .Y(n10241) );
  BUFX2 U10206 ( .A(fifo[991]), .Y(n10242) );
  INVX1 U10207 ( .A(n10245), .Y(n10243) );
  INVX1 U10208 ( .A(n10243), .Y(n10244) );
  BUFX2 U10209 ( .A(fifo[992]), .Y(n10245) );
  INVX1 U10210 ( .A(n10248), .Y(n10246) );
  INVX1 U10211 ( .A(n10246), .Y(n10247) );
  BUFX2 U10212 ( .A(fifo[993]), .Y(n10248) );
  INVX1 U10213 ( .A(n10251), .Y(n10249) );
  INVX1 U10214 ( .A(n10249), .Y(n10250) );
  BUFX2 U10215 ( .A(fifo[994]), .Y(n10251) );
  INVX1 U10216 ( .A(n10254), .Y(n10252) );
  INVX1 U10217 ( .A(n10252), .Y(n10253) );
  BUFX2 U10218 ( .A(fifo[995]), .Y(n10254) );
  INVX1 U10219 ( .A(n10257), .Y(n10255) );
  INVX1 U10220 ( .A(n10255), .Y(n10256) );
  BUFX2 U10221 ( .A(fifo[996]), .Y(n10257) );
  INVX1 U10222 ( .A(n10260), .Y(n10258) );
  INVX1 U10223 ( .A(n10258), .Y(n10259) );
  BUFX2 U10224 ( .A(fifo[997]), .Y(n10260) );
  INVX1 U10225 ( .A(n10263), .Y(n10261) );
  INVX1 U10226 ( .A(n10261), .Y(n10262) );
  BUFX2 U10227 ( .A(fifo[998]), .Y(n10263) );
  INVX1 U10228 ( .A(n10266), .Y(n10264) );
  INVX1 U10229 ( .A(n10264), .Y(n10265) );
  BUFX2 U10230 ( .A(fifo[999]), .Y(n10266) );
  INVX1 U10231 ( .A(n10269), .Y(n10267) );
  INVX1 U10232 ( .A(n10267), .Y(n10268) );
  BUFX2 U10233 ( .A(fifo[1000]), .Y(n10269) );
  INVX1 U10234 ( .A(n10272), .Y(n10270) );
  INVX1 U10235 ( .A(n10270), .Y(n10271) );
  BUFX2 U10236 ( .A(fifo[1001]), .Y(n10272) );
  INVX1 U10237 ( .A(n10275), .Y(n10273) );
  INVX1 U10238 ( .A(n10273), .Y(n10274) );
  BUFX2 U10239 ( .A(fifo[1002]), .Y(n10275) );
  INVX1 U10240 ( .A(n10278), .Y(n10276) );
  INVX1 U10241 ( .A(n10276), .Y(n10277) );
  BUFX2 U10242 ( .A(fifo[1003]), .Y(n10278) );
  INVX1 U10243 ( .A(n10281), .Y(n10279) );
  INVX1 U10244 ( .A(n10279), .Y(n10280) );
  BUFX2 U10245 ( .A(fifo[1004]), .Y(n10281) );
  INVX1 U10246 ( .A(n10284), .Y(n10282) );
  INVX1 U10247 ( .A(n10282), .Y(n10283) );
  BUFX2 U10248 ( .A(fifo[1005]), .Y(n10284) );
  INVX1 U10249 ( .A(n10287), .Y(n10285) );
  INVX1 U10250 ( .A(n10285), .Y(n10286) );
  BUFX2 U10251 ( .A(fifo[1006]), .Y(n10287) );
  INVX1 U10252 ( .A(n10290), .Y(n10288) );
  INVX1 U10253 ( .A(n10288), .Y(n10289) );
  BUFX2 U10254 ( .A(fifo[1007]), .Y(n10290) );
  INVX1 U10255 ( .A(n10293), .Y(n10291) );
  INVX1 U10256 ( .A(n10291), .Y(n10292) );
  BUFX2 U10257 ( .A(fifo[1050]), .Y(n10293) );
  INVX1 U10258 ( .A(n10296), .Y(n10294) );
  INVX1 U10259 ( .A(n10294), .Y(n10295) );
  BUFX2 U10260 ( .A(fifo[1051]), .Y(n10296) );
  INVX1 U10261 ( .A(n10299), .Y(n10297) );
  INVX1 U10262 ( .A(n10297), .Y(n10298) );
  BUFX2 U10263 ( .A(fifo[1052]), .Y(n10299) );
  INVX1 U10264 ( .A(n10302), .Y(n10300) );
  INVX1 U10265 ( .A(n10300), .Y(n10301) );
  BUFX2 U10266 ( .A(fifo[1053]), .Y(n10302) );
  INVX1 U10267 ( .A(n10305), .Y(n10303) );
  INVX1 U10268 ( .A(n10303), .Y(n10304) );
  BUFX2 U10269 ( .A(fifo[1054]), .Y(n10305) );
  INVX1 U10270 ( .A(n10308), .Y(n10306) );
  INVX1 U10271 ( .A(n10306), .Y(n10307) );
  BUFX2 U10272 ( .A(fifo[1055]), .Y(n10308) );
  INVX1 U10273 ( .A(n10311), .Y(n10309) );
  INVX1 U10274 ( .A(n10309), .Y(n10310) );
  BUFX2 U10275 ( .A(fifo[1056]), .Y(n10311) );
  INVX1 U10276 ( .A(n10314), .Y(n10312) );
  INVX1 U10277 ( .A(n10312), .Y(n10313) );
  BUFX2 U10278 ( .A(fifo[1057]), .Y(n10314) );
  INVX1 U10279 ( .A(n10317), .Y(n10315) );
  INVX1 U10280 ( .A(n10315), .Y(n10316) );
  BUFX2 U10281 ( .A(fifo[1058]), .Y(n10317) );
  INVX1 U10282 ( .A(n10320), .Y(n10318) );
  INVX1 U10283 ( .A(n10318), .Y(n10319) );
  BUFX2 U10284 ( .A(fifo[1059]), .Y(n10320) );
  INVX1 U10285 ( .A(n10323), .Y(n10321) );
  INVX1 U10286 ( .A(n10321), .Y(n10322) );
  BUFX2 U10287 ( .A(fifo[1060]), .Y(n10323) );
  INVX1 U10288 ( .A(n10326), .Y(n10324) );
  INVX1 U10289 ( .A(n10324), .Y(n10325) );
  BUFX2 U10290 ( .A(fifo[1061]), .Y(n10326) );
  INVX1 U10291 ( .A(n10329), .Y(n10327) );
  INVX1 U10292 ( .A(n10327), .Y(n10328) );
  BUFX2 U10293 ( .A(fifo[1062]), .Y(n10329) );
  INVX1 U10294 ( .A(n10332), .Y(n10330) );
  INVX1 U10295 ( .A(n10330), .Y(n10331) );
  BUFX2 U10296 ( .A(fifo[1063]), .Y(n10332) );
  INVX1 U10297 ( .A(n10335), .Y(n10333) );
  INVX1 U10298 ( .A(n10333), .Y(n10334) );
  BUFX2 U10299 ( .A(fifo[1064]), .Y(n10335) );
  INVX1 U10300 ( .A(n10338), .Y(n10336) );
  INVX1 U10301 ( .A(n10336), .Y(n10337) );
  BUFX2 U10302 ( .A(fifo[1065]), .Y(n10338) );
  INVX1 U10303 ( .A(n10341), .Y(n10339) );
  INVX1 U10304 ( .A(n10339), .Y(n10340) );
  BUFX2 U10305 ( .A(fifo[1066]), .Y(n10341) );
  INVX1 U10306 ( .A(n10344), .Y(n10342) );
  INVX1 U10307 ( .A(n10342), .Y(n10343) );
  BUFX2 U10308 ( .A(fifo[1067]), .Y(n10344) );
  INVX1 U10309 ( .A(n10347), .Y(n10345) );
  INVX1 U10310 ( .A(n10345), .Y(n10346) );
  BUFX2 U10311 ( .A(fifo[1068]), .Y(n10347) );
  INVX1 U10312 ( .A(n10350), .Y(n10348) );
  INVX1 U10313 ( .A(n10348), .Y(n10349) );
  BUFX2 U10314 ( .A(fifo[1069]), .Y(n10350) );
  INVX1 U10315 ( .A(n10353), .Y(n10351) );
  INVX1 U10316 ( .A(n10351), .Y(n10352) );
  BUFX2 U10317 ( .A(fifo[1070]), .Y(n10353) );
  INVX1 U10318 ( .A(n10356), .Y(n10354) );
  INVX1 U10319 ( .A(n10354), .Y(n10355) );
  BUFX2 U10320 ( .A(fifo[1071]), .Y(n10356) );
  INVX1 U10321 ( .A(n10359), .Y(n10357) );
  INVX1 U10322 ( .A(n10357), .Y(n10358) );
  BUFX2 U10323 ( .A(fifo[1072]), .Y(n10359) );
  INVX1 U10324 ( .A(n10362), .Y(n10360) );
  INVX1 U10325 ( .A(n10360), .Y(n10361) );
  BUFX2 U10326 ( .A(fifo[1073]), .Y(n10362) );
  INVX1 U10327 ( .A(n10365), .Y(n10363) );
  INVX1 U10328 ( .A(n10363), .Y(n10364) );
  BUFX2 U10329 ( .A(fifo[1074]), .Y(n10365) );
  INVX1 U10330 ( .A(n10368), .Y(n10366) );
  INVX1 U10331 ( .A(n10366), .Y(n10367) );
  BUFX2 U10332 ( .A(fifo[1075]), .Y(n10368) );
  INVX1 U10333 ( .A(n10371), .Y(n10369) );
  INVX1 U10334 ( .A(n10369), .Y(n10370) );
  BUFX2 U10335 ( .A(fifo[1076]), .Y(n10371) );
  INVX1 U10336 ( .A(n10374), .Y(n10372) );
  INVX1 U10337 ( .A(n10372), .Y(n10373) );
  BUFX2 U10338 ( .A(fifo[1077]), .Y(n10374) );
  INVX1 U10339 ( .A(n10377), .Y(n10375) );
  INVX1 U10340 ( .A(n10375), .Y(n10376) );
  BUFX2 U10341 ( .A(fifo[1078]), .Y(n10377) );
  INVX1 U10342 ( .A(n10380), .Y(n10378) );
  INVX1 U10343 ( .A(n10378), .Y(n10379) );
  BUFX2 U10344 ( .A(fifo[1079]), .Y(n10380) );
  INVX1 U10345 ( .A(n10383), .Y(n10381) );
  INVX1 U10346 ( .A(n10381), .Y(n10382) );
  BUFX2 U10347 ( .A(fifo[1080]), .Y(n10383) );
  INVX1 U10348 ( .A(n10386), .Y(n10384) );
  INVX1 U10349 ( .A(n10384), .Y(n10385) );
  BUFX2 U10350 ( .A(fifo[1081]), .Y(n10386) );
  INVX1 U10351 ( .A(n10389), .Y(n10387) );
  INVX1 U10352 ( .A(n10387), .Y(n10388) );
  BUFX2 U10353 ( .A(fifo[1082]), .Y(n10389) );
  INVX1 U10354 ( .A(n10392), .Y(n10390) );
  INVX1 U10355 ( .A(n10390), .Y(n10391) );
  BUFX2 U10356 ( .A(fifo[1083]), .Y(n10392) );
  INVX1 U10357 ( .A(n10395), .Y(n10393) );
  INVX1 U10358 ( .A(n10393), .Y(n10394) );
  BUFX2 U10359 ( .A(fifo[1084]), .Y(n10395) );
  INVX1 U10360 ( .A(n10398), .Y(n10396) );
  INVX1 U10361 ( .A(n10396), .Y(n10397) );
  BUFX2 U10362 ( .A(fifo[1085]), .Y(n10398) );
  INVX1 U10363 ( .A(n10401), .Y(n10399) );
  INVX1 U10364 ( .A(n10399), .Y(n10400) );
  BUFX2 U10365 ( .A(fifo[1086]), .Y(n10401) );
  INVX1 U10366 ( .A(n10404), .Y(n10402) );
  INVX1 U10367 ( .A(n10402), .Y(n10403) );
  BUFX2 U10368 ( .A(fifo[1087]), .Y(n10404) );
  INVX1 U10369 ( .A(n10407), .Y(n10405) );
  INVX1 U10370 ( .A(n10405), .Y(n10406) );
  BUFX2 U10371 ( .A(fifo[1088]), .Y(n10407) );
  INVX1 U10372 ( .A(n10410), .Y(n10408) );
  INVX1 U10373 ( .A(n10408), .Y(n10409) );
  BUFX2 U10374 ( .A(fifo[1089]), .Y(n10410) );
  INVX1 U10375 ( .A(n10413), .Y(n10411) );
  INVX1 U10376 ( .A(n10411), .Y(n10412) );
  BUFX2 U10377 ( .A(fifo[1090]), .Y(n10413) );
  INVX1 U10378 ( .A(n10416), .Y(n10414) );
  INVX1 U10379 ( .A(n10414), .Y(n10415) );
  BUFX2 U10380 ( .A(fifo[1091]), .Y(n10416) );
  INVX1 U10381 ( .A(n10419), .Y(n10417) );
  INVX1 U10382 ( .A(n10417), .Y(n10418) );
  BUFX2 U10383 ( .A(fifo[1134]), .Y(n10419) );
  INVX1 U10384 ( .A(n10422), .Y(n10420) );
  INVX1 U10385 ( .A(n10420), .Y(n10421) );
  BUFX2 U10386 ( .A(fifo[1135]), .Y(n10422) );
  INVX1 U10387 ( .A(n10425), .Y(n10423) );
  INVX1 U10388 ( .A(n10423), .Y(n10424) );
  BUFX2 U10389 ( .A(fifo[1136]), .Y(n10425) );
  INVX1 U10390 ( .A(n10428), .Y(n10426) );
  INVX1 U10391 ( .A(n10426), .Y(n10427) );
  BUFX2 U10392 ( .A(fifo[1137]), .Y(n10428) );
  INVX1 U10393 ( .A(n10431), .Y(n10429) );
  INVX1 U10394 ( .A(n10429), .Y(n10430) );
  BUFX2 U10395 ( .A(fifo[1138]), .Y(n10431) );
  INVX1 U10396 ( .A(n10434), .Y(n10432) );
  INVX1 U10397 ( .A(n10432), .Y(n10433) );
  BUFX2 U10398 ( .A(fifo[1139]), .Y(n10434) );
  INVX1 U10399 ( .A(n10437), .Y(n10435) );
  INVX1 U10400 ( .A(n10435), .Y(n10436) );
  BUFX2 U10401 ( .A(fifo[1140]), .Y(n10437) );
  INVX1 U10402 ( .A(n10440), .Y(n10438) );
  INVX1 U10403 ( .A(n10438), .Y(n10439) );
  BUFX2 U10404 ( .A(fifo[1141]), .Y(n10440) );
  INVX1 U10405 ( .A(n10443), .Y(n10441) );
  INVX1 U10406 ( .A(n10441), .Y(n10442) );
  BUFX2 U10407 ( .A(fifo[1142]), .Y(n10443) );
  INVX1 U10408 ( .A(n10446), .Y(n10444) );
  INVX1 U10409 ( .A(n10444), .Y(n10445) );
  BUFX2 U10410 ( .A(fifo[1143]), .Y(n10446) );
  INVX1 U10411 ( .A(n10449), .Y(n10447) );
  INVX1 U10412 ( .A(n10447), .Y(n10448) );
  BUFX2 U10413 ( .A(fifo[1144]), .Y(n10449) );
  INVX1 U10414 ( .A(n10452), .Y(n10450) );
  INVX1 U10415 ( .A(n10450), .Y(n10451) );
  BUFX2 U10416 ( .A(fifo[1145]), .Y(n10452) );
  INVX1 U10417 ( .A(n10455), .Y(n10453) );
  INVX1 U10418 ( .A(n10453), .Y(n10454) );
  BUFX2 U10419 ( .A(fifo[1146]), .Y(n10455) );
  INVX1 U10420 ( .A(n10458), .Y(n10456) );
  INVX1 U10421 ( .A(n10456), .Y(n10457) );
  BUFX2 U10422 ( .A(fifo[1147]), .Y(n10458) );
  INVX1 U10423 ( .A(n10461), .Y(n10459) );
  INVX1 U10424 ( .A(n10459), .Y(n10460) );
  BUFX2 U10425 ( .A(fifo[1148]), .Y(n10461) );
  INVX1 U10426 ( .A(n10464), .Y(n10462) );
  INVX1 U10427 ( .A(n10462), .Y(n10463) );
  BUFX2 U10428 ( .A(fifo[1149]), .Y(n10464) );
  INVX1 U10429 ( .A(n10467), .Y(n10465) );
  INVX1 U10430 ( .A(n10465), .Y(n10466) );
  BUFX2 U10431 ( .A(fifo[1150]), .Y(n10467) );
  INVX1 U10432 ( .A(n10470), .Y(n10468) );
  INVX1 U10433 ( .A(n10468), .Y(n10469) );
  BUFX2 U10434 ( .A(fifo[1151]), .Y(n10470) );
  INVX1 U10435 ( .A(n10473), .Y(n10471) );
  INVX1 U10436 ( .A(n10471), .Y(n10472) );
  BUFX2 U10437 ( .A(fifo[1152]), .Y(n10473) );
  INVX1 U10438 ( .A(n10476), .Y(n10474) );
  INVX1 U10439 ( .A(n10474), .Y(n10475) );
  BUFX2 U10440 ( .A(fifo[1153]), .Y(n10476) );
  INVX1 U10441 ( .A(n10479), .Y(n10477) );
  INVX1 U10442 ( .A(n10477), .Y(n10478) );
  BUFX2 U10443 ( .A(fifo[1154]), .Y(n10479) );
  INVX1 U10444 ( .A(n10482), .Y(n10480) );
  INVX1 U10445 ( .A(n10480), .Y(n10481) );
  BUFX2 U10446 ( .A(fifo[1155]), .Y(n10482) );
  INVX1 U10447 ( .A(n10485), .Y(n10483) );
  INVX1 U10448 ( .A(n10483), .Y(n10484) );
  BUFX2 U10449 ( .A(fifo[1156]), .Y(n10485) );
  INVX1 U10450 ( .A(n10488), .Y(n10486) );
  INVX1 U10451 ( .A(n10486), .Y(n10487) );
  BUFX2 U10452 ( .A(fifo[1157]), .Y(n10488) );
  INVX1 U10453 ( .A(n10491), .Y(n10489) );
  INVX1 U10454 ( .A(n10489), .Y(n10490) );
  BUFX2 U10455 ( .A(fifo[1158]), .Y(n10491) );
  INVX1 U10456 ( .A(n10494), .Y(n10492) );
  INVX1 U10457 ( .A(n10492), .Y(n10493) );
  BUFX2 U10458 ( .A(fifo[1159]), .Y(n10494) );
  INVX1 U10459 ( .A(n10497), .Y(n10495) );
  INVX1 U10460 ( .A(n10495), .Y(n10496) );
  BUFX2 U10461 ( .A(fifo[1160]), .Y(n10497) );
  INVX1 U10462 ( .A(n10500), .Y(n10498) );
  INVX1 U10463 ( .A(n10498), .Y(n10499) );
  BUFX2 U10464 ( .A(fifo[1161]), .Y(n10500) );
  INVX1 U10465 ( .A(n10503), .Y(n10501) );
  INVX1 U10466 ( .A(n10501), .Y(n10502) );
  BUFX2 U10467 ( .A(fifo[1162]), .Y(n10503) );
  INVX1 U10468 ( .A(n10506), .Y(n10504) );
  INVX1 U10469 ( .A(n10504), .Y(n10505) );
  BUFX2 U10470 ( .A(fifo[1163]), .Y(n10506) );
  INVX1 U10471 ( .A(n10509), .Y(n10507) );
  INVX1 U10472 ( .A(n10507), .Y(n10508) );
  BUFX2 U10473 ( .A(fifo[1164]), .Y(n10509) );
  INVX1 U10474 ( .A(n10512), .Y(n10510) );
  INVX1 U10475 ( .A(n10510), .Y(n10511) );
  BUFX2 U10476 ( .A(fifo[1165]), .Y(n10512) );
  INVX1 U10477 ( .A(n10515), .Y(n10513) );
  INVX1 U10478 ( .A(n10513), .Y(n10514) );
  BUFX2 U10479 ( .A(fifo[1166]), .Y(n10515) );
  INVX1 U10480 ( .A(n10518), .Y(n10516) );
  INVX1 U10481 ( .A(n10516), .Y(n10517) );
  BUFX2 U10482 ( .A(fifo[1167]), .Y(n10518) );
  INVX1 U10483 ( .A(n10521), .Y(n10519) );
  INVX1 U10484 ( .A(n10519), .Y(n10520) );
  BUFX2 U10485 ( .A(fifo[1168]), .Y(n10521) );
  INVX1 U10486 ( .A(n10524), .Y(n10522) );
  INVX1 U10487 ( .A(n10522), .Y(n10523) );
  BUFX2 U10488 ( .A(fifo[1169]), .Y(n10524) );
  INVX1 U10489 ( .A(n10527), .Y(n10525) );
  INVX1 U10490 ( .A(n10525), .Y(n10526) );
  BUFX2 U10491 ( .A(fifo[1170]), .Y(n10527) );
  INVX1 U10492 ( .A(n10530), .Y(n10528) );
  INVX1 U10493 ( .A(n10528), .Y(n10529) );
  BUFX2 U10494 ( .A(fifo[1171]), .Y(n10530) );
  INVX1 U10495 ( .A(n10533), .Y(n10531) );
  INVX1 U10496 ( .A(n10531), .Y(n10532) );
  BUFX2 U10497 ( .A(fifo[1172]), .Y(n10533) );
  INVX1 U10498 ( .A(n10536), .Y(n10534) );
  INVX1 U10499 ( .A(n10534), .Y(n10535) );
  BUFX2 U10500 ( .A(fifo[1173]), .Y(n10536) );
  INVX1 U10501 ( .A(n10539), .Y(n10537) );
  INVX1 U10502 ( .A(n10537), .Y(n10538) );
  BUFX2 U10503 ( .A(fifo[1174]), .Y(n10539) );
  INVX1 U10504 ( .A(n10542), .Y(n10540) );
  INVX1 U10505 ( .A(n10540), .Y(n10541) );
  BUFX2 U10506 ( .A(fifo[1175]), .Y(n10542) );
  INVX1 U10507 ( .A(n10545), .Y(n10543) );
  INVX1 U10508 ( .A(n10543), .Y(n10544) );
  BUFX2 U10509 ( .A(fifo[1218]), .Y(n10545) );
  INVX1 U10510 ( .A(n10548), .Y(n10546) );
  INVX1 U10511 ( .A(n10546), .Y(n10547) );
  BUFX2 U10512 ( .A(fifo[1219]), .Y(n10548) );
  INVX1 U10513 ( .A(n10551), .Y(n10549) );
  INVX1 U10514 ( .A(n10549), .Y(n10550) );
  BUFX2 U10515 ( .A(fifo[1220]), .Y(n10551) );
  INVX1 U10516 ( .A(n10554), .Y(n10552) );
  INVX1 U10517 ( .A(n10552), .Y(n10553) );
  BUFX2 U10518 ( .A(fifo[1221]), .Y(n10554) );
  INVX1 U10519 ( .A(n10557), .Y(n10555) );
  INVX1 U10520 ( .A(n10555), .Y(n10556) );
  BUFX2 U10521 ( .A(fifo[1222]), .Y(n10557) );
  INVX1 U10522 ( .A(n10560), .Y(n10558) );
  INVX1 U10523 ( .A(n10558), .Y(n10559) );
  BUFX2 U10524 ( .A(fifo[1223]), .Y(n10560) );
  INVX1 U10525 ( .A(n10563), .Y(n10561) );
  INVX1 U10526 ( .A(n10561), .Y(n10562) );
  BUFX2 U10527 ( .A(fifo[1224]), .Y(n10563) );
  INVX1 U10528 ( .A(n10566), .Y(n10564) );
  INVX1 U10529 ( .A(n10564), .Y(n10565) );
  BUFX2 U10530 ( .A(fifo[1225]), .Y(n10566) );
  INVX1 U10531 ( .A(n10569), .Y(n10567) );
  INVX1 U10532 ( .A(n10567), .Y(n10568) );
  BUFX2 U10533 ( .A(fifo[1226]), .Y(n10569) );
  INVX1 U10534 ( .A(n10572), .Y(n10570) );
  INVX1 U10535 ( .A(n10570), .Y(n10571) );
  BUFX2 U10536 ( .A(fifo[1227]), .Y(n10572) );
  INVX1 U10537 ( .A(n10575), .Y(n10573) );
  INVX1 U10538 ( .A(n10573), .Y(n10574) );
  BUFX2 U10539 ( .A(fifo[1228]), .Y(n10575) );
  INVX1 U10540 ( .A(n10578), .Y(n10576) );
  INVX1 U10541 ( .A(n10576), .Y(n10577) );
  BUFX2 U10542 ( .A(fifo[1229]), .Y(n10578) );
  INVX1 U10543 ( .A(n10581), .Y(n10579) );
  INVX1 U10544 ( .A(n10579), .Y(n10580) );
  BUFX2 U10545 ( .A(fifo[1230]), .Y(n10581) );
  INVX1 U10546 ( .A(n10584), .Y(n10582) );
  INVX1 U10547 ( .A(n10582), .Y(n10583) );
  BUFX2 U10548 ( .A(fifo[1231]), .Y(n10584) );
  INVX1 U10549 ( .A(n10587), .Y(n10585) );
  INVX1 U10550 ( .A(n10585), .Y(n10586) );
  BUFX2 U10551 ( .A(fifo[1232]), .Y(n10587) );
  INVX1 U10552 ( .A(n10590), .Y(n10588) );
  INVX1 U10553 ( .A(n10588), .Y(n10589) );
  BUFX2 U10554 ( .A(fifo[1233]), .Y(n10590) );
  INVX1 U10555 ( .A(n10593), .Y(n10591) );
  INVX1 U10556 ( .A(n10591), .Y(n10592) );
  BUFX2 U10557 ( .A(fifo[1234]), .Y(n10593) );
  INVX1 U10558 ( .A(n10596), .Y(n10594) );
  INVX1 U10559 ( .A(n10594), .Y(n10595) );
  BUFX2 U10560 ( .A(fifo[1235]), .Y(n10596) );
  INVX1 U10561 ( .A(n10599), .Y(n10597) );
  INVX1 U10562 ( .A(n10597), .Y(n10598) );
  BUFX2 U10563 ( .A(fifo[1236]), .Y(n10599) );
  INVX1 U10564 ( .A(n10602), .Y(n10600) );
  INVX1 U10565 ( .A(n10600), .Y(n10601) );
  BUFX2 U10566 ( .A(fifo[1237]), .Y(n10602) );
  INVX1 U10567 ( .A(n10605), .Y(n10603) );
  INVX1 U10568 ( .A(n10603), .Y(n10604) );
  BUFX2 U10569 ( .A(fifo[1238]), .Y(n10605) );
  INVX1 U10570 ( .A(n10608), .Y(n10606) );
  INVX1 U10571 ( .A(n10606), .Y(n10607) );
  BUFX2 U10572 ( .A(fifo[1239]), .Y(n10608) );
  INVX1 U10573 ( .A(n10611), .Y(n10609) );
  INVX1 U10574 ( .A(n10609), .Y(n10610) );
  BUFX2 U10575 ( .A(fifo[1240]), .Y(n10611) );
  INVX1 U10576 ( .A(n10614), .Y(n10612) );
  INVX1 U10577 ( .A(n10612), .Y(n10613) );
  BUFX2 U10578 ( .A(fifo[1241]), .Y(n10614) );
  INVX1 U10579 ( .A(n10617), .Y(n10615) );
  INVX1 U10580 ( .A(n10615), .Y(n10616) );
  BUFX2 U10581 ( .A(fifo[1242]), .Y(n10617) );
  INVX1 U10582 ( .A(n10620), .Y(n10618) );
  INVX1 U10583 ( .A(n10618), .Y(n10619) );
  BUFX2 U10584 ( .A(fifo[1243]), .Y(n10620) );
  INVX1 U10585 ( .A(n10623), .Y(n10621) );
  INVX1 U10586 ( .A(n10621), .Y(n10622) );
  BUFX2 U10587 ( .A(fifo[1244]), .Y(n10623) );
  INVX1 U10588 ( .A(n10626), .Y(n10624) );
  INVX1 U10589 ( .A(n10624), .Y(n10625) );
  BUFX2 U10590 ( .A(fifo[1245]), .Y(n10626) );
  INVX1 U10591 ( .A(n10629), .Y(n10627) );
  INVX1 U10592 ( .A(n10627), .Y(n10628) );
  BUFX2 U10593 ( .A(fifo[1246]), .Y(n10629) );
  INVX1 U10594 ( .A(n10632), .Y(n10630) );
  INVX1 U10595 ( .A(n10630), .Y(n10631) );
  BUFX2 U10596 ( .A(fifo[1247]), .Y(n10632) );
  INVX1 U10597 ( .A(n10635), .Y(n10633) );
  INVX1 U10598 ( .A(n10633), .Y(n10634) );
  BUFX2 U10599 ( .A(fifo[1248]), .Y(n10635) );
  INVX1 U10600 ( .A(n10638), .Y(n10636) );
  INVX1 U10601 ( .A(n10636), .Y(n10637) );
  BUFX2 U10602 ( .A(fifo[1249]), .Y(n10638) );
  INVX1 U10603 ( .A(n10641), .Y(n10639) );
  INVX1 U10604 ( .A(n10639), .Y(n10640) );
  BUFX2 U10605 ( .A(fifo[1250]), .Y(n10641) );
  INVX1 U10606 ( .A(n10644), .Y(n10642) );
  INVX1 U10607 ( .A(n10642), .Y(n10643) );
  BUFX2 U10608 ( .A(fifo[1251]), .Y(n10644) );
  INVX1 U10609 ( .A(n10647), .Y(n10645) );
  INVX1 U10610 ( .A(n10645), .Y(n10646) );
  BUFX2 U10611 ( .A(fifo[1252]), .Y(n10647) );
  INVX1 U10612 ( .A(n10650), .Y(n10648) );
  INVX1 U10613 ( .A(n10648), .Y(n10649) );
  BUFX2 U10614 ( .A(fifo[1253]), .Y(n10650) );
  INVX1 U10615 ( .A(n10653), .Y(n10651) );
  INVX1 U10616 ( .A(n10651), .Y(n10652) );
  BUFX2 U10617 ( .A(fifo[1254]), .Y(n10653) );
  INVX1 U10618 ( .A(n10656), .Y(n10654) );
  INVX1 U10619 ( .A(n10654), .Y(n10655) );
  BUFX2 U10620 ( .A(fifo[1255]), .Y(n10656) );
  INVX1 U10621 ( .A(n10659), .Y(n10657) );
  INVX1 U10622 ( .A(n10657), .Y(n10658) );
  BUFX2 U10623 ( .A(fifo[1256]), .Y(n10659) );
  INVX1 U10624 ( .A(n10662), .Y(n10660) );
  INVX1 U10625 ( .A(n10660), .Y(n10661) );
  BUFX2 U10626 ( .A(fifo[1257]), .Y(n10662) );
  INVX1 U10627 ( .A(n10665), .Y(n10663) );
  INVX1 U10628 ( .A(n10663), .Y(n10664) );
  BUFX2 U10629 ( .A(fifo[1258]), .Y(n10665) );
  INVX1 U10630 ( .A(n10668), .Y(n10666) );
  INVX1 U10631 ( .A(n10666), .Y(n10667) );
  BUFX2 U10632 ( .A(fifo[1259]), .Y(n10668) );
  INVX1 U10633 ( .A(n10671), .Y(n10669) );
  INVX1 U10634 ( .A(n10669), .Y(n10670) );
  BUFX2 U10635 ( .A(fifo[1302]), .Y(n10671) );
  INVX1 U10636 ( .A(n10674), .Y(n10672) );
  INVX1 U10637 ( .A(n10672), .Y(n10673) );
  BUFX2 U10638 ( .A(fifo[1303]), .Y(n10674) );
  INVX1 U10639 ( .A(n10677), .Y(n10675) );
  INVX1 U10640 ( .A(n10675), .Y(n10676) );
  BUFX2 U10641 ( .A(fifo[1304]), .Y(n10677) );
  INVX1 U10642 ( .A(n10680), .Y(n10678) );
  INVX1 U10643 ( .A(n10678), .Y(n10679) );
  BUFX2 U10644 ( .A(fifo[1305]), .Y(n10680) );
  INVX1 U10645 ( .A(n10683), .Y(n10681) );
  INVX1 U10646 ( .A(n10681), .Y(n10682) );
  BUFX2 U10647 ( .A(fifo[1306]), .Y(n10683) );
  INVX1 U10648 ( .A(n10686), .Y(n10684) );
  INVX1 U10649 ( .A(n10684), .Y(n10685) );
  BUFX2 U10650 ( .A(fifo[1307]), .Y(n10686) );
  INVX1 U10651 ( .A(n10689), .Y(n10687) );
  INVX1 U10652 ( .A(n10687), .Y(n10688) );
  BUFX2 U10653 ( .A(fifo[1308]), .Y(n10689) );
  INVX1 U10654 ( .A(n10692), .Y(n10690) );
  INVX1 U10655 ( .A(n10690), .Y(n10691) );
  BUFX2 U10656 ( .A(fifo[1309]), .Y(n10692) );
  INVX1 U10657 ( .A(n10695), .Y(n10693) );
  INVX1 U10658 ( .A(n10693), .Y(n10694) );
  BUFX2 U10659 ( .A(fifo[1310]), .Y(n10695) );
  INVX1 U10660 ( .A(n10698), .Y(n10696) );
  INVX1 U10661 ( .A(n10696), .Y(n10697) );
  BUFX2 U10662 ( .A(fifo[1311]), .Y(n10698) );
  INVX1 U10663 ( .A(n10701), .Y(n10699) );
  INVX1 U10664 ( .A(n10699), .Y(n10700) );
  BUFX2 U10665 ( .A(fifo[1312]), .Y(n10701) );
  INVX1 U10666 ( .A(n10704), .Y(n10702) );
  INVX1 U10667 ( .A(n10702), .Y(n10703) );
  BUFX2 U10668 ( .A(fifo[1313]), .Y(n10704) );
  INVX1 U10669 ( .A(n10707), .Y(n10705) );
  INVX1 U10670 ( .A(n10705), .Y(n10706) );
  BUFX2 U10671 ( .A(fifo[1314]), .Y(n10707) );
  INVX1 U10672 ( .A(n10710), .Y(n10708) );
  INVX1 U10673 ( .A(n10708), .Y(n10709) );
  BUFX2 U10674 ( .A(fifo[1315]), .Y(n10710) );
  INVX1 U10675 ( .A(n10713), .Y(n10711) );
  INVX1 U10676 ( .A(n10711), .Y(n10712) );
  BUFX2 U10677 ( .A(fifo[1316]), .Y(n10713) );
  INVX1 U10678 ( .A(n10716), .Y(n10714) );
  INVX1 U10679 ( .A(n10714), .Y(n10715) );
  BUFX2 U10680 ( .A(fifo[1317]), .Y(n10716) );
  INVX1 U10681 ( .A(n10719), .Y(n10717) );
  INVX1 U10682 ( .A(n10717), .Y(n10718) );
  BUFX2 U10683 ( .A(fifo[1318]), .Y(n10719) );
  INVX1 U10684 ( .A(n10722), .Y(n10720) );
  INVX1 U10685 ( .A(n10720), .Y(n10721) );
  BUFX2 U10686 ( .A(fifo[1319]), .Y(n10722) );
  INVX1 U10687 ( .A(n10725), .Y(n10723) );
  INVX1 U10688 ( .A(n10723), .Y(n10724) );
  BUFX2 U10689 ( .A(fifo[1320]), .Y(n10725) );
  INVX1 U10690 ( .A(n10728), .Y(n10726) );
  INVX1 U10691 ( .A(n10726), .Y(n10727) );
  BUFX2 U10692 ( .A(fifo[1321]), .Y(n10728) );
  INVX1 U10693 ( .A(n10731), .Y(n10729) );
  INVX1 U10694 ( .A(n10729), .Y(n10730) );
  BUFX2 U10695 ( .A(fifo[1322]), .Y(n10731) );
  INVX1 U10696 ( .A(n10734), .Y(n10732) );
  INVX1 U10697 ( .A(n10732), .Y(n10733) );
  BUFX2 U10698 ( .A(fifo[1323]), .Y(n10734) );
  INVX1 U10699 ( .A(n10737), .Y(n10735) );
  INVX1 U10700 ( .A(n10735), .Y(n10736) );
  BUFX2 U10701 ( .A(fifo[1324]), .Y(n10737) );
  INVX1 U10702 ( .A(n10740), .Y(n10738) );
  INVX1 U10703 ( .A(n10738), .Y(n10739) );
  BUFX2 U10704 ( .A(fifo[1325]), .Y(n10740) );
  INVX1 U10705 ( .A(n10743), .Y(n10741) );
  INVX1 U10706 ( .A(n10741), .Y(n10742) );
  BUFX2 U10707 ( .A(fifo[1326]), .Y(n10743) );
  INVX1 U10708 ( .A(n10746), .Y(n10744) );
  INVX1 U10709 ( .A(n10744), .Y(n10745) );
  BUFX2 U10710 ( .A(fifo[1327]), .Y(n10746) );
  INVX1 U10711 ( .A(n10749), .Y(n10747) );
  INVX1 U10712 ( .A(n10747), .Y(n10748) );
  BUFX2 U10713 ( .A(fifo[1328]), .Y(n10749) );
  INVX1 U10714 ( .A(n10752), .Y(n10750) );
  INVX1 U10715 ( .A(n10750), .Y(n10751) );
  BUFX2 U10716 ( .A(fifo[1329]), .Y(n10752) );
  INVX1 U10717 ( .A(n10755), .Y(n10753) );
  INVX1 U10718 ( .A(n10753), .Y(n10754) );
  BUFX2 U10719 ( .A(fifo[1330]), .Y(n10755) );
  INVX1 U10720 ( .A(n10758), .Y(n10756) );
  INVX1 U10721 ( .A(n10756), .Y(n10757) );
  BUFX2 U10722 ( .A(fifo[1331]), .Y(n10758) );
  INVX1 U10723 ( .A(n10761), .Y(n10759) );
  INVX1 U10724 ( .A(n10759), .Y(n10760) );
  BUFX2 U10725 ( .A(fifo[1332]), .Y(n10761) );
  INVX1 U10726 ( .A(n10764), .Y(n10762) );
  INVX1 U10727 ( .A(n10762), .Y(n10763) );
  BUFX2 U10728 ( .A(fifo[1333]), .Y(n10764) );
  INVX1 U10729 ( .A(n10767), .Y(n10765) );
  INVX1 U10730 ( .A(n10765), .Y(n10766) );
  BUFX2 U10731 ( .A(fifo[1334]), .Y(n10767) );
  INVX1 U10732 ( .A(n10770), .Y(n10768) );
  INVX1 U10733 ( .A(n10768), .Y(n10769) );
  BUFX2 U10734 ( .A(fifo[1335]), .Y(n10770) );
  INVX1 U10735 ( .A(n10773), .Y(n10771) );
  INVX1 U10736 ( .A(n10771), .Y(n10772) );
  BUFX2 U10737 ( .A(fifo[1336]), .Y(n10773) );
  INVX1 U10738 ( .A(n10776), .Y(n10774) );
  INVX1 U10739 ( .A(n10774), .Y(n10775) );
  BUFX2 U10740 ( .A(fifo[1337]), .Y(n10776) );
  INVX1 U10741 ( .A(n10779), .Y(n10777) );
  INVX1 U10742 ( .A(n10777), .Y(n10778) );
  BUFX2 U10743 ( .A(fifo[1338]), .Y(n10779) );
  INVX1 U10744 ( .A(n10782), .Y(n10780) );
  INVX1 U10745 ( .A(n10780), .Y(n10781) );
  BUFX2 U10746 ( .A(fifo[1339]), .Y(n10782) );
  INVX1 U10747 ( .A(n10785), .Y(n10783) );
  INVX1 U10748 ( .A(n10783), .Y(n10784) );
  BUFX2 U10749 ( .A(fifo[1340]), .Y(n10785) );
  INVX1 U10750 ( .A(n10788), .Y(n10786) );
  INVX1 U10751 ( .A(n10786), .Y(n10787) );
  BUFX2 U10752 ( .A(fifo[1341]), .Y(n10788) );
  INVX1 U10753 ( .A(n10791), .Y(n10789) );
  INVX1 U10754 ( .A(n10789), .Y(n10790) );
  BUFX2 U10755 ( .A(fifo[1342]), .Y(n10791) );
  INVX1 U10756 ( .A(n10794), .Y(n10792) );
  INVX1 U10757 ( .A(n10792), .Y(n10793) );
  BUFX2 U10758 ( .A(fifo[1343]), .Y(n10794) );
  INVX1 U10759 ( .A(n8762), .Y(n10795) );
  INVX1 U10760 ( .A(n10795), .Y(n10796) );
  INVX1 U10761 ( .A(n8770), .Y(n10797) );
  INVX1 U10762 ( .A(n10797), .Y(n10798) );
  INVX1 U10763 ( .A(n8746), .Y(n10799) );
  INVX1 U10764 ( .A(n10799), .Y(n10800) );
  INVX1 U10765 ( .A(n8748), .Y(n10801) );
  INVX1 U10766 ( .A(n10801), .Y(n10802) );
  INVX1 U10767 ( .A(n10805), .Y(n10803) );
  INVX1 U10768 ( .A(n10803), .Y(n10804) );
  BUFX2 U10769 ( .A(fifo[0]), .Y(n10805) );
  INVX1 U10770 ( .A(n10808), .Y(n10806) );
  INVX1 U10771 ( .A(n10806), .Y(n10807) );
  BUFX2 U10772 ( .A(fifo[1]), .Y(n10808) );
  INVX1 U10773 ( .A(n10811), .Y(n10809) );
  INVX1 U10774 ( .A(n10809), .Y(n10810) );
  BUFX2 U10775 ( .A(fifo[2]), .Y(n10811) );
  INVX1 U10776 ( .A(n10814), .Y(n10812) );
  INVX1 U10777 ( .A(n10812), .Y(n10813) );
  BUFX2 U10778 ( .A(fifo[3]), .Y(n10814) );
  INVX1 U10779 ( .A(n10817), .Y(n10815) );
  INVX1 U10780 ( .A(n10815), .Y(n10816) );
  BUFX2 U10781 ( .A(fifo[4]), .Y(n10817) );
  INVX1 U10782 ( .A(n10820), .Y(n10818) );
  INVX1 U10783 ( .A(n10818), .Y(n10819) );
  BUFX2 U10784 ( .A(fifo[5]), .Y(n10820) );
  INVX1 U10785 ( .A(n10823), .Y(n10821) );
  INVX1 U10786 ( .A(n10821), .Y(n10822) );
  BUFX2 U10787 ( .A(fifo[6]), .Y(n10823) );
  INVX1 U10788 ( .A(n10826), .Y(n10824) );
  INVX1 U10789 ( .A(n10824), .Y(n10825) );
  BUFX2 U10790 ( .A(fifo[7]), .Y(n10826) );
  INVX1 U10791 ( .A(n10829), .Y(n10827) );
  INVX1 U10792 ( .A(n10827), .Y(n10828) );
  BUFX2 U10793 ( .A(fifo[8]), .Y(n10829) );
  INVX1 U10794 ( .A(n10832), .Y(n10830) );
  INVX1 U10795 ( .A(n10830), .Y(n10831) );
  BUFX2 U10796 ( .A(fifo[9]), .Y(n10832) );
  INVX1 U10797 ( .A(n10835), .Y(n10833) );
  INVX1 U10798 ( .A(n10833), .Y(n10834) );
  BUFX2 U10799 ( .A(fifo[10]), .Y(n10835) );
  INVX1 U10800 ( .A(n10838), .Y(n10836) );
  INVX1 U10801 ( .A(n10836), .Y(n10837) );
  BUFX2 U10802 ( .A(fifo[11]), .Y(n10838) );
  INVX1 U10803 ( .A(n10841), .Y(n10839) );
  INVX1 U10804 ( .A(n10839), .Y(n10840) );
  BUFX2 U10805 ( .A(fifo[12]), .Y(n10841) );
  INVX1 U10806 ( .A(n10844), .Y(n10842) );
  INVX1 U10807 ( .A(n10842), .Y(n10843) );
  BUFX2 U10808 ( .A(fifo[13]), .Y(n10844) );
  INVX1 U10809 ( .A(n10847), .Y(n10845) );
  INVX1 U10810 ( .A(n10845), .Y(n10846) );
  BUFX2 U10811 ( .A(fifo[14]), .Y(n10847) );
  INVX1 U10812 ( .A(n10850), .Y(n10848) );
  INVX1 U10813 ( .A(n10848), .Y(n10849) );
  BUFX2 U10814 ( .A(fifo[15]), .Y(n10850) );
  INVX1 U10815 ( .A(n10853), .Y(n10851) );
  INVX1 U10816 ( .A(n10851), .Y(n10852) );
  BUFX2 U10817 ( .A(fifo[16]), .Y(n10853) );
  INVX1 U10818 ( .A(n10856), .Y(n10854) );
  INVX1 U10819 ( .A(n10854), .Y(n10855) );
  BUFX2 U10820 ( .A(fifo[17]), .Y(n10856) );
  INVX1 U10821 ( .A(n10859), .Y(n10857) );
  INVX1 U10822 ( .A(n10857), .Y(n10858) );
  BUFX2 U10823 ( .A(fifo[18]), .Y(n10859) );
  INVX1 U10824 ( .A(n10862), .Y(n10860) );
  INVX1 U10825 ( .A(n10860), .Y(n10861) );
  BUFX2 U10826 ( .A(fifo[19]), .Y(n10862) );
  INVX1 U10827 ( .A(n10865), .Y(n10863) );
  INVX1 U10828 ( .A(n10863), .Y(n10864) );
  BUFX2 U10829 ( .A(fifo[20]), .Y(n10865) );
  INVX1 U10830 ( .A(n10868), .Y(n10866) );
  INVX1 U10831 ( .A(n10866), .Y(n10867) );
  BUFX2 U10832 ( .A(fifo[21]), .Y(n10868) );
  INVX1 U10833 ( .A(n10871), .Y(n10869) );
  INVX1 U10834 ( .A(n10869), .Y(n10870) );
  BUFX2 U10835 ( .A(fifo[22]), .Y(n10871) );
  INVX1 U10836 ( .A(n10874), .Y(n10872) );
  INVX1 U10837 ( .A(n10872), .Y(n10873) );
  BUFX2 U10838 ( .A(fifo[23]), .Y(n10874) );
  INVX1 U10839 ( .A(n10877), .Y(n10875) );
  INVX1 U10840 ( .A(n10875), .Y(n10876) );
  BUFX2 U10841 ( .A(fifo[24]), .Y(n10877) );
  INVX1 U10842 ( .A(n10880), .Y(n10878) );
  INVX1 U10843 ( .A(n10878), .Y(n10879) );
  BUFX2 U10844 ( .A(fifo[25]), .Y(n10880) );
  INVX1 U10845 ( .A(n10883), .Y(n10881) );
  INVX1 U10846 ( .A(n10881), .Y(n10882) );
  BUFX2 U10847 ( .A(fifo[26]), .Y(n10883) );
  INVX1 U10848 ( .A(n10886), .Y(n10884) );
  INVX1 U10849 ( .A(n10884), .Y(n10885) );
  BUFX2 U10850 ( .A(fifo[27]), .Y(n10886) );
  INVX1 U10851 ( .A(n10889), .Y(n10887) );
  INVX1 U10852 ( .A(n10887), .Y(n10888) );
  BUFX2 U10853 ( .A(fifo[28]), .Y(n10889) );
  INVX1 U10854 ( .A(n10892), .Y(n10890) );
  INVX1 U10855 ( .A(n10890), .Y(n10891) );
  BUFX2 U10856 ( .A(fifo[29]), .Y(n10892) );
  INVX1 U10857 ( .A(n10895), .Y(n10893) );
  INVX1 U10858 ( .A(n10893), .Y(n10894) );
  BUFX2 U10859 ( .A(fifo[30]), .Y(n10895) );
  INVX1 U10860 ( .A(n10898), .Y(n10896) );
  INVX1 U10861 ( .A(n10896), .Y(n10897) );
  BUFX2 U10862 ( .A(fifo[31]), .Y(n10898) );
  INVX1 U10863 ( .A(n10901), .Y(n10899) );
  INVX1 U10864 ( .A(n10899), .Y(n10900) );
  BUFX2 U10865 ( .A(fifo[32]), .Y(n10901) );
  INVX1 U10866 ( .A(n10904), .Y(n10902) );
  INVX1 U10867 ( .A(n10902), .Y(n10903) );
  BUFX2 U10868 ( .A(fifo[33]), .Y(n10904) );
  INVX1 U10869 ( .A(n10907), .Y(n10905) );
  INVX1 U10870 ( .A(n10905), .Y(n10906) );
  BUFX2 U10871 ( .A(fifo[34]), .Y(n10907) );
  INVX1 U10872 ( .A(n10910), .Y(n10908) );
  INVX1 U10873 ( .A(n10908), .Y(n10909) );
  BUFX2 U10874 ( .A(fifo[35]), .Y(n10910) );
  INVX1 U10875 ( .A(n10913), .Y(n10911) );
  INVX1 U10876 ( .A(n10911), .Y(n10912) );
  BUFX2 U10877 ( .A(fifo[36]), .Y(n10913) );
  INVX1 U10878 ( .A(n10916), .Y(n10914) );
  INVX1 U10879 ( .A(n10914), .Y(n10915) );
  BUFX2 U10880 ( .A(fifo[37]), .Y(n10916) );
  INVX1 U10881 ( .A(n10919), .Y(n10917) );
  INVX1 U10882 ( .A(n10917), .Y(n10918) );
  BUFX2 U10883 ( .A(fifo[38]), .Y(n10919) );
  INVX1 U10884 ( .A(n10922), .Y(n10920) );
  INVX1 U10885 ( .A(n10920), .Y(n10921) );
  BUFX2 U10886 ( .A(fifo[39]), .Y(n10922) );
  INVX1 U10887 ( .A(n10925), .Y(n10923) );
  INVX1 U10888 ( .A(n10923), .Y(n10924) );
  BUFX2 U10889 ( .A(fifo[40]), .Y(n10925) );
  INVX1 U10890 ( .A(n10928), .Y(n10926) );
  INVX1 U10891 ( .A(n10926), .Y(n10927) );
  BUFX2 U10892 ( .A(fifo[41]), .Y(n10928) );
  INVX1 U10893 ( .A(n10931), .Y(n10929) );
  INVX1 U10894 ( .A(n10929), .Y(n10930) );
  BUFX2 U10895 ( .A(fifo[84]), .Y(n10931) );
  INVX1 U10896 ( .A(n10934), .Y(n10932) );
  INVX1 U10897 ( .A(n10932), .Y(n10933) );
  BUFX2 U10898 ( .A(fifo[85]), .Y(n10934) );
  INVX1 U10899 ( .A(n10937), .Y(n10935) );
  INVX1 U10900 ( .A(n10935), .Y(n10936) );
  BUFX2 U10901 ( .A(fifo[86]), .Y(n10937) );
  INVX1 U10902 ( .A(n10940), .Y(n10938) );
  INVX1 U10903 ( .A(n10938), .Y(n10939) );
  BUFX2 U10904 ( .A(fifo[87]), .Y(n10940) );
  INVX1 U10905 ( .A(n10943), .Y(n10941) );
  INVX1 U10906 ( .A(n10941), .Y(n10942) );
  BUFX2 U10907 ( .A(fifo[88]), .Y(n10943) );
  INVX1 U10908 ( .A(n10946), .Y(n10944) );
  INVX1 U10909 ( .A(n10944), .Y(n10945) );
  BUFX2 U10910 ( .A(fifo[89]), .Y(n10946) );
  INVX1 U10911 ( .A(n10949), .Y(n10947) );
  INVX1 U10912 ( .A(n10947), .Y(n10948) );
  BUFX2 U10913 ( .A(fifo[90]), .Y(n10949) );
  INVX1 U10914 ( .A(n10952), .Y(n10950) );
  INVX1 U10915 ( .A(n10950), .Y(n10951) );
  BUFX2 U10916 ( .A(fifo[91]), .Y(n10952) );
  INVX1 U10917 ( .A(n10955), .Y(n10953) );
  INVX1 U10918 ( .A(n10953), .Y(n10954) );
  BUFX2 U10919 ( .A(fifo[92]), .Y(n10955) );
  INVX1 U10920 ( .A(n10958), .Y(n10956) );
  INVX1 U10921 ( .A(n10956), .Y(n10957) );
  BUFX2 U10922 ( .A(fifo[93]), .Y(n10958) );
  INVX1 U10923 ( .A(n10961), .Y(n10959) );
  INVX1 U10924 ( .A(n10959), .Y(n10960) );
  BUFX2 U10925 ( .A(fifo[94]), .Y(n10961) );
  INVX1 U10926 ( .A(n10964), .Y(n10962) );
  INVX1 U10927 ( .A(n10962), .Y(n10963) );
  BUFX2 U10928 ( .A(fifo[95]), .Y(n10964) );
  INVX1 U10929 ( .A(n10967), .Y(n10965) );
  INVX1 U10930 ( .A(n10965), .Y(n10966) );
  BUFX2 U10931 ( .A(fifo[96]), .Y(n10967) );
  INVX1 U10932 ( .A(n10970), .Y(n10968) );
  INVX1 U10933 ( .A(n10968), .Y(n10969) );
  BUFX2 U10934 ( .A(fifo[97]), .Y(n10970) );
  INVX1 U10935 ( .A(n10973), .Y(n10971) );
  INVX1 U10936 ( .A(n10971), .Y(n10972) );
  BUFX2 U10937 ( .A(fifo[98]), .Y(n10973) );
  INVX1 U10938 ( .A(n10976), .Y(n10974) );
  INVX1 U10939 ( .A(n10974), .Y(n10975) );
  BUFX2 U10940 ( .A(fifo[99]), .Y(n10976) );
  INVX1 U10941 ( .A(n10979), .Y(n10977) );
  INVX1 U10942 ( .A(n10977), .Y(n10978) );
  BUFX2 U10943 ( .A(fifo[100]), .Y(n10979) );
  INVX1 U10944 ( .A(n10982), .Y(n10980) );
  INVX1 U10945 ( .A(n10980), .Y(n10981) );
  BUFX2 U10946 ( .A(fifo[101]), .Y(n10982) );
  INVX1 U10947 ( .A(n10985), .Y(n10983) );
  INVX1 U10948 ( .A(n10983), .Y(n10984) );
  BUFX2 U10949 ( .A(fifo[102]), .Y(n10985) );
  INVX1 U10950 ( .A(n10988), .Y(n10986) );
  INVX1 U10951 ( .A(n10986), .Y(n10987) );
  BUFX2 U10952 ( .A(fifo[103]), .Y(n10988) );
  INVX1 U10953 ( .A(n10991), .Y(n10989) );
  INVX1 U10954 ( .A(n10989), .Y(n10990) );
  BUFX2 U10955 ( .A(fifo[104]), .Y(n10991) );
  INVX1 U10956 ( .A(n10994), .Y(n10992) );
  INVX1 U10957 ( .A(n10992), .Y(n10993) );
  BUFX2 U10958 ( .A(fifo[105]), .Y(n10994) );
  INVX1 U10959 ( .A(n10997), .Y(n10995) );
  INVX1 U10960 ( .A(n10995), .Y(n10996) );
  BUFX2 U10961 ( .A(fifo[106]), .Y(n10997) );
  INVX1 U10962 ( .A(n11000), .Y(n10998) );
  INVX1 U10963 ( .A(n10998), .Y(n10999) );
  BUFX2 U10964 ( .A(fifo[107]), .Y(n11000) );
  INVX1 U10965 ( .A(n11003), .Y(n11001) );
  INVX1 U10966 ( .A(n11001), .Y(n11002) );
  BUFX2 U10967 ( .A(fifo[108]), .Y(n11003) );
  INVX1 U10968 ( .A(n11006), .Y(n11004) );
  INVX1 U10969 ( .A(n11004), .Y(n11005) );
  BUFX2 U10970 ( .A(fifo[109]), .Y(n11006) );
  INVX1 U10971 ( .A(n11009), .Y(n11007) );
  INVX1 U10972 ( .A(n11007), .Y(n11008) );
  BUFX2 U10973 ( .A(fifo[110]), .Y(n11009) );
  INVX1 U10974 ( .A(n11012), .Y(n11010) );
  INVX1 U10975 ( .A(n11010), .Y(n11011) );
  BUFX2 U10976 ( .A(fifo[111]), .Y(n11012) );
  INVX1 U10977 ( .A(n11015), .Y(n11013) );
  INVX1 U10978 ( .A(n11013), .Y(n11014) );
  BUFX2 U10979 ( .A(fifo[112]), .Y(n11015) );
  INVX1 U10980 ( .A(n11018), .Y(n11016) );
  INVX1 U10981 ( .A(n11016), .Y(n11017) );
  BUFX2 U10982 ( .A(fifo[113]), .Y(n11018) );
  INVX1 U10983 ( .A(n11021), .Y(n11019) );
  INVX1 U10984 ( .A(n11019), .Y(n11020) );
  BUFX2 U10985 ( .A(fifo[114]), .Y(n11021) );
  INVX1 U10986 ( .A(n11024), .Y(n11022) );
  INVX1 U10987 ( .A(n11022), .Y(n11023) );
  BUFX2 U10988 ( .A(fifo[115]), .Y(n11024) );
  INVX1 U10989 ( .A(n11027), .Y(n11025) );
  INVX1 U10990 ( .A(n11025), .Y(n11026) );
  BUFX2 U10991 ( .A(fifo[116]), .Y(n11027) );
  INVX1 U10992 ( .A(n11030), .Y(n11028) );
  INVX1 U10993 ( .A(n11028), .Y(n11029) );
  BUFX2 U10994 ( .A(fifo[117]), .Y(n11030) );
  INVX1 U10995 ( .A(n11033), .Y(n11031) );
  INVX1 U10996 ( .A(n11031), .Y(n11032) );
  BUFX2 U10997 ( .A(fifo[118]), .Y(n11033) );
  INVX1 U10998 ( .A(n11036), .Y(n11034) );
  INVX1 U10999 ( .A(n11034), .Y(n11035) );
  BUFX2 U11000 ( .A(fifo[119]), .Y(n11036) );
  INVX1 U11001 ( .A(n11039), .Y(n11037) );
  INVX1 U11002 ( .A(n11037), .Y(n11038) );
  BUFX2 U11003 ( .A(fifo[120]), .Y(n11039) );
  INVX1 U11004 ( .A(n11042), .Y(n11040) );
  INVX1 U11005 ( .A(n11040), .Y(n11041) );
  BUFX2 U11006 ( .A(fifo[121]), .Y(n11042) );
  INVX1 U11007 ( .A(n11045), .Y(n11043) );
  INVX1 U11008 ( .A(n11043), .Y(n11044) );
  BUFX2 U11009 ( .A(fifo[122]), .Y(n11045) );
  INVX1 U11010 ( .A(n11048), .Y(n11046) );
  INVX1 U11011 ( .A(n11046), .Y(n11047) );
  BUFX2 U11012 ( .A(fifo[123]), .Y(n11048) );
  INVX1 U11013 ( .A(n11051), .Y(n11049) );
  INVX1 U11014 ( .A(n11049), .Y(n11050) );
  BUFX2 U11015 ( .A(fifo[124]), .Y(n11051) );
  INVX1 U11016 ( .A(n11054), .Y(n11052) );
  INVX1 U11017 ( .A(n11052), .Y(n11053) );
  BUFX2 U11018 ( .A(fifo[125]), .Y(n11054) );
  INVX1 U11019 ( .A(n11057), .Y(n11055) );
  INVX1 U11020 ( .A(n11055), .Y(n11056) );
  BUFX2 U11021 ( .A(fifo[168]), .Y(n11057) );
  INVX1 U11022 ( .A(n11060), .Y(n11058) );
  INVX1 U11023 ( .A(n11058), .Y(n11059) );
  BUFX2 U11024 ( .A(fifo[169]), .Y(n11060) );
  INVX1 U11025 ( .A(n11063), .Y(n11061) );
  INVX1 U11026 ( .A(n11061), .Y(n11062) );
  BUFX2 U11027 ( .A(fifo[170]), .Y(n11063) );
  INVX1 U11028 ( .A(n11066), .Y(n11064) );
  INVX1 U11029 ( .A(n11064), .Y(n11065) );
  BUFX2 U11030 ( .A(fifo[171]), .Y(n11066) );
  INVX1 U11031 ( .A(n11069), .Y(n11067) );
  INVX1 U11032 ( .A(n11067), .Y(n11068) );
  BUFX2 U11033 ( .A(fifo[172]), .Y(n11069) );
  INVX1 U11034 ( .A(n11072), .Y(n11070) );
  INVX1 U11035 ( .A(n11070), .Y(n11071) );
  BUFX2 U11036 ( .A(fifo[173]), .Y(n11072) );
  INVX1 U11037 ( .A(n11075), .Y(n11073) );
  INVX1 U11038 ( .A(n11073), .Y(n11074) );
  BUFX2 U11039 ( .A(fifo[174]), .Y(n11075) );
  INVX1 U11040 ( .A(n11078), .Y(n11076) );
  INVX1 U11041 ( .A(n11076), .Y(n11077) );
  BUFX2 U11042 ( .A(fifo[175]), .Y(n11078) );
  INVX1 U11043 ( .A(n11081), .Y(n11079) );
  INVX1 U11044 ( .A(n11079), .Y(n11080) );
  BUFX2 U11045 ( .A(fifo[176]), .Y(n11081) );
  INVX1 U11046 ( .A(n11084), .Y(n11082) );
  INVX1 U11047 ( .A(n11082), .Y(n11083) );
  BUFX2 U11048 ( .A(fifo[177]), .Y(n11084) );
  INVX1 U11049 ( .A(n11087), .Y(n11085) );
  INVX1 U11050 ( .A(n11085), .Y(n11086) );
  BUFX2 U11051 ( .A(fifo[178]), .Y(n11087) );
  INVX1 U11052 ( .A(n11090), .Y(n11088) );
  INVX1 U11053 ( .A(n11088), .Y(n11089) );
  BUFX2 U11054 ( .A(fifo[179]), .Y(n11090) );
  INVX1 U11055 ( .A(n11093), .Y(n11091) );
  INVX1 U11056 ( .A(n11091), .Y(n11092) );
  BUFX2 U11057 ( .A(fifo[180]), .Y(n11093) );
  INVX1 U11058 ( .A(n11096), .Y(n11094) );
  INVX1 U11059 ( .A(n11094), .Y(n11095) );
  BUFX2 U11060 ( .A(fifo[181]), .Y(n11096) );
  INVX1 U11061 ( .A(n11099), .Y(n11097) );
  INVX1 U11062 ( .A(n11097), .Y(n11098) );
  BUFX2 U11063 ( .A(fifo[182]), .Y(n11099) );
  INVX1 U11064 ( .A(n11102), .Y(n11100) );
  INVX1 U11065 ( .A(n11100), .Y(n11101) );
  BUFX2 U11066 ( .A(fifo[183]), .Y(n11102) );
  INVX1 U11067 ( .A(n11105), .Y(n11103) );
  INVX1 U11068 ( .A(n11103), .Y(n11104) );
  BUFX2 U11069 ( .A(fifo[184]), .Y(n11105) );
  INVX1 U11070 ( .A(n11108), .Y(n11106) );
  INVX1 U11071 ( .A(n11106), .Y(n11107) );
  BUFX2 U11072 ( .A(fifo[185]), .Y(n11108) );
  INVX1 U11073 ( .A(n11111), .Y(n11109) );
  INVX1 U11074 ( .A(n11109), .Y(n11110) );
  BUFX2 U11075 ( .A(fifo[186]), .Y(n11111) );
  INVX1 U11076 ( .A(n11114), .Y(n11112) );
  INVX1 U11077 ( .A(n11112), .Y(n11113) );
  BUFX2 U11078 ( .A(fifo[187]), .Y(n11114) );
  INVX1 U11079 ( .A(n11117), .Y(n11115) );
  INVX1 U11080 ( .A(n11115), .Y(n11116) );
  BUFX2 U11081 ( .A(fifo[188]), .Y(n11117) );
  INVX1 U11082 ( .A(n11120), .Y(n11118) );
  INVX1 U11083 ( .A(n11118), .Y(n11119) );
  BUFX2 U11084 ( .A(fifo[189]), .Y(n11120) );
  INVX1 U11085 ( .A(n11123), .Y(n11121) );
  INVX1 U11086 ( .A(n11121), .Y(n11122) );
  BUFX2 U11087 ( .A(fifo[190]), .Y(n11123) );
  INVX1 U11088 ( .A(n11126), .Y(n11124) );
  INVX1 U11089 ( .A(n11124), .Y(n11125) );
  BUFX2 U11090 ( .A(fifo[191]), .Y(n11126) );
  INVX1 U11091 ( .A(n11129), .Y(n11127) );
  INVX1 U11092 ( .A(n11127), .Y(n11128) );
  BUFX2 U11093 ( .A(fifo[192]), .Y(n11129) );
  INVX1 U11094 ( .A(n11132), .Y(n11130) );
  INVX1 U11095 ( .A(n11130), .Y(n11131) );
  BUFX2 U11096 ( .A(fifo[193]), .Y(n11132) );
  INVX1 U11097 ( .A(n11135), .Y(n11133) );
  INVX1 U11098 ( .A(n11133), .Y(n11134) );
  BUFX2 U11099 ( .A(fifo[194]), .Y(n11135) );
  INVX1 U11100 ( .A(n11138), .Y(n11136) );
  INVX1 U11101 ( .A(n11136), .Y(n11137) );
  BUFX2 U11102 ( .A(fifo[195]), .Y(n11138) );
  INVX1 U11103 ( .A(n11141), .Y(n11139) );
  INVX1 U11104 ( .A(n11139), .Y(n11140) );
  BUFX2 U11105 ( .A(fifo[196]), .Y(n11141) );
  INVX1 U11106 ( .A(n11144), .Y(n11142) );
  INVX1 U11107 ( .A(n11142), .Y(n11143) );
  BUFX2 U11108 ( .A(fifo[197]), .Y(n11144) );
  INVX1 U11109 ( .A(n11147), .Y(n11145) );
  INVX1 U11110 ( .A(n11145), .Y(n11146) );
  BUFX2 U11111 ( .A(fifo[198]), .Y(n11147) );
  INVX1 U11112 ( .A(n11150), .Y(n11148) );
  INVX1 U11113 ( .A(n11148), .Y(n11149) );
  BUFX2 U11114 ( .A(fifo[199]), .Y(n11150) );
  INVX1 U11115 ( .A(n11153), .Y(n11151) );
  INVX1 U11116 ( .A(n11151), .Y(n11152) );
  BUFX2 U11117 ( .A(fifo[200]), .Y(n11153) );
  INVX1 U11118 ( .A(n11156), .Y(n11154) );
  INVX1 U11119 ( .A(n11154), .Y(n11155) );
  BUFX2 U11120 ( .A(fifo[201]), .Y(n11156) );
  INVX1 U11121 ( .A(n11159), .Y(n11157) );
  INVX1 U11122 ( .A(n11157), .Y(n11158) );
  BUFX2 U11123 ( .A(fifo[202]), .Y(n11159) );
  INVX1 U11124 ( .A(n11162), .Y(n11160) );
  INVX1 U11125 ( .A(n11160), .Y(n11161) );
  BUFX2 U11126 ( .A(fifo[203]), .Y(n11162) );
  INVX1 U11127 ( .A(n11165), .Y(n11163) );
  INVX1 U11128 ( .A(n11163), .Y(n11164) );
  BUFX2 U11129 ( .A(fifo[204]), .Y(n11165) );
  INVX1 U11130 ( .A(n11168), .Y(n11166) );
  INVX1 U11131 ( .A(n11166), .Y(n11167) );
  BUFX2 U11132 ( .A(fifo[205]), .Y(n11168) );
  INVX1 U11133 ( .A(n11171), .Y(n11169) );
  INVX1 U11134 ( .A(n11169), .Y(n11170) );
  BUFX2 U11135 ( .A(fifo[206]), .Y(n11171) );
  INVX1 U11136 ( .A(n11174), .Y(n11172) );
  INVX1 U11137 ( .A(n11172), .Y(n11173) );
  BUFX2 U11138 ( .A(fifo[207]), .Y(n11174) );
  INVX1 U11139 ( .A(n11177), .Y(n11175) );
  INVX1 U11140 ( .A(n11175), .Y(n11176) );
  BUFX2 U11141 ( .A(fifo[208]), .Y(n11177) );
  INVX1 U11142 ( .A(n11180), .Y(n11178) );
  INVX1 U11143 ( .A(n11178), .Y(n11179) );
  BUFX2 U11144 ( .A(fifo[209]), .Y(n11180) );
  INVX1 U11145 ( .A(n11183), .Y(n11181) );
  INVX1 U11146 ( .A(n11181), .Y(n11182) );
  BUFX2 U11147 ( .A(fifo[252]), .Y(n11183) );
  INVX1 U11148 ( .A(n11186), .Y(n11184) );
  INVX1 U11149 ( .A(n11184), .Y(n11185) );
  BUFX2 U11150 ( .A(fifo[253]), .Y(n11186) );
  INVX1 U11151 ( .A(n11189), .Y(n11187) );
  INVX1 U11152 ( .A(n11187), .Y(n11188) );
  BUFX2 U11153 ( .A(fifo[254]), .Y(n11189) );
  INVX1 U11154 ( .A(n11192), .Y(n11190) );
  INVX1 U11155 ( .A(n11190), .Y(n11191) );
  BUFX2 U11156 ( .A(fifo[255]), .Y(n11192) );
  INVX1 U11157 ( .A(n11195), .Y(n11193) );
  INVX1 U11158 ( .A(n11193), .Y(n11194) );
  BUFX2 U11159 ( .A(fifo[256]), .Y(n11195) );
  INVX1 U11160 ( .A(n11198), .Y(n11196) );
  INVX1 U11161 ( .A(n11196), .Y(n11197) );
  BUFX2 U11162 ( .A(fifo[257]), .Y(n11198) );
  INVX1 U11163 ( .A(n11201), .Y(n11199) );
  INVX1 U11164 ( .A(n11199), .Y(n11200) );
  BUFX2 U11165 ( .A(fifo[258]), .Y(n11201) );
  INVX1 U11166 ( .A(n11204), .Y(n11202) );
  INVX1 U11167 ( .A(n11202), .Y(n11203) );
  BUFX2 U11168 ( .A(fifo[259]), .Y(n11204) );
  INVX1 U11169 ( .A(n11207), .Y(n11205) );
  INVX1 U11170 ( .A(n11205), .Y(n11206) );
  BUFX2 U11171 ( .A(fifo[260]), .Y(n11207) );
  INVX1 U11172 ( .A(n11210), .Y(n11208) );
  INVX1 U11173 ( .A(n11208), .Y(n11209) );
  BUFX2 U11174 ( .A(fifo[261]), .Y(n11210) );
  INVX1 U11175 ( .A(n11213), .Y(n11211) );
  INVX1 U11176 ( .A(n11211), .Y(n11212) );
  BUFX2 U11177 ( .A(fifo[262]), .Y(n11213) );
  INVX1 U11178 ( .A(n11216), .Y(n11214) );
  INVX1 U11179 ( .A(n11214), .Y(n11215) );
  BUFX2 U11180 ( .A(fifo[263]), .Y(n11216) );
  INVX1 U11181 ( .A(n11219), .Y(n11217) );
  INVX1 U11182 ( .A(n11217), .Y(n11218) );
  BUFX2 U11183 ( .A(fifo[264]), .Y(n11219) );
  INVX1 U11184 ( .A(n11222), .Y(n11220) );
  INVX1 U11185 ( .A(n11220), .Y(n11221) );
  BUFX2 U11186 ( .A(fifo[265]), .Y(n11222) );
  INVX1 U11187 ( .A(n11225), .Y(n11223) );
  INVX1 U11188 ( .A(n11223), .Y(n11224) );
  BUFX2 U11189 ( .A(fifo[266]), .Y(n11225) );
  INVX1 U11190 ( .A(n11228), .Y(n11226) );
  INVX1 U11191 ( .A(n11226), .Y(n11227) );
  BUFX2 U11192 ( .A(fifo[267]), .Y(n11228) );
  INVX1 U11193 ( .A(n11231), .Y(n11229) );
  INVX1 U11194 ( .A(n11229), .Y(n11230) );
  BUFX2 U11195 ( .A(fifo[268]), .Y(n11231) );
  INVX1 U11196 ( .A(n11234), .Y(n11232) );
  INVX1 U11197 ( .A(n11232), .Y(n11233) );
  BUFX2 U11198 ( .A(fifo[269]), .Y(n11234) );
  INVX1 U11199 ( .A(n11237), .Y(n11235) );
  INVX1 U11200 ( .A(n11235), .Y(n11236) );
  BUFX2 U11201 ( .A(fifo[270]), .Y(n11237) );
  INVX1 U11202 ( .A(n11240), .Y(n11238) );
  INVX1 U11203 ( .A(n11238), .Y(n11239) );
  BUFX2 U11204 ( .A(fifo[271]), .Y(n11240) );
  INVX1 U11205 ( .A(n11243), .Y(n11241) );
  INVX1 U11206 ( .A(n11241), .Y(n11242) );
  BUFX2 U11207 ( .A(fifo[272]), .Y(n11243) );
  INVX1 U11208 ( .A(n11246), .Y(n11244) );
  INVX1 U11209 ( .A(n11244), .Y(n11245) );
  BUFX2 U11210 ( .A(fifo[273]), .Y(n11246) );
  INVX1 U11211 ( .A(n11249), .Y(n11247) );
  INVX1 U11212 ( .A(n11247), .Y(n11248) );
  BUFX2 U11213 ( .A(fifo[274]), .Y(n11249) );
  INVX1 U11214 ( .A(n11252), .Y(n11250) );
  INVX1 U11215 ( .A(n11250), .Y(n11251) );
  BUFX2 U11216 ( .A(fifo[275]), .Y(n11252) );
  INVX1 U11217 ( .A(n11255), .Y(n11253) );
  INVX1 U11218 ( .A(n11253), .Y(n11254) );
  BUFX2 U11219 ( .A(fifo[276]), .Y(n11255) );
  INVX1 U11220 ( .A(n11258), .Y(n11256) );
  INVX1 U11221 ( .A(n11256), .Y(n11257) );
  BUFX2 U11222 ( .A(fifo[277]), .Y(n11258) );
  INVX1 U11223 ( .A(n11261), .Y(n11259) );
  INVX1 U11224 ( .A(n11259), .Y(n11260) );
  BUFX2 U11225 ( .A(fifo[278]), .Y(n11261) );
  INVX1 U11226 ( .A(n11264), .Y(n11262) );
  INVX1 U11227 ( .A(n11262), .Y(n11263) );
  BUFX2 U11228 ( .A(fifo[279]), .Y(n11264) );
  INVX1 U11229 ( .A(n11267), .Y(n11265) );
  INVX1 U11230 ( .A(n11265), .Y(n11266) );
  BUFX2 U11231 ( .A(fifo[280]), .Y(n11267) );
  INVX1 U11232 ( .A(n11270), .Y(n11268) );
  INVX1 U11233 ( .A(n11268), .Y(n11269) );
  BUFX2 U11234 ( .A(fifo[281]), .Y(n11270) );
  INVX1 U11235 ( .A(n11273), .Y(n11271) );
  INVX1 U11236 ( .A(n11271), .Y(n11272) );
  BUFX2 U11237 ( .A(fifo[282]), .Y(n11273) );
  INVX1 U11238 ( .A(n11276), .Y(n11274) );
  INVX1 U11239 ( .A(n11274), .Y(n11275) );
  BUFX2 U11240 ( .A(fifo[283]), .Y(n11276) );
  INVX1 U11241 ( .A(n11279), .Y(n11277) );
  INVX1 U11242 ( .A(n11277), .Y(n11278) );
  BUFX2 U11243 ( .A(fifo[284]), .Y(n11279) );
  INVX1 U11244 ( .A(n11282), .Y(n11280) );
  INVX1 U11245 ( .A(n11280), .Y(n11281) );
  BUFX2 U11246 ( .A(fifo[285]), .Y(n11282) );
  INVX1 U11247 ( .A(n11285), .Y(n11283) );
  INVX1 U11248 ( .A(n11283), .Y(n11284) );
  BUFX2 U11249 ( .A(fifo[286]), .Y(n11285) );
  INVX1 U11250 ( .A(n11288), .Y(n11286) );
  INVX1 U11251 ( .A(n11286), .Y(n11287) );
  BUFX2 U11252 ( .A(fifo[287]), .Y(n11288) );
  INVX1 U11253 ( .A(n11291), .Y(n11289) );
  INVX1 U11254 ( .A(n11289), .Y(n11290) );
  BUFX2 U11255 ( .A(fifo[288]), .Y(n11291) );
  INVX1 U11256 ( .A(n11294), .Y(n11292) );
  INVX1 U11257 ( .A(n11292), .Y(n11293) );
  BUFX2 U11258 ( .A(fifo[289]), .Y(n11294) );
  INVX1 U11259 ( .A(n11297), .Y(n11295) );
  INVX1 U11260 ( .A(n11295), .Y(n11296) );
  BUFX2 U11261 ( .A(fifo[290]), .Y(n11297) );
  INVX1 U11262 ( .A(n11300), .Y(n11298) );
  INVX1 U11263 ( .A(n11298), .Y(n11299) );
  BUFX2 U11264 ( .A(fifo[291]), .Y(n11300) );
  INVX1 U11265 ( .A(n11303), .Y(n11301) );
  INVX1 U11266 ( .A(n11301), .Y(n11302) );
  BUFX2 U11267 ( .A(fifo[292]), .Y(n11303) );
  INVX1 U11268 ( .A(n11306), .Y(n11304) );
  INVX1 U11269 ( .A(n11304), .Y(n11305) );
  BUFX2 U11270 ( .A(fifo[293]), .Y(n11306) );
  INVX1 U11271 ( .A(n11309), .Y(n11307) );
  INVX1 U11272 ( .A(n11307), .Y(n11308) );
  BUFX2 U11273 ( .A(fifo[336]), .Y(n11309) );
  INVX1 U11274 ( .A(n11312), .Y(n11310) );
  INVX1 U11275 ( .A(n11310), .Y(n11311) );
  BUFX2 U11276 ( .A(fifo[337]), .Y(n11312) );
  INVX1 U11277 ( .A(n11315), .Y(n11313) );
  INVX1 U11278 ( .A(n11313), .Y(n11314) );
  BUFX2 U11279 ( .A(fifo[338]), .Y(n11315) );
  INVX1 U11280 ( .A(n11318), .Y(n11316) );
  INVX1 U11281 ( .A(n11316), .Y(n11317) );
  BUFX2 U11282 ( .A(fifo[339]), .Y(n11318) );
  INVX1 U11283 ( .A(n11321), .Y(n11319) );
  INVX1 U11284 ( .A(n11319), .Y(n11320) );
  BUFX2 U11285 ( .A(fifo[340]), .Y(n11321) );
  INVX1 U11286 ( .A(n11324), .Y(n11322) );
  INVX1 U11287 ( .A(n11322), .Y(n11323) );
  BUFX2 U11288 ( .A(fifo[341]), .Y(n11324) );
  INVX1 U11289 ( .A(n11327), .Y(n11325) );
  INVX1 U11290 ( .A(n11325), .Y(n11326) );
  BUFX2 U11291 ( .A(fifo[342]), .Y(n11327) );
  INVX1 U11292 ( .A(n11330), .Y(n11328) );
  INVX1 U11293 ( .A(n11328), .Y(n11329) );
  BUFX2 U11294 ( .A(fifo[343]), .Y(n11330) );
  INVX1 U11295 ( .A(n11333), .Y(n11331) );
  INVX1 U11296 ( .A(n11331), .Y(n11332) );
  BUFX2 U11297 ( .A(fifo[344]), .Y(n11333) );
  INVX1 U11298 ( .A(n11336), .Y(n11334) );
  INVX1 U11299 ( .A(n11334), .Y(n11335) );
  BUFX2 U11300 ( .A(fifo[345]), .Y(n11336) );
  INVX1 U11301 ( .A(n11339), .Y(n11337) );
  INVX1 U11302 ( .A(n11337), .Y(n11338) );
  BUFX2 U11303 ( .A(fifo[346]), .Y(n11339) );
  INVX1 U11304 ( .A(n11342), .Y(n11340) );
  INVX1 U11305 ( .A(n11340), .Y(n11341) );
  BUFX2 U11306 ( .A(fifo[347]), .Y(n11342) );
  INVX1 U11307 ( .A(n11345), .Y(n11343) );
  INVX1 U11308 ( .A(n11343), .Y(n11344) );
  BUFX2 U11309 ( .A(fifo[348]), .Y(n11345) );
  INVX1 U11310 ( .A(n11348), .Y(n11346) );
  INVX1 U11311 ( .A(n11346), .Y(n11347) );
  BUFX2 U11312 ( .A(fifo[349]), .Y(n11348) );
  INVX1 U11313 ( .A(n11351), .Y(n11349) );
  INVX1 U11314 ( .A(n11349), .Y(n11350) );
  BUFX2 U11315 ( .A(fifo[350]), .Y(n11351) );
  INVX1 U11316 ( .A(n11354), .Y(n11352) );
  INVX1 U11317 ( .A(n11352), .Y(n11353) );
  BUFX2 U11318 ( .A(fifo[351]), .Y(n11354) );
  INVX1 U11319 ( .A(n11357), .Y(n11355) );
  INVX1 U11320 ( .A(n11355), .Y(n11356) );
  BUFX2 U11321 ( .A(fifo[352]), .Y(n11357) );
  INVX1 U11322 ( .A(n11360), .Y(n11358) );
  INVX1 U11323 ( .A(n11358), .Y(n11359) );
  BUFX2 U11324 ( .A(fifo[353]), .Y(n11360) );
  INVX1 U11325 ( .A(n11363), .Y(n11361) );
  INVX1 U11326 ( .A(n11361), .Y(n11362) );
  BUFX2 U11327 ( .A(fifo[354]), .Y(n11363) );
  INVX1 U11328 ( .A(n11366), .Y(n11364) );
  INVX1 U11329 ( .A(n11364), .Y(n11365) );
  BUFX2 U11330 ( .A(fifo[355]), .Y(n11366) );
  INVX1 U11331 ( .A(n11369), .Y(n11367) );
  INVX1 U11332 ( .A(n11367), .Y(n11368) );
  BUFX2 U11333 ( .A(fifo[356]), .Y(n11369) );
  INVX1 U11334 ( .A(n11372), .Y(n11370) );
  INVX1 U11335 ( .A(n11370), .Y(n11371) );
  BUFX2 U11336 ( .A(fifo[357]), .Y(n11372) );
  INVX1 U11337 ( .A(n11375), .Y(n11373) );
  INVX1 U11338 ( .A(n11373), .Y(n11374) );
  BUFX2 U11339 ( .A(fifo[358]), .Y(n11375) );
  INVX1 U11340 ( .A(n11378), .Y(n11376) );
  INVX1 U11341 ( .A(n11376), .Y(n11377) );
  BUFX2 U11342 ( .A(fifo[359]), .Y(n11378) );
  INVX1 U11343 ( .A(n11381), .Y(n11379) );
  INVX1 U11344 ( .A(n11379), .Y(n11380) );
  BUFX2 U11345 ( .A(fifo[360]), .Y(n11381) );
  INVX1 U11346 ( .A(n11384), .Y(n11382) );
  INVX1 U11347 ( .A(n11382), .Y(n11383) );
  BUFX2 U11348 ( .A(fifo[361]), .Y(n11384) );
  INVX1 U11349 ( .A(n11387), .Y(n11385) );
  INVX1 U11350 ( .A(n11385), .Y(n11386) );
  BUFX2 U11351 ( .A(fifo[362]), .Y(n11387) );
  INVX1 U11352 ( .A(n11390), .Y(n11388) );
  INVX1 U11353 ( .A(n11388), .Y(n11389) );
  BUFX2 U11354 ( .A(fifo[363]), .Y(n11390) );
  INVX1 U11355 ( .A(n11393), .Y(n11391) );
  INVX1 U11356 ( .A(n11391), .Y(n11392) );
  BUFX2 U11357 ( .A(fifo[364]), .Y(n11393) );
  INVX1 U11358 ( .A(n11396), .Y(n11394) );
  INVX1 U11359 ( .A(n11394), .Y(n11395) );
  BUFX2 U11360 ( .A(fifo[365]), .Y(n11396) );
  INVX1 U11361 ( .A(n11399), .Y(n11397) );
  INVX1 U11362 ( .A(n11397), .Y(n11398) );
  BUFX2 U11363 ( .A(fifo[366]), .Y(n11399) );
  INVX1 U11364 ( .A(n11402), .Y(n11400) );
  INVX1 U11365 ( .A(n11400), .Y(n11401) );
  BUFX2 U11366 ( .A(fifo[367]), .Y(n11402) );
  INVX1 U11367 ( .A(n11405), .Y(n11403) );
  INVX1 U11368 ( .A(n11403), .Y(n11404) );
  BUFX2 U11369 ( .A(fifo[368]), .Y(n11405) );
  INVX1 U11370 ( .A(n11408), .Y(n11406) );
  INVX1 U11371 ( .A(n11406), .Y(n11407) );
  BUFX2 U11372 ( .A(fifo[369]), .Y(n11408) );
  INVX1 U11373 ( .A(n11411), .Y(n11409) );
  INVX1 U11374 ( .A(n11409), .Y(n11410) );
  BUFX2 U11375 ( .A(fifo[370]), .Y(n11411) );
  INVX1 U11376 ( .A(n11414), .Y(n11412) );
  INVX1 U11377 ( .A(n11412), .Y(n11413) );
  BUFX2 U11378 ( .A(fifo[371]), .Y(n11414) );
  INVX1 U11379 ( .A(n11417), .Y(n11415) );
  INVX1 U11380 ( .A(n11415), .Y(n11416) );
  BUFX2 U11381 ( .A(fifo[372]), .Y(n11417) );
  INVX1 U11382 ( .A(n11420), .Y(n11418) );
  INVX1 U11383 ( .A(n11418), .Y(n11419) );
  BUFX2 U11384 ( .A(fifo[373]), .Y(n11420) );
  INVX1 U11385 ( .A(n11423), .Y(n11421) );
  INVX1 U11386 ( .A(n11421), .Y(n11422) );
  BUFX2 U11387 ( .A(fifo[374]), .Y(n11423) );
  INVX1 U11388 ( .A(n11426), .Y(n11424) );
  INVX1 U11389 ( .A(n11424), .Y(n11425) );
  BUFX2 U11390 ( .A(fifo[375]), .Y(n11426) );
  INVX1 U11391 ( .A(n11429), .Y(n11427) );
  INVX1 U11392 ( .A(n11427), .Y(n11428) );
  BUFX2 U11393 ( .A(fifo[376]), .Y(n11429) );
  INVX1 U11394 ( .A(n11432), .Y(n11430) );
  INVX1 U11395 ( .A(n11430), .Y(n11431) );
  BUFX2 U11396 ( .A(fifo[377]), .Y(n11432) );
  INVX1 U11397 ( .A(n11435), .Y(n11433) );
  INVX1 U11398 ( .A(n11433), .Y(n11434) );
  BUFX2 U11399 ( .A(fifo[420]), .Y(n11435) );
  INVX1 U11400 ( .A(n11438), .Y(n11436) );
  INVX1 U11401 ( .A(n11436), .Y(n11437) );
  BUFX2 U11402 ( .A(fifo[421]), .Y(n11438) );
  INVX1 U11403 ( .A(n11441), .Y(n11439) );
  INVX1 U11404 ( .A(n11439), .Y(n11440) );
  BUFX2 U11405 ( .A(fifo[422]), .Y(n11441) );
  INVX1 U11406 ( .A(n11444), .Y(n11442) );
  INVX1 U11407 ( .A(n11442), .Y(n11443) );
  BUFX2 U11408 ( .A(fifo[423]), .Y(n11444) );
  INVX1 U11409 ( .A(n11447), .Y(n11445) );
  INVX1 U11410 ( .A(n11445), .Y(n11446) );
  BUFX2 U11411 ( .A(fifo[424]), .Y(n11447) );
  INVX1 U11412 ( .A(n11450), .Y(n11448) );
  INVX1 U11413 ( .A(n11448), .Y(n11449) );
  BUFX2 U11414 ( .A(fifo[425]), .Y(n11450) );
  INVX1 U11415 ( .A(n11453), .Y(n11451) );
  INVX1 U11416 ( .A(n11451), .Y(n11452) );
  BUFX2 U11417 ( .A(fifo[426]), .Y(n11453) );
  INVX1 U11418 ( .A(n11456), .Y(n11454) );
  INVX1 U11419 ( .A(n11454), .Y(n11455) );
  BUFX2 U11420 ( .A(fifo[427]), .Y(n11456) );
  INVX1 U11421 ( .A(n11459), .Y(n11457) );
  INVX1 U11422 ( .A(n11457), .Y(n11458) );
  BUFX2 U11423 ( .A(fifo[428]), .Y(n11459) );
  INVX1 U11424 ( .A(n11462), .Y(n11460) );
  INVX1 U11425 ( .A(n11460), .Y(n11461) );
  BUFX2 U11426 ( .A(fifo[429]), .Y(n11462) );
  INVX1 U11427 ( .A(n11465), .Y(n11463) );
  INVX1 U11428 ( .A(n11463), .Y(n11464) );
  BUFX2 U11429 ( .A(fifo[430]), .Y(n11465) );
  INVX1 U11430 ( .A(n11468), .Y(n11466) );
  INVX1 U11431 ( .A(n11466), .Y(n11467) );
  BUFX2 U11432 ( .A(fifo[431]), .Y(n11468) );
  INVX1 U11433 ( .A(n11471), .Y(n11469) );
  INVX1 U11434 ( .A(n11469), .Y(n11470) );
  BUFX2 U11435 ( .A(fifo[432]), .Y(n11471) );
  INVX1 U11436 ( .A(n11474), .Y(n11472) );
  INVX1 U11437 ( .A(n11472), .Y(n11473) );
  BUFX2 U11438 ( .A(fifo[433]), .Y(n11474) );
  INVX1 U11439 ( .A(n11477), .Y(n11475) );
  INVX1 U11440 ( .A(n11475), .Y(n11476) );
  BUFX2 U11441 ( .A(fifo[434]), .Y(n11477) );
  INVX1 U11442 ( .A(n11480), .Y(n11478) );
  INVX1 U11443 ( .A(n11478), .Y(n11479) );
  BUFX2 U11444 ( .A(fifo[435]), .Y(n11480) );
  INVX1 U11445 ( .A(n11483), .Y(n11481) );
  INVX1 U11446 ( .A(n11481), .Y(n11482) );
  BUFX2 U11447 ( .A(fifo[436]), .Y(n11483) );
  INVX1 U11448 ( .A(n11486), .Y(n11484) );
  INVX1 U11449 ( .A(n11484), .Y(n11485) );
  BUFX2 U11450 ( .A(fifo[437]), .Y(n11486) );
  INVX1 U11451 ( .A(n11489), .Y(n11487) );
  INVX1 U11452 ( .A(n11487), .Y(n11488) );
  BUFX2 U11453 ( .A(fifo[438]), .Y(n11489) );
  INVX1 U11454 ( .A(n11492), .Y(n11490) );
  INVX1 U11455 ( .A(n11490), .Y(n11491) );
  BUFX2 U11456 ( .A(fifo[439]), .Y(n11492) );
  INVX1 U11457 ( .A(n11495), .Y(n11493) );
  INVX1 U11458 ( .A(n11493), .Y(n11494) );
  BUFX2 U11459 ( .A(fifo[440]), .Y(n11495) );
  INVX1 U11460 ( .A(n11498), .Y(n11496) );
  INVX1 U11461 ( .A(n11496), .Y(n11497) );
  BUFX2 U11462 ( .A(fifo[441]), .Y(n11498) );
  INVX1 U11463 ( .A(n11501), .Y(n11499) );
  INVX1 U11464 ( .A(n11499), .Y(n11500) );
  BUFX2 U11465 ( .A(fifo[442]), .Y(n11501) );
  INVX1 U11466 ( .A(n11504), .Y(n11502) );
  INVX1 U11467 ( .A(n11502), .Y(n11503) );
  BUFX2 U11468 ( .A(fifo[443]), .Y(n11504) );
  INVX1 U11469 ( .A(n11507), .Y(n11505) );
  INVX1 U11470 ( .A(n11505), .Y(n11506) );
  BUFX2 U11471 ( .A(fifo[444]), .Y(n11507) );
  INVX1 U11472 ( .A(n11510), .Y(n11508) );
  INVX1 U11473 ( .A(n11508), .Y(n11509) );
  BUFX2 U11474 ( .A(fifo[445]), .Y(n11510) );
  INVX1 U11475 ( .A(n11513), .Y(n11511) );
  INVX1 U11476 ( .A(n11511), .Y(n11512) );
  BUFX2 U11477 ( .A(fifo[446]), .Y(n11513) );
  INVX1 U11478 ( .A(n11516), .Y(n11514) );
  INVX1 U11479 ( .A(n11514), .Y(n11515) );
  BUFX2 U11480 ( .A(fifo[447]), .Y(n11516) );
  INVX1 U11481 ( .A(n11519), .Y(n11517) );
  INVX1 U11482 ( .A(n11517), .Y(n11518) );
  BUFX2 U11483 ( .A(fifo[448]), .Y(n11519) );
  INVX1 U11484 ( .A(n11522), .Y(n11520) );
  INVX1 U11485 ( .A(n11520), .Y(n11521) );
  BUFX2 U11486 ( .A(fifo[449]), .Y(n11522) );
  INVX1 U11487 ( .A(n11525), .Y(n11523) );
  INVX1 U11488 ( .A(n11523), .Y(n11524) );
  BUFX2 U11489 ( .A(fifo[450]), .Y(n11525) );
  INVX1 U11490 ( .A(n11528), .Y(n11526) );
  INVX1 U11491 ( .A(n11526), .Y(n11527) );
  BUFX2 U11492 ( .A(fifo[451]), .Y(n11528) );
  INVX1 U11493 ( .A(n11531), .Y(n11529) );
  INVX1 U11494 ( .A(n11529), .Y(n11530) );
  BUFX2 U11495 ( .A(fifo[452]), .Y(n11531) );
  INVX1 U11496 ( .A(n11534), .Y(n11532) );
  INVX1 U11497 ( .A(n11532), .Y(n11533) );
  BUFX2 U11498 ( .A(fifo[453]), .Y(n11534) );
  INVX1 U11499 ( .A(n11537), .Y(n11535) );
  INVX1 U11500 ( .A(n11535), .Y(n11536) );
  BUFX2 U11501 ( .A(fifo[454]), .Y(n11537) );
  INVX1 U11502 ( .A(n11540), .Y(n11538) );
  INVX1 U11503 ( .A(n11538), .Y(n11539) );
  BUFX2 U11504 ( .A(fifo[455]), .Y(n11540) );
  INVX1 U11505 ( .A(n11543), .Y(n11541) );
  INVX1 U11506 ( .A(n11541), .Y(n11542) );
  BUFX2 U11507 ( .A(fifo[456]), .Y(n11543) );
  INVX1 U11508 ( .A(n11546), .Y(n11544) );
  INVX1 U11509 ( .A(n11544), .Y(n11545) );
  BUFX2 U11510 ( .A(fifo[457]), .Y(n11546) );
  INVX1 U11511 ( .A(n11549), .Y(n11547) );
  INVX1 U11512 ( .A(n11547), .Y(n11548) );
  BUFX2 U11513 ( .A(fifo[458]), .Y(n11549) );
  INVX1 U11514 ( .A(n11552), .Y(n11550) );
  INVX1 U11515 ( .A(n11550), .Y(n11551) );
  BUFX2 U11516 ( .A(fifo[459]), .Y(n11552) );
  INVX1 U11517 ( .A(n11555), .Y(n11553) );
  INVX1 U11518 ( .A(n11553), .Y(n11554) );
  BUFX2 U11519 ( .A(fifo[460]), .Y(n11555) );
  INVX1 U11520 ( .A(n11558), .Y(n11556) );
  INVX1 U11521 ( .A(n11556), .Y(n11557) );
  BUFX2 U11522 ( .A(fifo[461]), .Y(n11558) );
  INVX1 U11523 ( .A(n11561), .Y(n11559) );
  INVX1 U11524 ( .A(n11559), .Y(n11560) );
  BUFX2 U11525 ( .A(fifo[504]), .Y(n11561) );
  INVX1 U11526 ( .A(n11564), .Y(n11562) );
  INVX1 U11527 ( .A(n11562), .Y(n11563) );
  BUFX2 U11528 ( .A(fifo[505]), .Y(n11564) );
  INVX1 U11529 ( .A(n11567), .Y(n11565) );
  INVX1 U11530 ( .A(n11565), .Y(n11566) );
  BUFX2 U11531 ( .A(fifo[506]), .Y(n11567) );
  INVX1 U11532 ( .A(n11570), .Y(n11568) );
  INVX1 U11533 ( .A(n11568), .Y(n11569) );
  BUFX2 U11534 ( .A(fifo[507]), .Y(n11570) );
  INVX1 U11535 ( .A(n11573), .Y(n11571) );
  INVX1 U11536 ( .A(n11571), .Y(n11572) );
  BUFX2 U11537 ( .A(fifo[508]), .Y(n11573) );
  INVX1 U11538 ( .A(n11576), .Y(n11574) );
  INVX1 U11539 ( .A(n11574), .Y(n11575) );
  BUFX2 U11540 ( .A(fifo[509]), .Y(n11576) );
  INVX1 U11541 ( .A(n11579), .Y(n11577) );
  INVX1 U11542 ( .A(n11577), .Y(n11578) );
  BUFX2 U11543 ( .A(fifo[510]), .Y(n11579) );
  INVX1 U11544 ( .A(n11582), .Y(n11580) );
  INVX1 U11545 ( .A(n11580), .Y(n11581) );
  BUFX2 U11546 ( .A(fifo[511]), .Y(n11582) );
  INVX1 U11547 ( .A(n11585), .Y(n11583) );
  INVX1 U11548 ( .A(n11583), .Y(n11584) );
  BUFX2 U11549 ( .A(fifo[512]), .Y(n11585) );
  INVX1 U11550 ( .A(n11588), .Y(n11586) );
  INVX1 U11551 ( .A(n11586), .Y(n11587) );
  BUFX2 U11552 ( .A(fifo[513]), .Y(n11588) );
  INVX1 U11553 ( .A(n11591), .Y(n11589) );
  INVX1 U11554 ( .A(n11589), .Y(n11590) );
  BUFX2 U11555 ( .A(fifo[514]), .Y(n11591) );
  INVX1 U11556 ( .A(n11594), .Y(n11592) );
  INVX1 U11557 ( .A(n11592), .Y(n11593) );
  BUFX2 U11558 ( .A(fifo[515]), .Y(n11594) );
  INVX1 U11559 ( .A(n11597), .Y(n11595) );
  INVX1 U11560 ( .A(n11595), .Y(n11596) );
  BUFX2 U11561 ( .A(fifo[516]), .Y(n11597) );
  INVX1 U11562 ( .A(n11600), .Y(n11598) );
  INVX1 U11563 ( .A(n11598), .Y(n11599) );
  BUFX2 U11564 ( .A(fifo[517]), .Y(n11600) );
  INVX1 U11565 ( .A(n11603), .Y(n11601) );
  INVX1 U11566 ( .A(n11601), .Y(n11602) );
  BUFX2 U11567 ( .A(fifo[518]), .Y(n11603) );
  INVX1 U11568 ( .A(n11606), .Y(n11604) );
  INVX1 U11569 ( .A(n11604), .Y(n11605) );
  BUFX2 U11570 ( .A(fifo[519]), .Y(n11606) );
  INVX1 U11571 ( .A(n11609), .Y(n11607) );
  INVX1 U11572 ( .A(n11607), .Y(n11608) );
  BUFX2 U11573 ( .A(fifo[520]), .Y(n11609) );
  INVX1 U11574 ( .A(n11612), .Y(n11610) );
  INVX1 U11575 ( .A(n11610), .Y(n11611) );
  BUFX2 U11576 ( .A(fifo[521]), .Y(n11612) );
  INVX1 U11577 ( .A(n11615), .Y(n11613) );
  INVX1 U11578 ( .A(n11613), .Y(n11614) );
  BUFX2 U11579 ( .A(fifo[522]), .Y(n11615) );
  INVX1 U11580 ( .A(n11618), .Y(n11616) );
  INVX1 U11581 ( .A(n11616), .Y(n11617) );
  BUFX2 U11582 ( .A(fifo[523]), .Y(n11618) );
  INVX1 U11583 ( .A(n11621), .Y(n11619) );
  INVX1 U11584 ( .A(n11619), .Y(n11620) );
  BUFX2 U11585 ( .A(fifo[524]), .Y(n11621) );
  INVX1 U11586 ( .A(n11624), .Y(n11622) );
  INVX1 U11587 ( .A(n11622), .Y(n11623) );
  BUFX2 U11588 ( .A(fifo[525]), .Y(n11624) );
  INVX1 U11589 ( .A(n11627), .Y(n11625) );
  INVX1 U11590 ( .A(n11625), .Y(n11626) );
  BUFX2 U11591 ( .A(fifo[526]), .Y(n11627) );
  INVX1 U11592 ( .A(n11630), .Y(n11628) );
  INVX1 U11593 ( .A(n11628), .Y(n11629) );
  BUFX2 U11594 ( .A(fifo[527]), .Y(n11630) );
  INVX1 U11595 ( .A(n11633), .Y(n11631) );
  INVX1 U11596 ( .A(n11631), .Y(n11632) );
  BUFX2 U11597 ( .A(fifo[528]), .Y(n11633) );
  INVX1 U11598 ( .A(n11636), .Y(n11634) );
  INVX1 U11599 ( .A(n11634), .Y(n11635) );
  BUFX2 U11600 ( .A(fifo[529]), .Y(n11636) );
  INVX1 U11601 ( .A(n11639), .Y(n11637) );
  INVX1 U11602 ( .A(n11637), .Y(n11638) );
  BUFX2 U11603 ( .A(fifo[530]), .Y(n11639) );
  INVX1 U11604 ( .A(n11642), .Y(n11640) );
  INVX1 U11605 ( .A(n11640), .Y(n11641) );
  BUFX2 U11606 ( .A(fifo[531]), .Y(n11642) );
  INVX1 U11607 ( .A(n11645), .Y(n11643) );
  INVX1 U11608 ( .A(n11643), .Y(n11644) );
  BUFX2 U11609 ( .A(fifo[532]), .Y(n11645) );
  INVX1 U11610 ( .A(n11648), .Y(n11646) );
  INVX1 U11611 ( .A(n11646), .Y(n11647) );
  BUFX2 U11612 ( .A(fifo[533]), .Y(n11648) );
  INVX1 U11613 ( .A(n11651), .Y(n11649) );
  INVX1 U11614 ( .A(n11649), .Y(n11650) );
  BUFX2 U11615 ( .A(fifo[534]), .Y(n11651) );
  INVX1 U11616 ( .A(n11654), .Y(n11652) );
  INVX1 U11617 ( .A(n11652), .Y(n11653) );
  BUFX2 U11618 ( .A(fifo[535]), .Y(n11654) );
  INVX1 U11619 ( .A(n11657), .Y(n11655) );
  INVX1 U11620 ( .A(n11655), .Y(n11656) );
  BUFX2 U11621 ( .A(fifo[536]), .Y(n11657) );
  INVX1 U11622 ( .A(n11660), .Y(n11658) );
  INVX1 U11623 ( .A(n11658), .Y(n11659) );
  BUFX2 U11624 ( .A(fifo[537]), .Y(n11660) );
  INVX1 U11625 ( .A(n11663), .Y(n11661) );
  INVX1 U11626 ( .A(n11661), .Y(n11662) );
  BUFX2 U11627 ( .A(fifo[538]), .Y(n11663) );
  INVX1 U11628 ( .A(n11666), .Y(n11664) );
  INVX1 U11629 ( .A(n11664), .Y(n11665) );
  BUFX2 U11630 ( .A(fifo[539]), .Y(n11666) );
  INVX1 U11631 ( .A(n11669), .Y(n11667) );
  INVX1 U11632 ( .A(n11667), .Y(n11668) );
  BUFX2 U11633 ( .A(fifo[540]), .Y(n11669) );
  INVX1 U11634 ( .A(n11672), .Y(n11670) );
  INVX1 U11635 ( .A(n11670), .Y(n11671) );
  BUFX2 U11636 ( .A(fifo[541]), .Y(n11672) );
  INVX1 U11637 ( .A(n11675), .Y(n11673) );
  INVX1 U11638 ( .A(n11673), .Y(n11674) );
  BUFX2 U11639 ( .A(fifo[542]), .Y(n11675) );
  INVX1 U11640 ( .A(n11678), .Y(n11676) );
  INVX1 U11641 ( .A(n11676), .Y(n11677) );
  BUFX2 U11642 ( .A(fifo[543]), .Y(n11678) );
  INVX1 U11643 ( .A(n11681), .Y(n11679) );
  INVX1 U11644 ( .A(n11679), .Y(n11680) );
  BUFX2 U11645 ( .A(fifo[544]), .Y(n11681) );
  INVX1 U11646 ( .A(n11684), .Y(n11682) );
  INVX1 U11647 ( .A(n11682), .Y(n11683) );
  BUFX2 U11648 ( .A(fifo[545]), .Y(n11684) );
  INVX1 U11649 ( .A(n11687), .Y(n11685) );
  INVX1 U11650 ( .A(n11685), .Y(n11686) );
  BUFX2 U11651 ( .A(fifo[588]), .Y(n11687) );
  INVX1 U11652 ( .A(n11690), .Y(n11688) );
  INVX1 U11653 ( .A(n11688), .Y(n11689) );
  BUFX2 U11654 ( .A(fifo[589]), .Y(n11690) );
  INVX1 U11655 ( .A(n11693), .Y(n11691) );
  INVX1 U11656 ( .A(n11691), .Y(n11692) );
  BUFX2 U11657 ( .A(fifo[590]), .Y(n11693) );
  INVX1 U11658 ( .A(n11696), .Y(n11694) );
  INVX1 U11659 ( .A(n11694), .Y(n11695) );
  BUFX2 U11660 ( .A(fifo[591]), .Y(n11696) );
  INVX1 U11661 ( .A(n11699), .Y(n11697) );
  INVX1 U11662 ( .A(n11697), .Y(n11698) );
  BUFX2 U11663 ( .A(fifo[592]), .Y(n11699) );
  INVX1 U11664 ( .A(n11702), .Y(n11700) );
  INVX1 U11665 ( .A(n11700), .Y(n11701) );
  BUFX2 U11666 ( .A(fifo[593]), .Y(n11702) );
  INVX1 U11667 ( .A(n11705), .Y(n11703) );
  INVX1 U11668 ( .A(n11703), .Y(n11704) );
  BUFX2 U11669 ( .A(fifo[594]), .Y(n11705) );
  INVX1 U11670 ( .A(n11708), .Y(n11706) );
  INVX1 U11671 ( .A(n11706), .Y(n11707) );
  BUFX2 U11672 ( .A(fifo[595]), .Y(n11708) );
  INVX1 U11673 ( .A(n11711), .Y(n11709) );
  INVX1 U11674 ( .A(n11709), .Y(n11710) );
  BUFX2 U11675 ( .A(fifo[596]), .Y(n11711) );
  INVX1 U11676 ( .A(n11714), .Y(n11712) );
  INVX1 U11677 ( .A(n11712), .Y(n11713) );
  BUFX2 U11678 ( .A(fifo[597]), .Y(n11714) );
  INVX1 U11679 ( .A(n11717), .Y(n11715) );
  INVX1 U11680 ( .A(n11715), .Y(n11716) );
  BUFX2 U11681 ( .A(fifo[598]), .Y(n11717) );
  INVX1 U11682 ( .A(n11720), .Y(n11718) );
  INVX1 U11683 ( .A(n11718), .Y(n11719) );
  BUFX2 U11684 ( .A(fifo[599]), .Y(n11720) );
  INVX1 U11685 ( .A(n11723), .Y(n11721) );
  INVX1 U11686 ( .A(n11721), .Y(n11722) );
  BUFX2 U11687 ( .A(fifo[600]), .Y(n11723) );
  INVX1 U11688 ( .A(n11726), .Y(n11724) );
  INVX1 U11689 ( .A(n11724), .Y(n11725) );
  BUFX2 U11690 ( .A(fifo[601]), .Y(n11726) );
  INVX1 U11691 ( .A(n11729), .Y(n11727) );
  INVX1 U11692 ( .A(n11727), .Y(n11728) );
  BUFX2 U11693 ( .A(fifo[602]), .Y(n11729) );
  INVX1 U11694 ( .A(n11732), .Y(n11730) );
  INVX1 U11695 ( .A(n11730), .Y(n11731) );
  BUFX2 U11696 ( .A(fifo[603]), .Y(n11732) );
  INVX1 U11697 ( .A(n11735), .Y(n11733) );
  INVX1 U11698 ( .A(n11733), .Y(n11734) );
  BUFX2 U11699 ( .A(fifo[604]), .Y(n11735) );
  INVX1 U11700 ( .A(n11738), .Y(n11736) );
  INVX1 U11701 ( .A(n11736), .Y(n11737) );
  BUFX2 U11702 ( .A(fifo[605]), .Y(n11738) );
  INVX1 U11703 ( .A(n11741), .Y(n11739) );
  INVX1 U11704 ( .A(n11739), .Y(n11740) );
  BUFX2 U11705 ( .A(fifo[606]), .Y(n11741) );
  INVX1 U11706 ( .A(n11744), .Y(n11742) );
  INVX1 U11707 ( .A(n11742), .Y(n11743) );
  BUFX2 U11708 ( .A(fifo[607]), .Y(n11744) );
  INVX1 U11709 ( .A(n11747), .Y(n11745) );
  INVX1 U11710 ( .A(n11745), .Y(n11746) );
  BUFX2 U11711 ( .A(fifo[608]), .Y(n11747) );
  INVX1 U11712 ( .A(n11750), .Y(n11748) );
  INVX1 U11713 ( .A(n11748), .Y(n11749) );
  BUFX2 U11714 ( .A(fifo[609]), .Y(n11750) );
  INVX1 U11715 ( .A(n11753), .Y(n11751) );
  INVX1 U11716 ( .A(n11751), .Y(n11752) );
  BUFX2 U11717 ( .A(fifo[610]), .Y(n11753) );
  INVX1 U11718 ( .A(n11756), .Y(n11754) );
  INVX1 U11719 ( .A(n11754), .Y(n11755) );
  BUFX2 U11720 ( .A(fifo[611]), .Y(n11756) );
  INVX1 U11721 ( .A(n11759), .Y(n11757) );
  INVX1 U11722 ( .A(n11757), .Y(n11758) );
  BUFX2 U11723 ( .A(fifo[612]), .Y(n11759) );
  INVX1 U11724 ( .A(n11762), .Y(n11760) );
  INVX1 U11725 ( .A(n11760), .Y(n11761) );
  BUFX2 U11726 ( .A(fifo[613]), .Y(n11762) );
  INVX1 U11727 ( .A(n11765), .Y(n11763) );
  INVX1 U11728 ( .A(n11763), .Y(n11764) );
  BUFX2 U11729 ( .A(fifo[614]), .Y(n11765) );
  INVX1 U11730 ( .A(n11768), .Y(n11766) );
  INVX1 U11731 ( .A(n11766), .Y(n11767) );
  BUFX2 U11732 ( .A(fifo[615]), .Y(n11768) );
  INVX1 U11733 ( .A(n11771), .Y(n11769) );
  INVX1 U11734 ( .A(n11769), .Y(n11770) );
  BUFX2 U11735 ( .A(fifo[616]), .Y(n11771) );
  INVX1 U11736 ( .A(n11774), .Y(n11772) );
  INVX1 U11737 ( .A(n11772), .Y(n11773) );
  BUFX2 U11738 ( .A(fifo[617]), .Y(n11774) );
  INVX1 U11739 ( .A(n11777), .Y(n11775) );
  INVX1 U11740 ( .A(n11775), .Y(n11776) );
  BUFX2 U11741 ( .A(fifo[618]), .Y(n11777) );
  INVX1 U11742 ( .A(n11780), .Y(n11778) );
  INVX1 U11743 ( .A(n11778), .Y(n11779) );
  BUFX2 U11744 ( .A(fifo[619]), .Y(n11780) );
  INVX1 U11745 ( .A(n11783), .Y(n11781) );
  INVX1 U11746 ( .A(n11781), .Y(n11782) );
  BUFX2 U11747 ( .A(fifo[620]), .Y(n11783) );
  INVX1 U11748 ( .A(n11786), .Y(n11784) );
  INVX1 U11749 ( .A(n11784), .Y(n11785) );
  BUFX2 U11750 ( .A(fifo[621]), .Y(n11786) );
  INVX1 U11751 ( .A(n11789), .Y(n11787) );
  INVX1 U11752 ( .A(n11787), .Y(n11788) );
  BUFX2 U11753 ( .A(fifo[622]), .Y(n11789) );
  INVX1 U11754 ( .A(n11792), .Y(n11790) );
  INVX1 U11755 ( .A(n11790), .Y(n11791) );
  BUFX2 U11756 ( .A(fifo[623]), .Y(n11792) );
  INVX1 U11757 ( .A(n11795), .Y(n11793) );
  INVX1 U11758 ( .A(n11793), .Y(n11794) );
  BUFX2 U11759 ( .A(fifo[624]), .Y(n11795) );
  INVX1 U11760 ( .A(n11798), .Y(n11796) );
  INVX1 U11761 ( .A(n11796), .Y(n11797) );
  BUFX2 U11762 ( .A(fifo[625]), .Y(n11798) );
  INVX1 U11763 ( .A(n11801), .Y(n11799) );
  INVX1 U11764 ( .A(n11799), .Y(n11800) );
  BUFX2 U11765 ( .A(fifo[626]), .Y(n11801) );
  INVX1 U11766 ( .A(n11804), .Y(n11802) );
  INVX1 U11767 ( .A(n11802), .Y(n11803) );
  BUFX2 U11768 ( .A(fifo[627]), .Y(n11804) );
  INVX1 U11769 ( .A(n11807), .Y(n11805) );
  INVX1 U11770 ( .A(n11805), .Y(n11806) );
  BUFX2 U11771 ( .A(fifo[628]), .Y(n11807) );
  INVX1 U11772 ( .A(n11810), .Y(n11808) );
  INVX1 U11773 ( .A(n11808), .Y(n11809) );
  BUFX2 U11774 ( .A(fifo[629]), .Y(n11810) );
  INVX1 U11775 ( .A(n11813), .Y(n11811) );
  INVX1 U11776 ( .A(n11811), .Y(n11812) );
  BUFX2 U11777 ( .A(fifo[672]), .Y(n11813) );
  INVX1 U11778 ( .A(n11816), .Y(n11814) );
  INVX1 U11779 ( .A(n11814), .Y(n11815) );
  BUFX2 U11780 ( .A(fifo[673]), .Y(n11816) );
  INVX1 U11781 ( .A(n11819), .Y(n11817) );
  INVX1 U11782 ( .A(n11817), .Y(n11818) );
  BUFX2 U11783 ( .A(fifo[674]), .Y(n11819) );
  INVX1 U11784 ( .A(n11822), .Y(n11820) );
  INVX1 U11785 ( .A(n11820), .Y(n11821) );
  BUFX2 U11786 ( .A(fifo[675]), .Y(n11822) );
  INVX1 U11787 ( .A(n11825), .Y(n11823) );
  INVX1 U11788 ( .A(n11823), .Y(n11824) );
  BUFX2 U11789 ( .A(fifo[676]), .Y(n11825) );
  INVX1 U11790 ( .A(n11828), .Y(n11826) );
  INVX1 U11791 ( .A(n11826), .Y(n11827) );
  BUFX2 U11792 ( .A(fifo[677]), .Y(n11828) );
  INVX1 U11793 ( .A(n11831), .Y(n11829) );
  INVX1 U11794 ( .A(n11829), .Y(n11830) );
  BUFX2 U11795 ( .A(fifo[678]), .Y(n11831) );
  INVX1 U11796 ( .A(n11834), .Y(n11832) );
  INVX1 U11797 ( .A(n11832), .Y(n11833) );
  BUFX2 U11798 ( .A(fifo[679]), .Y(n11834) );
  INVX1 U11799 ( .A(n11837), .Y(n11835) );
  INVX1 U11800 ( .A(n11835), .Y(n11836) );
  BUFX2 U11801 ( .A(fifo[680]), .Y(n11837) );
  INVX1 U11802 ( .A(n11840), .Y(n11838) );
  INVX1 U11803 ( .A(n11838), .Y(n11839) );
  BUFX2 U11804 ( .A(fifo[681]), .Y(n11840) );
  INVX1 U11805 ( .A(n11843), .Y(n11841) );
  INVX1 U11806 ( .A(n11841), .Y(n11842) );
  BUFX2 U11807 ( .A(fifo[682]), .Y(n11843) );
  INVX1 U11808 ( .A(n11846), .Y(n11844) );
  INVX1 U11809 ( .A(n11844), .Y(n11845) );
  BUFX2 U11810 ( .A(fifo[683]), .Y(n11846) );
  INVX1 U11811 ( .A(n11849), .Y(n11847) );
  INVX1 U11812 ( .A(n11847), .Y(n11848) );
  BUFX2 U11813 ( .A(fifo[684]), .Y(n11849) );
  INVX1 U11814 ( .A(n11852), .Y(n11850) );
  INVX1 U11815 ( .A(n11850), .Y(n11851) );
  BUFX2 U11816 ( .A(fifo[685]), .Y(n11852) );
  INVX1 U11817 ( .A(n11855), .Y(n11853) );
  INVX1 U11818 ( .A(n11853), .Y(n11854) );
  BUFX2 U11819 ( .A(fifo[686]), .Y(n11855) );
  INVX1 U11820 ( .A(n11858), .Y(n11856) );
  INVX1 U11821 ( .A(n11856), .Y(n11857) );
  BUFX2 U11822 ( .A(fifo[687]), .Y(n11858) );
  INVX1 U11823 ( .A(n11861), .Y(n11859) );
  INVX1 U11824 ( .A(n11859), .Y(n11860) );
  BUFX2 U11825 ( .A(fifo[688]), .Y(n11861) );
  INVX1 U11826 ( .A(n11864), .Y(n11862) );
  INVX1 U11827 ( .A(n11862), .Y(n11863) );
  BUFX2 U11828 ( .A(fifo[689]), .Y(n11864) );
  INVX1 U11829 ( .A(n11867), .Y(n11865) );
  INVX1 U11830 ( .A(n11865), .Y(n11866) );
  BUFX2 U11831 ( .A(fifo[690]), .Y(n11867) );
  INVX1 U11832 ( .A(n11870), .Y(n11868) );
  INVX1 U11833 ( .A(n11868), .Y(n11869) );
  BUFX2 U11834 ( .A(fifo[691]), .Y(n11870) );
  INVX1 U11835 ( .A(n11873), .Y(n11871) );
  INVX1 U11836 ( .A(n11871), .Y(n11872) );
  BUFX2 U11837 ( .A(fifo[692]), .Y(n11873) );
  INVX1 U11838 ( .A(n11876), .Y(n11874) );
  INVX1 U11839 ( .A(n11874), .Y(n11875) );
  BUFX2 U11840 ( .A(fifo[693]), .Y(n11876) );
  INVX1 U11841 ( .A(n11879), .Y(n11877) );
  INVX1 U11842 ( .A(n11877), .Y(n11878) );
  BUFX2 U11843 ( .A(fifo[694]), .Y(n11879) );
  INVX1 U11844 ( .A(n11882), .Y(n11880) );
  INVX1 U11845 ( .A(n11880), .Y(n11881) );
  BUFX2 U11846 ( .A(fifo[695]), .Y(n11882) );
  INVX1 U11847 ( .A(n11885), .Y(n11883) );
  INVX1 U11848 ( .A(n11883), .Y(n11884) );
  BUFX2 U11849 ( .A(fifo[696]), .Y(n11885) );
  INVX1 U11850 ( .A(n11888), .Y(n11886) );
  INVX1 U11851 ( .A(n11886), .Y(n11887) );
  BUFX2 U11852 ( .A(fifo[697]), .Y(n11888) );
  INVX1 U11853 ( .A(n11891), .Y(n11889) );
  INVX1 U11854 ( .A(n11889), .Y(n11890) );
  BUFX2 U11855 ( .A(fifo[698]), .Y(n11891) );
  INVX1 U11856 ( .A(n11894), .Y(n11892) );
  INVX1 U11857 ( .A(n11892), .Y(n11893) );
  BUFX2 U11858 ( .A(fifo[699]), .Y(n11894) );
  INVX1 U11859 ( .A(n11897), .Y(n11895) );
  INVX1 U11860 ( .A(n11895), .Y(n11896) );
  BUFX2 U11861 ( .A(fifo[700]), .Y(n11897) );
  INVX1 U11862 ( .A(n11900), .Y(n11898) );
  INVX1 U11863 ( .A(n11898), .Y(n11899) );
  BUFX2 U11864 ( .A(fifo[701]), .Y(n11900) );
  INVX1 U11865 ( .A(n11903), .Y(n11901) );
  INVX1 U11866 ( .A(n11901), .Y(n11902) );
  BUFX2 U11867 ( .A(fifo[702]), .Y(n11903) );
  INVX1 U11868 ( .A(n11906), .Y(n11904) );
  INVX1 U11869 ( .A(n11904), .Y(n11905) );
  BUFX2 U11870 ( .A(fifo[703]), .Y(n11906) );
  INVX1 U11871 ( .A(n11909), .Y(n11907) );
  INVX1 U11872 ( .A(n11907), .Y(n11908) );
  BUFX2 U11873 ( .A(fifo[704]), .Y(n11909) );
  INVX1 U11874 ( .A(n11912), .Y(n11910) );
  INVX1 U11875 ( .A(n11910), .Y(n11911) );
  BUFX2 U11876 ( .A(fifo[705]), .Y(n11912) );
  INVX1 U11877 ( .A(n11915), .Y(n11913) );
  INVX1 U11878 ( .A(n11913), .Y(n11914) );
  BUFX2 U11879 ( .A(fifo[706]), .Y(n11915) );
  INVX1 U11880 ( .A(n11918), .Y(n11916) );
  INVX1 U11881 ( .A(n11916), .Y(n11917) );
  BUFX2 U11882 ( .A(fifo[707]), .Y(n11918) );
  INVX1 U11883 ( .A(n11921), .Y(n11919) );
  INVX1 U11884 ( .A(n11919), .Y(n11920) );
  BUFX2 U11885 ( .A(fifo[708]), .Y(n11921) );
  INVX1 U11886 ( .A(n11924), .Y(n11922) );
  INVX1 U11887 ( .A(n11922), .Y(n11923) );
  BUFX2 U11888 ( .A(fifo[709]), .Y(n11924) );
  INVX1 U11889 ( .A(n11927), .Y(n11925) );
  INVX1 U11890 ( .A(n11925), .Y(n11926) );
  BUFX2 U11891 ( .A(fifo[710]), .Y(n11927) );
  INVX1 U11892 ( .A(n11930), .Y(n11928) );
  INVX1 U11893 ( .A(n11928), .Y(n11929) );
  BUFX2 U11894 ( .A(fifo[711]), .Y(n11930) );
  INVX1 U11895 ( .A(n11933), .Y(n11931) );
  INVX1 U11896 ( .A(n11931), .Y(n11932) );
  BUFX2 U11897 ( .A(fifo[712]), .Y(n11933) );
  INVX1 U11898 ( .A(n11936), .Y(n11934) );
  INVX1 U11899 ( .A(n11934), .Y(n11935) );
  BUFX2 U11900 ( .A(fifo[713]), .Y(n11936) );
  INVX1 U11901 ( .A(n11939), .Y(n11937) );
  INVX1 U11902 ( .A(n11937), .Y(n11938) );
  BUFX2 U11903 ( .A(fifo[756]), .Y(n11939) );
  INVX1 U11904 ( .A(n11942), .Y(n11940) );
  INVX1 U11905 ( .A(n11940), .Y(n11941) );
  BUFX2 U11906 ( .A(fifo[757]), .Y(n11942) );
  INVX1 U11907 ( .A(n11945), .Y(n11943) );
  INVX1 U11908 ( .A(n11943), .Y(n11944) );
  BUFX2 U11909 ( .A(fifo[758]), .Y(n11945) );
  INVX1 U11910 ( .A(n11948), .Y(n11946) );
  INVX1 U11911 ( .A(n11946), .Y(n11947) );
  BUFX2 U11912 ( .A(fifo[759]), .Y(n11948) );
  INVX1 U11913 ( .A(n11951), .Y(n11949) );
  INVX1 U11914 ( .A(n11949), .Y(n11950) );
  BUFX2 U11915 ( .A(fifo[760]), .Y(n11951) );
  INVX1 U11916 ( .A(n11954), .Y(n11952) );
  INVX1 U11917 ( .A(n11952), .Y(n11953) );
  BUFX2 U11918 ( .A(fifo[761]), .Y(n11954) );
  INVX1 U11919 ( .A(n11957), .Y(n11955) );
  INVX1 U11920 ( .A(n11955), .Y(n11956) );
  BUFX2 U11921 ( .A(fifo[762]), .Y(n11957) );
  INVX1 U11922 ( .A(n11960), .Y(n11958) );
  INVX1 U11923 ( .A(n11958), .Y(n11959) );
  BUFX2 U11924 ( .A(fifo[763]), .Y(n11960) );
  INVX1 U11925 ( .A(n11963), .Y(n11961) );
  INVX1 U11926 ( .A(n11961), .Y(n11962) );
  BUFX2 U11927 ( .A(fifo[764]), .Y(n11963) );
  INVX1 U11928 ( .A(n11966), .Y(n11964) );
  INVX1 U11929 ( .A(n11964), .Y(n11965) );
  BUFX2 U11930 ( .A(fifo[765]), .Y(n11966) );
  INVX1 U11931 ( .A(n11969), .Y(n11967) );
  INVX1 U11932 ( .A(n11967), .Y(n11968) );
  BUFX2 U11933 ( .A(fifo[766]), .Y(n11969) );
  INVX1 U11934 ( .A(n11972), .Y(n11970) );
  INVX1 U11935 ( .A(n11970), .Y(n11971) );
  BUFX2 U11936 ( .A(fifo[767]), .Y(n11972) );
  INVX1 U11937 ( .A(n11975), .Y(n11973) );
  INVX1 U11938 ( .A(n11973), .Y(n11974) );
  BUFX2 U11939 ( .A(fifo[768]), .Y(n11975) );
  INVX1 U11940 ( .A(n11978), .Y(n11976) );
  INVX1 U11941 ( .A(n11976), .Y(n11977) );
  BUFX2 U11942 ( .A(fifo[769]), .Y(n11978) );
  INVX1 U11943 ( .A(n11981), .Y(n11979) );
  INVX1 U11944 ( .A(n11979), .Y(n11980) );
  BUFX2 U11945 ( .A(fifo[770]), .Y(n11981) );
  INVX1 U11946 ( .A(n11984), .Y(n11982) );
  INVX1 U11947 ( .A(n11982), .Y(n11983) );
  BUFX2 U11948 ( .A(fifo[771]), .Y(n11984) );
  INVX1 U11949 ( .A(n11987), .Y(n11985) );
  INVX1 U11950 ( .A(n11985), .Y(n11986) );
  BUFX2 U11951 ( .A(fifo[772]), .Y(n11987) );
  INVX1 U11952 ( .A(n11990), .Y(n11988) );
  INVX1 U11953 ( .A(n11988), .Y(n11989) );
  BUFX2 U11954 ( .A(fifo[773]), .Y(n11990) );
  INVX1 U11955 ( .A(n11993), .Y(n11991) );
  INVX1 U11956 ( .A(n11991), .Y(n11992) );
  BUFX2 U11957 ( .A(fifo[774]), .Y(n11993) );
  INVX1 U11958 ( .A(n11996), .Y(n11994) );
  INVX1 U11959 ( .A(n11994), .Y(n11995) );
  BUFX2 U11960 ( .A(fifo[775]), .Y(n11996) );
  INVX1 U11961 ( .A(n11999), .Y(n11997) );
  INVX1 U11962 ( .A(n11997), .Y(n11998) );
  BUFX2 U11963 ( .A(fifo[776]), .Y(n11999) );
  INVX1 U11964 ( .A(n12002), .Y(n12000) );
  INVX1 U11965 ( .A(n12000), .Y(n12001) );
  BUFX2 U11966 ( .A(fifo[777]), .Y(n12002) );
  INVX1 U11967 ( .A(n12005), .Y(n12003) );
  INVX1 U11968 ( .A(n12003), .Y(n12004) );
  BUFX2 U11969 ( .A(fifo[778]), .Y(n12005) );
  INVX1 U11970 ( .A(n12008), .Y(n12006) );
  INVX1 U11971 ( .A(n12006), .Y(n12007) );
  BUFX2 U11972 ( .A(fifo[779]), .Y(n12008) );
  INVX1 U11973 ( .A(n12011), .Y(n12009) );
  INVX1 U11974 ( .A(n12009), .Y(n12010) );
  BUFX2 U11975 ( .A(fifo[780]), .Y(n12011) );
  INVX1 U11976 ( .A(n12014), .Y(n12012) );
  INVX1 U11977 ( .A(n12012), .Y(n12013) );
  BUFX2 U11978 ( .A(fifo[781]), .Y(n12014) );
  INVX1 U11979 ( .A(n12017), .Y(n12015) );
  INVX1 U11980 ( .A(n12015), .Y(n12016) );
  BUFX2 U11981 ( .A(fifo[782]), .Y(n12017) );
  INVX1 U11982 ( .A(n12020), .Y(n12018) );
  INVX1 U11983 ( .A(n12018), .Y(n12019) );
  BUFX2 U11984 ( .A(fifo[783]), .Y(n12020) );
  INVX1 U11985 ( .A(n12023), .Y(n12021) );
  INVX1 U11986 ( .A(n12021), .Y(n12022) );
  BUFX2 U11987 ( .A(fifo[784]), .Y(n12023) );
  INVX1 U11988 ( .A(n12026), .Y(n12024) );
  INVX1 U11989 ( .A(n12024), .Y(n12025) );
  BUFX2 U11990 ( .A(fifo[785]), .Y(n12026) );
  INVX1 U11991 ( .A(n12029), .Y(n12027) );
  INVX1 U11992 ( .A(n12027), .Y(n12028) );
  BUFX2 U11993 ( .A(fifo[786]), .Y(n12029) );
  INVX1 U11994 ( .A(n12032), .Y(n12030) );
  INVX1 U11995 ( .A(n12030), .Y(n12031) );
  BUFX2 U11996 ( .A(fifo[787]), .Y(n12032) );
  INVX1 U11997 ( .A(n12035), .Y(n12033) );
  INVX1 U11998 ( .A(n12033), .Y(n12034) );
  BUFX2 U11999 ( .A(fifo[788]), .Y(n12035) );
  INVX1 U12000 ( .A(n12038), .Y(n12036) );
  INVX1 U12001 ( .A(n12036), .Y(n12037) );
  BUFX2 U12002 ( .A(fifo[789]), .Y(n12038) );
  INVX1 U12003 ( .A(n12041), .Y(n12039) );
  INVX1 U12004 ( .A(n12039), .Y(n12040) );
  BUFX2 U12005 ( .A(fifo[790]), .Y(n12041) );
  INVX1 U12006 ( .A(n12044), .Y(n12042) );
  INVX1 U12007 ( .A(n12042), .Y(n12043) );
  BUFX2 U12008 ( .A(fifo[791]), .Y(n12044) );
  INVX1 U12009 ( .A(n12047), .Y(n12045) );
  INVX1 U12010 ( .A(n12045), .Y(n12046) );
  BUFX2 U12011 ( .A(fifo[792]), .Y(n12047) );
  INVX1 U12012 ( .A(n12050), .Y(n12048) );
  INVX1 U12013 ( .A(n12048), .Y(n12049) );
  BUFX2 U12014 ( .A(fifo[793]), .Y(n12050) );
  INVX1 U12015 ( .A(n12053), .Y(n12051) );
  INVX1 U12016 ( .A(n12051), .Y(n12052) );
  BUFX2 U12017 ( .A(fifo[794]), .Y(n12053) );
  INVX1 U12018 ( .A(n12056), .Y(n12054) );
  INVX1 U12019 ( .A(n12054), .Y(n12055) );
  BUFX2 U12020 ( .A(fifo[795]), .Y(n12056) );
  INVX1 U12021 ( .A(n12059), .Y(n12057) );
  INVX1 U12022 ( .A(n12057), .Y(n12058) );
  BUFX2 U12023 ( .A(fifo[796]), .Y(n12059) );
  INVX1 U12024 ( .A(n12062), .Y(n12060) );
  INVX1 U12025 ( .A(n12060), .Y(n12061) );
  BUFX2 U12026 ( .A(fifo[797]), .Y(n12062) );
  INVX1 U12027 ( .A(n12065), .Y(n12063) );
  INVX1 U12028 ( .A(n12063), .Y(n12064) );
  BUFX2 U12029 ( .A(fifo[840]), .Y(n12065) );
  INVX1 U12030 ( .A(n12068), .Y(n12066) );
  INVX1 U12031 ( .A(n12066), .Y(n12067) );
  BUFX2 U12032 ( .A(fifo[841]), .Y(n12068) );
  INVX1 U12033 ( .A(n12071), .Y(n12069) );
  INVX1 U12034 ( .A(n12069), .Y(n12070) );
  BUFX2 U12035 ( .A(fifo[842]), .Y(n12071) );
  INVX1 U12036 ( .A(n12074), .Y(n12072) );
  INVX1 U12037 ( .A(n12072), .Y(n12073) );
  BUFX2 U12038 ( .A(fifo[843]), .Y(n12074) );
  INVX1 U12039 ( .A(n12077), .Y(n12075) );
  INVX1 U12040 ( .A(n12075), .Y(n12076) );
  BUFX2 U12041 ( .A(fifo[844]), .Y(n12077) );
  INVX1 U12042 ( .A(n12080), .Y(n12078) );
  INVX1 U12043 ( .A(n12078), .Y(n12079) );
  BUFX2 U12044 ( .A(fifo[845]), .Y(n12080) );
  INVX1 U12045 ( .A(n12083), .Y(n12081) );
  INVX1 U12046 ( .A(n12081), .Y(n12082) );
  BUFX2 U12047 ( .A(fifo[846]), .Y(n12083) );
  INVX1 U12048 ( .A(n12086), .Y(n12084) );
  INVX1 U12049 ( .A(n12084), .Y(n12085) );
  BUFX2 U12050 ( .A(fifo[847]), .Y(n12086) );
  INVX1 U12051 ( .A(n12089), .Y(n12087) );
  INVX1 U12052 ( .A(n12087), .Y(n12088) );
  BUFX2 U12053 ( .A(fifo[848]), .Y(n12089) );
  INVX1 U12054 ( .A(n12092), .Y(n12090) );
  INVX1 U12055 ( .A(n12090), .Y(n12091) );
  BUFX2 U12056 ( .A(fifo[849]), .Y(n12092) );
  INVX1 U12057 ( .A(n12095), .Y(n12093) );
  INVX1 U12058 ( .A(n12093), .Y(n12094) );
  BUFX2 U12059 ( .A(fifo[850]), .Y(n12095) );
  INVX1 U12060 ( .A(n12098), .Y(n12096) );
  INVX1 U12061 ( .A(n12096), .Y(n12097) );
  BUFX2 U12062 ( .A(fifo[851]), .Y(n12098) );
  INVX1 U12063 ( .A(n12101), .Y(n12099) );
  INVX1 U12064 ( .A(n12099), .Y(n12100) );
  BUFX2 U12065 ( .A(fifo[852]), .Y(n12101) );
  INVX1 U12066 ( .A(n12104), .Y(n12102) );
  INVX1 U12067 ( .A(n12102), .Y(n12103) );
  BUFX2 U12068 ( .A(fifo[853]), .Y(n12104) );
  INVX1 U12069 ( .A(n12107), .Y(n12105) );
  INVX1 U12070 ( .A(n12105), .Y(n12106) );
  BUFX2 U12071 ( .A(fifo[854]), .Y(n12107) );
  INVX1 U12072 ( .A(n12110), .Y(n12108) );
  INVX1 U12073 ( .A(n12108), .Y(n12109) );
  BUFX2 U12074 ( .A(fifo[855]), .Y(n12110) );
  INVX1 U12075 ( .A(n12113), .Y(n12111) );
  INVX1 U12076 ( .A(n12111), .Y(n12112) );
  BUFX2 U12077 ( .A(fifo[856]), .Y(n12113) );
  INVX1 U12078 ( .A(n12116), .Y(n12114) );
  INVX1 U12079 ( .A(n12114), .Y(n12115) );
  BUFX2 U12080 ( .A(fifo[857]), .Y(n12116) );
  INVX1 U12081 ( .A(n12119), .Y(n12117) );
  INVX1 U12082 ( .A(n12117), .Y(n12118) );
  BUFX2 U12083 ( .A(fifo[858]), .Y(n12119) );
  INVX1 U12084 ( .A(n12122), .Y(n12120) );
  INVX1 U12085 ( .A(n12120), .Y(n12121) );
  BUFX2 U12086 ( .A(fifo[859]), .Y(n12122) );
  INVX1 U12087 ( .A(n12125), .Y(n12123) );
  INVX1 U12088 ( .A(n12123), .Y(n12124) );
  BUFX2 U12089 ( .A(fifo[860]), .Y(n12125) );
  INVX1 U12090 ( .A(n12128), .Y(n12126) );
  INVX1 U12091 ( .A(n12126), .Y(n12127) );
  BUFX2 U12092 ( .A(fifo[861]), .Y(n12128) );
  INVX1 U12093 ( .A(n12131), .Y(n12129) );
  INVX1 U12094 ( .A(n12129), .Y(n12130) );
  BUFX2 U12095 ( .A(fifo[862]), .Y(n12131) );
  INVX1 U12096 ( .A(n12134), .Y(n12132) );
  INVX1 U12097 ( .A(n12132), .Y(n12133) );
  BUFX2 U12098 ( .A(fifo[863]), .Y(n12134) );
  INVX1 U12099 ( .A(n12137), .Y(n12135) );
  INVX1 U12100 ( .A(n12135), .Y(n12136) );
  BUFX2 U12101 ( .A(fifo[864]), .Y(n12137) );
  INVX1 U12102 ( .A(n12140), .Y(n12138) );
  INVX1 U12103 ( .A(n12138), .Y(n12139) );
  BUFX2 U12104 ( .A(fifo[865]), .Y(n12140) );
  INVX1 U12105 ( .A(n12143), .Y(n12141) );
  INVX1 U12106 ( .A(n12141), .Y(n12142) );
  BUFX2 U12107 ( .A(fifo[866]), .Y(n12143) );
  INVX1 U12108 ( .A(n12146), .Y(n12144) );
  INVX1 U12109 ( .A(n12144), .Y(n12145) );
  BUFX2 U12110 ( .A(fifo[867]), .Y(n12146) );
  INVX1 U12111 ( .A(n12149), .Y(n12147) );
  INVX1 U12112 ( .A(n12147), .Y(n12148) );
  BUFX2 U12113 ( .A(fifo[868]), .Y(n12149) );
  INVX1 U12114 ( .A(n12152), .Y(n12150) );
  INVX1 U12115 ( .A(n12150), .Y(n12151) );
  BUFX2 U12116 ( .A(fifo[869]), .Y(n12152) );
  INVX1 U12117 ( .A(n12155), .Y(n12153) );
  INVX1 U12118 ( .A(n12153), .Y(n12154) );
  BUFX2 U12119 ( .A(fifo[870]), .Y(n12155) );
  INVX1 U12120 ( .A(n12158), .Y(n12156) );
  INVX1 U12121 ( .A(n12156), .Y(n12157) );
  BUFX2 U12122 ( .A(fifo[871]), .Y(n12158) );
  INVX1 U12123 ( .A(n12161), .Y(n12159) );
  INVX1 U12124 ( .A(n12159), .Y(n12160) );
  BUFX2 U12125 ( .A(fifo[872]), .Y(n12161) );
  INVX1 U12126 ( .A(n12164), .Y(n12162) );
  INVX1 U12127 ( .A(n12162), .Y(n12163) );
  BUFX2 U12128 ( .A(fifo[873]), .Y(n12164) );
  INVX1 U12129 ( .A(n12167), .Y(n12165) );
  INVX1 U12130 ( .A(n12165), .Y(n12166) );
  BUFX2 U12131 ( .A(fifo[874]), .Y(n12167) );
  INVX1 U12132 ( .A(n12170), .Y(n12168) );
  INVX1 U12133 ( .A(n12168), .Y(n12169) );
  BUFX2 U12134 ( .A(fifo[875]), .Y(n12170) );
  INVX1 U12135 ( .A(n12173), .Y(n12171) );
  INVX1 U12136 ( .A(n12171), .Y(n12172) );
  BUFX2 U12137 ( .A(fifo[876]), .Y(n12173) );
  INVX1 U12138 ( .A(n12176), .Y(n12174) );
  INVX1 U12139 ( .A(n12174), .Y(n12175) );
  BUFX2 U12140 ( .A(fifo[877]), .Y(n12176) );
  INVX1 U12141 ( .A(n12179), .Y(n12177) );
  INVX1 U12142 ( .A(n12177), .Y(n12178) );
  BUFX2 U12143 ( .A(fifo[878]), .Y(n12179) );
  INVX1 U12144 ( .A(n12182), .Y(n12180) );
  INVX1 U12145 ( .A(n12180), .Y(n12181) );
  BUFX2 U12146 ( .A(fifo[879]), .Y(n12182) );
  INVX1 U12147 ( .A(n12185), .Y(n12183) );
  INVX1 U12148 ( .A(n12183), .Y(n12184) );
  BUFX2 U12149 ( .A(fifo[880]), .Y(n12185) );
  INVX1 U12150 ( .A(n12188), .Y(n12186) );
  INVX1 U12151 ( .A(n12186), .Y(n12187) );
  BUFX2 U12152 ( .A(fifo[881]), .Y(n12188) );
  INVX1 U12153 ( .A(n12191), .Y(n12189) );
  INVX1 U12154 ( .A(n12189), .Y(n12190) );
  BUFX2 U12155 ( .A(fifo[924]), .Y(n12191) );
  INVX1 U12156 ( .A(n12194), .Y(n12192) );
  INVX1 U12157 ( .A(n12192), .Y(n12193) );
  BUFX2 U12158 ( .A(fifo[925]), .Y(n12194) );
  INVX1 U12159 ( .A(n12197), .Y(n12195) );
  INVX1 U12160 ( .A(n12195), .Y(n12196) );
  BUFX2 U12161 ( .A(fifo[926]), .Y(n12197) );
  INVX1 U12162 ( .A(n12200), .Y(n12198) );
  INVX1 U12163 ( .A(n12198), .Y(n12199) );
  BUFX2 U12164 ( .A(fifo[927]), .Y(n12200) );
  INVX1 U12165 ( .A(n12203), .Y(n12201) );
  INVX1 U12166 ( .A(n12201), .Y(n12202) );
  BUFX2 U12167 ( .A(fifo[928]), .Y(n12203) );
  INVX1 U12168 ( .A(n12206), .Y(n12204) );
  INVX1 U12169 ( .A(n12204), .Y(n12205) );
  BUFX2 U12170 ( .A(fifo[929]), .Y(n12206) );
  INVX1 U12171 ( .A(n12209), .Y(n12207) );
  INVX1 U12172 ( .A(n12207), .Y(n12208) );
  BUFX2 U12173 ( .A(fifo[930]), .Y(n12209) );
  INVX1 U12174 ( .A(n12212), .Y(n12210) );
  INVX1 U12175 ( .A(n12210), .Y(n12211) );
  BUFX2 U12176 ( .A(fifo[931]), .Y(n12212) );
  INVX1 U12177 ( .A(n12215), .Y(n12213) );
  INVX1 U12178 ( .A(n12213), .Y(n12214) );
  BUFX2 U12179 ( .A(fifo[932]), .Y(n12215) );
  INVX1 U12180 ( .A(n12218), .Y(n12216) );
  INVX1 U12181 ( .A(n12216), .Y(n12217) );
  BUFX2 U12182 ( .A(fifo[933]), .Y(n12218) );
  INVX1 U12183 ( .A(n12221), .Y(n12219) );
  INVX1 U12184 ( .A(n12219), .Y(n12220) );
  BUFX2 U12185 ( .A(fifo[934]), .Y(n12221) );
  INVX1 U12186 ( .A(n12224), .Y(n12222) );
  INVX1 U12187 ( .A(n12222), .Y(n12223) );
  BUFX2 U12188 ( .A(fifo[935]), .Y(n12224) );
  INVX1 U12189 ( .A(n12227), .Y(n12225) );
  INVX1 U12190 ( .A(n12225), .Y(n12226) );
  BUFX2 U12191 ( .A(fifo[936]), .Y(n12227) );
  INVX1 U12192 ( .A(n12230), .Y(n12228) );
  INVX1 U12193 ( .A(n12228), .Y(n12229) );
  BUFX2 U12194 ( .A(fifo[937]), .Y(n12230) );
  INVX1 U12195 ( .A(n12233), .Y(n12231) );
  INVX1 U12196 ( .A(n12231), .Y(n12232) );
  BUFX2 U12197 ( .A(fifo[938]), .Y(n12233) );
  INVX1 U12198 ( .A(n12236), .Y(n12234) );
  INVX1 U12199 ( .A(n12234), .Y(n12235) );
  BUFX2 U12200 ( .A(fifo[939]), .Y(n12236) );
  INVX1 U12201 ( .A(n12239), .Y(n12237) );
  INVX1 U12202 ( .A(n12237), .Y(n12238) );
  BUFX2 U12203 ( .A(fifo[940]), .Y(n12239) );
  INVX1 U12204 ( .A(n12242), .Y(n12240) );
  INVX1 U12205 ( .A(n12240), .Y(n12241) );
  BUFX2 U12206 ( .A(fifo[941]), .Y(n12242) );
  INVX1 U12207 ( .A(n12245), .Y(n12243) );
  INVX1 U12208 ( .A(n12243), .Y(n12244) );
  BUFX2 U12209 ( .A(fifo[942]), .Y(n12245) );
  INVX1 U12210 ( .A(n12248), .Y(n12246) );
  INVX1 U12211 ( .A(n12246), .Y(n12247) );
  BUFX2 U12212 ( .A(fifo[943]), .Y(n12248) );
  INVX1 U12213 ( .A(n12251), .Y(n12249) );
  INVX1 U12214 ( .A(n12249), .Y(n12250) );
  BUFX2 U12215 ( .A(fifo[944]), .Y(n12251) );
  INVX1 U12216 ( .A(n12254), .Y(n12252) );
  INVX1 U12217 ( .A(n12252), .Y(n12253) );
  BUFX2 U12218 ( .A(fifo[945]), .Y(n12254) );
  INVX1 U12219 ( .A(n12257), .Y(n12255) );
  INVX1 U12220 ( .A(n12255), .Y(n12256) );
  BUFX2 U12221 ( .A(fifo[946]), .Y(n12257) );
  INVX1 U12222 ( .A(n12260), .Y(n12258) );
  INVX1 U12223 ( .A(n12258), .Y(n12259) );
  BUFX2 U12224 ( .A(fifo[947]), .Y(n12260) );
  INVX1 U12225 ( .A(n12263), .Y(n12261) );
  INVX1 U12226 ( .A(n12261), .Y(n12262) );
  BUFX2 U12227 ( .A(fifo[948]), .Y(n12263) );
  INVX1 U12228 ( .A(n12266), .Y(n12264) );
  INVX1 U12229 ( .A(n12264), .Y(n12265) );
  BUFX2 U12230 ( .A(fifo[949]), .Y(n12266) );
  INVX1 U12231 ( .A(n12269), .Y(n12267) );
  INVX1 U12232 ( .A(n12267), .Y(n12268) );
  BUFX2 U12233 ( .A(fifo[950]), .Y(n12269) );
  INVX1 U12234 ( .A(n12272), .Y(n12270) );
  INVX1 U12235 ( .A(n12270), .Y(n12271) );
  BUFX2 U12236 ( .A(fifo[951]), .Y(n12272) );
  INVX1 U12237 ( .A(n12275), .Y(n12273) );
  INVX1 U12238 ( .A(n12273), .Y(n12274) );
  BUFX2 U12239 ( .A(fifo[952]), .Y(n12275) );
  INVX1 U12240 ( .A(n12278), .Y(n12276) );
  INVX1 U12241 ( .A(n12276), .Y(n12277) );
  BUFX2 U12242 ( .A(fifo[953]), .Y(n12278) );
  INVX1 U12243 ( .A(n12281), .Y(n12279) );
  INVX1 U12244 ( .A(n12279), .Y(n12280) );
  BUFX2 U12245 ( .A(fifo[954]), .Y(n12281) );
  INVX1 U12246 ( .A(n12284), .Y(n12282) );
  INVX1 U12247 ( .A(n12282), .Y(n12283) );
  BUFX2 U12248 ( .A(fifo[955]), .Y(n12284) );
  INVX1 U12249 ( .A(n12287), .Y(n12285) );
  INVX1 U12250 ( .A(n12285), .Y(n12286) );
  BUFX2 U12251 ( .A(fifo[956]), .Y(n12287) );
  INVX1 U12252 ( .A(n12290), .Y(n12288) );
  INVX1 U12253 ( .A(n12288), .Y(n12289) );
  BUFX2 U12254 ( .A(fifo[957]), .Y(n12290) );
  INVX1 U12255 ( .A(n12293), .Y(n12291) );
  INVX1 U12256 ( .A(n12291), .Y(n12292) );
  BUFX2 U12257 ( .A(fifo[958]), .Y(n12293) );
  INVX1 U12258 ( .A(n12296), .Y(n12294) );
  INVX1 U12259 ( .A(n12294), .Y(n12295) );
  BUFX2 U12260 ( .A(fifo[959]), .Y(n12296) );
  INVX1 U12261 ( .A(n12299), .Y(n12297) );
  INVX1 U12262 ( .A(n12297), .Y(n12298) );
  BUFX2 U12263 ( .A(fifo[960]), .Y(n12299) );
  INVX1 U12264 ( .A(n12302), .Y(n12300) );
  INVX1 U12265 ( .A(n12300), .Y(n12301) );
  BUFX2 U12266 ( .A(fifo[961]), .Y(n12302) );
  INVX1 U12267 ( .A(n12305), .Y(n12303) );
  INVX1 U12268 ( .A(n12303), .Y(n12304) );
  BUFX2 U12269 ( .A(fifo[962]), .Y(n12305) );
  INVX1 U12270 ( .A(n12308), .Y(n12306) );
  INVX1 U12271 ( .A(n12306), .Y(n12307) );
  BUFX2 U12272 ( .A(fifo[963]), .Y(n12308) );
  INVX1 U12273 ( .A(n12311), .Y(n12309) );
  INVX1 U12274 ( .A(n12309), .Y(n12310) );
  BUFX2 U12275 ( .A(fifo[964]), .Y(n12311) );
  INVX1 U12276 ( .A(n12314), .Y(n12312) );
  INVX1 U12277 ( .A(n12312), .Y(n12313) );
  BUFX2 U12278 ( .A(fifo[965]), .Y(n12314) );
  INVX1 U12279 ( .A(n12317), .Y(n12315) );
  INVX1 U12280 ( .A(n12315), .Y(n12316) );
  BUFX2 U12281 ( .A(fifo[1008]), .Y(n12317) );
  INVX1 U12282 ( .A(n12320), .Y(n12318) );
  INVX1 U12283 ( .A(n12318), .Y(n12319) );
  BUFX2 U12284 ( .A(fifo[1009]), .Y(n12320) );
  INVX1 U12285 ( .A(n12323), .Y(n12321) );
  INVX1 U12286 ( .A(n12321), .Y(n12322) );
  BUFX2 U12287 ( .A(fifo[1010]), .Y(n12323) );
  INVX1 U12288 ( .A(n12326), .Y(n12324) );
  INVX1 U12289 ( .A(n12324), .Y(n12325) );
  BUFX2 U12290 ( .A(fifo[1011]), .Y(n12326) );
  INVX1 U12291 ( .A(n12329), .Y(n12327) );
  INVX1 U12292 ( .A(n12327), .Y(n12328) );
  BUFX2 U12293 ( .A(fifo[1012]), .Y(n12329) );
  INVX1 U12294 ( .A(n12332), .Y(n12330) );
  INVX1 U12295 ( .A(n12330), .Y(n12331) );
  BUFX2 U12296 ( .A(fifo[1013]), .Y(n12332) );
  INVX1 U12297 ( .A(n12335), .Y(n12333) );
  INVX1 U12298 ( .A(n12333), .Y(n12334) );
  BUFX2 U12299 ( .A(fifo[1014]), .Y(n12335) );
  INVX1 U12300 ( .A(n12338), .Y(n12336) );
  INVX1 U12301 ( .A(n12336), .Y(n12337) );
  BUFX2 U12302 ( .A(fifo[1015]), .Y(n12338) );
  INVX1 U12303 ( .A(n12341), .Y(n12339) );
  INVX1 U12304 ( .A(n12339), .Y(n12340) );
  BUFX2 U12305 ( .A(fifo[1016]), .Y(n12341) );
  INVX1 U12306 ( .A(n12344), .Y(n12342) );
  INVX1 U12307 ( .A(n12342), .Y(n12343) );
  BUFX2 U12308 ( .A(fifo[1017]), .Y(n12344) );
  INVX1 U12309 ( .A(n12347), .Y(n12345) );
  INVX1 U12310 ( .A(n12345), .Y(n12346) );
  BUFX2 U12311 ( .A(fifo[1018]), .Y(n12347) );
  INVX1 U12312 ( .A(n12350), .Y(n12348) );
  INVX1 U12313 ( .A(n12348), .Y(n12349) );
  BUFX2 U12314 ( .A(fifo[1019]), .Y(n12350) );
  INVX1 U12315 ( .A(n12353), .Y(n12351) );
  INVX1 U12316 ( .A(n12351), .Y(n12352) );
  BUFX2 U12317 ( .A(fifo[1020]), .Y(n12353) );
  INVX1 U12318 ( .A(n12356), .Y(n12354) );
  INVX1 U12319 ( .A(n12354), .Y(n12355) );
  BUFX2 U12320 ( .A(fifo[1021]), .Y(n12356) );
  INVX1 U12321 ( .A(n12359), .Y(n12357) );
  INVX1 U12322 ( .A(n12357), .Y(n12358) );
  BUFX2 U12323 ( .A(fifo[1022]), .Y(n12359) );
  INVX1 U12324 ( .A(n12362), .Y(n12360) );
  INVX1 U12325 ( .A(n12360), .Y(n12361) );
  BUFX2 U12326 ( .A(fifo[1023]), .Y(n12362) );
  INVX1 U12327 ( .A(n12365), .Y(n12363) );
  INVX1 U12328 ( .A(n12363), .Y(n12364) );
  BUFX2 U12329 ( .A(fifo[1024]), .Y(n12365) );
  INVX1 U12330 ( .A(n12368), .Y(n12366) );
  INVX1 U12331 ( .A(n12366), .Y(n12367) );
  BUFX2 U12332 ( .A(fifo[1025]), .Y(n12368) );
  INVX1 U12333 ( .A(n12371), .Y(n12369) );
  INVX1 U12334 ( .A(n12369), .Y(n12370) );
  BUFX2 U12335 ( .A(fifo[1026]), .Y(n12371) );
  INVX1 U12336 ( .A(n12374), .Y(n12372) );
  INVX1 U12337 ( .A(n12372), .Y(n12373) );
  BUFX2 U12338 ( .A(fifo[1027]), .Y(n12374) );
  INVX1 U12339 ( .A(n12377), .Y(n12375) );
  INVX1 U12340 ( .A(n12375), .Y(n12376) );
  BUFX2 U12341 ( .A(fifo[1028]), .Y(n12377) );
  INVX1 U12342 ( .A(n12380), .Y(n12378) );
  INVX1 U12343 ( .A(n12378), .Y(n12379) );
  BUFX2 U12344 ( .A(fifo[1029]), .Y(n12380) );
  INVX1 U12345 ( .A(n12383), .Y(n12381) );
  INVX1 U12346 ( .A(n12381), .Y(n12382) );
  BUFX2 U12347 ( .A(fifo[1030]), .Y(n12383) );
  INVX1 U12348 ( .A(n12386), .Y(n12384) );
  INVX1 U12349 ( .A(n12384), .Y(n12385) );
  BUFX2 U12350 ( .A(fifo[1031]), .Y(n12386) );
  INVX1 U12351 ( .A(n12389), .Y(n12387) );
  INVX1 U12352 ( .A(n12387), .Y(n12388) );
  BUFX2 U12353 ( .A(fifo[1032]), .Y(n12389) );
  INVX1 U12354 ( .A(n12392), .Y(n12390) );
  INVX1 U12355 ( .A(n12390), .Y(n12391) );
  BUFX2 U12356 ( .A(fifo[1033]), .Y(n12392) );
  INVX1 U12357 ( .A(n12395), .Y(n12393) );
  INVX1 U12358 ( .A(n12393), .Y(n12394) );
  BUFX2 U12359 ( .A(fifo[1034]), .Y(n12395) );
  INVX1 U12360 ( .A(n12398), .Y(n12396) );
  INVX1 U12361 ( .A(n12396), .Y(n12397) );
  BUFX2 U12362 ( .A(fifo[1035]), .Y(n12398) );
  INVX1 U12363 ( .A(n12401), .Y(n12399) );
  INVX1 U12364 ( .A(n12399), .Y(n12400) );
  BUFX2 U12365 ( .A(fifo[1036]), .Y(n12401) );
  INVX1 U12366 ( .A(n12404), .Y(n12402) );
  INVX1 U12367 ( .A(n12402), .Y(n12403) );
  BUFX2 U12368 ( .A(fifo[1037]), .Y(n12404) );
  INVX1 U12369 ( .A(n12407), .Y(n12405) );
  INVX1 U12370 ( .A(n12405), .Y(n12406) );
  BUFX2 U12371 ( .A(fifo[1038]), .Y(n12407) );
  INVX1 U12372 ( .A(n12410), .Y(n12408) );
  INVX1 U12373 ( .A(n12408), .Y(n12409) );
  BUFX2 U12374 ( .A(fifo[1039]), .Y(n12410) );
  INVX1 U12375 ( .A(n12413), .Y(n12411) );
  INVX1 U12376 ( .A(n12411), .Y(n12412) );
  BUFX2 U12377 ( .A(fifo[1040]), .Y(n12413) );
  INVX1 U12378 ( .A(n12416), .Y(n12414) );
  INVX1 U12379 ( .A(n12414), .Y(n12415) );
  BUFX2 U12380 ( .A(fifo[1041]), .Y(n12416) );
  INVX1 U12381 ( .A(n12419), .Y(n12417) );
  INVX1 U12382 ( .A(n12417), .Y(n12418) );
  BUFX2 U12383 ( .A(fifo[1042]), .Y(n12419) );
  INVX1 U12384 ( .A(n12422), .Y(n12420) );
  INVX1 U12385 ( .A(n12420), .Y(n12421) );
  BUFX2 U12386 ( .A(fifo[1043]), .Y(n12422) );
  INVX1 U12387 ( .A(n12425), .Y(n12423) );
  INVX1 U12388 ( .A(n12423), .Y(n12424) );
  BUFX2 U12389 ( .A(fifo[1044]), .Y(n12425) );
  INVX1 U12390 ( .A(n12428), .Y(n12426) );
  INVX1 U12391 ( .A(n12426), .Y(n12427) );
  BUFX2 U12392 ( .A(fifo[1045]), .Y(n12428) );
  INVX1 U12393 ( .A(n12431), .Y(n12429) );
  INVX1 U12394 ( .A(n12429), .Y(n12430) );
  BUFX2 U12395 ( .A(fifo[1046]), .Y(n12431) );
  INVX1 U12396 ( .A(n12434), .Y(n12432) );
  INVX1 U12397 ( .A(n12432), .Y(n12433) );
  BUFX2 U12398 ( .A(fifo[1047]), .Y(n12434) );
  INVX1 U12399 ( .A(n12437), .Y(n12435) );
  INVX1 U12400 ( .A(n12435), .Y(n12436) );
  BUFX2 U12401 ( .A(fifo[1048]), .Y(n12437) );
  INVX1 U12402 ( .A(n12440), .Y(n12438) );
  INVX1 U12403 ( .A(n12438), .Y(n12439) );
  BUFX2 U12404 ( .A(fifo[1049]), .Y(n12440) );
  INVX1 U12405 ( .A(n12443), .Y(n12441) );
  INVX1 U12406 ( .A(n12441), .Y(n12442) );
  BUFX2 U12407 ( .A(fifo[1092]), .Y(n12443) );
  INVX1 U12408 ( .A(n12446), .Y(n12444) );
  INVX1 U12409 ( .A(n12444), .Y(n12445) );
  BUFX2 U12410 ( .A(fifo[1093]), .Y(n12446) );
  INVX1 U12411 ( .A(n12449), .Y(n12447) );
  INVX1 U12412 ( .A(n12447), .Y(n12448) );
  BUFX2 U12413 ( .A(fifo[1094]), .Y(n12449) );
  INVX1 U12414 ( .A(n12452), .Y(n12450) );
  INVX1 U12415 ( .A(n12450), .Y(n12451) );
  BUFX2 U12416 ( .A(fifo[1095]), .Y(n12452) );
  INVX1 U12417 ( .A(n12455), .Y(n12453) );
  INVX1 U12418 ( .A(n12453), .Y(n12454) );
  BUFX2 U12419 ( .A(fifo[1096]), .Y(n12455) );
  INVX1 U12420 ( .A(n12458), .Y(n12456) );
  INVX1 U12421 ( .A(n12456), .Y(n12457) );
  BUFX2 U12422 ( .A(fifo[1097]), .Y(n12458) );
  INVX1 U12423 ( .A(n12461), .Y(n12459) );
  INVX1 U12424 ( .A(n12459), .Y(n12460) );
  BUFX2 U12425 ( .A(fifo[1098]), .Y(n12461) );
  INVX1 U12426 ( .A(n12464), .Y(n12462) );
  INVX1 U12427 ( .A(n12462), .Y(n12463) );
  BUFX2 U12428 ( .A(fifo[1099]), .Y(n12464) );
  INVX1 U12429 ( .A(n12467), .Y(n12465) );
  INVX1 U12430 ( .A(n12465), .Y(n12466) );
  BUFX2 U12431 ( .A(fifo[1100]), .Y(n12467) );
  INVX1 U12432 ( .A(n12470), .Y(n12468) );
  INVX1 U12433 ( .A(n12468), .Y(n12469) );
  BUFX2 U12434 ( .A(fifo[1101]), .Y(n12470) );
  INVX1 U12435 ( .A(n12473), .Y(n12471) );
  INVX1 U12436 ( .A(n12471), .Y(n12472) );
  BUFX2 U12437 ( .A(fifo[1102]), .Y(n12473) );
  INVX1 U12438 ( .A(n12476), .Y(n12474) );
  INVX1 U12439 ( .A(n12474), .Y(n12475) );
  BUFX2 U12440 ( .A(fifo[1103]), .Y(n12476) );
  INVX1 U12441 ( .A(n12479), .Y(n12477) );
  INVX1 U12442 ( .A(n12477), .Y(n12478) );
  BUFX2 U12443 ( .A(fifo[1104]), .Y(n12479) );
  INVX1 U12444 ( .A(n12482), .Y(n12480) );
  INVX1 U12445 ( .A(n12480), .Y(n12481) );
  BUFX2 U12446 ( .A(fifo[1105]), .Y(n12482) );
  INVX1 U12447 ( .A(n12485), .Y(n12483) );
  INVX1 U12448 ( .A(n12483), .Y(n12484) );
  BUFX2 U12449 ( .A(fifo[1106]), .Y(n12485) );
  INVX1 U12450 ( .A(n12488), .Y(n12486) );
  INVX1 U12451 ( .A(n12486), .Y(n12487) );
  BUFX2 U12452 ( .A(fifo[1107]), .Y(n12488) );
  INVX1 U12453 ( .A(n12491), .Y(n12489) );
  INVX1 U12454 ( .A(n12489), .Y(n12490) );
  BUFX2 U12455 ( .A(fifo[1108]), .Y(n12491) );
  INVX1 U12456 ( .A(n12494), .Y(n12492) );
  INVX1 U12457 ( .A(n12492), .Y(n12493) );
  BUFX2 U12458 ( .A(fifo[1109]), .Y(n12494) );
  INVX1 U12459 ( .A(n12497), .Y(n12495) );
  INVX1 U12460 ( .A(n12495), .Y(n12496) );
  BUFX2 U12461 ( .A(fifo[1110]), .Y(n12497) );
  INVX1 U12462 ( .A(n12500), .Y(n12498) );
  INVX1 U12463 ( .A(n12498), .Y(n12499) );
  BUFX2 U12464 ( .A(fifo[1111]), .Y(n12500) );
  INVX1 U12465 ( .A(n12503), .Y(n12501) );
  INVX1 U12466 ( .A(n12501), .Y(n12502) );
  BUFX2 U12467 ( .A(fifo[1112]), .Y(n12503) );
  INVX1 U12468 ( .A(n12506), .Y(n12504) );
  INVX1 U12469 ( .A(n12504), .Y(n12505) );
  BUFX2 U12470 ( .A(fifo[1113]), .Y(n12506) );
  INVX1 U12471 ( .A(n12509), .Y(n12507) );
  INVX1 U12472 ( .A(n12507), .Y(n12508) );
  BUFX2 U12473 ( .A(fifo[1114]), .Y(n12509) );
  INVX1 U12474 ( .A(n12512), .Y(n12510) );
  INVX1 U12475 ( .A(n12510), .Y(n12511) );
  BUFX2 U12476 ( .A(fifo[1115]), .Y(n12512) );
  INVX1 U12477 ( .A(n12515), .Y(n12513) );
  INVX1 U12478 ( .A(n12513), .Y(n12514) );
  BUFX2 U12479 ( .A(fifo[1116]), .Y(n12515) );
  INVX1 U12480 ( .A(n12518), .Y(n12516) );
  INVX1 U12481 ( .A(n12516), .Y(n12517) );
  BUFX2 U12482 ( .A(fifo[1117]), .Y(n12518) );
  INVX1 U12483 ( .A(n12521), .Y(n12519) );
  INVX1 U12484 ( .A(n12519), .Y(n12520) );
  BUFX2 U12485 ( .A(fifo[1118]), .Y(n12521) );
  INVX1 U12486 ( .A(n12524), .Y(n12522) );
  INVX1 U12487 ( .A(n12522), .Y(n12523) );
  BUFX2 U12488 ( .A(fifo[1119]), .Y(n12524) );
  INVX1 U12489 ( .A(n12527), .Y(n12525) );
  INVX1 U12490 ( .A(n12525), .Y(n12526) );
  BUFX2 U12491 ( .A(fifo[1120]), .Y(n12527) );
  INVX1 U12492 ( .A(n12530), .Y(n12528) );
  INVX1 U12493 ( .A(n12528), .Y(n12529) );
  BUFX2 U12494 ( .A(fifo[1121]), .Y(n12530) );
  INVX1 U12495 ( .A(n12533), .Y(n12531) );
  INVX1 U12496 ( .A(n12531), .Y(n12532) );
  BUFX2 U12497 ( .A(fifo[1122]), .Y(n12533) );
  INVX1 U12498 ( .A(n12536), .Y(n12534) );
  INVX1 U12499 ( .A(n12534), .Y(n12535) );
  BUFX2 U12500 ( .A(fifo[1123]), .Y(n12536) );
  INVX1 U12501 ( .A(n12539), .Y(n12537) );
  INVX1 U12502 ( .A(n12537), .Y(n12538) );
  BUFX2 U12503 ( .A(fifo[1124]), .Y(n12539) );
  INVX1 U12504 ( .A(n12542), .Y(n12540) );
  INVX1 U12505 ( .A(n12540), .Y(n12541) );
  BUFX2 U12506 ( .A(fifo[1125]), .Y(n12542) );
  INVX1 U12507 ( .A(n12545), .Y(n12543) );
  INVX1 U12508 ( .A(n12543), .Y(n12544) );
  BUFX2 U12509 ( .A(fifo[1126]), .Y(n12545) );
  INVX1 U12510 ( .A(n12548), .Y(n12546) );
  INVX1 U12511 ( .A(n12546), .Y(n12547) );
  BUFX2 U12512 ( .A(fifo[1127]), .Y(n12548) );
  INVX1 U12513 ( .A(n12551), .Y(n12549) );
  INVX1 U12514 ( .A(n12549), .Y(n12550) );
  BUFX2 U12515 ( .A(fifo[1128]), .Y(n12551) );
  INVX1 U12516 ( .A(n12554), .Y(n12552) );
  INVX1 U12517 ( .A(n12552), .Y(n12553) );
  BUFX2 U12518 ( .A(fifo[1129]), .Y(n12554) );
  INVX1 U12519 ( .A(n12557), .Y(n12555) );
  INVX1 U12520 ( .A(n12555), .Y(n12556) );
  BUFX2 U12521 ( .A(fifo[1130]), .Y(n12557) );
  INVX1 U12522 ( .A(n12560), .Y(n12558) );
  INVX1 U12523 ( .A(n12558), .Y(n12559) );
  BUFX2 U12524 ( .A(fifo[1131]), .Y(n12560) );
  INVX1 U12525 ( .A(n12563), .Y(n12561) );
  INVX1 U12526 ( .A(n12561), .Y(n12562) );
  BUFX2 U12527 ( .A(fifo[1132]), .Y(n12563) );
  INVX1 U12528 ( .A(n12566), .Y(n12564) );
  INVX1 U12529 ( .A(n12564), .Y(n12565) );
  BUFX2 U12530 ( .A(fifo[1133]), .Y(n12566) );
  INVX1 U12531 ( .A(n12569), .Y(n12567) );
  INVX1 U12532 ( .A(n12567), .Y(n12568) );
  BUFX2 U12533 ( .A(fifo[1176]), .Y(n12569) );
  INVX1 U12534 ( .A(n12572), .Y(n12570) );
  INVX1 U12535 ( .A(n12570), .Y(n12571) );
  BUFX2 U12536 ( .A(fifo[1177]), .Y(n12572) );
  INVX1 U12537 ( .A(n12575), .Y(n12573) );
  INVX1 U12538 ( .A(n12573), .Y(n12574) );
  BUFX2 U12539 ( .A(fifo[1178]), .Y(n12575) );
  INVX1 U12540 ( .A(n12578), .Y(n12576) );
  INVX1 U12541 ( .A(n12576), .Y(n12577) );
  BUFX2 U12542 ( .A(fifo[1179]), .Y(n12578) );
  INVX1 U12543 ( .A(n12581), .Y(n12579) );
  INVX1 U12544 ( .A(n12579), .Y(n12580) );
  BUFX2 U12545 ( .A(fifo[1180]), .Y(n12581) );
  INVX1 U12546 ( .A(n12584), .Y(n12582) );
  INVX1 U12547 ( .A(n12582), .Y(n12583) );
  BUFX2 U12548 ( .A(fifo[1181]), .Y(n12584) );
  INVX1 U12549 ( .A(n12587), .Y(n12585) );
  INVX1 U12550 ( .A(n12585), .Y(n12586) );
  BUFX2 U12551 ( .A(fifo[1182]), .Y(n12587) );
  INVX1 U12552 ( .A(n12590), .Y(n12588) );
  INVX1 U12553 ( .A(n12588), .Y(n12589) );
  BUFX2 U12554 ( .A(fifo[1183]), .Y(n12590) );
  INVX1 U12555 ( .A(n12593), .Y(n12591) );
  INVX1 U12556 ( .A(n12591), .Y(n12592) );
  BUFX2 U12557 ( .A(fifo[1184]), .Y(n12593) );
  INVX1 U12558 ( .A(n12596), .Y(n12594) );
  INVX1 U12559 ( .A(n12594), .Y(n12595) );
  BUFX2 U12560 ( .A(fifo[1185]), .Y(n12596) );
  INVX1 U12561 ( .A(n12599), .Y(n12597) );
  INVX1 U12562 ( .A(n12597), .Y(n12598) );
  BUFX2 U12563 ( .A(fifo[1186]), .Y(n12599) );
  INVX1 U12564 ( .A(n12602), .Y(n12600) );
  INVX1 U12565 ( .A(n12600), .Y(n12601) );
  BUFX2 U12566 ( .A(fifo[1187]), .Y(n12602) );
  INVX1 U12567 ( .A(n12605), .Y(n12603) );
  INVX1 U12568 ( .A(n12603), .Y(n12604) );
  BUFX2 U12569 ( .A(fifo[1188]), .Y(n12605) );
  INVX1 U12570 ( .A(n12608), .Y(n12606) );
  INVX1 U12571 ( .A(n12606), .Y(n12607) );
  BUFX2 U12572 ( .A(fifo[1189]), .Y(n12608) );
  INVX1 U12573 ( .A(n12611), .Y(n12609) );
  INVX1 U12574 ( .A(n12609), .Y(n12610) );
  BUFX2 U12575 ( .A(fifo[1190]), .Y(n12611) );
  INVX1 U12576 ( .A(n12614), .Y(n12612) );
  INVX1 U12577 ( .A(n12612), .Y(n12613) );
  BUFX2 U12578 ( .A(fifo[1191]), .Y(n12614) );
  INVX1 U12579 ( .A(n12617), .Y(n12615) );
  INVX1 U12580 ( .A(n12615), .Y(n12616) );
  BUFX2 U12581 ( .A(fifo[1192]), .Y(n12617) );
  INVX1 U12582 ( .A(n12620), .Y(n12618) );
  INVX1 U12583 ( .A(n12618), .Y(n12619) );
  BUFX2 U12584 ( .A(fifo[1193]), .Y(n12620) );
  INVX1 U12585 ( .A(n12623), .Y(n12621) );
  INVX1 U12586 ( .A(n12621), .Y(n12622) );
  BUFX2 U12587 ( .A(fifo[1194]), .Y(n12623) );
  INVX1 U12588 ( .A(n12626), .Y(n12624) );
  INVX1 U12589 ( .A(n12624), .Y(n12625) );
  BUFX2 U12590 ( .A(fifo[1195]), .Y(n12626) );
  INVX1 U12591 ( .A(n12629), .Y(n12627) );
  INVX1 U12592 ( .A(n12627), .Y(n12628) );
  BUFX2 U12593 ( .A(fifo[1196]), .Y(n12629) );
  INVX1 U12594 ( .A(n12632), .Y(n12630) );
  INVX1 U12595 ( .A(n12630), .Y(n12631) );
  BUFX2 U12596 ( .A(fifo[1197]), .Y(n12632) );
  INVX1 U12597 ( .A(n12635), .Y(n12633) );
  INVX1 U12598 ( .A(n12633), .Y(n12634) );
  BUFX2 U12599 ( .A(fifo[1198]), .Y(n12635) );
  INVX1 U12600 ( .A(n12638), .Y(n12636) );
  INVX1 U12601 ( .A(n12636), .Y(n12637) );
  BUFX2 U12602 ( .A(fifo[1199]), .Y(n12638) );
  INVX1 U12603 ( .A(n12641), .Y(n12639) );
  INVX1 U12604 ( .A(n12639), .Y(n12640) );
  BUFX2 U12605 ( .A(fifo[1200]), .Y(n12641) );
  INVX1 U12606 ( .A(n12644), .Y(n12642) );
  INVX1 U12607 ( .A(n12642), .Y(n12643) );
  BUFX2 U12608 ( .A(fifo[1201]), .Y(n12644) );
  INVX1 U12609 ( .A(n12647), .Y(n12645) );
  INVX1 U12610 ( .A(n12645), .Y(n12646) );
  BUFX2 U12611 ( .A(fifo[1202]), .Y(n12647) );
  INVX1 U12612 ( .A(n12650), .Y(n12648) );
  INVX1 U12613 ( .A(n12648), .Y(n12649) );
  BUFX2 U12614 ( .A(fifo[1203]), .Y(n12650) );
  INVX1 U12615 ( .A(n12653), .Y(n12651) );
  INVX1 U12616 ( .A(n12651), .Y(n12652) );
  BUFX2 U12617 ( .A(fifo[1204]), .Y(n12653) );
  INVX1 U12618 ( .A(n12656), .Y(n12654) );
  INVX1 U12619 ( .A(n12654), .Y(n12655) );
  BUFX2 U12620 ( .A(fifo[1205]), .Y(n12656) );
  INVX1 U12621 ( .A(n12659), .Y(n12657) );
  INVX1 U12622 ( .A(n12657), .Y(n12658) );
  BUFX2 U12623 ( .A(fifo[1206]), .Y(n12659) );
  INVX1 U12624 ( .A(n12662), .Y(n12660) );
  INVX1 U12625 ( .A(n12660), .Y(n12661) );
  BUFX2 U12626 ( .A(fifo[1207]), .Y(n12662) );
  INVX1 U12627 ( .A(n12665), .Y(n12663) );
  INVX1 U12628 ( .A(n12663), .Y(n12664) );
  BUFX2 U12629 ( .A(fifo[1208]), .Y(n12665) );
  INVX1 U12630 ( .A(n12668), .Y(n12666) );
  INVX1 U12631 ( .A(n12666), .Y(n12667) );
  BUFX2 U12632 ( .A(fifo[1209]), .Y(n12668) );
  INVX1 U12633 ( .A(n12671), .Y(n12669) );
  INVX1 U12634 ( .A(n12669), .Y(n12670) );
  BUFX2 U12635 ( .A(fifo[1210]), .Y(n12671) );
  INVX1 U12636 ( .A(n12674), .Y(n12672) );
  INVX1 U12637 ( .A(n12672), .Y(n12673) );
  BUFX2 U12638 ( .A(fifo[1211]), .Y(n12674) );
  INVX1 U12639 ( .A(n12677), .Y(n12675) );
  INVX1 U12640 ( .A(n12675), .Y(n12676) );
  BUFX2 U12641 ( .A(fifo[1212]), .Y(n12677) );
  INVX1 U12642 ( .A(n12680), .Y(n12678) );
  INVX1 U12643 ( .A(n12678), .Y(n12679) );
  BUFX2 U12644 ( .A(fifo[1213]), .Y(n12680) );
  INVX1 U12645 ( .A(n12683), .Y(n12681) );
  INVX1 U12646 ( .A(n12681), .Y(n12682) );
  BUFX2 U12647 ( .A(fifo[1214]), .Y(n12683) );
  INVX1 U12648 ( .A(n12686), .Y(n12684) );
  INVX1 U12649 ( .A(n12684), .Y(n12685) );
  BUFX2 U12650 ( .A(fifo[1215]), .Y(n12686) );
  INVX1 U12651 ( .A(n12689), .Y(n12687) );
  INVX1 U12652 ( .A(n12687), .Y(n12688) );
  BUFX2 U12653 ( .A(fifo[1216]), .Y(n12689) );
  INVX1 U12654 ( .A(n12692), .Y(n12690) );
  INVX1 U12655 ( .A(n12690), .Y(n12691) );
  BUFX2 U12656 ( .A(fifo[1217]), .Y(n12692) );
  INVX1 U12657 ( .A(n12695), .Y(n12693) );
  INVX1 U12658 ( .A(n12693), .Y(n12694) );
  BUFX2 U12659 ( .A(fifo[1260]), .Y(n12695) );
  INVX1 U12660 ( .A(n12698), .Y(n12696) );
  INVX1 U12661 ( .A(n12696), .Y(n12697) );
  BUFX2 U12662 ( .A(fifo[1261]), .Y(n12698) );
  INVX1 U12663 ( .A(n12701), .Y(n12699) );
  INVX1 U12664 ( .A(n12699), .Y(n12700) );
  BUFX2 U12665 ( .A(fifo[1262]), .Y(n12701) );
  INVX1 U12666 ( .A(n12704), .Y(n12702) );
  INVX1 U12667 ( .A(n12702), .Y(n12703) );
  BUFX2 U12668 ( .A(fifo[1263]), .Y(n12704) );
  INVX1 U12669 ( .A(n12707), .Y(n12705) );
  INVX1 U12670 ( .A(n12705), .Y(n12706) );
  BUFX2 U12671 ( .A(fifo[1264]), .Y(n12707) );
  INVX1 U12672 ( .A(n12710), .Y(n12708) );
  INVX1 U12673 ( .A(n12708), .Y(n12709) );
  BUFX2 U12674 ( .A(fifo[1265]), .Y(n12710) );
  INVX1 U12675 ( .A(n12713), .Y(n12711) );
  INVX1 U12676 ( .A(n12711), .Y(n12712) );
  BUFX2 U12677 ( .A(fifo[1266]), .Y(n12713) );
  INVX1 U12678 ( .A(n12716), .Y(n12714) );
  INVX1 U12679 ( .A(n12714), .Y(n12715) );
  BUFX2 U12680 ( .A(fifo[1267]), .Y(n12716) );
  INVX1 U12681 ( .A(n12719), .Y(n12717) );
  INVX1 U12682 ( .A(n12717), .Y(n12718) );
  BUFX2 U12683 ( .A(fifo[1268]), .Y(n12719) );
  INVX1 U12684 ( .A(n12722), .Y(n12720) );
  INVX1 U12685 ( .A(n12720), .Y(n12721) );
  BUFX2 U12686 ( .A(fifo[1269]), .Y(n12722) );
  INVX1 U12687 ( .A(n12725), .Y(n12723) );
  INVX1 U12688 ( .A(n12723), .Y(n12724) );
  BUFX2 U12689 ( .A(fifo[1270]), .Y(n12725) );
  INVX1 U12690 ( .A(n12728), .Y(n12726) );
  INVX1 U12691 ( .A(n12726), .Y(n12727) );
  BUFX2 U12692 ( .A(fifo[1271]), .Y(n12728) );
  INVX1 U12693 ( .A(n12731), .Y(n12729) );
  INVX1 U12694 ( .A(n12729), .Y(n12730) );
  BUFX2 U12695 ( .A(fifo[1272]), .Y(n12731) );
  INVX1 U12696 ( .A(n12734), .Y(n12732) );
  INVX1 U12697 ( .A(n12732), .Y(n12733) );
  BUFX2 U12698 ( .A(fifo[1273]), .Y(n12734) );
  INVX1 U12699 ( .A(n12737), .Y(n12735) );
  INVX1 U12700 ( .A(n12735), .Y(n12736) );
  BUFX2 U12701 ( .A(fifo[1274]), .Y(n12737) );
  INVX1 U12702 ( .A(n12740), .Y(n12738) );
  INVX1 U12703 ( .A(n12738), .Y(n12739) );
  BUFX2 U12704 ( .A(fifo[1275]), .Y(n12740) );
  INVX1 U12705 ( .A(n12743), .Y(n12741) );
  INVX1 U12706 ( .A(n12741), .Y(n12742) );
  BUFX2 U12707 ( .A(fifo[1276]), .Y(n12743) );
  INVX1 U12708 ( .A(n12746), .Y(n12744) );
  INVX1 U12709 ( .A(n12744), .Y(n12745) );
  BUFX2 U12710 ( .A(fifo[1277]), .Y(n12746) );
  INVX1 U12711 ( .A(n12749), .Y(n12747) );
  INVX1 U12712 ( .A(n12747), .Y(n12748) );
  BUFX2 U12713 ( .A(fifo[1278]), .Y(n12749) );
  INVX1 U12714 ( .A(n12752), .Y(n12750) );
  INVX1 U12715 ( .A(n12750), .Y(n12751) );
  BUFX2 U12716 ( .A(fifo[1279]), .Y(n12752) );
  INVX1 U12717 ( .A(n12755), .Y(n12753) );
  INVX1 U12718 ( .A(n12753), .Y(n12754) );
  BUFX2 U12719 ( .A(fifo[1280]), .Y(n12755) );
  INVX1 U12720 ( .A(n12758), .Y(n12756) );
  INVX1 U12721 ( .A(n12756), .Y(n12757) );
  BUFX2 U12722 ( .A(fifo[1281]), .Y(n12758) );
  INVX1 U12723 ( .A(n12761), .Y(n12759) );
  INVX1 U12724 ( .A(n12759), .Y(n12760) );
  BUFX2 U12725 ( .A(fifo[1282]), .Y(n12761) );
  INVX1 U12726 ( .A(n12764), .Y(n12762) );
  INVX1 U12727 ( .A(n12762), .Y(n12763) );
  BUFX2 U12728 ( .A(fifo[1283]), .Y(n12764) );
  INVX1 U12729 ( .A(n12767), .Y(n12765) );
  INVX1 U12730 ( .A(n12765), .Y(n12766) );
  BUFX2 U12731 ( .A(fifo[1284]), .Y(n12767) );
  INVX1 U12732 ( .A(n12770), .Y(n12768) );
  INVX1 U12733 ( .A(n12768), .Y(n12769) );
  BUFX2 U12734 ( .A(fifo[1285]), .Y(n12770) );
  INVX1 U12735 ( .A(n12773), .Y(n12771) );
  INVX1 U12736 ( .A(n12771), .Y(n12772) );
  BUFX2 U12737 ( .A(fifo[1286]), .Y(n12773) );
  INVX1 U12738 ( .A(n12776), .Y(n12774) );
  INVX1 U12739 ( .A(n12774), .Y(n12775) );
  BUFX2 U12740 ( .A(fifo[1287]), .Y(n12776) );
  INVX1 U12741 ( .A(n12779), .Y(n12777) );
  INVX1 U12742 ( .A(n12777), .Y(n12778) );
  BUFX2 U12743 ( .A(fifo[1288]), .Y(n12779) );
  INVX1 U12744 ( .A(n12782), .Y(n12780) );
  INVX1 U12745 ( .A(n12780), .Y(n12781) );
  BUFX2 U12746 ( .A(fifo[1289]), .Y(n12782) );
  INVX1 U12747 ( .A(n12785), .Y(n12783) );
  INVX1 U12748 ( .A(n12783), .Y(n12784) );
  BUFX2 U12749 ( .A(fifo[1290]), .Y(n12785) );
  INVX1 U12750 ( .A(n12788), .Y(n12786) );
  INVX1 U12751 ( .A(n12786), .Y(n12787) );
  BUFX2 U12752 ( .A(fifo[1291]), .Y(n12788) );
  INVX1 U12753 ( .A(n12791), .Y(n12789) );
  INVX1 U12754 ( .A(n12789), .Y(n12790) );
  BUFX2 U12755 ( .A(fifo[1292]), .Y(n12791) );
  INVX1 U12756 ( .A(n12794), .Y(n12792) );
  INVX1 U12757 ( .A(n12792), .Y(n12793) );
  BUFX2 U12758 ( .A(fifo[1293]), .Y(n12794) );
  INVX1 U12759 ( .A(n12797), .Y(n12795) );
  INVX1 U12760 ( .A(n12795), .Y(n12796) );
  BUFX2 U12761 ( .A(fifo[1294]), .Y(n12797) );
  INVX1 U12762 ( .A(n12800), .Y(n12798) );
  INVX1 U12763 ( .A(n12798), .Y(n12799) );
  BUFX2 U12764 ( .A(fifo[1295]), .Y(n12800) );
  INVX1 U12765 ( .A(n12803), .Y(n12801) );
  INVX1 U12766 ( .A(n12801), .Y(n12802) );
  BUFX2 U12767 ( .A(fifo[1296]), .Y(n12803) );
  INVX1 U12768 ( .A(n12806), .Y(n12804) );
  INVX1 U12769 ( .A(n12804), .Y(n12805) );
  BUFX2 U12770 ( .A(fifo[1297]), .Y(n12806) );
  INVX1 U12771 ( .A(n12809), .Y(n12807) );
  INVX1 U12772 ( .A(n12807), .Y(n12808) );
  BUFX2 U12773 ( .A(fifo[1298]), .Y(n12809) );
  INVX1 U12774 ( .A(n12812), .Y(n12810) );
  INVX1 U12775 ( .A(n12810), .Y(n12811) );
  BUFX2 U12776 ( .A(fifo[1299]), .Y(n12812) );
  INVX1 U12777 ( .A(n12815), .Y(n12813) );
  INVX1 U12778 ( .A(n12813), .Y(n12814) );
  BUFX2 U12779 ( .A(fifo[1300]), .Y(n12815) );
  INVX1 U12780 ( .A(n12818), .Y(n12816) );
  INVX1 U12781 ( .A(n12816), .Y(n12817) );
  BUFX2 U12782 ( .A(fifo[1301]), .Y(n12818) );
  INVX1 U12783 ( .A(n12821), .Y(n12819) );
  INVX1 U12784 ( .A(n12819), .Y(data_out[0]) );
  BUFX2 U12785 ( .A(n14723), .Y(n12821) );
  BUFX2 U12786 ( .A(n12), .Y(n12822) );
  INVX1 U12787 ( .A(n12822), .Y(n13282) );
  BUFX2 U12788 ( .A(n11), .Y(n12823) );
  INVX1 U12789 ( .A(n12823), .Y(n13315) );
  BUFX2 U12790 ( .A(n10), .Y(n12824) );
  INVX1 U12791 ( .A(n12824), .Y(n13378) );
  INVX1 U12792 ( .A(n12827), .Y(n12825) );
  INVX1 U12793 ( .A(n12825), .Y(data_out[41]) );
  BUFX2 U12794 ( .A(n14682), .Y(n12827) );
  INVX1 U12795 ( .A(n12830), .Y(n12828) );
  INVX1 U12796 ( .A(n12828), .Y(data_out[40]) );
  BUFX2 U12797 ( .A(n14683), .Y(n12830) );
  INVX1 U12798 ( .A(n12833), .Y(n12831) );
  INVX1 U12799 ( .A(n12831), .Y(data_out[39]) );
  BUFX2 U12800 ( .A(n14684), .Y(n12833) );
  INVX1 U12801 ( .A(n12836), .Y(n12834) );
  INVX1 U12802 ( .A(n12834), .Y(data_out[38]) );
  BUFX2 U12803 ( .A(n14685), .Y(n12836) );
  INVX1 U12804 ( .A(n12839), .Y(n12837) );
  INVX1 U12805 ( .A(n12837), .Y(data_out[37]) );
  BUFX2 U12806 ( .A(n14686), .Y(n12839) );
  INVX1 U12807 ( .A(n12842), .Y(n12840) );
  INVX1 U12808 ( .A(n12840), .Y(data_out[36]) );
  BUFX2 U12809 ( .A(n14687), .Y(n12842) );
  INVX1 U12810 ( .A(n12845), .Y(n12843) );
  INVX1 U12811 ( .A(n12843), .Y(data_out[35]) );
  BUFX2 U12812 ( .A(n14688), .Y(n12845) );
  INVX1 U12813 ( .A(n12848), .Y(n12846) );
  INVX1 U12814 ( .A(n12846), .Y(data_out[34]) );
  BUFX2 U12815 ( .A(n14689), .Y(n12848) );
  INVX1 U12816 ( .A(n12851), .Y(n12849) );
  INVX1 U12817 ( .A(n12849), .Y(data_out[33]) );
  BUFX2 U12818 ( .A(n14690), .Y(n12851) );
  INVX1 U12819 ( .A(n12854), .Y(n12852) );
  INVX1 U12820 ( .A(n12852), .Y(data_out[32]) );
  BUFX2 U12821 ( .A(n14691), .Y(n12854) );
  INVX1 U12822 ( .A(n12857), .Y(n12855) );
  INVX1 U12823 ( .A(n12855), .Y(data_out[31]) );
  BUFX2 U12824 ( .A(n14692), .Y(n12857) );
  INVX1 U12825 ( .A(n12860), .Y(n12858) );
  INVX1 U12826 ( .A(n12858), .Y(data_out[30]) );
  BUFX2 U12827 ( .A(n14693), .Y(n12860) );
  INVX1 U12828 ( .A(n12863), .Y(n12861) );
  INVX1 U12829 ( .A(n12861), .Y(data_out[29]) );
  BUFX2 U12830 ( .A(n14694), .Y(n12863) );
  INVX1 U12831 ( .A(n12866), .Y(n12864) );
  INVX1 U12832 ( .A(n12864), .Y(data_out[28]) );
  BUFX2 U12833 ( .A(n14695), .Y(n12866) );
  INVX1 U12834 ( .A(n12869), .Y(n12867) );
  INVX1 U12835 ( .A(n12867), .Y(data_out[27]) );
  BUFX2 U12836 ( .A(n14696), .Y(n12869) );
  INVX1 U12837 ( .A(n12872), .Y(n12870) );
  INVX1 U12838 ( .A(n12870), .Y(data_out[26]) );
  BUFX2 U12839 ( .A(n14697), .Y(n12872) );
  INVX1 U12840 ( .A(n12875), .Y(n12873) );
  INVX1 U12841 ( .A(n12873), .Y(data_out[25]) );
  BUFX2 U12842 ( .A(n14698), .Y(n12875) );
  INVX1 U12843 ( .A(n12878), .Y(n12876) );
  INVX1 U12844 ( .A(n12876), .Y(data_out[24]) );
  BUFX2 U12845 ( .A(n14699), .Y(n12878) );
  INVX1 U12846 ( .A(n12881), .Y(n12879) );
  INVX1 U12847 ( .A(n12879), .Y(data_out[23]) );
  BUFX2 U12848 ( .A(n14700), .Y(n12881) );
  INVX1 U12849 ( .A(n12884), .Y(n12882) );
  INVX1 U12850 ( .A(n12882), .Y(data_out[22]) );
  BUFX2 U12851 ( .A(n14701), .Y(n12884) );
  INVX1 U12852 ( .A(n12887), .Y(n12885) );
  INVX1 U12853 ( .A(n12885), .Y(data_out[21]) );
  BUFX2 U12854 ( .A(n14702), .Y(n12887) );
  INVX1 U12855 ( .A(n12890), .Y(n12888) );
  INVX1 U12856 ( .A(n12888), .Y(data_out[20]) );
  BUFX2 U12857 ( .A(n14703), .Y(n12890) );
  INVX1 U12858 ( .A(n12893), .Y(n12891) );
  INVX1 U12859 ( .A(n12891), .Y(data_out[19]) );
  BUFX2 U12860 ( .A(n14704), .Y(n12893) );
  INVX1 U12861 ( .A(n12896), .Y(n12894) );
  INVX1 U12862 ( .A(n12894), .Y(data_out[18]) );
  BUFX2 U12863 ( .A(n14705), .Y(n12896) );
  INVX1 U12864 ( .A(n12899), .Y(n12897) );
  INVX1 U12865 ( .A(n12897), .Y(data_out[17]) );
  BUFX2 U12866 ( .A(n14706), .Y(n12899) );
  INVX1 U12867 ( .A(n12902), .Y(n12900) );
  INVX1 U12868 ( .A(n12900), .Y(data_out[16]) );
  BUFX2 U12869 ( .A(n14707), .Y(n12902) );
  INVX1 U12870 ( .A(n12905), .Y(n12903) );
  INVX1 U12871 ( .A(n12903), .Y(data_out[15]) );
  BUFX2 U12872 ( .A(n14708), .Y(n12905) );
  INVX1 U12873 ( .A(n12908), .Y(n12906) );
  INVX1 U12874 ( .A(n12906), .Y(data_out[14]) );
  BUFX2 U12875 ( .A(n14709), .Y(n12908) );
  INVX1 U12876 ( .A(n12911), .Y(n12909) );
  INVX1 U12877 ( .A(n12909), .Y(data_out[13]) );
  BUFX2 U12878 ( .A(n14710), .Y(n12911) );
  INVX1 U12879 ( .A(n12914), .Y(n12912) );
  INVX1 U12880 ( .A(n12912), .Y(data_out[12]) );
  BUFX2 U12881 ( .A(n14711), .Y(n12914) );
  INVX1 U12882 ( .A(n12917), .Y(n12915) );
  INVX1 U12883 ( .A(n12915), .Y(data_out[11]) );
  BUFX2 U12884 ( .A(n14712), .Y(n12917) );
  INVX1 U12885 ( .A(n12920), .Y(n12918) );
  INVX1 U12886 ( .A(n12918), .Y(data_out[10]) );
  BUFX2 U12887 ( .A(n14713), .Y(n12920) );
  INVX1 U12888 ( .A(n12923), .Y(n12921) );
  INVX1 U12889 ( .A(n12921), .Y(data_out[9]) );
  BUFX2 U12890 ( .A(n14714), .Y(n12923) );
  INVX1 U12891 ( .A(n12926), .Y(n12924) );
  INVX1 U12892 ( .A(n12924), .Y(data_out[8]) );
  BUFX2 U12893 ( .A(n14715), .Y(n12926) );
  INVX1 U12894 ( .A(n12929), .Y(n12927) );
  INVX1 U12895 ( .A(n12927), .Y(data_out[7]) );
  BUFX2 U12896 ( .A(n14716), .Y(n12929) );
  INVX1 U12897 ( .A(n12932), .Y(n12930) );
  INVX1 U12898 ( .A(n12930), .Y(data_out[6]) );
  BUFX2 U12899 ( .A(n14717), .Y(n12932) );
  INVX1 U12900 ( .A(n12935), .Y(n12933) );
  INVX1 U12901 ( .A(n12933), .Y(data_out[5]) );
  BUFX2 U12902 ( .A(n14718), .Y(n12935) );
  INVX1 U12903 ( .A(n12938), .Y(n12936) );
  INVX1 U12904 ( .A(n12936), .Y(data_out[4]) );
  BUFX2 U12905 ( .A(n14719), .Y(n12938) );
  INVX1 U12906 ( .A(n12941), .Y(n12939) );
  INVX1 U12907 ( .A(n12939), .Y(data_out[3]) );
  BUFX2 U12908 ( .A(n14720), .Y(n12941) );
  INVX1 U12909 ( .A(n12944), .Y(n12942) );
  INVX1 U12910 ( .A(n12942), .Y(data_out[2]) );
  BUFX2 U12911 ( .A(n14721), .Y(n12944) );
  INVX1 U12912 ( .A(n12947), .Y(n12945) );
  INVX1 U12913 ( .A(n12945), .Y(data_out[1]) );
  BUFX2 U12914 ( .A(n14722), .Y(n12947) );
  INVX1 U12915 ( .A(n12969), .Y(n12948) );
  INVX1 U12916 ( .A(n12948), .Y(n12949) );
  AND2X2 U12917 ( .A(net91816), .B(n68), .Y(net91712) );
  INVX1 U12918 ( .A(net91712), .Y(n12950) );
  INVX1 U12919 ( .A(net91712), .Y(n12951) );
  INVX1 U12920 ( .A(net95822), .Y(n12952) );
  INVX1 U12921 ( .A(n28), .Y(n12953) );
  INVX1 U12922 ( .A(n12956), .Y(n12954) );
  INVX1 U12923 ( .A(n12954), .Y(n12955) );
  AND2X2 U12924 ( .A(n13015), .B(n258), .Y(n1488) );
  INVX1 U12925 ( .A(n1488), .Y(n12956) );
  INVX1 U12926 ( .A(n12959), .Y(n12957) );
  INVX1 U12927 ( .A(n12957), .Y(n12958) );
  AND2X2 U12928 ( .A(n68), .B(n260), .Y(n1575) );
  INVX1 U12929 ( .A(n1575), .Y(n12959) );
  INVX1 U12930 ( .A(n12970), .Y(n12960) );
  INVX1 U12931 ( .A(n12972), .Y(n12961) );
  INVX1 U12932 ( .A(n12974), .Y(n12962) );
  INVX1 U12933 ( .A(n12965), .Y(n12963) );
  INVX1 U12934 ( .A(n12963), .Y(n12964) );
  BUFX2 U12935 ( .A(wr_ptr_gray_ss[5]), .Y(n12965) );
  INVX1 U12936 ( .A(net94528), .Y(n12966) );
  INVX1 U12937 ( .A(n41), .Y(net94528) );
  INVX1 U12938 ( .A(n10795), .Y(n12967) );
  INVX1 U12939 ( .A(n12990), .Y(n12968) );
  INVX1 U12940 ( .A(n12968), .Y(n12969) );
  INVX1 U12941 ( .A(n8752), .Y(n12970) );
  INVX1 U12942 ( .A(n12970), .Y(n12971) );
  INVX1 U12943 ( .A(n665), .Y(n356) );
  INVX1 U12944 ( .A(n8775), .Y(n12972) );
  INVX1 U12945 ( .A(n12972), .Y(n12973) );
  INVX1 U12946 ( .A(n1011), .Y(n709) );
  INVX1 U12947 ( .A(n8772), .Y(n12974) );
  INVX1 U12948 ( .A(n12974), .Y(n12975) );
  INVX1 U12949 ( .A(n1357), .Y(n1055) );
  INVX1 U12950 ( .A(n12979), .Y(n12977) );
  INVX1 U12951 ( .A(n12977), .Y(n12978) );
  BUFX2 U12952 ( .A(wr_ptr_gray_ss[1]), .Y(n12979) );
  INVX1 U12953 ( .A(n12982), .Y(n12980) );
  INVX1 U12954 ( .A(n12980), .Y(n12981) );
  BUFX2 U12955 ( .A(rd_ptr_bin_5_), .Y(n12982) );
  INVX1 U12956 ( .A(n8754), .Y(n12983) );
  INVX1 U12957 ( .A(n12983), .Y(n12984) );
  INVX1 U12958 ( .A(n8756), .Y(n12985) );
  INVX1 U12959 ( .A(n12985), .Y(n12986) );
  INVX1 U12960 ( .A(n1706), .Y(n12987) );
  INVX1 U12961 ( .A(n12987), .Y(n12988) );
  INVX1 U12962 ( .A(n12967), .Y(n12989) );
  INVX1 U12963 ( .A(n12989), .Y(n12990) );
  INVX1 U12964 ( .A(n13032), .Y(n12991) );
  INVX1 U12965 ( .A(n12991), .Y(n12992) );
  INVX1 U12966 ( .A(n12996), .Y(n12993) );
  INVX1 U12967 ( .A(n12993), .Y(n12994) );
  INVX1 U12968 ( .A(n12993), .Y(n12995) );
  BUFX2 U12969 ( .A(wr_ptr_bin[5]), .Y(n12996) );
  INVX1 U12970 ( .A(n12999), .Y(n12997) );
  INVX1 U12971 ( .A(n12997), .Y(n12998) );
  OR2X2 U12972 ( .A(n12958), .B(n13030), .Y(n532) );
  INVX1 U12973 ( .A(n532), .Y(n12999) );
  INVX1 U12974 ( .A(n13002), .Y(n13000) );
  INVX1 U12975 ( .A(n13000), .Y(n13001) );
  OR2X2 U12976 ( .A(n12958), .B(n262), .Y(n576) );
  INVX1 U12977 ( .A(n576), .Y(n13002) );
  INVX1 U12978 ( .A(n13005), .Y(n13003) );
  INVX1 U12979 ( .A(n13003), .Y(n13004) );
  OR2X2 U12980 ( .A(n12955), .B(n262), .Y(n488) );
  INVX1 U12981 ( .A(n488), .Y(n13005) );
  INVX1 U12982 ( .A(n13008), .Y(n13006) );
  INVX1 U12983 ( .A(n13006), .Y(n13007) );
  OR2X2 U12984 ( .A(n12955), .B(n13030), .Y(n444) );
  INVX1 U12985 ( .A(n444), .Y(n13008) );
  INVX1 U12986 ( .A(n13012), .Y(n13009) );
  INVX1 U12987 ( .A(n13009), .Y(n13010) );
  INVX1 U12988 ( .A(n13009), .Y(n13011) );
  BUFX2 U12989 ( .A(wr_ptr_bin[3]), .Y(n13012) );
  INVX1 U12990 ( .A(n13017), .Y(n13013) );
  INVX1 U12991 ( .A(n13013), .Y(n13014) );
  INVX1 U12992 ( .A(n13013), .Y(n13015) );
  INVX1 U12993 ( .A(n13013), .Y(n13016) );
  BUFX2 U12994 ( .A(wr_ptr_bin[1]), .Y(n13017) );
  INVX1 U12995 ( .A(n13023), .Y(n13018) );
  INVX1 U12996 ( .A(n13018), .Y(n13019) );
  INVX1 U12997 ( .A(n13018), .Y(n13020) );
  INVX1 U12998 ( .A(n13018), .Y(n13021) );
  INVX1 U12999 ( .A(n13018), .Y(n13022) );
  BUFX2 U13000 ( .A(wr_ptr_bin[4]), .Y(n13023) );
  INVX1 U13001 ( .A(n13041), .Y(n13024) );
  INVX1 U13002 ( .A(n13037), .Y(n13025) );
  INVX1 U13003 ( .A(n13033), .Y(n13026) );
  INVX1 U13004 ( .A(n13031), .Y(n13027) );
  INVX1 U13005 ( .A(n13027), .Y(n13028) );
  INVX1 U13006 ( .A(n13027), .Y(n13029) );
  INVX1 U13007 ( .A(n13027), .Y(n13030) );
  BUFX2 U13008 ( .A(wr_ptr_bin[0]), .Y(n13031) );
  INVX1 U13009 ( .A(n12989), .Y(n13032) );
  INVX1 U13010 ( .A(n12984), .Y(n13033) );
  INVX1 U13011 ( .A(n13033), .Y(n13034) );
  BUFX2 U13012 ( .A(n8754), .Y(n13035) );
  BUFX2 U13013 ( .A(n8748), .Y(n13036) );
  INVX1 U13014 ( .A(n12986), .Y(n13037) );
  INVX1 U13015 ( .A(n13037), .Y(n13038) );
  BUFX2 U13016 ( .A(n8756), .Y(n13039) );
  BUFX2 U13017 ( .A(n8746), .Y(n13040) );
  INVX1 U13018 ( .A(n12988), .Y(n13041) );
  INVX1 U13019 ( .A(n13041), .Y(n13042) );
  BUFX2 U13020 ( .A(n8750), .Y(n13043) );
  INVX1 U13021 ( .A(n1228), .Y(n13044) );
  INVX1 U13022 ( .A(n13048), .Y(n13046) );
  INVX2 U13023 ( .A(n13046), .Y(n13047) );
  AND2X2 U13024 ( .A(re), .B(empty_bar), .Y(n211) );
  INVX1 U13025 ( .A(n211), .Y(n13048) );
  FAX1 U13026 ( .A(n29), .B(n13050), .C(n13051), .YC(), .YS(n13049) );
  INVX4 U13027 ( .A(net95813), .Y(n13050) );
  INVX1 U13028 ( .A(net95817), .Y(n13051) );
  INVX1 U13029 ( .A(n12953), .Y(net95817) );
  AND2X2 U13030 ( .A(n69), .B(n12951), .Y(n13055) );
  INVX1 U13031 ( .A(net91679), .Y(n13057) );
  INVX1 U13032 ( .A(n13028), .Y(net91711) );
  XOR2X1 U13033 ( .A(net89699), .B(net82058), .Y(fillcount[1]) );
  OAI21X1 U13034 ( .A(net91757), .B(n68), .C(net84771), .Y(net91679) );
  OAI21X1 U13035 ( .A(n12976), .B(n12966), .C(n49), .Y(net84770) );
  OR2X2 U13036 ( .A(fillcount[1]), .B(fillcount[0]), .Y(net92930) );
  AOI21X1 U13037 ( .A(n5), .B(n1), .C(net91715), .Y(net84760) );
  INVX1 U13038 ( .A(net91731), .Y(net91715) );
  NAND3X1 U13039 ( .A(n13055), .B(n63), .C(n61), .Y(net91731) );
  INVX2 U13040 ( .A(net82274), .Y(r301_B_not_0_) );
  INVX1 U13041 ( .A(r301_B_not_0_), .Y(net94575) );
  OR2X2 U13042 ( .A(r301_B_not_0_), .B(n13030), .Y(net89699) );
  INVX8 U13043 ( .A(net80615), .Y(net82259) );
  INVX1 U13044 ( .A(net94575), .Y(net93027) );
  AND2X2 U13045 ( .A(net80615), .B(net84761), .Y(net84769) );
  XNOR2X1 U13046 ( .A(net89715), .B(net84737), .Y(net82058) );
  INVX1 U13047 ( .A(n32), .Y(net84864) );
  INVX1 U13048 ( .A(net84864), .Y(net92912) );
  INVX2 U13049 ( .A(n13014), .Y(net84737) );
  AND2X2 U13050 ( .A(net82274), .B(net91711), .Y(net84723) );
  AOI22X1 U13051 ( .A(net94517), .B(net94519), .C(n8778), .D(net94527), .Y(
        net94530) );
  INVX1 U13052 ( .A(n12950), .Y(net94515) );
  INVX1 U13053 ( .A(n13060), .Y(fillcount[2]) );
  XNOR2X1 U13054 ( .A(net82074), .B(net82060), .Y(n13060) );
  XNOR2X1 U13055 ( .A(net91757), .B(n68), .Y(net82060) );
  INVX1 U13056 ( .A(net91756), .Y(net91757) );
  INVX1 U13057 ( .A(net94543), .Y(net91756) );
  INVX1 U13058 ( .A(net91756), .Y(net91816) );
  OR2X2 U13059 ( .A(net94543), .B(n68), .Y(net91739) );
  INVX1 U13060 ( .A(net82246), .Y(net82074) );
  AOI21X1 U13061 ( .A(net94487), .B(net84723), .C(net92910), .Y(net82246) );
  INVX1 U13062 ( .A(net94574), .Y(net94487) );
  INVX1 U13063 ( .A(net94487), .Y(net94546) );
  OR2X2 U13064 ( .A(n12976), .B(n12966), .Y(net84761) );
  XNOR2X1 U13065 ( .A(net98077), .B(n65), .Y(net98087) );
  BUFX2 U13066 ( .A(n59), .Y(net80878) );
  XNOR2X1 U13067 ( .A(net82107), .B(n12994), .Y(net84863) );
  INVX1 U13068 ( .A(net95813), .Y(net82107) );
  XNOR2X1 U13069 ( .A(net82107), .B(net95818), .Y(net94541) );
  NAND3X1 U13070 ( .A(n196), .B(n8729), .C(n56), .Y(n13064) );
  AOI21X1 U13071 ( .A(net94546), .B(net94553), .C(n13062), .Y(n13061) );
  BUFX2 U13072 ( .A(net91739), .Y(net94553) );
  INVX2 U13073 ( .A(n13049), .Y(net82457) );
  INVX1 U13074 ( .A(net95817), .Y(net95818) );
  AND2X2 U13075 ( .A(net84864), .B(n13015), .Y(net94574) );
  INVX2 U13076 ( .A(n13021), .Y(net94517) );
  INVX2 U13077 ( .A(net94541), .Y(net94519) );
  XNOR2X1 U13078 ( .A(net94541), .B(n13019), .Y(net80615) );
  AND2X2 U13079 ( .A(net94528), .B(n8777), .Y(net94527) );
  INVX1 U13080 ( .A(net84723), .Y(net94521) );
  INVX1 U13081 ( .A(net94515), .Y(net94407) );
  INVX1 U13082 ( .A(n13068), .Y(net82055) );
  OAI21X1 U13083 ( .A(net84723), .B(n55), .C(n13067), .Y(n13068) );
  INVX1 U13084 ( .A(net84771), .Y(net91760) );
  INVX1 U13085 ( .A(net82062), .Y(net82512) );
  XNOR2X1 U13086 ( .A(net82062), .B(net82038), .Y(net82056) );
  INVX1 U13087 ( .A(net82038), .Y(net82147) );
  INVX2 U13088 ( .A(n13010), .Y(net82038) );
  INVX1 U13089 ( .A(n13010), .Y(net82511) );
  INVX1 U13090 ( .A(n4), .Y(net89715) );
  AND2X1 U13091 ( .A(n355), .B(n356), .Y(n13069) );
  INVX8 U13092 ( .A(n13069), .Y(n270) );
  INVX8 U13093 ( .A(n13070), .Y(n577) );
  INVX8 U13094 ( .A(n13071), .Y(n621) );
  INVX8 U13095 ( .A(n13072), .Y(n357) );
  INVX8 U13096 ( .A(n13073), .Y(n445) );
  INVX8 U13097 ( .A(n13074), .Y(n533) );
  INVX8 U13098 ( .A(n13075), .Y(n489) );
  AND2X1 U13099 ( .A(n1401), .B(n355), .Y(n13076) );
  INVX8 U13100 ( .A(n13076), .Y(n1358) );
  AND2X2 U13101 ( .A(n1401), .B(n400), .Y(n13077) );
  INVX8 U13102 ( .A(n13077), .Y(n1402) );
  INVX8 U13103 ( .A(n13078), .Y(n1619) );
  AND2X2 U13104 ( .A(n1401), .B(n664), .Y(n13079) );
  INVX8 U13105 ( .A(n13079), .Y(n1662) );
  INVX8 U13106 ( .A(n13080), .Y(n1445) );
  INVX8 U13107 ( .A(n13081), .Y(n1489) );
  INVX8 U13108 ( .A(n13082), .Y(n1576) );
  AND2X1 U13109 ( .A(n709), .B(n355), .Y(n13083) );
  INVX8 U13110 ( .A(n13083), .Y(n666) );
  AND2X1 U13111 ( .A(n1055), .B(n355), .Y(n13084) );
  INVX8 U13112 ( .A(n13084), .Y(n1012) );
  INVX8 U13113 ( .A(n13085), .Y(n710) );
  INVX8 U13114 ( .A(n13086), .Y(n1056) );
  INVX8 U13115 ( .A(n13087), .Y(n925) );
  INVX8 U13116 ( .A(n13088), .Y(n1271) );
  INVX8 U13117 ( .A(n13089), .Y(n968) );
  INVX8 U13118 ( .A(n13090), .Y(n1314) );
  INVX8 U13119 ( .A(n13091), .Y(n753) );
  INVX8 U13120 ( .A(n13092), .Y(n1099) );
  INVX8 U13121 ( .A(n13093), .Y(n882) );
  INVX8 U13122 ( .A(n13094), .Y(n1142) );
  INVX8 U13123 ( .A(n13095), .Y(n839) );
  INVX8 U13124 ( .A(n13096), .Y(n1185) );
  AND2X2 U13125 ( .A(net84864), .B(n13016), .Y(net84771) );
  XNOR2X1 U13126 ( .A(net93027), .B(n13029), .Y(fillcount[0]) );
  INVX8 U13127 ( .A(net82056), .Y(net84855) );
  INVX1 U13128 ( .A(n14), .Y(n13099) );
  INVX1 U13129 ( .A(n13099), .Y(n13100) );
  INVX1 U13130 ( .A(n13099), .Y(n13101) );
  INVX1 U13131 ( .A(n13030), .Y(net82004) );
  INVX1 U13132 ( .A(net80878), .Y(net80702) );
  INVX1 U13133 ( .A(net80702), .Y(net80703) );
  AND2X2 U13134 ( .A(net80703), .B(we), .Y(n253) );
  INVX1 U13135 ( .A(n13), .Y(n13102) );
  INVX1 U13136 ( .A(n13102), .Y(n13103) );
  INVX2 U13137 ( .A(n13102), .Y(n13104) );
  BUFX4 U13138 ( .A(n13264), .Y(n13105) );
  BUFX4 U13139 ( .A(n13264), .Y(n13106) );
  BUFX4 U13140 ( .A(n13264), .Y(n13107) );
  BUFX4 U13141 ( .A(n13263), .Y(n13108) );
  BUFX4 U13142 ( .A(n13263), .Y(n13109) );
  BUFX4 U13143 ( .A(n13263), .Y(n13110) );
  BUFX4 U13144 ( .A(n13262), .Y(n13111) );
  BUFX4 U13145 ( .A(n13262), .Y(n13112) );
  BUFX4 U13146 ( .A(n13262), .Y(n13113) );
  BUFX4 U13147 ( .A(n13261), .Y(n13114) );
  BUFX4 U13148 ( .A(n13261), .Y(n13115) );
  BUFX4 U13149 ( .A(n13261), .Y(n13116) );
  BUFX4 U13150 ( .A(n13260), .Y(n13117) );
  BUFX4 U13151 ( .A(n13260), .Y(n13118) );
  BUFX4 U13152 ( .A(n13260), .Y(n13119) );
  BUFX4 U13153 ( .A(n13259), .Y(n13120) );
  BUFX4 U13154 ( .A(n13259), .Y(n13121) );
  BUFX4 U13155 ( .A(n13259), .Y(n13122) );
  BUFX4 U13156 ( .A(n13258), .Y(n13123) );
  BUFX4 U13157 ( .A(n13258), .Y(n13124) );
  BUFX4 U13158 ( .A(n13258), .Y(n13125) );
  BUFX4 U13159 ( .A(n13257), .Y(n13126) );
  BUFX4 U13160 ( .A(n13257), .Y(n13127) );
  BUFX4 U13161 ( .A(n13257), .Y(n13128) );
  BUFX4 U13162 ( .A(n13256), .Y(n13129) );
  BUFX4 U13163 ( .A(n13256), .Y(n13130) );
  BUFX4 U13164 ( .A(n13256), .Y(n13131) );
  BUFX4 U13165 ( .A(n13255), .Y(n13132) );
  BUFX4 U13166 ( .A(n13255), .Y(n13133) );
  BUFX4 U13167 ( .A(n13255), .Y(n13134) );
  BUFX4 U13168 ( .A(n13254), .Y(n13135) );
  BUFX4 U13169 ( .A(n13254), .Y(n13136) );
  BUFX4 U13170 ( .A(n13254), .Y(n13137) );
  BUFX4 U13171 ( .A(n13253), .Y(n13138) );
  BUFX4 U13172 ( .A(n13253), .Y(n13139) );
  BUFX4 U13173 ( .A(n13253), .Y(n13140) );
  BUFX4 U13174 ( .A(n13252), .Y(n13141) );
  BUFX4 U13175 ( .A(n13252), .Y(n13142) );
  BUFX4 U13176 ( .A(n13252), .Y(n13143) );
  BUFX4 U13177 ( .A(n13251), .Y(n13144) );
  BUFX4 U13178 ( .A(n13251), .Y(n13145) );
  BUFX4 U13179 ( .A(n13251), .Y(n13146) );
  BUFX4 U13180 ( .A(n13250), .Y(n13147) );
  BUFX4 U13181 ( .A(n13250), .Y(n13148) );
  BUFX4 U13182 ( .A(n13250), .Y(n13149) );
  BUFX4 U13183 ( .A(n13249), .Y(n13150) );
  BUFX4 U13184 ( .A(n13249), .Y(n13151) );
  BUFX4 U13185 ( .A(n13249), .Y(n13152) );
  BUFX4 U13186 ( .A(n13248), .Y(n13153) );
  BUFX4 U13187 ( .A(n13248), .Y(n13154) );
  BUFX4 U13188 ( .A(n13248), .Y(n13155) );
  BUFX4 U13189 ( .A(n13247), .Y(n13156) );
  BUFX4 U13190 ( .A(n13247), .Y(n13157) );
  BUFX4 U13191 ( .A(n13247), .Y(n13158) );
  BUFX4 U13192 ( .A(n13246), .Y(n13159) );
  BUFX4 U13193 ( .A(n13246), .Y(n13160) );
  BUFX4 U13194 ( .A(n13246), .Y(n13161) );
  BUFX4 U13195 ( .A(n13245), .Y(n13162) );
  BUFX4 U13196 ( .A(n13245), .Y(n13163) );
  BUFX4 U13197 ( .A(n13245), .Y(n13164) );
  BUFX4 U13198 ( .A(n13244), .Y(n13165) );
  BUFX4 U13199 ( .A(n13244), .Y(n13166) );
  BUFX4 U13200 ( .A(n13244), .Y(n13167) );
  BUFX4 U13201 ( .A(n13243), .Y(n13168) );
  BUFX4 U13202 ( .A(n13243), .Y(n13169) );
  BUFX4 U13203 ( .A(n13243), .Y(n13170) );
  BUFX4 U13204 ( .A(n13242), .Y(n13171) );
  BUFX4 U13205 ( .A(n13242), .Y(n13172) );
  BUFX4 U13206 ( .A(n13242), .Y(n13173) );
  BUFX4 U13207 ( .A(n13241), .Y(n13174) );
  BUFX4 U13208 ( .A(n13241), .Y(n13175) );
  BUFX4 U13209 ( .A(n13241), .Y(n13176) );
  BUFX4 U13210 ( .A(n13240), .Y(n13177) );
  BUFX4 U13211 ( .A(n13240), .Y(n13178) );
  BUFX4 U13212 ( .A(n13240), .Y(n13179) );
  BUFX4 U13213 ( .A(n13239), .Y(n13180) );
  BUFX4 U13214 ( .A(n13239), .Y(n13181) );
  BUFX4 U13215 ( .A(n13239), .Y(n13182) );
  BUFX4 U13216 ( .A(n13238), .Y(n13183) );
  BUFX4 U13217 ( .A(n13238), .Y(n13184) );
  BUFX4 U13218 ( .A(n13238), .Y(n13185) );
  BUFX4 U13219 ( .A(n13237), .Y(n13186) );
  BUFX4 U13220 ( .A(n13237), .Y(n13187) );
  BUFX4 U13221 ( .A(n13237), .Y(n13188) );
  BUFX4 U13222 ( .A(n13236), .Y(n13189) );
  BUFX4 U13223 ( .A(n13236), .Y(n13190) );
  BUFX4 U13224 ( .A(n13236), .Y(n13191) );
  BUFX4 U13225 ( .A(n13235), .Y(n13192) );
  BUFX4 U13226 ( .A(n13235), .Y(n13193) );
  BUFX4 U13227 ( .A(n13235), .Y(n13194) );
  BUFX4 U13228 ( .A(n13234), .Y(n13195) );
  BUFX4 U13229 ( .A(n13234), .Y(n13196) );
  BUFX4 U13230 ( .A(n13234), .Y(n13197) );
  BUFX4 U13231 ( .A(n13233), .Y(n13198) );
  BUFX4 U13232 ( .A(n13233), .Y(n13199) );
  BUFX4 U13233 ( .A(n13233), .Y(n13200) );
  BUFX4 U13234 ( .A(n13232), .Y(n13201) );
  BUFX4 U13235 ( .A(n13232), .Y(n13202) );
  BUFX4 U13236 ( .A(n13232), .Y(n13203) );
  BUFX4 U13237 ( .A(n13231), .Y(n13204) );
  BUFX4 U13238 ( .A(n13231), .Y(n13205) );
  BUFX4 U13239 ( .A(n13231), .Y(n13206) );
  BUFX4 U13240 ( .A(n13230), .Y(n13207) );
  BUFX4 U13241 ( .A(n13230), .Y(n13208) );
  BUFX4 U13242 ( .A(n13230), .Y(n13209) );
  BUFX4 U13243 ( .A(n13229), .Y(n13210) );
  BUFX4 U13244 ( .A(n13229), .Y(n13211) );
  BUFX4 U13245 ( .A(n13229), .Y(n13212) );
  BUFX4 U13246 ( .A(n13228), .Y(n13213) );
  BUFX4 U13247 ( .A(n13228), .Y(n13214) );
  BUFX4 U13248 ( .A(n13228), .Y(n13215) );
  BUFX4 U13249 ( .A(n13227), .Y(n13216) );
  BUFX4 U13250 ( .A(n13227), .Y(n13217) );
  BUFX4 U13251 ( .A(n13227), .Y(n13218) );
  BUFX4 U13252 ( .A(n13226), .Y(n13219) );
  BUFX4 U13253 ( .A(n13226), .Y(n13220) );
  BUFX4 U13254 ( .A(n13226), .Y(n13221) );
  BUFX4 U13255 ( .A(n13225), .Y(n13222) );
  BUFX4 U13256 ( .A(n13225), .Y(n13223) );
  BUFX4 U13257 ( .A(n13225), .Y(n13224) );
  BUFX4 U13258 ( .A(n3210), .Y(n13225) );
  BUFX4 U13259 ( .A(n3210), .Y(n13226) );
  BUFX4 U13260 ( .A(n3210), .Y(n13227) );
  BUFX4 U13261 ( .A(n3210), .Y(n13228) );
  BUFX4 U13262 ( .A(n3210), .Y(n13229) );
  BUFX4 U13263 ( .A(n3210), .Y(n13230) );
  BUFX4 U13264 ( .A(n3210), .Y(n13231) );
  BUFX4 U13265 ( .A(n3210), .Y(n13232) );
  BUFX4 U13266 ( .A(n3210), .Y(n13233) );
  BUFX4 U13267 ( .A(n3210), .Y(n13234) );
  BUFX4 U13268 ( .A(n3210), .Y(n13235) );
  BUFX4 U13269 ( .A(n3210), .Y(n13236) );
  BUFX4 U13270 ( .A(n3210), .Y(n13237) );
  BUFX4 U13271 ( .A(n3210), .Y(n13238) );
  BUFX4 U13272 ( .A(n3210), .Y(n13239) );
  BUFX4 U13273 ( .A(n3210), .Y(n13240) );
  BUFX4 U13274 ( .A(n3210), .Y(n13241) );
  BUFX4 U13275 ( .A(n3210), .Y(n13242) );
  BUFX4 U13276 ( .A(n3210), .Y(n13243) );
  BUFX4 U13277 ( .A(n3210), .Y(n13244) );
  BUFX4 U13278 ( .A(n3210), .Y(n13245) );
  BUFX4 U13279 ( .A(n3210), .Y(n13246) );
  BUFX4 U13280 ( .A(n3210), .Y(n13247) );
  BUFX4 U13281 ( .A(n3210), .Y(n13248) );
  BUFX4 U13282 ( .A(n3210), .Y(n13249) );
  BUFX4 U13283 ( .A(n3210), .Y(n13250) );
  BUFX4 U13284 ( .A(n3210), .Y(n13251) );
  BUFX4 U13285 ( .A(n3210), .Y(n13252) );
  BUFX4 U13286 ( .A(n3210), .Y(n13253) );
  BUFX4 U13287 ( .A(n3210), .Y(n13254) );
  BUFX4 U13288 ( .A(n3210), .Y(n13255) );
  BUFX4 U13289 ( .A(n3210), .Y(n13256) );
  BUFX4 U13290 ( .A(n3210), .Y(n13257) );
  BUFX4 U13291 ( .A(n3210), .Y(n13258) );
  BUFX4 U13292 ( .A(n3210), .Y(n13259) );
  BUFX4 U13293 ( .A(n3210), .Y(n13260) );
  BUFX4 U13294 ( .A(n3210), .Y(n13261) );
  BUFX4 U13295 ( .A(n3210), .Y(n13262) );
  BUFX4 U13296 ( .A(n3210), .Y(n13263) );
  BUFX4 U13297 ( .A(n3210), .Y(n13264) );
  INVX8 U13298 ( .A(n13276), .Y(n13265) );
  INVX8 U13299 ( .A(n13276), .Y(n13266) );
  INVX8 U13300 ( .A(n13276), .Y(n13267) );
  INVX8 U13301 ( .A(n13277), .Y(n13268) );
  INVX8 U13302 ( .A(n13277), .Y(n13269) );
  INVX8 U13303 ( .A(n13278), .Y(n13270) );
  INVX8 U13304 ( .A(n13278), .Y(n13271) );
  INVX8 U13305 ( .A(n13278), .Y(n13272) );
  INVX8 U13306 ( .A(n13279), .Y(n13273) );
  INVX8 U13307 ( .A(n13279), .Y(n13274) );
  INVX8 U13308 ( .A(n13277), .Y(n13275) );
  INVX8 U13309 ( .A(n13281), .Y(n13276) );
  INVX8 U13310 ( .A(n13280), .Y(n13277) );
  INVX8 U13311 ( .A(n13280), .Y(n13278) );
  INVX8 U13312 ( .A(n13280), .Y(n13279) );
  INVX8 U13313 ( .A(n13282), .Y(n13280) );
  INVX8 U13314 ( .A(n13282), .Y(n13281) );
  INVX8 U13315 ( .A(n13310), .Y(n13283) );
  INVX8 U13316 ( .A(n13310), .Y(n13284) );
  INVX8 U13317 ( .A(n13310), .Y(n13285) );
  INVX8 U13318 ( .A(n13309), .Y(n13286) );
  INVX8 U13319 ( .A(n13309), .Y(n13287) );
  INVX8 U13320 ( .A(n13309), .Y(n13288) );
  INVX8 U13321 ( .A(n13308), .Y(n13289) );
  INVX8 U13322 ( .A(n13308), .Y(n13290) );
  INVX8 U13323 ( .A(n13308), .Y(n13291) );
  INVX8 U13324 ( .A(n13307), .Y(n13292) );
  INVX8 U13325 ( .A(n13307), .Y(n13293) );
  INVX8 U13326 ( .A(n13307), .Y(n13294) );
  INVX8 U13327 ( .A(n13306), .Y(n13295) );
  INVX8 U13328 ( .A(n13306), .Y(n13296) );
  INVX8 U13329 ( .A(n13306), .Y(n13297) );
  INVX8 U13330 ( .A(n13305), .Y(n13298) );
  INVX8 U13331 ( .A(n13305), .Y(n13299) );
  INVX8 U13332 ( .A(n13305), .Y(n13300) );
  INVX8 U13333 ( .A(n13304), .Y(n13301) );
  INVX8 U13334 ( .A(n13304), .Y(n13302) );
  INVX8 U13335 ( .A(n13304), .Y(n13303) );
  INVX8 U13336 ( .A(n13314), .Y(n13304) );
  INVX8 U13337 ( .A(n13314), .Y(n13305) );
  INVX8 U13338 ( .A(n13313), .Y(n13306) );
  INVX8 U13339 ( .A(n13313), .Y(n13307) );
  INVX8 U13340 ( .A(n13313), .Y(n13308) );
  INVX8 U13341 ( .A(n13312), .Y(n13309) );
  INVX8 U13342 ( .A(n13312), .Y(n13310) );
  INVX8 U13343 ( .A(n13312), .Y(n13311) );
  INVX8 U13344 ( .A(n13315), .Y(n13312) );
  INVX8 U13345 ( .A(n13315), .Y(n13313) );
  INVX8 U13346 ( .A(n13315), .Y(n13314) );
  INVX8 U13347 ( .A(n13356), .Y(n13316) );
  INVX8 U13348 ( .A(n13356), .Y(n13317) );
  INVX8 U13349 ( .A(n13357), .Y(n13318) );
  INVX8 U13350 ( .A(n13357), .Y(n13319) );
  INVX8 U13351 ( .A(n13357), .Y(n13320) );
  INVX8 U13352 ( .A(n13358), .Y(n13321) );
  INVX8 U13353 ( .A(n13358), .Y(n13322) );
  INVX8 U13354 ( .A(n13362), .Y(n13323) );
  INVX8 U13355 ( .A(n13358), .Y(n13324) );
  INVX8 U13356 ( .A(n13359), .Y(n13325) );
  INVX8 U13357 ( .A(n13359), .Y(n13326) );
  INVX8 U13358 ( .A(n13359), .Y(n13327) );
  INVX8 U13359 ( .A(n13360), .Y(n13328) );
  INVX8 U13360 ( .A(n13360), .Y(n13329) );
  INVX8 U13361 ( .A(n13360), .Y(n13330) );
  INVX8 U13362 ( .A(n13361), .Y(n13331) );
  INVX8 U13363 ( .A(n13361), .Y(n13332) );
  INVX8 U13364 ( .A(n13361), .Y(n13333) );
  INVX8 U13365 ( .A(n13362), .Y(n13334) );
  INVX8 U13366 ( .A(n13362), .Y(n13335) );
  INVX8 U13367 ( .A(n13363), .Y(n13336) );
  INVX8 U13368 ( .A(n13363), .Y(n13337) );
  INVX8 U13369 ( .A(n13363), .Y(n13338) );
  INVX8 U13370 ( .A(n13364), .Y(n13339) );
  INVX8 U13371 ( .A(n13364), .Y(n13340) );
  INVX8 U13372 ( .A(n13364), .Y(n13341) );
  INVX8 U13373 ( .A(n13365), .Y(n13342) );
  INVX8 U13374 ( .A(n13365), .Y(n13343) );
  INVX8 U13375 ( .A(n13365), .Y(n13344) );
  INVX8 U13376 ( .A(n13366), .Y(n13345) );
  INVX8 U13377 ( .A(n13366), .Y(n13346) );
  INVX8 U13378 ( .A(n13367), .Y(n13347) );
  INVX8 U13379 ( .A(n13367), .Y(n13348) );
  INVX8 U13380 ( .A(n13367), .Y(n13349) );
  INVX8 U13381 ( .A(n13368), .Y(n13350) );
  INVX8 U13382 ( .A(n13368), .Y(n13351) );
  INVX8 U13383 ( .A(n13368), .Y(n13352) );
  INVX8 U13384 ( .A(n13369), .Y(n13353) );
  INVX8 U13385 ( .A(n13366), .Y(n13354) );
  INVX8 U13386 ( .A(n13356), .Y(n13355) );
  INVX8 U13387 ( .A(n13374), .Y(n13356) );
  INVX8 U13388 ( .A(n13374), .Y(n13357) );
  INVX8 U13389 ( .A(n13373), .Y(n13358) );
  INVX8 U13390 ( .A(n13373), .Y(n13359) );
  INVX8 U13391 ( .A(n13373), .Y(n13360) );
  INVX8 U13392 ( .A(n13372), .Y(n13361) );
  INVX8 U13393 ( .A(n13372), .Y(n13362) );
  INVX8 U13394 ( .A(n13372), .Y(n13363) );
  INVX8 U13395 ( .A(n13371), .Y(n13364) );
  INVX8 U13396 ( .A(n13371), .Y(n13365) );
  INVX8 U13397 ( .A(n13371), .Y(n13366) );
  INVX8 U13398 ( .A(n13370), .Y(n13367) );
  INVX8 U13399 ( .A(n13370), .Y(n13368) );
  INVX8 U13400 ( .A(n13370), .Y(n13369) );
  INVX8 U13401 ( .A(n13376), .Y(n13370) );
  INVX8 U13402 ( .A(n13376), .Y(n13371) );
  INVX8 U13403 ( .A(n13375), .Y(n13372) );
  INVX8 U13404 ( .A(n13375), .Y(n13373) );
  INVX8 U13405 ( .A(n13375), .Y(n13374) );
  INVX8 U13406 ( .A(n13377), .Y(n13375) );
  INVX8 U13407 ( .A(n13377), .Y(n13376) );
  INVX8 U13408 ( .A(n13378), .Y(n13377) );
  MUX2X1 U13409 ( .B(n13380), .A(n13381), .S(n13303), .Y(n13379) );
  MUX2X1 U13410 ( .B(n13383), .A(n13384), .S(n13302), .Y(n13382) );
  MUX2X1 U13411 ( .B(n13386), .A(n13387), .S(n13302), .Y(n13385) );
  MUX2X1 U13412 ( .B(n13389), .A(n13390), .S(n13302), .Y(n13388) );
  MUX2X1 U13413 ( .B(n13392), .A(n13393), .S(n13104), .Y(n13391) );
  MUX2X1 U13414 ( .B(n13395), .A(n13396), .S(n13302), .Y(n13394) );
  MUX2X1 U13415 ( .B(n13398), .A(n13399), .S(n13302), .Y(n13397) );
  MUX2X1 U13416 ( .B(n13401), .A(n13402), .S(n13302), .Y(n13400) );
  MUX2X1 U13417 ( .B(n13404), .A(n13405), .S(n13302), .Y(n13403) );
  MUX2X1 U13418 ( .B(n13407), .A(n13408), .S(n13104), .Y(n13406) );
  MUX2X1 U13419 ( .B(n13410), .A(n13411), .S(n13302), .Y(n13409) );
  MUX2X1 U13420 ( .B(n13413), .A(n13414), .S(n13302), .Y(n13412) );
  MUX2X1 U13421 ( .B(n13416), .A(n13417), .S(n13302), .Y(n13415) );
  MUX2X1 U13422 ( .B(n13419), .A(n13420), .S(n13302), .Y(n13418) );
  MUX2X1 U13423 ( .B(n13422), .A(n13423), .S(n13104), .Y(n13421) );
  MUX2X1 U13424 ( .B(n13425), .A(n13426), .S(n13302), .Y(n13424) );
  MUX2X1 U13425 ( .B(n13428), .A(n13429), .S(n13302), .Y(n13427) );
  MUX2X1 U13426 ( .B(n13431), .A(n13432), .S(n13302), .Y(n13430) );
  MUX2X1 U13427 ( .B(n13434), .A(n13435), .S(n13302), .Y(n13433) );
  MUX2X1 U13428 ( .B(n13437), .A(n13438), .S(n13104), .Y(n13436) );
  MUX2X1 U13429 ( .B(n13440), .A(n13441), .S(n13302), .Y(n13439) );
  MUX2X1 U13430 ( .B(n13443), .A(n13444), .S(n13302), .Y(n13442) );
  MUX2X1 U13431 ( .B(n13446), .A(n13447), .S(n13301), .Y(n13445) );
  MUX2X1 U13432 ( .B(n13449), .A(n13450), .S(n13301), .Y(n13448) );
  MUX2X1 U13433 ( .B(n13452), .A(n13453), .S(n13104), .Y(n13451) );
  MUX2X1 U13434 ( .B(n13455), .A(n13456), .S(n13301), .Y(n13454) );
  MUX2X1 U13435 ( .B(n13458), .A(n13459), .S(n13301), .Y(n13457) );
  MUX2X1 U13436 ( .B(n13461), .A(n13462), .S(n13301), .Y(n13460) );
  MUX2X1 U13437 ( .B(n13464), .A(n13465), .S(n13301), .Y(n13463) );
  MUX2X1 U13438 ( .B(n13467), .A(n13468), .S(n13104), .Y(n13466) );
  MUX2X1 U13439 ( .B(n13470), .A(n13471), .S(n13301), .Y(n13469) );
  MUX2X1 U13440 ( .B(n13473), .A(n13474), .S(n13301), .Y(n13472) );
  MUX2X1 U13441 ( .B(n13476), .A(n13477), .S(n13301), .Y(n13475) );
  MUX2X1 U13442 ( .B(n13479), .A(n13480), .S(n13301), .Y(n13478) );
  MUX2X1 U13443 ( .B(n13482), .A(n13483), .S(n13104), .Y(n13481) );
  MUX2X1 U13444 ( .B(n13485), .A(n13486), .S(n13301), .Y(n13484) );
  MUX2X1 U13445 ( .B(n13488), .A(n13489), .S(n13301), .Y(n13487) );
  MUX2X1 U13446 ( .B(n13491), .A(n13492), .S(n13301), .Y(n13490) );
  MUX2X1 U13447 ( .B(n13494), .A(n13495), .S(n13301), .Y(n13493) );
  MUX2X1 U13448 ( .B(n13497), .A(n13498), .S(n13104), .Y(n13496) );
  MUX2X1 U13449 ( .B(n13500), .A(n13501), .S(n13301), .Y(n13499) );
  MUX2X1 U13450 ( .B(n13503), .A(n13504), .S(n13301), .Y(n13502) );
  MUX2X1 U13451 ( .B(n13506), .A(n13507), .S(n13301), .Y(n13505) );
  MUX2X1 U13452 ( .B(n13509), .A(n13510), .S(n13300), .Y(n13508) );
  MUX2X1 U13453 ( .B(n13512), .A(n13513), .S(n13104), .Y(n13511) );
  MUX2X1 U13454 ( .B(n13515), .A(n13516), .S(n13300), .Y(n13514) );
  MUX2X1 U13455 ( .B(n13518), .A(n13519), .S(n13300), .Y(n13517) );
  MUX2X1 U13456 ( .B(n13521), .A(n13522), .S(n13300), .Y(n13520) );
  MUX2X1 U13457 ( .B(n13524), .A(n13525), .S(n13300), .Y(n13523) );
  MUX2X1 U13458 ( .B(n13527), .A(n13528), .S(n13104), .Y(n13526) );
  MUX2X1 U13459 ( .B(n13530), .A(n13531), .S(n13300), .Y(n13529) );
  MUX2X1 U13460 ( .B(n13533), .A(n13534), .S(n13300), .Y(n13532) );
  MUX2X1 U13461 ( .B(n13536), .A(n13537), .S(n13300), .Y(n13535) );
  MUX2X1 U13462 ( .B(n13539), .A(n13540), .S(n13300), .Y(n13538) );
  MUX2X1 U13463 ( .B(n13542), .A(n13543), .S(n13104), .Y(n13541) );
  MUX2X1 U13464 ( .B(n13545), .A(n13546), .S(n13300), .Y(n13544) );
  MUX2X1 U13465 ( .B(n13548), .A(n13549), .S(n13300), .Y(n13547) );
  MUX2X1 U13466 ( .B(n13551), .A(n13552), .S(n13300), .Y(n13550) );
  MUX2X1 U13467 ( .B(n13554), .A(n13555), .S(n13300), .Y(n13553) );
  MUX2X1 U13468 ( .B(n13557), .A(n13558), .S(n13104), .Y(n13556) );
  MUX2X1 U13469 ( .B(n13560), .A(n13561), .S(n13300), .Y(n13559) );
  MUX2X1 U13470 ( .B(n13563), .A(n13564), .S(n13300), .Y(n13562) );
  MUX2X1 U13471 ( .B(n13566), .A(n13567), .S(n13300), .Y(n13565) );
  MUX2X1 U13472 ( .B(n13569), .A(n13570), .S(n13300), .Y(n13568) );
  MUX2X1 U13473 ( .B(n13572), .A(n13573), .S(n13104), .Y(n13571) );
  MUX2X1 U13474 ( .B(n13575), .A(n13576), .S(n13299), .Y(n13574) );
  MUX2X1 U13475 ( .B(n13578), .A(n13579), .S(n13299), .Y(n13577) );
  MUX2X1 U13476 ( .B(n13581), .A(n13582), .S(n13299), .Y(n13580) );
  MUX2X1 U13477 ( .B(n13584), .A(n13585), .S(n13299), .Y(n13583) );
  MUX2X1 U13478 ( .B(n13587), .A(n13588), .S(n13104), .Y(n13586) );
  MUX2X1 U13479 ( .B(n13590), .A(n13591), .S(n13299), .Y(n13589) );
  MUX2X1 U13480 ( .B(n13593), .A(n13594), .S(n13299), .Y(n13592) );
  MUX2X1 U13481 ( .B(n13596), .A(n13597), .S(n13299), .Y(n13595) );
  MUX2X1 U13482 ( .B(n13599), .A(n13600), .S(n13299), .Y(n13598) );
  MUX2X1 U13483 ( .B(n13602), .A(n13603), .S(n13104), .Y(n13601) );
  MUX2X1 U13484 ( .B(n13605), .A(n13606), .S(n13299), .Y(n13604) );
  MUX2X1 U13485 ( .B(n13608), .A(n13609), .S(n13299), .Y(n13607) );
  MUX2X1 U13486 ( .B(n13611), .A(n13612), .S(n13299), .Y(n13610) );
  MUX2X1 U13487 ( .B(n13614), .A(n13615), .S(n13299), .Y(n13613) );
  MUX2X1 U13488 ( .B(n13617), .A(n13618), .S(n13104), .Y(n13616) );
  MUX2X1 U13489 ( .B(n13620), .A(n13621), .S(n13299), .Y(n13619) );
  MUX2X1 U13490 ( .B(n13623), .A(n13624), .S(n13299), .Y(n13622) );
  MUX2X1 U13491 ( .B(n13626), .A(n13627), .S(n13299), .Y(n13625) );
  MUX2X1 U13492 ( .B(n13629), .A(n13630), .S(n13299), .Y(n13628) );
  MUX2X1 U13493 ( .B(n13632), .A(n13633), .S(n13104), .Y(n13631) );
  MUX2X1 U13494 ( .B(n13635), .A(n13636), .S(n13299), .Y(n13634) );
  MUX2X1 U13495 ( .B(n13638), .A(n13639), .S(n13298), .Y(n13637) );
  MUX2X1 U13496 ( .B(n13641), .A(n13642), .S(n13298), .Y(n13640) );
  MUX2X1 U13497 ( .B(n13644), .A(n13645), .S(n13298), .Y(n13643) );
  MUX2X1 U13498 ( .B(n13647), .A(n13648), .S(n13104), .Y(n13646) );
  MUX2X1 U13499 ( .B(n13650), .A(n13651), .S(n13298), .Y(n13649) );
  MUX2X1 U13500 ( .B(n13653), .A(n13654), .S(n13298), .Y(n13652) );
  MUX2X1 U13501 ( .B(n13656), .A(n13657), .S(n13298), .Y(n13655) );
  MUX2X1 U13502 ( .B(n13659), .A(n13660), .S(n13298), .Y(n13658) );
  MUX2X1 U13503 ( .B(n13662), .A(n13663), .S(n13104), .Y(n13661) );
  MUX2X1 U13504 ( .B(n13665), .A(n13666), .S(n13298), .Y(n13664) );
  MUX2X1 U13505 ( .B(n13668), .A(n13669), .S(n13298), .Y(n13667) );
  MUX2X1 U13506 ( .B(n13671), .A(n13672), .S(n13298), .Y(n13670) );
  MUX2X1 U13507 ( .B(n13674), .A(n13675), .S(n13298), .Y(n13673) );
  MUX2X1 U13508 ( .B(n13677), .A(n13678), .S(n13104), .Y(n13676) );
  MUX2X1 U13509 ( .B(n13680), .A(n13681), .S(n13298), .Y(n13679) );
  MUX2X1 U13510 ( .B(n13683), .A(n13684), .S(n13298), .Y(n13682) );
  MUX2X1 U13511 ( .B(n13686), .A(n13687), .S(n13298), .Y(n13685) );
  MUX2X1 U13512 ( .B(n13689), .A(n13690), .S(n13298), .Y(n13688) );
  MUX2X1 U13513 ( .B(n13692), .A(n13693), .S(n13104), .Y(n13691) );
  MUX2X1 U13514 ( .B(n13695), .A(n13696), .S(n13298), .Y(n13694) );
  MUX2X1 U13515 ( .B(n13698), .A(n13699), .S(n13298), .Y(n13697) );
  MUX2X1 U13516 ( .B(n13701), .A(n13702), .S(n13297), .Y(n13700) );
  MUX2X1 U13517 ( .B(n13704), .A(n13705), .S(n13297), .Y(n13703) );
  MUX2X1 U13518 ( .B(n13707), .A(n13708), .S(n13104), .Y(n13706) );
  MUX2X1 U13519 ( .B(n13710), .A(n13711), .S(n13297), .Y(n13709) );
  MUX2X1 U13520 ( .B(n13713), .A(n13714), .S(n13297), .Y(n13712) );
  MUX2X1 U13521 ( .B(n13716), .A(n13717), .S(n13297), .Y(n13715) );
  MUX2X1 U13522 ( .B(n13719), .A(n13720), .S(n13297), .Y(n13718) );
  MUX2X1 U13523 ( .B(n13722), .A(n13723), .S(n13104), .Y(n13721) );
  MUX2X1 U13524 ( .B(n13725), .A(n13726), .S(n13297), .Y(n13724) );
  MUX2X1 U13525 ( .B(n13728), .A(n13729), .S(n13297), .Y(n13727) );
  MUX2X1 U13526 ( .B(n13731), .A(n13732), .S(n13297), .Y(n13730) );
  MUX2X1 U13527 ( .B(n13734), .A(n13735), .S(n13297), .Y(n13733) );
  MUX2X1 U13528 ( .B(n13737), .A(n13738), .S(n13104), .Y(n13736) );
  MUX2X1 U13529 ( .B(n13740), .A(n13741), .S(n13297), .Y(n13739) );
  MUX2X1 U13530 ( .B(n13743), .A(n13744), .S(n13297), .Y(n13742) );
  MUX2X1 U13531 ( .B(n13746), .A(n13747), .S(n13297), .Y(n13745) );
  MUX2X1 U13532 ( .B(n13749), .A(n13750), .S(n13297), .Y(n13748) );
  MUX2X1 U13533 ( .B(n13752), .A(n13753), .S(n13104), .Y(n13751) );
  MUX2X1 U13534 ( .B(n13755), .A(n13756), .S(n13297), .Y(n13754) );
  MUX2X1 U13535 ( .B(n13758), .A(n13759), .S(n13297), .Y(n13757) );
  MUX2X1 U13536 ( .B(n13761), .A(n13762), .S(n13297), .Y(n13760) );
  MUX2X1 U13537 ( .B(n13764), .A(n13765), .S(n13296), .Y(n13763) );
  MUX2X1 U13538 ( .B(n13767), .A(n13768), .S(n13104), .Y(n13766) );
  MUX2X1 U13539 ( .B(n13770), .A(n13771), .S(n13296), .Y(n13769) );
  MUX2X1 U13540 ( .B(n13773), .A(n13774), .S(n13296), .Y(n13772) );
  MUX2X1 U13541 ( .B(n13776), .A(n13777), .S(n13296), .Y(n13775) );
  MUX2X1 U13542 ( .B(n13779), .A(n13780), .S(n13296), .Y(n13778) );
  MUX2X1 U13543 ( .B(n13782), .A(n13783), .S(n13104), .Y(n13781) );
  MUX2X1 U13544 ( .B(n13785), .A(n13786), .S(n13296), .Y(n13784) );
  MUX2X1 U13545 ( .B(n13788), .A(n13789), .S(n13296), .Y(n13787) );
  MUX2X1 U13546 ( .B(n13791), .A(n13792), .S(n13296), .Y(n13790) );
  MUX2X1 U13547 ( .B(n13794), .A(n13795), .S(n13296), .Y(n13793) );
  MUX2X1 U13548 ( .B(n13797), .A(n13798), .S(n13104), .Y(n13796) );
  MUX2X1 U13549 ( .B(n13800), .A(n13801), .S(n13296), .Y(n13799) );
  MUX2X1 U13550 ( .B(n13803), .A(n13804), .S(n13296), .Y(n13802) );
  MUX2X1 U13551 ( .B(n13806), .A(n13807), .S(n13296), .Y(n13805) );
  MUX2X1 U13552 ( .B(n13809), .A(n13810), .S(n13296), .Y(n13808) );
  MUX2X1 U13553 ( .B(n13812), .A(n13813), .S(n13104), .Y(n13811) );
  MUX2X1 U13554 ( .B(n13815), .A(n13816), .S(n13296), .Y(n13814) );
  MUX2X1 U13555 ( .B(n13818), .A(n13819), .S(n13296), .Y(n13817) );
  MUX2X1 U13556 ( .B(n13821), .A(n13822), .S(n13296), .Y(n13820) );
  MUX2X1 U13557 ( .B(n13824), .A(n13825), .S(n13296), .Y(n13823) );
  MUX2X1 U13558 ( .B(n13827), .A(n13828), .S(n13104), .Y(n13826) );
  MUX2X1 U13559 ( .B(n13830), .A(n13831), .S(n13295), .Y(n13829) );
  MUX2X1 U13560 ( .B(n13833), .A(n13834), .S(n13295), .Y(n13832) );
  MUX2X1 U13561 ( .B(n13836), .A(n13837), .S(n13295), .Y(n13835) );
  MUX2X1 U13562 ( .B(n13839), .A(n13840), .S(n13295), .Y(n13838) );
  MUX2X1 U13563 ( .B(n13842), .A(n13843), .S(n13104), .Y(n13841) );
  MUX2X1 U13564 ( .B(n13845), .A(n13846), .S(n13295), .Y(n13844) );
  MUX2X1 U13565 ( .B(n13848), .A(n13849), .S(n13295), .Y(n13847) );
  MUX2X1 U13566 ( .B(n13851), .A(n13852), .S(n13295), .Y(n13850) );
  MUX2X1 U13567 ( .B(n13854), .A(n13855), .S(n13295), .Y(n13853) );
  MUX2X1 U13568 ( .B(n13857), .A(n13858), .S(n13104), .Y(n13856) );
  MUX2X1 U13569 ( .B(n13860), .A(n13861), .S(n13295), .Y(n13859) );
  MUX2X1 U13570 ( .B(n13863), .A(n13864), .S(n13295), .Y(n13862) );
  MUX2X1 U13571 ( .B(n13866), .A(n13867), .S(n13295), .Y(n13865) );
  MUX2X1 U13572 ( .B(n13869), .A(n13870), .S(n13295), .Y(n13868) );
  MUX2X1 U13573 ( .B(n13872), .A(n13873), .S(n13104), .Y(n13871) );
  MUX2X1 U13574 ( .B(n13875), .A(n13876), .S(n13295), .Y(n13874) );
  MUX2X1 U13575 ( .B(n13878), .A(n13879), .S(n13295), .Y(n13877) );
  MUX2X1 U13576 ( .B(n13881), .A(n13882), .S(n13295), .Y(n13880) );
  MUX2X1 U13577 ( .B(n13884), .A(n13885), .S(n13295), .Y(n13883) );
  MUX2X1 U13578 ( .B(n13887), .A(n13888), .S(n13104), .Y(n13886) );
  MUX2X1 U13579 ( .B(n13890), .A(n13891), .S(n13295), .Y(n13889) );
  MUX2X1 U13580 ( .B(n13893), .A(n13894), .S(n13294), .Y(n13892) );
  MUX2X1 U13581 ( .B(n13896), .A(n13897), .S(n13294), .Y(n13895) );
  MUX2X1 U13582 ( .B(n13899), .A(n13900), .S(n13294), .Y(n13898) );
  MUX2X1 U13583 ( .B(n13902), .A(n13903), .S(n13104), .Y(n13901) );
  MUX2X1 U13584 ( .B(n13905), .A(n13906), .S(n13294), .Y(n13904) );
  MUX2X1 U13585 ( .B(n13908), .A(n13909), .S(n13294), .Y(n13907) );
  MUX2X1 U13586 ( .B(n13911), .A(n13912), .S(n13294), .Y(n13910) );
  MUX2X1 U13587 ( .B(n13914), .A(n13915), .S(n13294), .Y(n13913) );
  MUX2X1 U13588 ( .B(n13917), .A(n13918), .S(n13104), .Y(n13916) );
  MUX2X1 U13589 ( .B(n13920), .A(n13921), .S(n13294), .Y(n13919) );
  MUX2X1 U13590 ( .B(n13923), .A(n13924), .S(n13294), .Y(n13922) );
  MUX2X1 U13591 ( .B(n13926), .A(n13927), .S(n13294), .Y(n13925) );
  MUX2X1 U13592 ( .B(n13929), .A(n13930), .S(n13294), .Y(n13928) );
  MUX2X1 U13593 ( .B(n13932), .A(n13933), .S(n13104), .Y(n13931) );
  MUX2X1 U13594 ( .B(n13935), .A(n13936), .S(n13294), .Y(n13934) );
  MUX2X1 U13595 ( .B(n13938), .A(n13939), .S(n13294), .Y(n13937) );
  MUX2X1 U13596 ( .B(n13941), .A(n13942), .S(n13294), .Y(n13940) );
  MUX2X1 U13597 ( .B(n13944), .A(n13945), .S(n13294), .Y(n13943) );
  MUX2X1 U13598 ( .B(n13947), .A(n13948), .S(n13104), .Y(n13946) );
  MUX2X1 U13599 ( .B(n13950), .A(n13951), .S(n13294), .Y(n13949) );
  MUX2X1 U13600 ( .B(n13953), .A(n13954), .S(n13294), .Y(n13952) );
  MUX2X1 U13601 ( .B(n13956), .A(n13957), .S(n13293), .Y(n13955) );
  MUX2X1 U13602 ( .B(n13959), .A(n13960), .S(n13293), .Y(n13958) );
  MUX2X1 U13603 ( .B(n13962), .A(n13963), .S(n13104), .Y(n13961) );
  MUX2X1 U13604 ( .B(n13965), .A(n13966), .S(n13293), .Y(n13964) );
  MUX2X1 U13605 ( .B(n13968), .A(n13969), .S(n13293), .Y(n13967) );
  MUX2X1 U13606 ( .B(n13971), .A(n13972), .S(n13293), .Y(n13970) );
  MUX2X1 U13607 ( .B(n13974), .A(n13975), .S(n13293), .Y(n13973) );
  MUX2X1 U13608 ( .B(n13977), .A(n13978), .S(n13104), .Y(n13976) );
  MUX2X1 U13609 ( .B(n13980), .A(n13981), .S(n13293), .Y(n13979) );
  MUX2X1 U13610 ( .B(n13983), .A(n13984), .S(n13293), .Y(n13982) );
  MUX2X1 U13611 ( .B(n13986), .A(n13987), .S(n13293), .Y(n13985) );
  MUX2X1 U13612 ( .B(n13989), .A(n13990), .S(n13293), .Y(n13988) );
  MUX2X1 U13613 ( .B(n13992), .A(n13993), .S(n13104), .Y(n13991) );
  MUX2X1 U13614 ( .B(n13995), .A(n13996), .S(n13293), .Y(n13994) );
  MUX2X1 U13615 ( .B(n13998), .A(n13999), .S(n13293), .Y(n13997) );
  MUX2X1 U13616 ( .B(n14001), .A(n14002), .S(n13293), .Y(n14000) );
  MUX2X1 U13617 ( .B(n14004), .A(n14005), .S(n13293), .Y(n14003) );
  MUX2X1 U13618 ( .B(n14007), .A(n14008), .S(n13104), .Y(n14006) );
  MUX2X1 U13619 ( .B(n14010), .A(n14011), .S(n13293), .Y(n14009) );
  MUX2X1 U13620 ( .B(n14013), .A(n14014), .S(n13293), .Y(n14012) );
  MUX2X1 U13621 ( .B(n14016), .A(n14017), .S(n13293), .Y(n14015) );
  MUX2X1 U13622 ( .B(n14019), .A(n14020), .S(n13292), .Y(n14018) );
  MUX2X1 U13623 ( .B(n14022), .A(n14023), .S(n13104), .Y(n14021) );
  MUX2X1 U13624 ( .B(n14025), .A(n14026), .S(n13292), .Y(n14024) );
  MUX2X1 U13625 ( .B(n14028), .A(n14029), .S(n13292), .Y(n14027) );
  MUX2X1 U13626 ( .B(n14031), .A(n14032), .S(n13292), .Y(n14030) );
  MUX2X1 U13627 ( .B(n14034), .A(n14035), .S(n13292), .Y(n14033) );
  MUX2X1 U13628 ( .B(n14037), .A(n14038), .S(n13104), .Y(n14036) );
  MUX2X1 U13629 ( .B(n14040), .A(n14041), .S(n13292), .Y(n14039) );
  MUX2X1 U13630 ( .B(n14043), .A(n14044), .S(n13292), .Y(n14042) );
  MUX2X1 U13631 ( .B(n14046), .A(n14047), .S(n13292), .Y(n14045) );
  MUX2X1 U13632 ( .B(n14049), .A(n14050), .S(n13292), .Y(n14048) );
  MUX2X1 U13633 ( .B(n14052), .A(n14053), .S(n13104), .Y(n14051) );
  MUX2X1 U13634 ( .B(n14055), .A(n14056), .S(n13292), .Y(n14054) );
  MUX2X1 U13635 ( .B(n14058), .A(n14059), .S(n13292), .Y(n14057) );
  MUX2X1 U13636 ( .B(n14061), .A(n14062), .S(n13292), .Y(n14060) );
  MUX2X1 U13637 ( .B(n14064), .A(n14065), .S(n13292), .Y(n14063) );
  MUX2X1 U13638 ( .B(n14067), .A(n14068), .S(n13104), .Y(n14066) );
  MUX2X1 U13639 ( .B(n14070), .A(n14071), .S(n13292), .Y(n14069) );
  MUX2X1 U13640 ( .B(n14073), .A(n14074), .S(n13292), .Y(n14072) );
  MUX2X1 U13641 ( .B(n14076), .A(n14077), .S(n13292), .Y(n14075) );
  MUX2X1 U13642 ( .B(n14079), .A(n14080), .S(n13292), .Y(n14078) );
  MUX2X1 U13643 ( .B(n14082), .A(n14083), .S(n13104), .Y(n14081) );
  MUX2X1 U13644 ( .B(n14085), .A(n14086), .S(n13291), .Y(n14084) );
  MUX2X1 U13645 ( .B(n14088), .A(n14089), .S(n13291), .Y(n14087) );
  MUX2X1 U13646 ( .B(n14091), .A(n14092), .S(n13291), .Y(n14090) );
  MUX2X1 U13647 ( .B(n14094), .A(n14095), .S(n13291), .Y(n14093) );
  MUX2X1 U13648 ( .B(n14097), .A(n14098), .S(n13104), .Y(n14096) );
  MUX2X1 U13649 ( .B(n14100), .A(n14101), .S(n13291), .Y(n14099) );
  MUX2X1 U13650 ( .B(n14103), .A(n14104), .S(n13291), .Y(n14102) );
  MUX2X1 U13651 ( .B(n14106), .A(n14107), .S(n13291), .Y(n14105) );
  MUX2X1 U13652 ( .B(n14109), .A(n14110), .S(n13291), .Y(n14108) );
  MUX2X1 U13653 ( .B(n14112), .A(n14113), .S(n13104), .Y(n14111) );
  MUX2X1 U13654 ( .B(n14115), .A(n14116), .S(n13291), .Y(n14114) );
  MUX2X1 U13655 ( .B(n14118), .A(n14119), .S(n13291), .Y(n14117) );
  MUX2X1 U13656 ( .B(n14121), .A(n14122), .S(n13291), .Y(n14120) );
  MUX2X1 U13657 ( .B(n14124), .A(n14125), .S(n13291), .Y(n14123) );
  MUX2X1 U13658 ( .B(n14127), .A(n14128), .S(n13104), .Y(n14126) );
  MUX2X1 U13659 ( .B(n14130), .A(n14131), .S(n13291), .Y(n14129) );
  MUX2X1 U13660 ( .B(n14133), .A(n14134), .S(n13291), .Y(n14132) );
  MUX2X1 U13661 ( .B(n14136), .A(n14137), .S(n13291), .Y(n14135) );
  MUX2X1 U13662 ( .B(n14139), .A(n14140), .S(n13291), .Y(n14138) );
  MUX2X1 U13663 ( .B(n14142), .A(n14143), .S(n13104), .Y(n14141) );
  MUX2X1 U13664 ( .B(n14145), .A(n14146), .S(n13291), .Y(n14144) );
  MUX2X1 U13665 ( .B(n14148), .A(n14149), .S(n13290), .Y(n14147) );
  MUX2X1 U13666 ( .B(n14151), .A(n14152), .S(n13290), .Y(n14150) );
  MUX2X1 U13667 ( .B(n14154), .A(n14155), .S(n13290), .Y(n14153) );
  MUX2X1 U13668 ( .B(n14157), .A(n14158), .S(n13104), .Y(n14156) );
  MUX2X1 U13669 ( .B(n14160), .A(n14161), .S(n13290), .Y(n14159) );
  MUX2X1 U13670 ( .B(n14163), .A(n14164), .S(n13290), .Y(n14162) );
  MUX2X1 U13671 ( .B(n14166), .A(n14167), .S(n13290), .Y(n14165) );
  MUX2X1 U13672 ( .B(n14169), .A(n14170), .S(n13290), .Y(n14168) );
  MUX2X1 U13673 ( .B(n14172), .A(n14173), .S(n13104), .Y(n14171) );
  MUX2X1 U13674 ( .B(n14175), .A(n14176), .S(n13290), .Y(n14174) );
  MUX2X1 U13675 ( .B(n14178), .A(n14179), .S(n13290), .Y(n14177) );
  MUX2X1 U13676 ( .B(n14181), .A(n14182), .S(n13290), .Y(n14180) );
  MUX2X1 U13677 ( .B(n14184), .A(n14185), .S(n13290), .Y(n14183) );
  MUX2X1 U13678 ( .B(n14187), .A(n14188), .S(n13104), .Y(n14186) );
  MUX2X1 U13679 ( .B(n14190), .A(n14191), .S(n13290), .Y(n14189) );
  MUX2X1 U13680 ( .B(n14193), .A(n14194), .S(n13290), .Y(n14192) );
  MUX2X1 U13681 ( .B(n14196), .A(n14197), .S(n13290), .Y(n14195) );
  MUX2X1 U13682 ( .B(n14199), .A(n14200), .S(n13290), .Y(n14198) );
  MUX2X1 U13683 ( .B(n14202), .A(n14203), .S(n13104), .Y(n14201) );
  MUX2X1 U13684 ( .B(n14205), .A(n14206), .S(n13290), .Y(n14204) );
  MUX2X1 U13685 ( .B(n14208), .A(n14209), .S(n13290), .Y(n14207) );
  MUX2X1 U13686 ( .B(n14211), .A(n14212), .S(n13289), .Y(n14210) );
  MUX2X1 U13687 ( .B(n14214), .A(n14215), .S(n13289), .Y(n14213) );
  MUX2X1 U13688 ( .B(n14217), .A(n14218), .S(n13104), .Y(n14216) );
  MUX2X1 U13689 ( .B(n14220), .A(n14221), .S(n13289), .Y(n14219) );
  MUX2X1 U13690 ( .B(n14223), .A(n14224), .S(n13289), .Y(n14222) );
  MUX2X1 U13691 ( .B(n14226), .A(n14227), .S(n13289), .Y(n14225) );
  MUX2X1 U13692 ( .B(n14229), .A(n14230), .S(n13289), .Y(n14228) );
  MUX2X1 U13693 ( .B(n14232), .A(n14233), .S(n13104), .Y(n14231) );
  MUX2X1 U13694 ( .B(n14235), .A(n14236), .S(n13289), .Y(n14234) );
  MUX2X1 U13695 ( .B(n14238), .A(n14239), .S(n13289), .Y(n14237) );
  MUX2X1 U13696 ( .B(n14241), .A(n14242), .S(n13289), .Y(n14240) );
  MUX2X1 U13697 ( .B(n14244), .A(n14245), .S(n13289), .Y(n14243) );
  MUX2X1 U13698 ( .B(n14247), .A(n14248), .S(n13104), .Y(n14246) );
  MUX2X1 U13699 ( .B(n14250), .A(n14251), .S(n13289), .Y(n14249) );
  MUX2X1 U13700 ( .B(n14253), .A(n14254), .S(n13289), .Y(n14252) );
  MUX2X1 U13701 ( .B(n14256), .A(n14257), .S(n13289), .Y(n14255) );
  MUX2X1 U13702 ( .B(n14259), .A(n14260), .S(n13289), .Y(n14258) );
  MUX2X1 U13703 ( .B(n14262), .A(n14263), .S(n13104), .Y(n14261) );
  MUX2X1 U13704 ( .B(n14265), .A(n14266), .S(n13289), .Y(n14264) );
  MUX2X1 U13705 ( .B(n14268), .A(n14269), .S(n13289), .Y(n14267) );
  MUX2X1 U13706 ( .B(n14271), .A(n14272), .S(n13289), .Y(n14270) );
  MUX2X1 U13707 ( .B(n14274), .A(n14275), .S(n13288), .Y(n14273) );
  MUX2X1 U13708 ( .B(n14277), .A(n14278), .S(n13104), .Y(n14276) );
  MUX2X1 U13709 ( .B(n14280), .A(n14281), .S(n13288), .Y(n14279) );
  MUX2X1 U13710 ( .B(n14283), .A(n14284), .S(n13288), .Y(n14282) );
  MUX2X1 U13711 ( .B(n14286), .A(n14287), .S(n13288), .Y(n14285) );
  MUX2X1 U13712 ( .B(n14289), .A(n14290), .S(n13288), .Y(n14288) );
  MUX2X1 U13713 ( .B(n14292), .A(n14293), .S(n13104), .Y(n14291) );
  MUX2X1 U13714 ( .B(n14295), .A(n14296), .S(n13288), .Y(n14294) );
  MUX2X1 U13715 ( .B(n14298), .A(n14299), .S(n13288), .Y(n14297) );
  MUX2X1 U13716 ( .B(n14301), .A(n14302), .S(n13288), .Y(n14300) );
  MUX2X1 U13717 ( .B(n14304), .A(n14305), .S(n13288), .Y(n14303) );
  MUX2X1 U13718 ( .B(n14307), .A(n14308), .S(n13104), .Y(n14306) );
  MUX2X1 U13719 ( .B(n14310), .A(n14311), .S(n13288), .Y(n14309) );
  MUX2X1 U13720 ( .B(n14313), .A(n14314), .S(n13288), .Y(n14312) );
  MUX2X1 U13721 ( .B(n14316), .A(n14317), .S(n13288), .Y(n14315) );
  MUX2X1 U13722 ( .B(n14319), .A(n14320), .S(n13288), .Y(n14318) );
  MUX2X1 U13723 ( .B(n14322), .A(n14323), .S(n13104), .Y(n14321) );
  MUX2X1 U13724 ( .B(n14325), .A(n14326), .S(n13288), .Y(n14324) );
  MUX2X1 U13725 ( .B(n14328), .A(n14329), .S(n13288), .Y(n14327) );
  MUX2X1 U13726 ( .B(n14331), .A(n14332), .S(n13288), .Y(n14330) );
  MUX2X1 U13727 ( .B(n14334), .A(n14335), .S(n13288), .Y(n14333) );
  MUX2X1 U13728 ( .B(n14337), .A(n14338), .S(n13104), .Y(n14336) );
  MUX2X1 U13729 ( .B(n14340), .A(n14341), .S(n13287), .Y(n14339) );
  MUX2X1 U13730 ( .B(n14343), .A(n14344), .S(n13287), .Y(n14342) );
  MUX2X1 U13731 ( .B(n14346), .A(n14347), .S(n13287), .Y(n14345) );
  MUX2X1 U13732 ( .B(n14349), .A(n14350), .S(n13287), .Y(n14348) );
  MUX2X1 U13733 ( .B(n14352), .A(n14353), .S(n13104), .Y(n14351) );
  MUX2X1 U13734 ( .B(n14355), .A(n14356), .S(n13287), .Y(n14354) );
  MUX2X1 U13735 ( .B(n14358), .A(n14359), .S(n13287), .Y(n14357) );
  MUX2X1 U13736 ( .B(n14361), .A(n14362), .S(n13287), .Y(n14360) );
  MUX2X1 U13737 ( .B(n14364), .A(n14365), .S(n13287), .Y(n14363) );
  MUX2X1 U13738 ( .B(n14367), .A(n14368), .S(n13104), .Y(n14366) );
  MUX2X1 U13739 ( .B(n14370), .A(n14371), .S(n13287), .Y(n14369) );
  MUX2X1 U13740 ( .B(n14373), .A(n14374), .S(n13287), .Y(n14372) );
  MUX2X1 U13741 ( .B(n14376), .A(n14377), .S(n13287), .Y(n14375) );
  MUX2X1 U13742 ( .B(n14379), .A(n14380), .S(n13287), .Y(n14378) );
  MUX2X1 U13743 ( .B(n14382), .A(n14383), .S(n13104), .Y(n14381) );
  MUX2X1 U13744 ( .B(n14385), .A(n14386), .S(n13287), .Y(n14384) );
  MUX2X1 U13745 ( .B(n14388), .A(n14389), .S(n13287), .Y(n14387) );
  MUX2X1 U13746 ( .B(n14391), .A(n14392), .S(n13287), .Y(n14390) );
  MUX2X1 U13747 ( .B(n14394), .A(n14395), .S(n13287), .Y(n14393) );
  MUX2X1 U13748 ( .B(n14397), .A(n14398), .S(n13104), .Y(n14396) );
  MUX2X1 U13749 ( .B(n14400), .A(n14401), .S(n13287), .Y(n14399) );
  MUX2X1 U13750 ( .B(n14403), .A(n14404), .S(n13286), .Y(n14402) );
  MUX2X1 U13751 ( .B(n14406), .A(n14407), .S(n13286), .Y(n14405) );
  MUX2X1 U13752 ( .B(n14409), .A(n14410), .S(n13286), .Y(n14408) );
  MUX2X1 U13753 ( .B(n14412), .A(n14413), .S(n13104), .Y(n14411) );
  MUX2X1 U13754 ( .B(n14415), .A(n14416), .S(n13286), .Y(n14414) );
  MUX2X1 U13755 ( .B(n14418), .A(n14419), .S(n13286), .Y(n14417) );
  MUX2X1 U13756 ( .B(n14421), .A(n14422), .S(n13286), .Y(n14420) );
  MUX2X1 U13757 ( .B(n14424), .A(n14425), .S(n13286), .Y(n14423) );
  MUX2X1 U13758 ( .B(n14427), .A(n14428), .S(n13104), .Y(n14426) );
  MUX2X1 U13759 ( .B(n14430), .A(n14431), .S(n13286), .Y(n14429) );
  MUX2X1 U13760 ( .B(n14433), .A(n14434), .S(n13286), .Y(n14432) );
  MUX2X1 U13761 ( .B(n14436), .A(n14437), .S(n13286), .Y(n14435) );
  MUX2X1 U13762 ( .B(n14439), .A(n14440), .S(n13286), .Y(n14438) );
  MUX2X1 U13763 ( .B(n14442), .A(n14443), .S(n13104), .Y(n14441) );
  MUX2X1 U13764 ( .B(n14445), .A(n14446), .S(n13286), .Y(n14444) );
  MUX2X1 U13765 ( .B(n14448), .A(n14449), .S(n13286), .Y(n14447) );
  MUX2X1 U13766 ( .B(n14451), .A(n14452), .S(n13286), .Y(n14450) );
  MUX2X1 U13767 ( .B(n14454), .A(n14455), .S(n13286), .Y(n14453) );
  MUX2X1 U13768 ( .B(n14457), .A(n14458), .S(n13104), .Y(n14456) );
  MUX2X1 U13769 ( .B(n14460), .A(n14461), .S(n13286), .Y(n14459) );
  MUX2X1 U13770 ( .B(n14463), .A(n14464), .S(n13286), .Y(n14462) );
  MUX2X1 U13771 ( .B(n14466), .A(n14467), .S(n13285), .Y(n14465) );
  MUX2X1 U13772 ( .B(n14469), .A(n14470), .S(n13285), .Y(n14468) );
  MUX2X1 U13773 ( .B(n14472), .A(n14473), .S(n13104), .Y(n14471) );
  MUX2X1 U13774 ( .B(n14475), .A(n14476), .S(n13285), .Y(n14474) );
  MUX2X1 U13775 ( .B(n14478), .A(n14479), .S(n13285), .Y(n14477) );
  MUX2X1 U13776 ( .B(n14481), .A(n14482), .S(n13285), .Y(n14480) );
  MUX2X1 U13777 ( .B(n14484), .A(n14485), .S(n13285), .Y(n14483) );
  MUX2X1 U13778 ( .B(n14487), .A(n14488), .S(n13104), .Y(n14486) );
  MUX2X1 U13779 ( .B(n14490), .A(n14491), .S(n13285), .Y(n14489) );
  MUX2X1 U13780 ( .B(n14493), .A(n14494), .S(n13285), .Y(n14492) );
  MUX2X1 U13781 ( .B(n14496), .A(n14497), .S(n13285), .Y(n14495) );
  MUX2X1 U13782 ( .B(n14499), .A(n14500), .S(n13285), .Y(n14498) );
  MUX2X1 U13783 ( .B(n14502), .A(n14503), .S(n13104), .Y(n14501) );
  MUX2X1 U13784 ( .B(n14505), .A(n14506), .S(n13285), .Y(n14504) );
  MUX2X1 U13785 ( .B(n14508), .A(n14509), .S(n13285), .Y(n14507) );
  MUX2X1 U13786 ( .B(n14511), .A(n14512), .S(n13285), .Y(n14510) );
  MUX2X1 U13787 ( .B(n14514), .A(n14515), .S(n13285), .Y(n14513) );
  MUX2X1 U13788 ( .B(n14517), .A(n14518), .S(n13104), .Y(n14516) );
  MUX2X1 U13789 ( .B(n14520), .A(n14521), .S(n13285), .Y(n14519) );
  MUX2X1 U13790 ( .B(n14523), .A(n14524), .S(n13285), .Y(n14522) );
  MUX2X1 U13791 ( .B(n14526), .A(n14527), .S(n13285), .Y(n14525) );
  MUX2X1 U13792 ( .B(n14529), .A(n14530), .S(n13284), .Y(n14528) );
  MUX2X1 U13793 ( .B(n14532), .A(n14533), .S(n13104), .Y(n14531) );
  MUX2X1 U13794 ( .B(n14535), .A(n14536), .S(n13284), .Y(n14534) );
  MUX2X1 U13795 ( .B(n14538), .A(n14539), .S(n13284), .Y(n14537) );
  MUX2X1 U13796 ( .B(n14541), .A(n14542), .S(n13284), .Y(n14540) );
  MUX2X1 U13797 ( .B(n14544), .A(n14545), .S(n13284), .Y(n14543) );
  MUX2X1 U13798 ( .B(n14547), .A(n14548), .S(n13104), .Y(n14546) );
  MUX2X1 U13799 ( .B(n14550), .A(n14551), .S(n13284), .Y(n14549) );
  MUX2X1 U13800 ( .B(n14553), .A(n14554), .S(n13284), .Y(n14552) );
  MUX2X1 U13801 ( .B(n14556), .A(n14557), .S(n13284), .Y(n14555) );
  MUX2X1 U13802 ( .B(n14559), .A(n14560), .S(n13284), .Y(n14558) );
  MUX2X1 U13803 ( .B(n14562), .A(n14563), .S(n13104), .Y(n14561) );
  MUX2X1 U13804 ( .B(n14565), .A(n14566), .S(n13284), .Y(n14564) );
  MUX2X1 U13805 ( .B(n14568), .A(n14569), .S(n13284), .Y(n14567) );
  MUX2X1 U13806 ( .B(n14571), .A(n14572), .S(n13284), .Y(n14570) );
  MUX2X1 U13807 ( .B(n14574), .A(n14575), .S(n13284), .Y(n14573) );
  MUX2X1 U13808 ( .B(n14577), .A(n14578), .S(n13104), .Y(n14576) );
  MUX2X1 U13809 ( .B(n14580), .A(n14581), .S(n13284), .Y(n14579) );
  MUX2X1 U13810 ( .B(n14583), .A(n14584), .S(n13284), .Y(n14582) );
  MUX2X1 U13811 ( .B(n14586), .A(n14587), .S(n13284), .Y(n14585) );
  MUX2X1 U13812 ( .B(n14589), .A(n14590), .S(n13284), .Y(n14588) );
  MUX2X1 U13813 ( .B(n14592), .A(n14593), .S(n13104), .Y(n14591) );
  MUX2X1 U13814 ( .B(n14595), .A(n14596), .S(n13283), .Y(n14594) );
  MUX2X1 U13815 ( .B(n14598), .A(n14599), .S(n13283), .Y(n14597) );
  MUX2X1 U13816 ( .B(n14601), .A(n14602), .S(n13283), .Y(n14600) );
  MUX2X1 U13817 ( .B(n14604), .A(n14605), .S(n13283), .Y(n14603) );
  MUX2X1 U13818 ( .B(n14607), .A(n14608), .S(n13104), .Y(n14606) );
  MUX2X1 U13819 ( .B(n14610), .A(n14611), .S(n13283), .Y(n14609) );
  MUX2X1 U13820 ( .B(n14613), .A(n14614), .S(n13283), .Y(n14612) );
  MUX2X1 U13821 ( .B(n14616), .A(n14617), .S(n13283), .Y(n14615) );
  MUX2X1 U13822 ( .B(n14619), .A(n14620), .S(n13283), .Y(n14618) );
  MUX2X1 U13823 ( .B(n14622), .A(n14623), .S(n13104), .Y(n14621) );
  MUX2X1 U13824 ( .B(n14625), .A(n14626), .S(n13283), .Y(n14624) );
  MUX2X1 U13825 ( .B(n14628), .A(n14629), .S(n13283), .Y(n14627) );
  MUX2X1 U13826 ( .B(n14631), .A(n14632), .S(n13283), .Y(n14630) );
  MUX2X1 U13827 ( .B(n14634), .A(n14635), .S(n13283), .Y(n14633) );
  MUX2X1 U13828 ( .B(n14637), .A(n14638), .S(n13104), .Y(n14636) );
  MUX2X1 U13829 ( .B(n8780), .A(n10804), .S(n13316), .Y(n13381) );
  MUX2X1 U13830 ( .B(n8906), .A(n10930), .S(n13345), .Y(n13380) );
  MUX2X1 U13831 ( .B(n9032), .A(n11056), .S(n13345), .Y(n13384) );
  MUX2X1 U13832 ( .B(n9158), .A(n11182), .S(n13345), .Y(n13383) );
  MUX2X1 U13833 ( .B(n13382), .A(n13379), .S(n13265), .Y(n13393) );
  MUX2X1 U13834 ( .B(n9284), .A(n11308), .S(n13345), .Y(n13387) );
  MUX2X1 U13835 ( .B(n9410), .A(n11434), .S(n13345), .Y(n13386) );
  MUX2X1 U13836 ( .B(n9536), .A(n11560), .S(n13345), .Y(n13390) );
  MUX2X1 U13837 ( .B(n9662), .A(n11686), .S(n13345), .Y(n13389) );
  MUX2X1 U13838 ( .B(n13388), .A(n13385), .S(n13274), .Y(n13392) );
  MUX2X1 U13839 ( .B(n9788), .A(n11812), .S(n13345), .Y(n13396) );
  MUX2X1 U13840 ( .B(n9914), .A(n11938), .S(n13345), .Y(n13395) );
  MUX2X1 U13841 ( .B(n10040), .A(n12064), .S(n13345), .Y(n13399) );
  MUX2X1 U13842 ( .B(n10166), .A(n12190), .S(n13345), .Y(n13398) );
  MUX2X1 U13843 ( .B(n13397), .A(n13394), .S(n13275), .Y(n13408) );
  MUX2X1 U13844 ( .B(n10292), .A(n12316), .S(n13345), .Y(n13402) );
  MUX2X1 U13845 ( .B(n10418), .A(n12442), .S(n13345), .Y(n13401) );
  MUX2X1 U13846 ( .B(n10544), .A(n12568), .S(n13345), .Y(n13405) );
  MUX2X1 U13847 ( .B(n10670), .A(n12694), .S(n13344), .Y(n13404) );
  MUX2X1 U13848 ( .B(n13403), .A(n13400), .S(n13275), .Y(n13407) );
  MUX2X1 U13849 ( .B(n13406), .A(n13391), .S(n13101), .Y(n14639) );
  INVX2 U13850 ( .A(n14639), .Y(n112) );
  MUX2X1 U13851 ( .B(n8783), .A(n10807), .S(n13344), .Y(n13411) );
  MUX2X1 U13852 ( .B(n8909), .A(n10933), .S(n13344), .Y(n13410) );
  MUX2X1 U13853 ( .B(n9035), .A(n11059), .S(n13344), .Y(n13414) );
  MUX2X1 U13854 ( .B(n9161), .A(n11185), .S(n13344), .Y(n13413) );
  MUX2X1 U13855 ( .B(n13412), .A(n13409), .S(n13274), .Y(n13423) );
  MUX2X1 U13856 ( .B(n9287), .A(n11311), .S(n13344), .Y(n13417) );
  MUX2X1 U13857 ( .B(n9413), .A(n11437), .S(n13344), .Y(n13416) );
  MUX2X1 U13858 ( .B(n9539), .A(n11563), .S(n13344), .Y(n13420) );
  MUX2X1 U13859 ( .B(n9665), .A(n11689), .S(n13344), .Y(n13419) );
  MUX2X1 U13860 ( .B(n13418), .A(n13415), .S(n13274), .Y(n13422) );
  MUX2X1 U13861 ( .B(n9791), .A(n11815), .S(n13344), .Y(n13426) );
  MUX2X1 U13862 ( .B(n9917), .A(n11941), .S(n13344), .Y(n13425) );
  MUX2X1 U13863 ( .B(n10043), .A(n12067), .S(n13344), .Y(n13429) );
  MUX2X1 U13864 ( .B(n10169), .A(n12193), .S(n13344), .Y(n13428) );
  MUX2X1 U13865 ( .B(n13427), .A(n13424), .S(n13274), .Y(n13438) );
  MUX2X1 U13866 ( .B(n10295), .A(n12319), .S(n13344), .Y(n13432) );
  MUX2X1 U13867 ( .B(n10421), .A(n12445), .S(n13344), .Y(n13431) );
  MUX2X1 U13868 ( .B(n10547), .A(n12571), .S(n13344), .Y(n13435) );
  MUX2X1 U13869 ( .B(n10673), .A(n12697), .S(n13344), .Y(n13434) );
  MUX2X1 U13870 ( .B(n13433), .A(n13430), .S(n13274), .Y(n13437) );
  MUX2X1 U13871 ( .B(n13436), .A(n13421), .S(n13101), .Y(n14640) );
  INVX2 U13872 ( .A(n14640), .Y(n111) );
  MUX2X1 U13873 ( .B(n8786), .A(n10810), .S(n13343), .Y(n13441) );
  MUX2X1 U13874 ( .B(n8912), .A(n10936), .S(n13343), .Y(n13440) );
  MUX2X1 U13875 ( .B(n9038), .A(n11062), .S(n13343), .Y(n13444) );
  MUX2X1 U13876 ( .B(n9164), .A(n11188), .S(n13343), .Y(n13443) );
  MUX2X1 U13877 ( .B(n13442), .A(n13439), .S(n13274), .Y(n13453) );
  MUX2X1 U13878 ( .B(n9290), .A(n11314), .S(n13343), .Y(n13447) );
  MUX2X1 U13879 ( .B(n9416), .A(n11440), .S(n13343), .Y(n13446) );
  MUX2X1 U13880 ( .B(n9542), .A(n11566), .S(n13343), .Y(n13450) );
  MUX2X1 U13881 ( .B(n9668), .A(n11692), .S(n13343), .Y(n13449) );
  MUX2X1 U13882 ( .B(n13448), .A(n13445), .S(n13274), .Y(n13452) );
  MUX2X1 U13883 ( .B(n9794), .A(n11818), .S(n13343), .Y(n13456) );
  MUX2X1 U13884 ( .B(n9920), .A(n11944), .S(n13343), .Y(n13455) );
  MUX2X1 U13885 ( .B(n10046), .A(n12070), .S(n13343), .Y(n13459) );
  MUX2X1 U13886 ( .B(n10172), .A(n12196), .S(n13343), .Y(n13458) );
  MUX2X1 U13887 ( .B(n13457), .A(n13454), .S(n13274), .Y(n13468) );
  MUX2X1 U13888 ( .B(n10298), .A(n12322), .S(n13343), .Y(n13462) );
  MUX2X1 U13889 ( .B(n10424), .A(n12448), .S(n13343), .Y(n13461) );
  MUX2X1 U13890 ( .B(n10550), .A(n12574), .S(n13343), .Y(n13465) );
  MUX2X1 U13891 ( .B(n10676), .A(n12700), .S(n13343), .Y(n13464) );
  MUX2X1 U13892 ( .B(n13463), .A(n13460), .S(n13274), .Y(n13467) );
  MUX2X1 U13893 ( .B(n13466), .A(n13451), .S(n13101), .Y(n14641) );
  INVX2 U13894 ( .A(n14641), .Y(n110) );
  MUX2X1 U13895 ( .B(n8789), .A(n10813), .S(n13343), .Y(n13471) );
  MUX2X1 U13896 ( .B(n8915), .A(n10939), .S(n13342), .Y(n13470) );
  MUX2X1 U13897 ( .B(n9041), .A(n11065), .S(n13342), .Y(n13474) );
  MUX2X1 U13898 ( .B(n9167), .A(n11191), .S(n13342), .Y(n13473) );
  MUX2X1 U13899 ( .B(n13472), .A(n13469), .S(n13274), .Y(n13483) );
  MUX2X1 U13900 ( .B(n9293), .A(n11317), .S(n13342), .Y(n13477) );
  MUX2X1 U13901 ( .B(n9419), .A(n11443), .S(n13342), .Y(n13476) );
  MUX2X1 U13902 ( .B(n9545), .A(n11569), .S(n13342), .Y(n13480) );
  MUX2X1 U13903 ( .B(n9671), .A(n11695), .S(n13342), .Y(n13479) );
  MUX2X1 U13904 ( .B(n13478), .A(n13475), .S(n13274), .Y(n13482) );
  MUX2X1 U13905 ( .B(n9797), .A(n11821), .S(n13342), .Y(n13486) );
  MUX2X1 U13906 ( .B(n9923), .A(n11947), .S(n13342), .Y(n13485) );
  MUX2X1 U13907 ( .B(n10049), .A(n12073), .S(n13342), .Y(n13489) );
  MUX2X1 U13908 ( .B(n10175), .A(n12199), .S(n13342), .Y(n13488) );
  MUX2X1 U13909 ( .B(n13487), .A(n13484), .S(n13274), .Y(n13498) );
  MUX2X1 U13910 ( .B(n10301), .A(n12325), .S(n13342), .Y(n13492) );
  MUX2X1 U13911 ( .B(n10427), .A(n12451), .S(n13342), .Y(n13491) );
  MUX2X1 U13912 ( .B(n10553), .A(n12577), .S(n13342), .Y(n13495) );
  MUX2X1 U13913 ( .B(n10679), .A(n12703), .S(n13342), .Y(n13494) );
  MUX2X1 U13914 ( .B(n13493), .A(n13490), .S(n13273), .Y(n13497) );
  MUX2X1 U13915 ( .B(n13496), .A(n13481), .S(n13101), .Y(n14642) );
  INVX2 U13916 ( .A(n14642), .Y(n109) );
  MUX2X1 U13917 ( .B(n8792), .A(n10816), .S(n13342), .Y(n13501) );
  MUX2X1 U13918 ( .B(n8918), .A(n10942), .S(n13342), .Y(n13500) );
  MUX2X1 U13919 ( .B(n9044), .A(n11068), .S(n13341), .Y(n13504) );
  MUX2X1 U13920 ( .B(n9170), .A(n11194), .S(n13341), .Y(n13503) );
  MUX2X1 U13921 ( .B(n13502), .A(n13499), .S(n13274), .Y(n13513) );
  MUX2X1 U13922 ( .B(n9296), .A(n11320), .S(n13341), .Y(n13507) );
  MUX2X1 U13923 ( .B(n9422), .A(n11446), .S(n13341), .Y(n13506) );
  MUX2X1 U13924 ( .B(n9548), .A(n11572), .S(n13341), .Y(n13510) );
  MUX2X1 U13925 ( .B(n9674), .A(n11698), .S(n13341), .Y(n13509) );
  MUX2X1 U13926 ( .B(n13508), .A(n13505), .S(n13274), .Y(n13512) );
  MUX2X1 U13927 ( .B(n9800), .A(n11824), .S(n13341), .Y(n13516) );
  MUX2X1 U13928 ( .B(n9926), .A(n11950), .S(n13341), .Y(n13515) );
  MUX2X1 U13929 ( .B(n10052), .A(n12076), .S(n13341), .Y(n13519) );
  MUX2X1 U13930 ( .B(n10178), .A(n12202), .S(n13341), .Y(n13518) );
  MUX2X1 U13931 ( .B(n13517), .A(n13514), .S(n13274), .Y(n13528) );
  MUX2X1 U13932 ( .B(n10304), .A(n12328), .S(n13341), .Y(n13522) );
  MUX2X1 U13933 ( .B(n10430), .A(n12454), .S(n13341), .Y(n13521) );
  MUX2X1 U13934 ( .B(n10556), .A(n12580), .S(n13341), .Y(n13525) );
  MUX2X1 U13935 ( .B(n10682), .A(n12706), .S(n13341), .Y(n13524) );
  MUX2X1 U13936 ( .B(n13523), .A(n13520), .S(n13274), .Y(n13527) );
  MUX2X1 U13937 ( .B(n13526), .A(n13511), .S(n13101), .Y(n14643) );
  INVX2 U13938 ( .A(n14643), .Y(n108) );
  MUX2X1 U13939 ( .B(n8795), .A(n10819), .S(n13341), .Y(n13531) );
  MUX2X1 U13940 ( .B(n8921), .A(n10945), .S(n13341), .Y(n13530) );
  MUX2X1 U13941 ( .B(n9047), .A(n11071), .S(n13341), .Y(n13534) );
  MUX2X1 U13942 ( .B(n9173), .A(n11197), .S(n13340), .Y(n13533) );
  MUX2X1 U13943 ( .B(n13532), .A(n13529), .S(n13274), .Y(n13543) );
  MUX2X1 U13944 ( .B(n9299), .A(n11323), .S(n13340), .Y(n13537) );
  MUX2X1 U13945 ( .B(n9425), .A(n11449), .S(n13340), .Y(n13536) );
  MUX2X1 U13946 ( .B(n9551), .A(n11575), .S(n13340), .Y(n13540) );
  MUX2X1 U13947 ( .B(n9677), .A(n11701), .S(n13340), .Y(n13539) );
  MUX2X1 U13948 ( .B(n13538), .A(n13535), .S(n13273), .Y(n13542) );
  MUX2X1 U13949 ( .B(n9803), .A(n11827), .S(n13340), .Y(n13546) );
  MUX2X1 U13950 ( .B(n9929), .A(n11953), .S(n13340), .Y(n13545) );
  MUX2X1 U13951 ( .B(n10055), .A(n12079), .S(n13340), .Y(n13549) );
  MUX2X1 U13952 ( .B(n10181), .A(n12205), .S(n13340), .Y(n13548) );
  MUX2X1 U13953 ( .B(n13547), .A(n13544), .S(n13273), .Y(n13558) );
  MUX2X1 U13954 ( .B(n10307), .A(n12331), .S(n13340), .Y(n13552) );
  MUX2X1 U13955 ( .B(n10433), .A(n12457), .S(n13340), .Y(n13551) );
  MUX2X1 U13956 ( .B(n10559), .A(n12583), .S(n13340), .Y(n13555) );
  MUX2X1 U13957 ( .B(n10685), .A(n12709), .S(n13340), .Y(n13554) );
  MUX2X1 U13958 ( .B(n13553), .A(n13550), .S(n13273), .Y(n13557) );
  MUX2X1 U13959 ( .B(n13556), .A(n13541), .S(n13101), .Y(n14644) );
  INVX2 U13960 ( .A(n14644), .Y(n107) );
  MUX2X1 U13961 ( .B(n8798), .A(n10822), .S(n13340), .Y(n13561) );
  MUX2X1 U13962 ( .B(n8924), .A(n10948), .S(n13340), .Y(n13560) );
  MUX2X1 U13963 ( .B(n9050), .A(n11074), .S(n13340), .Y(n13564) );
  MUX2X1 U13964 ( .B(n9176), .A(n11200), .S(n13339), .Y(n13563) );
  MUX2X1 U13965 ( .B(n13562), .A(n13559), .S(n13273), .Y(n13573) );
  MUX2X1 U13966 ( .B(n9302), .A(n11326), .S(n13339), .Y(n13567) );
  MUX2X1 U13967 ( .B(n9428), .A(n11452), .S(n13339), .Y(n13566) );
  MUX2X1 U13968 ( .B(n9554), .A(n11578), .S(n13339), .Y(n13570) );
  MUX2X1 U13969 ( .B(n9680), .A(n11704), .S(n13339), .Y(n13569) );
  MUX2X1 U13970 ( .B(n13568), .A(n13565), .S(n13273), .Y(n13572) );
  MUX2X1 U13971 ( .B(n9806), .A(n11830), .S(n13339), .Y(n13576) );
  MUX2X1 U13972 ( .B(n9932), .A(n11956), .S(n13339), .Y(n13575) );
  MUX2X1 U13973 ( .B(n10058), .A(n12082), .S(n13339), .Y(n13579) );
  MUX2X1 U13974 ( .B(n10184), .A(n12208), .S(n13339), .Y(n13578) );
  MUX2X1 U13975 ( .B(n13577), .A(n13574), .S(n13273), .Y(n13588) );
  MUX2X1 U13976 ( .B(n10310), .A(n12334), .S(n13339), .Y(n13582) );
  MUX2X1 U13977 ( .B(n10436), .A(n12460), .S(n13339), .Y(n13581) );
  MUX2X1 U13978 ( .B(n10562), .A(n12586), .S(n13339), .Y(n13585) );
  MUX2X1 U13979 ( .B(n10688), .A(n12712), .S(n13339), .Y(n13584) );
  MUX2X1 U13980 ( .B(n13583), .A(n13580), .S(n13273), .Y(n13587) );
  MUX2X1 U13981 ( .B(n13586), .A(n13571), .S(n13101), .Y(n14645) );
  INVX2 U13982 ( .A(n14645), .Y(n106) );
  MUX2X1 U13983 ( .B(n8801), .A(n10825), .S(n13339), .Y(n13591) );
  MUX2X1 U13984 ( .B(n8927), .A(n10951), .S(n13339), .Y(n13590) );
  MUX2X1 U13985 ( .B(n9053), .A(n11077), .S(n13339), .Y(n13594) );
  MUX2X1 U13986 ( .B(n9179), .A(n11203), .S(n13339), .Y(n13593) );
  MUX2X1 U13987 ( .B(n13592), .A(n13589), .S(n13273), .Y(n13603) );
  MUX2X1 U13988 ( .B(n9305), .A(n11329), .S(n13338), .Y(n13597) );
  MUX2X1 U13989 ( .B(n9431), .A(n11455), .S(n13338), .Y(n13596) );
  MUX2X1 U13990 ( .B(n9557), .A(n11581), .S(n13338), .Y(n13600) );
  MUX2X1 U13991 ( .B(n9683), .A(n11707), .S(n13338), .Y(n13599) );
  MUX2X1 U13992 ( .B(n13598), .A(n13595), .S(n13273), .Y(n13602) );
  MUX2X1 U13993 ( .B(n9809), .A(n11833), .S(n13338), .Y(n13606) );
  MUX2X1 U13994 ( .B(n9935), .A(n11959), .S(n13338), .Y(n13605) );
  MUX2X1 U13995 ( .B(n10061), .A(n12085), .S(n13338), .Y(n13609) );
  MUX2X1 U13996 ( .B(n10187), .A(n12211), .S(n13338), .Y(n13608) );
  MUX2X1 U13997 ( .B(n13607), .A(n13604), .S(n13273), .Y(n13618) );
  MUX2X1 U13998 ( .B(n10313), .A(n12337), .S(n13338), .Y(n13612) );
  MUX2X1 U13999 ( .B(n10439), .A(n12463), .S(n13338), .Y(n13611) );
  MUX2X1 U14000 ( .B(n10565), .A(n12589), .S(n13338), .Y(n13615) );
  MUX2X1 U14001 ( .B(n10691), .A(n12715), .S(n13338), .Y(n13614) );
  MUX2X1 U14002 ( .B(n13613), .A(n13610), .S(n13273), .Y(n13617) );
  MUX2X1 U14003 ( .B(n13616), .A(n13601), .S(n13101), .Y(n14646) );
  INVX2 U14004 ( .A(n14646), .Y(n105) );
  MUX2X1 U14005 ( .B(n8804), .A(n10828), .S(n13338), .Y(n13621) );
  MUX2X1 U14006 ( .B(n8930), .A(n10954), .S(n13338), .Y(n13620) );
  MUX2X1 U14007 ( .B(n9056), .A(n11080), .S(n13338), .Y(n13624) );
  MUX2X1 U14008 ( .B(n9182), .A(n11206), .S(n13338), .Y(n13623) );
  MUX2X1 U14009 ( .B(n13622), .A(n13619), .S(n13273), .Y(n13633) );
  MUX2X1 U14010 ( .B(n9308), .A(n11332), .S(n13338), .Y(n13627) );
  MUX2X1 U14011 ( .B(n9434), .A(n11458), .S(n13337), .Y(n13626) );
  MUX2X1 U14012 ( .B(n9560), .A(n11584), .S(n13337), .Y(n13630) );
  MUX2X1 U14013 ( .B(n9686), .A(n11710), .S(n13337), .Y(n13629) );
  MUX2X1 U14014 ( .B(n13628), .A(n13625), .S(n13273), .Y(n13632) );
  MUX2X1 U14015 ( .B(n9812), .A(n11836), .S(n13337), .Y(n13636) );
  MUX2X1 U14016 ( .B(n9938), .A(n11962), .S(n13337), .Y(n13635) );
  MUX2X1 U14017 ( .B(n10064), .A(n12088), .S(n13337), .Y(n13639) );
  MUX2X1 U14018 ( .B(n10190), .A(n12214), .S(n13337), .Y(n13638) );
  MUX2X1 U14019 ( .B(n13637), .A(n13634), .S(n13273), .Y(n13648) );
  MUX2X1 U14020 ( .B(n10316), .A(n12340), .S(n13337), .Y(n13642) );
  MUX2X1 U14021 ( .B(n10442), .A(n12466), .S(n13337), .Y(n13641) );
  MUX2X1 U14022 ( .B(n10568), .A(n12592), .S(n13337), .Y(n13645) );
  MUX2X1 U14023 ( .B(n10694), .A(n12718), .S(n13337), .Y(n13644) );
  MUX2X1 U14024 ( .B(n13643), .A(n13640), .S(n13273), .Y(n13647) );
  MUX2X1 U14025 ( .B(n13646), .A(n13631), .S(n13101), .Y(n14647) );
  INVX2 U14026 ( .A(n14647), .Y(n104) );
  MUX2X1 U14027 ( .B(n8807), .A(n10831), .S(n13337), .Y(n13651) );
  MUX2X1 U14028 ( .B(n8933), .A(n10957), .S(n13337), .Y(n13650) );
  MUX2X1 U14029 ( .B(n9059), .A(n11083), .S(n13337), .Y(n13654) );
  MUX2X1 U14030 ( .B(n9185), .A(n11209), .S(n13337), .Y(n13653) );
  MUX2X1 U14031 ( .B(n13652), .A(n13649), .S(n13272), .Y(n13663) );
  MUX2X1 U14032 ( .B(n9311), .A(n11335), .S(n13337), .Y(n13657) );
  MUX2X1 U14033 ( .B(n9437), .A(n11461), .S(n13337), .Y(n13656) );
  MUX2X1 U14034 ( .B(n9563), .A(n11587), .S(n13336), .Y(n13660) );
  MUX2X1 U14035 ( .B(n9689), .A(n11713), .S(n13336), .Y(n13659) );
  MUX2X1 U14036 ( .B(n13658), .A(n13655), .S(n13273), .Y(n13662) );
  MUX2X1 U14037 ( .B(n9815), .A(n11839), .S(n13336), .Y(n13666) );
  MUX2X1 U14038 ( .B(n9941), .A(n11965), .S(n13336), .Y(n13665) );
  MUX2X1 U14039 ( .B(n10067), .A(n12091), .S(n13336), .Y(n13669) );
  MUX2X1 U14040 ( .B(n10193), .A(n12217), .S(n13336), .Y(n13668) );
  MUX2X1 U14041 ( .B(n13667), .A(n13664), .S(n13272), .Y(n13678) );
  MUX2X1 U14042 ( .B(n10319), .A(n12343), .S(n13336), .Y(n13672) );
  MUX2X1 U14043 ( .B(n10445), .A(n12469), .S(n13336), .Y(n13671) );
  MUX2X1 U14044 ( .B(n10571), .A(n12595), .S(n13336), .Y(n13675) );
  MUX2X1 U14045 ( .B(n10697), .A(n12721), .S(n13336), .Y(n13674) );
  MUX2X1 U14046 ( .B(n13673), .A(n13670), .S(n13272), .Y(n13677) );
  MUX2X1 U14047 ( .B(n13676), .A(n13661), .S(n13101), .Y(n14648) );
  INVX2 U14048 ( .A(n14648), .Y(n103) );
  MUX2X1 U14049 ( .B(n8810), .A(n10834), .S(n13336), .Y(n13681) );
  MUX2X1 U14050 ( .B(n8936), .A(n10960), .S(n13336), .Y(n13680) );
  MUX2X1 U14051 ( .B(n9062), .A(n11086), .S(n13336), .Y(n13684) );
  MUX2X1 U14052 ( .B(n9188), .A(n11212), .S(n13336), .Y(n13683) );
  MUX2X1 U14053 ( .B(n13682), .A(n13679), .S(n13272), .Y(n13693) );
  MUX2X1 U14054 ( .B(n9314), .A(n11338), .S(n13336), .Y(n13687) );
  MUX2X1 U14055 ( .B(n9440), .A(n11464), .S(n13336), .Y(n13686) );
  MUX2X1 U14056 ( .B(n9566), .A(n11590), .S(n13336), .Y(n13690) );
  MUX2X1 U14057 ( .B(n9692), .A(n11716), .S(n13335), .Y(n13689) );
  MUX2X1 U14058 ( .B(n13688), .A(n13685), .S(n13272), .Y(n13692) );
  MUX2X1 U14059 ( .B(n9818), .A(n11842), .S(n13340), .Y(n13696) );
  MUX2X1 U14060 ( .B(n9944), .A(n11968), .S(n13355), .Y(n13695) );
  MUX2X1 U14061 ( .B(n10070), .A(n12094), .S(n13355), .Y(n13699) );
  MUX2X1 U14062 ( .B(n10196), .A(n12220), .S(n13355), .Y(n13698) );
  MUX2X1 U14063 ( .B(n13697), .A(n13694), .S(n13272), .Y(n13708) );
  MUX2X1 U14064 ( .B(n10322), .A(n12346), .S(n13355), .Y(n13702) );
  MUX2X1 U14065 ( .B(n10448), .A(n12472), .S(n13355), .Y(n13701) );
  MUX2X1 U14066 ( .B(n10574), .A(n12598), .S(n13355), .Y(n13705) );
  MUX2X1 U14067 ( .B(n10700), .A(n12724), .S(n13355), .Y(n13704) );
  MUX2X1 U14068 ( .B(n13703), .A(n13700), .S(n13272), .Y(n13707) );
  MUX2X1 U14069 ( .B(n13706), .A(n13691), .S(n13101), .Y(n14649) );
  INVX2 U14070 ( .A(n14649), .Y(n102) );
  MUX2X1 U14071 ( .B(n8813), .A(n10837), .S(n13355), .Y(n13711) );
  MUX2X1 U14072 ( .B(n8939), .A(n10963), .S(n13355), .Y(n13710) );
  MUX2X1 U14073 ( .B(n9065), .A(n11089), .S(n13355), .Y(n13714) );
  MUX2X1 U14074 ( .B(n9191), .A(n11215), .S(n13355), .Y(n13713) );
  MUX2X1 U14075 ( .B(n13712), .A(n13709), .S(n13272), .Y(n13723) );
  MUX2X1 U14076 ( .B(n9317), .A(n11341), .S(n13355), .Y(n13717) );
  MUX2X1 U14077 ( .B(n9443), .A(n11467), .S(n13354), .Y(n13716) );
  MUX2X1 U14078 ( .B(n9569), .A(n11593), .S(n13354), .Y(n13720) );
  MUX2X1 U14079 ( .B(n9695), .A(n11719), .S(n13354), .Y(n13719) );
  MUX2X1 U14080 ( .B(n13718), .A(n13715), .S(n13272), .Y(n13722) );
  MUX2X1 U14081 ( .B(n9821), .A(n11845), .S(n13354), .Y(n13726) );
  MUX2X1 U14082 ( .B(n9947), .A(n11971), .S(n13354), .Y(n13725) );
  MUX2X1 U14083 ( .B(n10073), .A(n12097), .S(n13354), .Y(n13729) );
  MUX2X1 U14084 ( .B(n10199), .A(n12223), .S(n13354), .Y(n13728) );
  MUX2X1 U14085 ( .B(n13727), .A(n13724), .S(n13272), .Y(n13738) );
  MUX2X1 U14086 ( .B(n10325), .A(n12349), .S(n13354), .Y(n13732) );
  MUX2X1 U14087 ( .B(n10451), .A(n12475), .S(n13354), .Y(n13731) );
  MUX2X1 U14088 ( .B(n10577), .A(n12601), .S(n13354), .Y(n13735) );
  MUX2X1 U14089 ( .B(n10703), .A(n12727), .S(n13354), .Y(n13734) );
  MUX2X1 U14090 ( .B(n13733), .A(n13730), .S(n13272), .Y(n13737) );
  MUX2X1 U14091 ( .B(n13736), .A(n13721), .S(n13101), .Y(n14650) );
  INVX2 U14092 ( .A(n14650), .Y(n101) );
  MUX2X1 U14093 ( .B(n8816), .A(n10840), .S(n13354), .Y(n13741) );
  MUX2X1 U14094 ( .B(n8942), .A(n10966), .S(n13354), .Y(n13740) );
  MUX2X1 U14095 ( .B(n9068), .A(n11092), .S(n13354), .Y(n13744) );
  MUX2X1 U14096 ( .B(n9194), .A(n11218), .S(n13354), .Y(n13743) );
  MUX2X1 U14097 ( .B(n13742), .A(n13739), .S(n13272), .Y(n13753) );
  MUX2X1 U14098 ( .B(n9320), .A(n11344), .S(n13354), .Y(n13747) );
  MUX2X1 U14099 ( .B(n9446), .A(n11470), .S(n13354), .Y(n13746) );
  MUX2X1 U14100 ( .B(n9572), .A(n11596), .S(n13353), .Y(n13750) );
  MUX2X1 U14101 ( .B(n9698), .A(n11722), .S(n13353), .Y(n13749) );
  MUX2X1 U14102 ( .B(n13748), .A(n13745), .S(n13272), .Y(n13752) );
  MUX2X1 U14103 ( .B(n9824), .A(n11848), .S(n13353), .Y(n13756) );
  MUX2X1 U14104 ( .B(n9950), .A(n11974), .S(n13353), .Y(n13755) );
  MUX2X1 U14105 ( .B(n10076), .A(n12100), .S(n13353), .Y(n13759) );
  MUX2X1 U14106 ( .B(n10202), .A(n12226), .S(n13353), .Y(n13758) );
  MUX2X1 U14107 ( .B(n13757), .A(n13754), .S(n13272), .Y(n13768) );
  MUX2X1 U14108 ( .B(n10328), .A(n12352), .S(n13353), .Y(n13762) );
  MUX2X1 U14109 ( .B(n10454), .A(n12478), .S(n13353), .Y(n13761) );
  MUX2X1 U14110 ( .B(n10580), .A(n12604), .S(n13353), .Y(n13765) );
  MUX2X1 U14111 ( .B(n10706), .A(n12730), .S(n13353), .Y(n13764) );
  MUX2X1 U14112 ( .B(n13763), .A(n13760), .S(n13272), .Y(n13767) );
  MUX2X1 U14113 ( .B(n13766), .A(n13751), .S(n13101), .Y(n14651) );
  INVX2 U14114 ( .A(n14651), .Y(n100) );
  MUX2X1 U14115 ( .B(n8819), .A(n10843), .S(n13353), .Y(n13771) );
  MUX2X1 U14116 ( .B(n8945), .A(n10969), .S(n13353), .Y(n13770) );
  MUX2X1 U14117 ( .B(n9071), .A(n11095), .S(n13353), .Y(n13774) );
  MUX2X1 U14118 ( .B(n9197), .A(n11221), .S(n13353), .Y(n13773) );
  MUX2X1 U14119 ( .B(n13772), .A(n13769), .S(n13272), .Y(n13783) );
  MUX2X1 U14120 ( .B(n9323), .A(n11347), .S(n13353), .Y(n13777) );
  MUX2X1 U14121 ( .B(n9449), .A(n11473), .S(n13353), .Y(n13776) );
  MUX2X1 U14122 ( .B(n9575), .A(n11599), .S(n13353), .Y(n13780) );
  MUX2X1 U14123 ( .B(n9701), .A(n11725), .S(n13352), .Y(n13779) );
  MUX2X1 U14124 ( .B(n13778), .A(n13775), .S(n13272), .Y(n13782) );
  MUX2X1 U14125 ( .B(n9827), .A(n11851), .S(n13352), .Y(n13786) );
  MUX2X1 U14126 ( .B(n9953), .A(n11977), .S(n13352), .Y(n13785) );
  MUX2X1 U14127 ( .B(n10079), .A(n12103), .S(n13352), .Y(n13789) );
  MUX2X1 U14128 ( .B(n10205), .A(n12229), .S(n13352), .Y(n13788) );
  MUX2X1 U14129 ( .B(n13787), .A(n13784), .S(n13271), .Y(n13798) );
  MUX2X1 U14130 ( .B(n10331), .A(n12355), .S(n13352), .Y(n13792) );
  MUX2X1 U14131 ( .B(n10457), .A(n12481), .S(n13352), .Y(n13791) );
  MUX2X1 U14132 ( .B(n10583), .A(n12607), .S(n13352), .Y(n13795) );
  MUX2X1 U14133 ( .B(n10709), .A(n12733), .S(n13352), .Y(n13794) );
  MUX2X1 U14134 ( .B(n13793), .A(n13790), .S(n13271), .Y(n13797) );
  MUX2X1 U14135 ( .B(n13796), .A(n13781), .S(n13101), .Y(n14652) );
  INVX2 U14136 ( .A(n14652), .Y(n99) );
  MUX2X1 U14137 ( .B(n8822), .A(n10846), .S(n13352), .Y(n13801) );
  MUX2X1 U14138 ( .B(n8948), .A(n10972), .S(n13352), .Y(n13800) );
  MUX2X1 U14139 ( .B(n9074), .A(n11098), .S(n13352), .Y(n13804) );
  MUX2X1 U14140 ( .B(n9200), .A(n11224), .S(n13352), .Y(n13803) );
  MUX2X1 U14141 ( .B(n13802), .A(n13799), .S(n13271), .Y(n13813) );
  MUX2X1 U14142 ( .B(n9326), .A(n11350), .S(n13352), .Y(n13807) );
  MUX2X1 U14143 ( .B(n9452), .A(n11476), .S(n13352), .Y(n13806) );
  MUX2X1 U14144 ( .B(n9578), .A(n11602), .S(n13352), .Y(n13810) );
  MUX2X1 U14145 ( .B(n9704), .A(n11728), .S(n13352), .Y(n13809) );
  MUX2X1 U14146 ( .B(n13808), .A(n13805), .S(n13271), .Y(n13812) );
  MUX2X1 U14147 ( .B(n9830), .A(n11854), .S(n13351), .Y(n13816) );
  MUX2X1 U14148 ( .B(n9956), .A(n11980), .S(n13351), .Y(n13815) );
  MUX2X1 U14149 ( .B(n10082), .A(n12106), .S(n13351), .Y(n13819) );
  MUX2X1 U14150 ( .B(n10208), .A(n12232), .S(n13351), .Y(n13818) );
  MUX2X1 U14151 ( .B(n13817), .A(n13814), .S(n13271), .Y(n13828) );
  MUX2X1 U14152 ( .B(n10334), .A(n12358), .S(n13351), .Y(n13822) );
  MUX2X1 U14153 ( .B(n10460), .A(n12484), .S(n13351), .Y(n13821) );
  MUX2X1 U14154 ( .B(n10586), .A(n12610), .S(n13351), .Y(n13825) );
  MUX2X1 U14155 ( .B(n10712), .A(n12736), .S(n13351), .Y(n13824) );
  MUX2X1 U14156 ( .B(n13823), .A(n13820), .S(n13271), .Y(n13827) );
  MUX2X1 U14157 ( .B(n13826), .A(n13811), .S(n13101), .Y(n14653) );
  INVX2 U14158 ( .A(n14653), .Y(n98) );
  MUX2X1 U14159 ( .B(n8825), .A(n10849), .S(n13351), .Y(n13831) );
  MUX2X1 U14160 ( .B(n8951), .A(n10975), .S(n13351), .Y(n13830) );
  MUX2X1 U14161 ( .B(n9077), .A(n11101), .S(n13351), .Y(n13834) );
  MUX2X1 U14162 ( .B(n9203), .A(n11227), .S(n13351), .Y(n13833) );
  MUX2X1 U14163 ( .B(n13832), .A(n13829), .S(n13271), .Y(n13843) );
  MUX2X1 U14164 ( .B(n9329), .A(n11353), .S(n13351), .Y(n13837) );
  MUX2X1 U14165 ( .B(n9455), .A(n11479), .S(n13351), .Y(n13836) );
  MUX2X1 U14166 ( .B(n9581), .A(n11605), .S(n13351), .Y(n13840) );
  MUX2X1 U14167 ( .B(n9707), .A(n11731), .S(n13351), .Y(n13839) );
  MUX2X1 U14168 ( .B(n13838), .A(n13835), .S(n13271), .Y(n13842) );
  MUX2X1 U14169 ( .B(n9833), .A(n11857), .S(n13351), .Y(n13846) );
  MUX2X1 U14170 ( .B(n9959), .A(n11983), .S(n13350), .Y(n13845) );
  MUX2X1 U14171 ( .B(n10085), .A(n12109), .S(n13350), .Y(n13849) );
  MUX2X1 U14172 ( .B(n10211), .A(n12235), .S(n13350), .Y(n13848) );
  MUX2X1 U14173 ( .B(n13847), .A(n13844), .S(n13271), .Y(n13858) );
  MUX2X1 U14174 ( .B(n10337), .A(n12361), .S(n13350), .Y(n13852) );
  MUX2X1 U14175 ( .B(n10463), .A(n12487), .S(n13350), .Y(n13851) );
  MUX2X1 U14176 ( .B(n10589), .A(n12613), .S(n13350), .Y(n13855) );
  MUX2X1 U14177 ( .B(n10715), .A(n12739), .S(n13350), .Y(n13854) );
  MUX2X1 U14178 ( .B(n13853), .A(n13850), .S(n13271), .Y(n13857) );
  MUX2X1 U14179 ( .B(n13856), .A(n13841), .S(n13101), .Y(n14654) );
  INVX2 U14180 ( .A(n14654), .Y(n97) );
  MUX2X1 U14181 ( .B(n8828), .A(n10852), .S(n13350), .Y(n13861) );
  MUX2X1 U14182 ( .B(n8954), .A(n10978), .S(n13350), .Y(n13860) );
  MUX2X1 U14183 ( .B(n9080), .A(n11104), .S(n13350), .Y(n13864) );
  MUX2X1 U14184 ( .B(n9206), .A(n11230), .S(n13350), .Y(n13863) );
  MUX2X1 U14185 ( .B(n13862), .A(n13859), .S(n13271), .Y(n13873) );
  MUX2X1 U14186 ( .B(n9332), .A(n11356), .S(n13350), .Y(n13867) );
  MUX2X1 U14187 ( .B(n9458), .A(n11482), .S(n13350), .Y(n13866) );
  MUX2X1 U14188 ( .B(n9584), .A(n11608), .S(n13350), .Y(n13870) );
  MUX2X1 U14189 ( .B(n9710), .A(n11734), .S(n13350), .Y(n13869) );
  MUX2X1 U14190 ( .B(n13868), .A(n13865), .S(n13271), .Y(n13872) );
  MUX2X1 U14191 ( .B(n9836), .A(n11860), .S(n13350), .Y(n13876) );
  MUX2X1 U14192 ( .B(n9962), .A(n11986), .S(n13349), .Y(n13875) );
  MUX2X1 U14193 ( .B(n10088), .A(n12112), .S(n13349), .Y(n13879) );
  MUX2X1 U14194 ( .B(n10214), .A(n12238), .S(n13349), .Y(n13878) );
  MUX2X1 U14195 ( .B(n13877), .A(n13874), .S(n13271), .Y(n13888) );
  MUX2X1 U14196 ( .B(n10340), .A(n12364), .S(n13349), .Y(n13882) );
  MUX2X1 U14197 ( .B(n10466), .A(n12490), .S(n13349), .Y(n13881) );
  MUX2X1 U14198 ( .B(n10592), .A(n12616), .S(n13349), .Y(n13885) );
  MUX2X1 U14199 ( .B(n10718), .A(n12742), .S(n13349), .Y(n13884) );
  MUX2X1 U14200 ( .B(n13883), .A(n13880), .S(n13271), .Y(n13887) );
  MUX2X1 U14201 ( .B(n13886), .A(n13871), .S(n13101), .Y(n14655) );
  INVX2 U14202 ( .A(n14655), .Y(n96) );
  MUX2X1 U14203 ( .B(n8831), .A(n10855), .S(n13349), .Y(n13891) );
  MUX2X1 U14204 ( .B(n8957), .A(n10981), .S(n13349), .Y(n13890) );
  MUX2X1 U14205 ( .B(n9083), .A(n11107), .S(n13349), .Y(n13894) );
  MUX2X1 U14206 ( .B(n9209), .A(n11233), .S(n13349), .Y(n13893) );
  MUX2X1 U14207 ( .B(n13892), .A(n13889), .S(n13271), .Y(n13903) );
  MUX2X1 U14208 ( .B(n9335), .A(n11359), .S(n13349), .Y(n13897) );
  MUX2X1 U14209 ( .B(n9461), .A(n11485), .S(n13349), .Y(n13896) );
  MUX2X1 U14210 ( .B(n9587), .A(n11611), .S(n13349), .Y(n13900) );
  MUX2X1 U14211 ( .B(n9713), .A(n11737), .S(n13349), .Y(n13899) );
  MUX2X1 U14212 ( .B(n13898), .A(n13895), .S(n13271), .Y(n13902) );
  MUX2X1 U14213 ( .B(n9839), .A(n11863), .S(n13349), .Y(n13906) );
  MUX2X1 U14214 ( .B(n9965), .A(n11989), .S(n13349), .Y(n13905) );
  MUX2X1 U14215 ( .B(n10091), .A(n12115), .S(n13348), .Y(n13909) );
  MUX2X1 U14216 ( .B(n10217), .A(n12241), .S(n13348), .Y(n13908) );
  MUX2X1 U14217 ( .B(n13907), .A(n13904), .S(n13271), .Y(n13918) );
  MUX2X1 U14218 ( .B(n10343), .A(n12367), .S(n13348), .Y(n13912) );
  MUX2X1 U14219 ( .B(n10469), .A(n12493), .S(n13348), .Y(n13911) );
  MUX2X1 U14220 ( .B(n10595), .A(n12619), .S(n13348), .Y(n13915) );
  MUX2X1 U14221 ( .B(n10721), .A(n12745), .S(n13348), .Y(n13914) );
  MUX2X1 U14222 ( .B(n13913), .A(n13910), .S(n13270), .Y(n13917) );
  MUX2X1 U14223 ( .B(n13916), .A(n13901), .S(n13101), .Y(n14656) );
  INVX2 U14224 ( .A(n14656), .Y(n95) );
  MUX2X1 U14225 ( .B(n8834), .A(n10858), .S(n13348), .Y(n13921) );
  MUX2X1 U14226 ( .B(n8960), .A(n10984), .S(n13348), .Y(n13920) );
  MUX2X1 U14227 ( .B(n9086), .A(n11110), .S(n13348), .Y(n13924) );
  MUX2X1 U14228 ( .B(n9212), .A(n11236), .S(n13348), .Y(n13923) );
  MUX2X1 U14229 ( .B(n13922), .A(n13919), .S(n13270), .Y(n13933) );
  MUX2X1 U14230 ( .B(n9338), .A(n11362), .S(n13348), .Y(n13927) );
  MUX2X1 U14231 ( .B(n9464), .A(n11488), .S(n13348), .Y(n13926) );
  MUX2X1 U14232 ( .B(n9590), .A(n11614), .S(n13348), .Y(n13930) );
  MUX2X1 U14233 ( .B(n9716), .A(n11740), .S(n13348), .Y(n13929) );
  MUX2X1 U14234 ( .B(n13928), .A(n13925), .S(n13270), .Y(n13932) );
  MUX2X1 U14235 ( .B(n9842), .A(n11866), .S(n13348), .Y(n13936) );
  MUX2X1 U14236 ( .B(n9968), .A(n11992), .S(n13348), .Y(n13935) );
  MUX2X1 U14237 ( .B(n10094), .A(n12118), .S(n13348), .Y(n13939) );
  MUX2X1 U14238 ( .B(n10220), .A(n12244), .S(n13347), .Y(n13938) );
  MUX2X1 U14239 ( .B(n13937), .A(n13934), .S(n13270), .Y(n13948) );
  MUX2X1 U14240 ( .B(n10346), .A(n12370), .S(n13347), .Y(n13942) );
  MUX2X1 U14241 ( .B(n10472), .A(n12496), .S(n13347), .Y(n13941) );
  MUX2X1 U14242 ( .B(n10598), .A(n12622), .S(n13347), .Y(n13945) );
  MUX2X1 U14243 ( .B(n10724), .A(n12748), .S(n13347), .Y(n13944) );
  MUX2X1 U14244 ( .B(n13943), .A(n13940), .S(n13270), .Y(n13947) );
  MUX2X1 U14245 ( .B(n13946), .A(n13931), .S(n13101), .Y(n14657) );
  INVX2 U14246 ( .A(n14657), .Y(n94) );
  MUX2X1 U14247 ( .B(n8837), .A(n10861), .S(n13347), .Y(n13951) );
  MUX2X1 U14248 ( .B(n8963), .A(n10987), .S(n13347), .Y(n13950) );
  MUX2X1 U14249 ( .B(n9089), .A(n11113), .S(n13347), .Y(n13954) );
  MUX2X1 U14250 ( .B(n9215), .A(n11239), .S(n13347), .Y(n13953) );
  MUX2X1 U14251 ( .B(n13952), .A(n13949), .S(n13270), .Y(n13963) );
  MUX2X1 U14252 ( .B(n9341), .A(n11365), .S(n13347), .Y(n13957) );
  MUX2X1 U14253 ( .B(n9467), .A(n11491), .S(n13347), .Y(n13956) );
  MUX2X1 U14254 ( .B(n9593), .A(n11617), .S(n13347), .Y(n13960) );
  MUX2X1 U14255 ( .B(n9719), .A(n11743), .S(n13347), .Y(n13959) );
  MUX2X1 U14256 ( .B(n13958), .A(n13955), .S(n13270), .Y(n13962) );
  MUX2X1 U14257 ( .B(n9845), .A(n11869), .S(n13347), .Y(n13966) );
  MUX2X1 U14258 ( .B(n9971), .A(n11995), .S(n13347), .Y(n13965) );
  MUX2X1 U14259 ( .B(n10097), .A(n12121), .S(n13347), .Y(n13969) );
  MUX2X1 U14260 ( .B(n10223), .A(n12247), .S(n13347), .Y(n13968) );
  MUX2X1 U14261 ( .B(n13967), .A(n13964), .S(n13270), .Y(n13978) );
  MUX2X1 U14262 ( .B(n10349), .A(n12373), .S(n13346), .Y(n13972) );
  MUX2X1 U14263 ( .B(n10475), .A(n12499), .S(n13346), .Y(n13971) );
  MUX2X1 U14264 ( .B(n10601), .A(n12625), .S(n13346), .Y(n13975) );
  MUX2X1 U14265 ( .B(n10727), .A(n12751), .S(n13346), .Y(n13974) );
  MUX2X1 U14266 ( .B(n13973), .A(n13970), .S(n13270), .Y(n13977) );
  MUX2X1 U14267 ( .B(n13976), .A(n13961), .S(n13101), .Y(n14658) );
  INVX2 U14268 ( .A(n14658), .Y(n93) );
  MUX2X1 U14269 ( .B(n8840), .A(n10864), .S(n13346), .Y(n13981) );
  MUX2X1 U14270 ( .B(n8966), .A(n10990), .S(n13346), .Y(n13980) );
  MUX2X1 U14271 ( .B(n9092), .A(n11116), .S(n13346), .Y(n13984) );
  MUX2X1 U14272 ( .B(n9218), .A(n11242), .S(n13346), .Y(n13983) );
  MUX2X1 U14273 ( .B(n13982), .A(n13979), .S(n13270), .Y(n13993) );
  MUX2X1 U14274 ( .B(n9344), .A(n11368), .S(n13346), .Y(n13987) );
  MUX2X1 U14275 ( .B(n9470), .A(n11494), .S(n13346), .Y(n13986) );
  MUX2X1 U14276 ( .B(n9596), .A(n11620), .S(n13346), .Y(n13990) );
  MUX2X1 U14277 ( .B(n9722), .A(n11746), .S(n13346), .Y(n13989) );
  MUX2X1 U14278 ( .B(n13988), .A(n13985), .S(n13270), .Y(n13992) );
  MUX2X1 U14279 ( .B(n9848), .A(n11872), .S(n13346), .Y(n13996) );
  MUX2X1 U14280 ( .B(n9974), .A(n11998), .S(n13346), .Y(n13995) );
  MUX2X1 U14281 ( .B(n10100), .A(n12124), .S(n13346), .Y(n13999) );
  MUX2X1 U14282 ( .B(n10226), .A(n12250), .S(n13346), .Y(n13998) );
  MUX2X1 U14283 ( .B(n13997), .A(n13994), .S(n13270), .Y(n14008) );
  MUX2X1 U14284 ( .B(n10352), .A(n12376), .S(n13346), .Y(n14002) );
  MUX2X1 U14285 ( .B(n10478), .A(n12502), .S(n13345), .Y(n14001) );
  MUX2X1 U14286 ( .B(n10604), .A(n12628), .S(n13345), .Y(n14005) );
  MUX2X1 U14287 ( .B(n10730), .A(n12754), .S(n13345), .Y(n14004) );
  MUX2X1 U14288 ( .B(n14003), .A(n14000), .S(n13270), .Y(n14007) );
  MUX2X1 U14289 ( .B(n14006), .A(n13991), .S(n13101), .Y(n14659) );
  INVX2 U14290 ( .A(n14659), .Y(n92) );
  MUX2X1 U14291 ( .B(n8843), .A(n10867), .S(n13350), .Y(n14011) );
  MUX2X1 U14292 ( .B(n8969), .A(n10993), .S(n13326), .Y(n14010) );
  MUX2X1 U14293 ( .B(n9095), .A(n11119), .S(n13325), .Y(n14014) );
  MUX2X1 U14294 ( .B(n9221), .A(n11245), .S(n13325), .Y(n14013) );
  MUX2X1 U14295 ( .B(n14012), .A(n14009), .S(n13270), .Y(n14023) );
  MUX2X1 U14296 ( .B(n9347), .A(n11371), .S(n13325), .Y(n14017) );
  MUX2X1 U14297 ( .B(n9473), .A(n11497), .S(n13325), .Y(n14016) );
  MUX2X1 U14298 ( .B(n9599), .A(n11623), .S(n13325), .Y(n14020) );
  MUX2X1 U14299 ( .B(n9725), .A(n11749), .S(n13325), .Y(n14019) );
  MUX2X1 U14300 ( .B(n14018), .A(n14015), .S(n13270), .Y(n14022) );
  MUX2X1 U14301 ( .B(n9851), .A(n11875), .S(n13325), .Y(n14026) );
  MUX2X1 U14302 ( .B(n9977), .A(n12001), .S(n13325), .Y(n14025) );
  MUX2X1 U14303 ( .B(n10103), .A(n12127), .S(n13325), .Y(n14029) );
  MUX2X1 U14304 ( .B(n10229), .A(n12253), .S(n13325), .Y(n14028) );
  MUX2X1 U14305 ( .B(n14027), .A(n14024), .S(n13270), .Y(n14038) );
  MUX2X1 U14306 ( .B(n10355), .A(n12379), .S(n13325), .Y(n14032) );
  MUX2X1 U14307 ( .B(n10481), .A(n12505), .S(n13325), .Y(n14031) );
  MUX2X1 U14308 ( .B(n10607), .A(n12631), .S(n13325), .Y(n14035) );
  MUX2X1 U14309 ( .B(n10733), .A(n12757), .S(n13325), .Y(n14034) );
  MUX2X1 U14310 ( .B(n14033), .A(n14030), .S(n13269), .Y(n14037) );
  MUX2X1 U14311 ( .B(n14036), .A(n14021), .S(n13101), .Y(n14660) );
  INVX2 U14312 ( .A(n14660), .Y(n91) );
  MUX2X1 U14313 ( .B(n8846), .A(n10870), .S(n13325), .Y(n14041) );
  MUX2X1 U14314 ( .B(n8972), .A(n10996), .S(n13325), .Y(n14040) );
  MUX2X1 U14315 ( .B(n9098), .A(n11122), .S(n13325), .Y(n14044) );
  MUX2X1 U14316 ( .B(n9224), .A(n11248), .S(n13324), .Y(n14043) );
  MUX2X1 U14317 ( .B(n14042), .A(n14039), .S(n13269), .Y(n14053) );
  MUX2X1 U14318 ( .B(n9350), .A(n11374), .S(n13324), .Y(n14047) );
  MUX2X1 U14319 ( .B(n9476), .A(n11500), .S(n13324), .Y(n14046) );
  MUX2X1 U14320 ( .B(n9602), .A(n11626), .S(n13324), .Y(n14050) );
  MUX2X1 U14321 ( .B(n9728), .A(n11752), .S(n13324), .Y(n14049) );
  MUX2X1 U14322 ( .B(n14048), .A(n14045), .S(n13269), .Y(n14052) );
  MUX2X1 U14323 ( .B(n9854), .A(n11878), .S(n13324), .Y(n14056) );
  MUX2X1 U14324 ( .B(n9980), .A(n12004), .S(n13324), .Y(n14055) );
  MUX2X1 U14325 ( .B(n10106), .A(n12130), .S(n13324), .Y(n14059) );
  MUX2X1 U14326 ( .B(n10232), .A(n12256), .S(n13324), .Y(n14058) );
  MUX2X1 U14327 ( .B(n14057), .A(n14054), .S(n13269), .Y(n14068) );
  MUX2X1 U14328 ( .B(n10358), .A(n12382), .S(n13324), .Y(n14062) );
  MUX2X1 U14329 ( .B(n10484), .A(n12508), .S(n13324), .Y(n14061) );
  MUX2X1 U14330 ( .B(n10610), .A(n12634), .S(n13324), .Y(n14065) );
  MUX2X1 U14331 ( .B(n10736), .A(n12760), .S(n13324), .Y(n14064) );
  MUX2X1 U14332 ( .B(n14063), .A(n14060), .S(n13269), .Y(n14067) );
  MUX2X1 U14333 ( .B(n14066), .A(n14051), .S(n13101), .Y(n14661) );
  INVX2 U14334 ( .A(n14661), .Y(n90) );
  MUX2X1 U14335 ( .B(n8849), .A(n10873), .S(n13324), .Y(n14071) );
  MUX2X1 U14336 ( .B(n8975), .A(n10999), .S(n13324), .Y(n14070) );
  MUX2X1 U14337 ( .B(n9101), .A(n11125), .S(n13324), .Y(n14074) );
  MUX2X1 U14338 ( .B(n9227), .A(n11251), .S(n13324), .Y(n14073) );
  MUX2X1 U14339 ( .B(n14072), .A(n14069), .S(n13269), .Y(n14083) );
  MUX2X1 U14340 ( .B(n9353), .A(n11377), .S(n13323), .Y(n14077) );
  MUX2X1 U14341 ( .B(n9479), .A(n11503), .S(n13323), .Y(n14076) );
  MUX2X1 U14342 ( .B(n9605), .A(n11629), .S(n13323), .Y(n14080) );
  MUX2X1 U14343 ( .B(n9731), .A(n11755), .S(n13323), .Y(n14079) );
  MUX2X1 U14344 ( .B(n14078), .A(n14075), .S(n13269), .Y(n14082) );
  MUX2X1 U14345 ( .B(n9857), .A(n11881), .S(n13323), .Y(n14086) );
  MUX2X1 U14346 ( .B(n9983), .A(n12007), .S(n13323), .Y(n14085) );
  MUX2X1 U14347 ( .B(n10109), .A(n12133), .S(n13323), .Y(n14089) );
  MUX2X1 U14348 ( .B(n10235), .A(n12259), .S(n13323), .Y(n14088) );
  MUX2X1 U14349 ( .B(n14087), .A(n14084), .S(n13269), .Y(n14098) );
  MUX2X1 U14350 ( .B(n10361), .A(n12385), .S(n13323), .Y(n14092) );
  MUX2X1 U14351 ( .B(n10487), .A(n12511), .S(n13323), .Y(n14091) );
  MUX2X1 U14352 ( .B(n10613), .A(n12637), .S(n13323), .Y(n14095) );
  MUX2X1 U14353 ( .B(n10739), .A(n12763), .S(n13323), .Y(n14094) );
  MUX2X1 U14354 ( .B(n14093), .A(n14090), .S(n13269), .Y(n14097) );
  MUX2X1 U14355 ( .B(n14096), .A(n14081), .S(n13101), .Y(n14662) );
  INVX2 U14356 ( .A(n14662), .Y(n89) );
  MUX2X1 U14357 ( .B(n8852), .A(n10876), .S(n13323), .Y(n14101) );
  MUX2X1 U14358 ( .B(n8978), .A(n11002), .S(n13323), .Y(n14100) );
  MUX2X1 U14359 ( .B(n9104), .A(n11128), .S(n13323), .Y(n14104) );
  MUX2X1 U14360 ( .B(n9230), .A(n11254), .S(n13323), .Y(n14103) );
  MUX2X1 U14361 ( .B(n14102), .A(n14099), .S(n13269), .Y(n14113) );
  MUX2X1 U14362 ( .B(n9356), .A(n11380), .S(n13323), .Y(n14107) );
  MUX2X1 U14363 ( .B(n9482), .A(n11506), .S(n13322), .Y(n14106) );
  MUX2X1 U14364 ( .B(n9608), .A(n11632), .S(n13322), .Y(n14110) );
  MUX2X1 U14365 ( .B(n9734), .A(n11758), .S(n13322), .Y(n14109) );
  MUX2X1 U14366 ( .B(n14108), .A(n14105), .S(n13269), .Y(n14112) );
  MUX2X1 U14367 ( .B(n9860), .A(n11884), .S(n13322), .Y(n14116) );
  MUX2X1 U14368 ( .B(n9986), .A(n12010), .S(n13322), .Y(n14115) );
  MUX2X1 U14369 ( .B(n10112), .A(n12136), .S(n13322), .Y(n14119) );
  MUX2X1 U14370 ( .B(n10238), .A(n12262), .S(n13322), .Y(n14118) );
  MUX2X1 U14371 ( .B(n14117), .A(n14114), .S(n13269), .Y(n14128) );
  MUX2X1 U14372 ( .B(n10364), .A(n12388), .S(n13322), .Y(n14122) );
  MUX2X1 U14373 ( .B(n10490), .A(n12514), .S(n13322), .Y(n14121) );
  MUX2X1 U14374 ( .B(n10616), .A(n12640), .S(n13322), .Y(n14125) );
  MUX2X1 U14375 ( .B(n10742), .A(n12766), .S(n13322), .Y(n14124) );
  MUX2X1 U14376 ( .B(n14123), .A(n14120), .S(n13269), .Y(n14127) );
  MUX2X1 U14377 ( .B(n14126), .A(n14111), .S(n13101), .Y(n14663) );
  INVX2 U14378 ( .A(n14663), .Y(n88) );
  MUX2X1 U14379 ( .B(n8855), .A(n10879), .S(n13322), .Y(n14131) );
  MUX2X1 U14380 ( .B(n8981), .A(n11005), .S(n13322), .Y(n14130) );
  MUX2X1 U14381 ( .B(n9107), .A(n11131), .S(n13322), .Y(n14134) );
  MUX2X1 U14382 ( .B(n9233), .A(n11257), .S(n13322), .Y(n14133) );
  MUX2X1 U14383 ( .B(n14132), .A(n14129), .S(n13269), .Y(n14143) );
  MUX2X1 U14384 ( .B(n9359), .A(n11383), .S(n13322), .Y(n14137) );
  MUX2X1 U14385 ( .B(n9485), .A(n11509), .S(n13322), .Y(n14136) );
  MUX2X1 U14386 ( .B(n9611), .A(n11635), .S(n13321), .Y(n14140) );
  MUX2X1 U14387 ( .B(n9737), .A(n11761), .S(n13321), .Y(n14139) );
  MUX2X1 U14388 ( .B(n14138), .A(n14135), .S(n13269), .Y(n14142) );
  MUX2X1 U14389 ( .B(n9863), .A(n11887), .S(n13321), .Y(n14146) );
  MUX2X1 U14390 ( .B(n9989), .A(n12013), .S(n13321), .Y(n14145) );
  MUX2X1 U14391 ( .B(n10115), .A(n12139), .S(n13321), .Y(n14149) );
  MUX2X1 U14392 ( .B(n10241), .A(n12265), .S(n13321), .Y(n14148) );
  MUX2X1 U14393 ( .B(n14147), .A(n14144), .S(n13269), .Y(n14158) );
  MUX2X1 U14394 ( .B(n10367), .A(n12391), .S(n13321), .Y(n14152) );
  MUX2X1 U14395 ( .B(n10493), .A(n12517), .S(n13321), .Y(n14151) );
  MUX2X1 U14396 ( .B(n10619), .A(n12643), .S(n13321), .Y(n14155) );
  MUX2X1 U14397 ( .B(n10745), .A(n12769), .S(n13321), .Y(n14154) );
  MUX2X1 U14398 ( .B(n14153), .A(n14150), .S(n13269), .Y(n14157) );
  MUX2X1 U14399 ( .B(n14156), .A(n14141), .S(n13101), .Y(n14664) );
  INVX2 U14400 ( .A(n14664), .Y(n87) );
  MUX2X1 U14401 ( .B(n8858), .A(n10882), .S(n13321), .Y(n14161) );
  MUX2X1 U14402 ( .B(n8984), .A(n11008), .S(n13321), .Y(n14160) );
  MUX2X1 U14403 ( .B(n9110), .A(n11134), .S(n13321), .Y(n14164) );
  MUX2X1 U14404 ( .B(n9236), .A(n11260), .S(n13321), .Y(n14163) );
  MUX2X1 U14405 ( .B(n14162), .A(n14159), .S(n13268), .Y(n14173) );
  MUX2X1 U14406 ( .B(n9362), .A(n11386), .S(n13321), .Y(n14167) );
  MUX2X1 U14407 ( .B(n9488), .A(n11512), .S(n13321), .Y(n14166) );
  MUX2X1 U14408 ( .B(n9614), .A(n11638), .S(n13320), .Y(n14170) );
  MUX2X1 U14409 ( .B(n9740), .A(n11764), .S(n13320), .Y(n14169) );
  MUX2X1 U14410 ( .B(n14168), .A(n14165), .S(n13268), .Y(n14172) );
  MUX2X1 U14411 ( .B(n9866), .A(n11890), .S(n13320), .Y(n14176) );
  MUX2X1 U14412 ( .B(n9992), .A(n12016), .S(n13320), .Y(n14175) );
  MUX2X1 U14413 ( .B(n10118), .A(n12142), .S(n13320), .Y(n14179) );
  MUX2X1 U14414 ( .B(n10244), .A(n12268), .S(n13320), .Y(n14178) );
  MUX2X1 U14415 ( .B(n14177), .A(n14174), .S(n13268), .Y(n14188) );
  MUX2X1 U14416 ( .B(n10370), .A(n12394), .S(n13320), .Y(n14182) );
  MUX2X1 U14417 ( .B(n10496), .A(n12520), .S(n13320), .Y(n14181) );
  MUX2X1 U14418 ( .B(n10622), .A(n12646), .S(n13320), .Y(n14185) );
  MUX2X1 U14419 ( .B(n10748), .A(n12772), .S(n13320), .Y(n14184) );
  MUX2X1 U14420 ( .B(n14183), .A(n14180), .S(n13268), .Y(n14187) );
  MUX2X1 U14421 ( .B(n14186), .A(n14171), .S(n13101), .Y(n14665) );
  INVX2 U14422 ( .A(n14665), .Y(n86) );
  MUX2X1 U14423 ( .B(n8861), .A(n10885), .S(n13320), .Y(n14191) );
  MUX2X1 U14424 ( .B(n8987), .A(n11011), .S(n13320), .Y(n14190) );
  MUX2X1 U14425 ( .B(n9113), .A(n11137), .S(n13320), .Y(n14194) );
  MUX2X1 U14426 ( .B(n9239), .A(n11263), .S(n13320), .Y(n14193) );
  MUX2X1 U14427 ( .B(n14192), .A(n14189), .S(n13268), .Y(n14203) );
  MUX2X1 U14428 ( .B(n9365), .A(n11389), .S(n13320), .Y(n14197) );
  MUX2X1 U14429 ( .B(n9491), .A(n11515), .S(n13320), .Y(n14196) );
  MUX2X1 U14430 ( .B(n9617), .A(n11641), .S(n13320), .Y(n14200) );
  MUX2X1 U14431 ( .B(n9743), .A(n11767), .S(n13319), .Y(n14199) );
  MUX2X1 U14432 ( .B(n14198), .A(n14195), .S(n13268), .Y(n14202) );
  MUX2X1 U14433 ( .B(n9869), .A(n11893), .S(n13319), .Y(n14206) );
  MUX2X1 U14434 ( .B(n9995), .A(n12019), .S(n13319), .Y(n14205) );
  MUX2X1 U14435 ( .B(n10121), .A(n12145), .S(n13319), .Y(n14209) );
  MUX2X1 U14436 ( .B(n10247), .A(n12271), .S(n13319), .Y(n14208) );
  MUX2X1 U14437 ( .B(n14207), .A(n14204), .S(n13268), .Y(n14218) );
  MUX2X1 U14438 ( .B(n10373), .A(n12397), .S(n13319), .Y(n14212) );
  MUX2X1 U14439 ( .B(n10499), .A(n12523), .S(n13319), .Y(n14211) );
  MUX2X1 U14440 ( .B(n10625), .A(n12649), .S(n13319), .Y(n14215) );
  MUX2X1 U14441 ( .B(n10751), .A(n12775), .S(n13319), .Y(n14214) );
  MUX2X1 U14442 ( .B(n14213), .A(n14210), .S(n13268), .Y(n14217) );
  MUX2X1 U14443 ( .B(n14216), .A(n14201), .S(n13101), .Y(n14666) );
  INVX2 U14444 ( .A(n14666), .Y(n85) );
  MUX2X1 U14445 ( .B(n8864), .A(n10888), .S(n13319), .Y(n14221) );
  MUX2X1 U14446 ( .B(n8990), .A(n11014), .S(n13319), .Y(n14220) );
  MUX2X1 U14447 ( .B(n9116), .A(n11140), .S(n13319), .Y(n14224) );
  MUX2X1 U14448 ( .B(n9242), .A(n11266), .S(n13319), .Y(n14223) );
  MUX2X1 U14449 ( .B(n14222), .A(n14219), .S(n13268), .Y(n14233) );
  MUX2X1 U14450 ( .B(n9368), .A(n11392), .S(n13319), .Y(n14227) );
  MUX2X1 U14451 ( .B(n9494), .A(n11518), .S(n13319), .Y(n14226) );
  MUX2X1 U14452 ( .B(n9620), .A(n11644), .S(n13319), .Y(n14230) );
  MUX2X1 U14453 ( .B(n9746), .A(n11770), .S(n13319), .Y(n14229) );
  MUX2X1 U14454 ( .B(n14228), .A(n14225), .S(n13268), .Y(n14232) );
  MUX2X1 U14455 ( .B(n9872), .A(n11896), .S(n13318), .Y(n14236) );
  MUX2X1 U14456 ( .B(n9998), .A(n12022), .S(n13318), .Y(n14235) );
  MUX2X1 U14457 ( .B(n10124), .A(n12148), .S(n13318), .Y(n14239) );
  MUX2X1 U14458 ( .B(n10250), .A(n12274), .S(n13318), .Y(n14238) );
  MUX2X1 U14459 ( .B(n14237), .A(n14234), .S(n13268), .Y(n14248) );
  MUX2X1 U14460 ( .B(n10376), .A(n12400), .S(n13318), .Y(n14242) );
  MUX2X1 U14461 ( .B(n10502), .A(n12526), .S(n13318), .Y(n14241) );
  MUX2X1 U14462 ( .B(n10628), .A(n12652), .S(n13318), .Y(n14245) );
  MUX2X1 U14463 ( .B(n10754), .A(n12778), .S(n13318), .Y(n14244) );
  MUX2X1 U14464 ( .B(n14243), .A(n14240), .S(n13268), .Y(n14247) );
  MUX2X1 U14465 ( .B(n14246), .A(n14231), .S(n13101), .Y(n14667) );
  INVX2 U14466 ( .A(n14667), .Y(n84) );
  MUX2X1 U14467 ( .B(n8867), .A(n10891), .S(n13318), .Y(n14251) );
  MUX2X1 U14468 ( .B(n8993), .A(n11017), .S(n13318), .Y(n14250) );
  MUX2X1 U14469 ( .B(n9119), .A(n11143), .S(n13318), .Y(n14254) );
  MUX2X1 U14470 ( .B(n9245), .A(n11269), .S(n13318), .Y(n14253) );
  MUX2X1 U14471 ( .B(n14252), .A(n14249), .S(n13268), .Y(n14263) );
  MUX2X1 U14472 ( .B(n9371), .A(n11395), .S(n13318), .Y(n14257) );
  MUX2X1 U14473 ( .B(n9497), .A(n11521), .S(n13318), .Y(n14256) );
  MUX2X1 U14474 ( .B(n9623), .A(n11647), .S(n13318), .Y(n14260) );
  MUX2X1 U14475 ( .B(n9749), .A(n11773), .S(n13318), .Y(n14259) );
  MUX2X1 U14476 ( .B(n14258), .A(n14255), .S(n13268), .Y(n14262) );
  MUX2X1 U14477 ( .B(n9875), .A(n11899), .S(n13318), .Y(n14266) );
  MUX2X1 U14478 ( .B(n10001), .A(n12025), .S(n13317), .Y(n14265) );
  MUX2X1 U14479 ( .B(n10127), .A(n12151), .S(n13317), .Y(n14269) );
  MUX2X1 U14480 ( .B(n10253), .A(n12277), .S(n13317), .Y(n14268) );
  MUX2X1 U14481 ( .B(n14267), .A(n14264), .S(n13268), .Y(n14278) );
  MUX2X1 U14482 ( .B(n10379), .A(n12403), .S(n13317), .Y(n14272) );
  MUX2X1 U14483 ( .B(n10505), .A(n12529), .S(n13317), .Y(n14271) );
  MUX2X1 U14484 ( .B(n10631), .A(n12655), .S(n13317), .Y(n14275) );
  MUX2X1 U14485 ( .B(n10757), .A(n12781), .S(n13317), .Y(n14274) );
  MUX2X1 U14486 ( .B(n14273), .A(n14270), .S(n13268), .Y(n14277) );
  MUX2X1 U14487 ( .B(n14276), .A(n14261), .S(n13101), .Y(n14668) );
  INVX2 U14488 ( .A(n14668), .Y(n83) );
  MUX2X1 U14489 ( .B(n8870), .A(n10894), .S(n13317), .Y(n14281) );
  MUX2X1 U14490 ( .B(n8996), .A(n11020), .S(n13317), .Y(n14280) );
  MUX2X1 U14491 ( .B(n9122), .A(n11146), .S(n13317), .Y(n14284) );
  MUX2X1 U14492 ( .B(n9248), .A(n11272), .S(n13317), .Y(n14283) );
  MUX2X1 U14493 ( .B(n14282), .A(n14279), .S(n13268), .Y(n14293) );
  MUX2X1 U14494 ( .B(n9374), .A(n11398), .S(n13317), .Y(n14287) );
  MUX2X1 U14495 ( .B(n9500), .A(n11524), .S(n13317), .Y(n14286) );
  MUX2X1 U14496 ( .B(n9626), .A(n11650), .S(n13317), .Y(n14290) );
  MUX2X1 U14497 ( .B(n9752), .A(n11776), .S(n13317), .Y(n14289) );
  MUX2X1 U14498 ( .B(n14288), .A(n14285), .S(n13267), .Y(n14292) );
  MUX2X1 U14499 ( .B(n9878), .A(n11902), .S(n13317), .Y(n14296) );
  MUX2X1 U14500 ( .B(n10004), .A(n12028), .S(n13317), .Y(n14295) );
  MUX2X1 U14501 ( .B(n10130), .A(n12154), .S(n13316), .Y(n14299) );
  MUX2X1 U14502 ( .B(n10256), .A(n12280), .S(n13316), .Y(n14298) );
  MUX2X1 U14503 ( .B(n14297), .A(n14294), .S(n13267), .Y(n14308) );
  MUX2X1 U14504 ( .B(n10382), .A(n12406), .S(n13316), .Y(n14302) );
  MUX2X1 U14505 ( .B(n10508), .A(n12532), .S(n13316), .Y(n14301) );
  MUX2X1 U14506 ( .B(n10634), .A(n12658), .S(n13316), .Y(n14305) );
  MUX2X1 U14507 ( .B(n10760), .A(n12784), .S(n13316), .Y(n14304) );
  MUX2X1 U14508 ( .B(n14303), .A(n14300), .S(n13267), .Y(n14307) );
  MUX2X1 U14509 ( .B(n14306), .A(n14291), .S(n13101), .Y(n14669) );
  INVX2 U14510 ( .A(n14669), .Y(n82) );
  MUX2X1 U14511 ( .B(n8873), .A(n10897), .S(n13316), .Y(n14311) );
  MUX2X1 U14512 ( .B(n8999), .A(n11023), .S(n13316), .Y(n14310) );
  MUX2X1 U14513 ( .B(n9125), .A(n11149), .S(n13316), .Y(n14314) );
  MUX2X1 U14514 ( .B(n9251), .A(n11275), .S(n13316), .Y(n14313) );
  MUX2X1 U14515 ( .B(n14312), .A(n14309), .S(n13267), .Y(n14323) );
  MUX2X1 U14516 ( .B(n9377), .A(n11401), .S(n13316), .Y(n14317) );
  MUX2X1 U14517 ( .B(n9503), .A(n11527), .S(n13316), .Y(n14316) );
  MUX2X1 U14518 ( .B(n9629), .A(n11653), .S(n13316), .Y(n14320) );
  MUX2X1 U14519 ( .B(n9755), .A(n11779), .S(n13321), .Y(n14319) );
  MUX2X1 U14520 ( .B(n14318), .A(n14315), .S(n13267), .Y(n14322) );
  MUX2X1 U14521 ( .B(n9881), .A(n11905), .S(n13335), .Y(n14326) );
  MUX2X1 U14522 ( .B(n10007), .A(n12031), .S(n13335), .Y(n14325) );
  MUX2X1 U14523 ( .B(n10133), .A(n12157), .S(n13335), .Y(n14329) );
  MUX2X1 U14524 ( .B(n10259), .A(n12283), .S(n13335), .Y(n14328) );
  MUX2X1 U14525 ( .B(n14327), .A(n14324), .S(n13267), .Y(n14338) );
  MUX2X1 U14526 ( .B(n10385), .A(n12409), .S(n13335), .Y(n14332) );
  MUX2X1 U14527 ( .B(n10511), .A(n12535), .S(n13335), .Y(n14331) );
  MUX2X1 U14528 ( .B(n10637), .A(n12661), .S(n13335), .Y(n14335) );
  MUX2X1 U14529 ( .B(n10763), .A(n12787), .S(n13335), .Y(n14334) );
  MUX2X1 U14530 ( .B(n14333), .A(n14330), .S(n13267), .Y(n14337) );
  MUX2X1 U14531 ( .B(n14336), .A(n14321), .S(n13101), .Y(n14670) );
  INVX2 U14532 ( .A(n14670), .Y(n81) );
  MUX2X1 U14533 ( .B(n8876), .A(n10900), .S(n13335), .Y(n14341) );
  MUX2X1 U14534 ( .B(n9002), .A(n11026), .S(n13335), .Y(n14340) );
  MUX2X1 U14535 ( .B(n9128), .A(n11152), .S(n13335), .Y(n14344) );
  MUX2X1 U14536 ( .B(n9254), .A(n11278), .S(n13335), .Y(n14343) );
  MUX2X1 U14537 ( .B(n14342), .A(n14339), .S(n13267), .Y(n14353) );
  MUX2X1 U14538 ( .B(n9380), .A(n11404), .S(n13335), .Y(n14347) );
  MUX2X1 U14539 ( .B(n9506), .A(n11530), .S(n13335), .Y(n14346) );
  MUX2X1 U14540 ( .B(n9632), .A(n11656), .S(n13335), .Y(n14350) );
  MUX2X1 U14541 ( .B(n9758), .A(n11782), .S(n13335), .Y(n14349) );
  MUX2X1 U14542 ( .B(n14348), .A(n14345), .S(n13270), .Y(n14352) );
  MUX2X1 U14543 ( .B(n9884), .A(n11908), .S(n13334), .Y(n14356) );
  MUX2X1 U14544 ( .B(n10010), .A(n12034), .S(n13334), .Y(n14355) );
  MUX2X1 U14545 ( .B(n10136), .A(n12160), .S(n13334), .Y(n14359) );
  MUX2X1 U14546 ( .B(n10262), .A(n12286), .S(n13334), .Y(n14358) );
  MUX2X1 U14547 ( .B(n14357), .A(n14354), .S(n13267), .Y(n14368) );
  MUX2X1 U14548 ( .B(n10388), .A(n12412), .S(n13334), .Y(n14362) );
  MUX2X1 U14549 ( .B(n10514), .A(n12538), .S(n13334), .Y(n14361) );
  MUX2X1 U14550 ( .B(n10640), .A(n12664), .S(n13334), .Y(n14365) );
  MUX2X1 U14551 ( .B(n10766), .A(n12790), .S(n13334), .Y(n14364) );
  MUX2X1 U14552 ( .B(n14363), .A(n14360), .S(n13267), .Y(n14367) );
  MUX2X1 U14553 ( .B(n14366), .A(n14351), .S(n13101), .Y(n14671) );
  INVX2 U14554 ( .A(n14671), .Y(n80) );
  MUX2X1 U14555 ( .B(n8879), .A(n10903), .S(n13334), .Y(n14371) );
  MUX2X1 U14556 ( .B(n9005), .A(n11029), .S(n13334), .Y(n14370) );
  MUX2X1 U14557 ( .B(n9131), .A(n11155), .S(n13334), .Y(n14374) );
  MUX2X1 U14558 ( .B(n9257), .A(n11281), .S(n13334), .Y(n14373) );
  MUX2X1 U14559 ( .B(n14372), .A(n14369), .S(n13267), .Y(n14383) );
  MUX2X1 U14560 ( .B(n9383), .A(n11407), .S(n13334), .Y(n14377) );
  MUX2X1 U14561 ( .B(n9509), .A(n11533), .S(n13334), .Y(n14376) );
  MUX2X1 U14562 ( .B(n9635), .A(n11659), .S(n13334), .Y(n14380) );
  MUX2X1 U14563 ( .B(n9761), .A(n11785), .S(n13334), .Y(n14379) );
  MUX2X1 U14564 ( .B(n14378), .A(n14375), .S(n13267), .Y(n14382) );
  MUX2X1 U14565 ( .B(n9887), .A(n11911), .S(n13334), .Y(n14386) );
  MUX2X1 U14566 ( .B(n10013), .A(n12037), .S(n13333), .Y(n14385) );
  MUX2X1 U14567 ( .B(n10139), .A(n12163), .S(n13333), .Y(n14389) );
  MUX2X1 U14568 ( .B(n10265), .A(n12289), .S(n13333), .Y(n14388) );
  MUX2X1 U14569 ( .B(n14387), .A(n14384), .S(n13267), .Y(n14398) );
  MUX2X1 U14570 ( .B(n10391), .A(n12415), .S(n13333), .Y(n14392) );
  MUX2X1 U14571 ( .B(n10517), .A(n12541), .S(n13333), .Y(n14391) );
  MUX2X1 U14572 ( .B(n10643), .A(n12667), .S(n13333), .Y(n14395) );
  MUX2X1 U14573 ( .B(n10769), .A(n12793), .S(n13333), .Y(n14394) );
  MUX2X1 U14574 ( .B(n14393), .A(n14390), .S(n13267), .Y(n14397) );
  MUX2X1 U14575 ( .B(n14396), .A(n14381), .S(n13101), .Y(n14672) );
  INVX2 U14576 ( .A(n14672), .Y(n79) );
  MUX2X1 U14577 ( .B(n8882), .A(n10906), .S(n13333), .Y(n14401) );
  MUX2X1 U14578 ( .B(n9008), .A(n11032), .S(n13333), .Y(n14400) );
  MUX2X1 U14579 ( .B(n9134), .A(n11158), .S(n13333), .Y(n14404) );
  MUX2X1 U14580 ( .B(n9260), .A(n11284), .S(n13333), .Y(n14403) );
  MUX2X1 U14581 ( .B(n14402), .A(n14399), .S(n13267), .Y(n14413) );
  MUX2X1 U14582 ( .B(n9386), .A(n11410), .S(n13333), .Y(n14407) );
  MUX2X1 U14583 ( .B(n9512), .A(n11536), .S(n13333), .Y(n14406) );
  MUX2X1 U14584 ( .B(n9638), .A(n11662), .S(n13333), .Y(n14410) );
  MUX2X1 U14585 ( .B(n9764), .A(n11788), .S(n13333), .Y(n14409) );
  MUX2X1 U14586 ( .B(n14408), .A(n14405), .S(n13267), .Y(n14412) );
  MUX2X1 U14587 ( .B(n9890), .A(n11914), .S(n13333), .Y(n14416) );
  MUX2X1 U14588 ( .B(n10016), .A(n12040), .S(n13333), .Y(n14415) );
  MUX2X1 U14589 ( .B(n10142), .A(n12166), .S(n13332), .Y(n14419) );
  MUX2X1 U14590 ( .B(n10268), .A(n12292), .S(n13332), .Y(n14418) );
  MUX2X1 U14591 ( .B(n14417), .A(n14414), .S(n13267), .Y(n14428) );
  MUX2X1 U14592 ( .B(n10394), .A(n12418), .S(n13332), .Y(n14422) );
  MUX2X1 U14593 ( .B(n10520), .A(n12544), .S(n13332), .Y(n14421) );
  MUX2X1 U14594 ( .B(n10646), .A(n12670), .S(n13332), .Y(n14425) );
  MUX2X1 U14595 ( .B(n10772), .A(n12796), .S(n13332), .Y(n14424) );
  MUX2X1 U14596 ( .B(n14423), .A(n14420), .S(n13266), .Y(n14427) );
  MUX2X1 U14597 ( .B(n14426), .A(n14411), .S(n13101), .Y(n14673) );
  INVX2 U14598 ( .A(n14673), .Y(n78) );
  MUX2X1 U14599 ( .B(n8885), .A(n10909), .S(n13332), .Y(n14431) );
  MUX2X1 U14600 ( .B(n9011), .A(n11035), .S(n13332), .Y(n14430) );
  MUX2X1 U14601 ( .B(n9137), .A(n11161), .S(n13332), .Y(n14434) );
  MUX2X1 U14602 ( .B(n9263), .A(n11287), .S(n13332), .Y(n14433) );
  MUX2X1 U14603 ( .B(n14432), .A(n14429), .S(n13266), .Y(n14443) );
  MUX2X1 U14604 ( .B(n9389), .A(n11413), .S(n13332), .Y(n14437) );
  MUX2X1 U14605 ( .B(n9515), .A(n11539), .S(n13332), .Y(n14436) );
  MUX2X1 U14606 ( .B(n9641), .A(n11665), .S(n13332), .Y(n14440) );
  MUX2X1 U14607 ( .B(n9767), .A(n11791), .S(n13332), .Y(n14439) );
  MUX2X1 U14608 ( .B(n14438), .A(n14435), .S(n13266), .Y(n14442) );
  MUX2X1 U14609 ( .B(n9893), .A(n11917), .S(n13332), .Y(n14446) );
  MUX2X1 U14610 ( .B(n10019), .A(n12043), .S(n13332), .Y(n14445) );
  MUX2X1 U14611 ( .B(n10145), .A(n12169), .S(n13332), .Y(n14449) );
  MUX2X1 U14612 ( .B(n10271), .A(n12295), .S(n13331), .Y(n14448) );
  MUX2X1 U14613 ( .B(n14447), .A(n14444), .S(n13266), .Y(n14458) );
  MUX2X1 U14614 ( .B(n10397), .A(n12421), .S(n13331), .Y(n14452) );
  MUX2X1 U14615 ( .B(n10523), .A(n12547), .S(n13331), .Y(n14451) );
  MUX2X1 U14616 ( .B(n10649), .A(n12673), .S(n13331), .Y(n14455) );
  MUX2X1 U14617 ( .B(n10775), .A(n12799), .S(n13331), .Y(n14454) );
  MUX2X1 U14618 ( .B(n14453), .A(n14450), .S(n13266), .Y(n14457) );
  MUX2X1 U14619 ( .B(n14456), .A(n14441), .S(n13101), .Y(n14674) );
  INVX2 U14620 ( .A(n14674), .Y(n77) );
  MUX2X1 U14621 ( .B(n8888), .A(n10912), .S(n13331), .Y(n14461) );
  MUX2X1 U14622 ( .B(n9014), .A(n11038), .S(n13331), .Y(n14460) );
  MUX2X1 U14623 ( .B(n9140), .A(n11164), .S(n13331), .Y(n14464) );
  MUX2X1 U14624 ( .B(n9266), .A(n11290), .S(n13331), .Y(n14463) );
  MUX2X1 U14625 ( .B(n14462), .A(n14459), .S(n13266), .Y(n14473) );
  MUX2X1 U14626 ( .B(n9392), .A(n11416), .S(n13331), .Y(n14467) );
  MUX2X1 U14627 ( .B(n9518), .A(n11542), .S(n13331), .Y(n14466) );
  MUX2X1 U14628 ( .B(n9644), .A(n11668), .S(n13331), .Y(n14470) );
  MUX2X1 U14629 ( .B(n9770), .A(n11794), .S(n13331), .Y(n14469) );
  MUX2X1 U14630 ( .B(n14468), .A(n14465), .S(n13266), .Y(n14472) );
  MUX2X1 U14631 ( .B(n9896), .A(n11920), .S(n13331), .Y(n14476) );
  MUX2X1 U14632 ( .B(n10022), .A(n12046), .S(n13331), .Y(n14475) );
  MUX2X1 U14633 ( .B(n10148), .A(n12172), .S(n13331), .Y(n14479) );
  MUX2X1 U14634 ( .B(n10274), .A(n12298), .S(n13331), .Y(n14478) );
  MUX2X1 U14635 ( .B(n14477), .A(n14474), .S(n13266), .Y(n14488) );
  MUX2X1 U14636 ( .B(n10400), .A(n12424), .S(n13330), .Y(n14482) );
  MUX2X1 U14637 ( .B(n10526), .A(n12550), .S(n13330), .Y(n14481) );
  MUX2X1 U14638 ( .B(n10652), .A(n12676), .S(n13330), .Y(n14485) );
  MUX2X1 U14639 ( .B(n10778), .A(n12802), .S(n13330), .Y(n14484) );
  MUX2X1 U14640 ( .B(n14483), .A(n14480), .S(n13266), .Y(n14487) );
  MUX2X1 U14641 ( .B(n14486), .A(n14471), .S(n13101), .Y(n14675) );
  INVX2 U14642 ( .A(n14675), .Y(n76) );
  MUX2X1 U14643 ( .B(n8891), .A(n10915), .S(n13330), .Y(n14491) );
  MUX2X1 U14644 ( .B(n9017), .A(n11041), .S(n13330), .Y(n14490) );
  MUX2X1 U14645 ( .B(n9143), .A(n11167), .S(n13330), .Y(n14494) );
  MUX2X1 U14646 ( .B(n9269), .A(n11293), .S(n13330), .Y(n14493) );
  MUX2X1 U14647 ( .B(n14492), .A(n14489), .S(n13266), .Y(n14503) );
  MUX2X1 U14648 ( .B(n9395), .A(n11419), .S(n13330), .Y(n14497) );
  MUX2X1 U14649 ( .B(n9521), .A(n11545), .S(n13330), .Y(n14496) );
  MUX2X1 U14650 ( .B(n9647), .A(n11671), .S(n13330), .Y(n14500) );
  MUX2X1 U14651 ( .B(n9773), .A(n11797), .S(n13330), .Y(n14499) );
  MUX2X1 U14652 ( .B(n14498), .A(n14495), .S(n13266), .Y(n14502) );
  MUX2X1 U14653 ( .B(n9899), .A(n11923), .S(n13330), .Y(n14506) );
  MUX2X1 U14654 ( .B(n10025), .A(n12049), .S(n13330), .Y(n14505) );
  MUX2X1 U14655 ( .B(n10151), .A(n12175), .S(n13330), .Y(n14509) );
  MUX2X1 U14656 ( .B(n10277), .A(n12301), .S(n13330), .Y(n14508) );
  MUX2X1 U14657 ( .B(n14507), .A(n14504), .S(n13266), .Y(n14518) );
  MUX2X1 U14658 ( .B(n10403), .A(n12427), .S(n13329), .Y(n14512) );
  MUX2X1 U14659 ( .B(n10529), .A(n12553), .S(n13329), .Y(n14511) );
  MUX2X1 U14660 ( .B(n10655), .A(n12679), .S(n13329), .Y(n14515) );
  MUX2X1 U14661 ( .B(n10781), .A(n12805), .S(n13329), .Y(n14514) );
  MUX2X1 U14662 ( .B(n14513), .A(n14510), .S(n13266), .Y(n14517) );
  MUX2X1 U14663 ( .B(n14516), .A(n14501), .S(n13101), .Y(n14676) );
  INVX2 U14664 ( .A(n14676), .Y(n75) );
  MUX2X1 U14665 ( .B(n8894), .A(n10918), .S(n13329), .Y(n14521) );
  MUX2X1 U14666 ( .B(n9020), .A(n11044), .S(n13329), .Y(n14520) );
  MUX2X1 U14667 ( .B(n9146), .A(n11170), .S(n13329), .Y(n14524) );
  MUX2X1 U14668 ( .B(n9272), .A(n11296), .S(n13329), .Y(n14523) );
  MUX2X1 U14669 ( .B(n14522), .A(n14519), .S(n13266), .Y(n14533) );
  MUX2X1 U14670 ( .B(n9398), .A(n11422), .S(n13329), .Y(n14527) );
  MUX2X1 U14671 ( .B(n9524), .A(n11548), .S(n13329), .Y(n14526) );
  MUX2X1 U14672 ( .B(n9650), .A(n11674), .S(n13329), .Y(n14530) );
  MUX2X1 U14673 ( .B(n9776), .A(n11800), .S(n13329), .Y(n14529) );
  MUX2X1 U14674 ( .B(n14528), .A(n14525), .S(n13266), .Y(n14532) );
  MUX2X1 U14675 ( .B(n9902), .A(n11926), .S(n13329), .Y(n14536) );
  MUX2X1 U14676 ( .B(n10028), .A(n12052), .S(n13329), .Y(n14535) );
  MUX2X1 U14677 ( .B(n10154), .A(n12178), .S(n13329), .Y(n14539) );
  MUX2X1 U14678 ( .B(n10280), .A(n12304), .S(n13329), .Y(n14538) );
  MUX2X1 U14679 ( .B(n14537), .A(n14534), .S(n13266), .Y(n14548) );
  MUX2X1 U14680 ( .B(n10406), .A(n12430), .S(n13329), .Y(n14542) );
  MUX2X1 U14681 ( .B(n10532), .A(n12556), .S(n13328), .Y(n14541) );
  MUX2X1 U14682 ( .B(n10658), .A(n12682), .S(n13328), .Y(n14545) );
  MUX2X1 U14683 ( .B(n10784), .A(n12808), .S(n13328), .Y(n14544) );
  MUX2X1 U14684 ( .B(n14543), .A(n14540), .S(n13266), .Y(n14547) );
  MUX2X1 U14685 ( .B(n14546), .A(n14531), .S(n13101), .Y(n14677) );
  INVX2 U14686 ( .A(n14677), .Y(n74) );
  MUX2X1 U14687 ( .B(n8897), .A(n10921), .S(n13328), .Y(n14551) );
  MUX2X1 U14688 ( .B(n9023), .A(n11047), .S(n13328), .Y(n14550) );
  MUX2X1 U14689 ( .B(n9149), .A(n11173), .S(n13328), .Y(n14554) );
  MUX2X1 U14690 ( .B(n9275), .A(n11299), .S(n13328), .Y(n14553) );
  MUX2X1 U14691 ( .B(n14552), .A(n14549), .S(n13265), .Y(n14563) );
  MUX2X1 U14692 ( .B(n9401), .A(n11425), .S(n13328), .Y(n14557) );
  MUX2X1 U14693 ( .B(n9527), .A(n11551), .S(n13328), .Y(n14556) );
  MUX2X1 U14694 ( .B(n9653), .A(n11677), .S(n13328), .Y(n14560) );
  MUX2X1 U14695 ( .B(n9779), .A(n11803), .S(n13328), .Y(n14559) );
  MUX2X1 U14696 ( .B(n14558), .A(n14555), .S(n13265), .Y(n14562) );
  MUX2X1 U14697 ( .B(n9905), .A(n11929), .S(n13328), .Y(n14566) );
  MUX2X1 U14698 ( .B(n10031), .A(n12055), .S(n13328), .Y(n14565) );
  MUX2X1 U14699 ( .B(n10157), .A(n12181), .S(n13328), .Y(n14569) );
  MUX2X1 U14700 ( .B(n10283), .A(n12307), .S(n13328), .Y(n14568) );
  MUX2X1 U14701 ( .B(n14567), .A(n14564), .S(n13265), .Y(n14578) );
  MUX2X1 U14702 ( .B(n10409), .A(n12433), .S(n13328), .Y(n14572) );
  MUX2X1 U14703 ( .B(n10535), .A(n12559), .S(n13328), .Y(n14571) );
  MUX2X1 U14704 ( .B(n10661), .A(n12685), .S(n13327), .Y(n14575) );
  MUX2X1 U14705 ( .B(n10787), .A(n12811), .S(n13327), .Y(n14574) );
  MUX2X1 U14706 ( .B(n14573), .A(n14570), .S(n13265), .Y(n14577) );
  MUX2X1 U14707 ( .B(n14576), .A(n14561), .S(n13101), .Y(n14678) );
  INVX2 U14708 ( .A(n14678), .Y(n73) );
  MUX2X1 U14709 ( .B(n8900), .A(n10924), .S(n13327), .Y(n14581) );
  MUX2X1 U14710 ( .B(n9026), .A(n11050), .S(n13327), .Y(n14580) );
  MUX2X1 U14711 ( .B(n9152), .A(n11176), .S(n13327), .Y(n14584) );
  MUX2X1 U14712 ( .B(n9278), .A(n11302), .S(n13327), .Y(n14583) );
  MUX2X1 U14713 ( .B(n14582), .A(n14579), .S(n13265), .Y(n14593) );
  MUX2X1 U14714 ( .B(n9404), .A(n11428), .S(n13327), .Y(n14587) );
  MUX2X1 U14715 ( .B(n9530), .A(n11554), .S(n13327), .Y(n14586) );
  MUX2X1 U14716 ( .B(n9656), .A(n11680), .S(n13327), .Y(n14590) );
  MUX2X1 U14717 ( .B(n9782), .A(n11806), .S(n13327), .Y(n14589) );
  MUX2X1 U14718 ( .B(n14588), .A(n14585), .S(n13265), .Y(n14592) );
  MUX2X1 U14719 ( .B(n9908), .A(n11932), .S(n13327), .Y(n14596) );
  MUX2X1 U14720 ( .B(n10034), .A(n12058), .S(n13327), .Y(n14595) );
  MUX2X1 U14721 ( .B(n10160), .A(n12184), .S(n13327), .Y(n14599) );
  MUX2X1 U14722 ( .B(n10286), .A(n12310), .S(n13327), .Y(n14598) );
  MUX2X1 U14723 ( .B(n14597), .A(n14594), .S(n13265), .Y(n14608) );
  MUX2X1 U14724 ( .B(n10412), .A(n12436), .S(n13327), .Y(n14602) );
  MUX2X1 U14725 ( .B(n10538), .A(n12562), .S(n13327), .Y(n14601) );
  MUX2X1 U14726 ( .B(n10664), .A(n12688), .S(n13327), .Y(n14605) );
  MUX2X1 U14727 ( .B(n10790), .A(n12814), .S(n13326), .Y(n14604) );
  MUX2X1 U14728 ( .B(n14603), .A(n14600), .S(n13265), .Y(n14607) );
  MUX2X1 U14729 ( .B(n14606), .A(n14591), .S(n13101), .Y(n14679) );
  INVX2 U14730 ( .A(n14679), .Y(n72) );
  MUX2X1 U14731 ( .B(n8903), .A(n10927), .S(n13326), .Y(n14611) );
  MUX2X1 U14732 ( .B(n9029), .A(n11053), .S(n13326), .Y(n14610) );
  MUX2X1 U14733 ( .B(n9155), .A(n11179), .S(n13326), .Y(n14614) );
  MUX2X1 U14734 ( .B(n9281), .A(n11305), .S(n13326), .Y(n14613) );
  MUX2X1 U14735 ( .B(n14612), .A(n14609), .S(n13265), .Y(n14623) );
  MUX2X1 U14736 ( .B(n9407), .A(n11431), .S(n13326), .Y(n14617) );
  MUX2X1 U14737 ( .B(n9533), .A(n11557), .S(n13326), .Y(n14616) );
  MUX2X1 U14738 ( .B(n9659), .A(n11683), .S(n13326), .Y(n14620) );
  MUX2X1 U14739 ( .B(n9785), .A(n11809), .S(n13326), .Y(n14619) );
  MUX2X1 U14740 ( .B(n14618), .A(n14615), .S(n13265), .Y(n14622) );
  MUX2X1 U14741 ( .B(n9911), .A(n11935), .S(n13326), .Y(n14626) );
  MUX2X1 U14742 ( .B(n10037), .A(n12061), .S(n13326), .Y(n14625) );
  MUX2X1 U14743 ( .B(n10163), .A(n12187), .S(n13326), .Y(n14629) );
  MUX2X1 U14744 ( .B(n10289), .A(n12313), .S(n13326), .Y(n14628) );
  MUX2X1 U14745 ( .B(n14627), .A(n14624), .S(n13265), .Y(n14638) );
  MUX2X1 U14746 ( .B(n10415), .A(n12439), .S(n13326), .Y(n14632) );
  MUX2X1 U14747 ( .B(n10541), .A(n12565), .S(n13326), .Y(n14631) );
  MUX2X1 U14748 ( .B(n10667), .A(n12691), .S(n13326), .Y(n14635) );
  MUX2X1 U14749 ( .B(n10793), .A(n12817), .S(n13330), .Y(n14634) );
  MUX2X1 U14750 ( .B(n14633), .A(n14630), .S(n13265), .Y(n14637) );
  MUX2X1 U14751 ( .B(n14636), .A(n14621), .S(n13101), .Y(n14680) );
  INVX2 U14752 ( .A(n14680), .Y(n71) );
  XOR2X1 U14753 ( .A(add_158_carry[5]), .B(n12995), .Y(n38) );
  XOR2X1 U14754 ( .A(add_176_carry[5]), .B(n12981), .Y(n118) );
endmodule


module ddr3_init_engine_DW01_inc_0 ( A, SUM );
  input [18:0] A;
  output [18:0] SUM;

  wire   [18:2] carry;

  HAX1 U1_1_17 ( .A(A[17]), .B(carry[17]), .YC(carry[18]), .YS(SUM[17]) );
  HAX1 U1_1_16 ( .A(A[16]), .B(carry[16]), .YC(carry[17]), .YS(SUM[16]) );
  HAX1 U1_1_15 ( .A(A[15]), .B(carry[15]), .YC(carry[16]), .YS(SUM[15]) );
  HAX1 U1_1_14 ( .A(A[14]), .B(carry[14]), .YC(carry[15]), .YS(SUM[14]) );
  HAX1 U1_1_13 ( .A(A[13]), .B(carry[13]), .YC(carry[14]), .YS(SUM[13]) );
  HAX1 U1_1_12 ( .A(A[12]), .B(carry[12]), .YC(carry[13]), .YS(SUM[12]) );
  HAX1 U1_1_11 ( .A(A[11]), .B(carry[11]), .YC(carry[12]), .YS(SUM[11]) );
  HAX1 U1_1_10 ( .A(A[10]), .B(carry[10]), .YC(carry[11]), .YS(SUM[10]) );
  HAX1 U1_1_9 ( .A(A[9]), .B(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  HAX1 U1_1_8 ( .A(A[8]), .B(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  HAX1 U1_1_7 ( .A(A[7]), .B(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  HAX1 U1_1_6 ( .A(A[6]), .B(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  HAX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry[2]), .YS(SUM[1]) );
  XOR2X1 U1 ( .A(carry[18]), .B(A[18]), .Y(SUM[18]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module ddr3_init_engine ( ready, csbar, rasbar, casbar, webar, ba, a, odt, 
        ts_con, cke, clk, reset, init, ck, reset_out );
  output [2:0] ba;
  output [12:0] a;
  input clk, reset, init, ck;
  output ready, csbar, rasbar, casbar, webar, odt, ts_con, cke, reset_out;
  wire   flag, RESET, INIT, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n326, n327, n332, n335,
         n1, n2, n3, n4, n5, n6, n7, n8, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n328, n329, n330, n331, n333, n334, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396;
  wire   [18:0] counter;
  assign csbar = 1'b0;
  assign ba[2] = 1'b0;
  assign a[12] = 1'b0;
  assign a[11] = 1'b0;
  assign a[9] = 1'b0;
  assign a[7] = 1'b0;
  assign a[6] = 1'b0;
  assign a[5] = 1'b0;
  assign a[3] = 1'b0;
  assign a[2] = 1'b0;
  assign a[1] = 1'b0;
  assign a[0] = 1'b0;
  assign odt = 1'b0;
  assign ts_con = 1'b0;

  DFFPOSX1 RESET_reg ( .D(reset), .CLK(clk), .Q(RESET) );
  DFFPOSX1 INIT_reg ( .D(init), .CLK(clk), .Q(INIT) );
  DFFPOSX1 flag_reg ( .D(n179), .CLK(clk), .Q(flag) );
  DFFPOSX1 counter_reg_17_ ( .D(n160), .CLK(clk), .Q(counter[17]) );
  DFFPOSX1 counter_reg_0_ ( .D(n177), .CLK(clk), .Q(counter[0]) );
  DFFPOSX1 counter_reg_1_ ( .D(n176), .CLK(clk), .Q(counter[1]) );
  DFFPOSX1 counter_reg_2_ ( .D(n175), .CLK(clk), .Q(counter[2]) );
  DFFPOSX1 counter_reg_3_ ( .D(n174), .CLK(clk), .Q(counter[3]) );
  DFFPOSX1 counter_reg_4_ ( .D(n173), .CLK(clk), .Q(counter[4]) );
  DFFPOSX1 counter_reg_5_ ( .D(n172), .CLK(clk), .Q(counter[5]) );
  DFFPOSX1 counter_reg_6_ ( .D(n171), .CLK(clk), .Q(counter[6]) );
  DFFPOSX1 counter_reg_7_ ( .D(n170), .CLK(clk), .Q(counter[7]) );
  DFFPOSX1 counter_reg_8_ ( .D(n169), .CLK(clk), .Q(counter[8]) );
  DFFPOSX1 counter_reg_9_ ( .D(n168), .CLK(clk), .Q(counter[9]) );
  DFFPOSX1 counter_reg_10_ ( .D(n167), .CLK(clk), .Q(counter[10]) );
  DFFPOSX1 counter_reg_11_ ( .D(n166), .CLK(clk), .Q(counter[11]) );
  DFFPOSX1 counter_reg_12_ ( .D(n165), .CLK(clk), .Q(counter[12]) );
  DFFPOSX1 counter_reg_13_ ( .D(n164), .CLK(clk), .Q(counter[13]) );
  DFFPOSX1 counter_reg_14_ ( .D(n163), .CLK(clk), .Q(counter[14]) );
  DFFPOSX1 counter_reg_15_ ( .D(n162), .CLK(clk), .Q(counter[15]) );
  DFFPOSX1 counter_reg_16_ ( .D(n161), .CLK(clk), .Q(counter[16]) );
  DFFPOSX1 counter_reg_18_ ( .D(n178), .CLK(clk), .Q(counter[18]) );
  DFFPOSX1 ready_reg ( .D(n156), .CLK(clk), .Q(ready) );
  DFFPOSX1 rasbar_reg ( .D(n220), .CLK(clk), .Q(rasbar) );
  DFFPOSX1 casbar_reg ( .D(n217), .CLK(clk), .Q(casbar) );
  DFFPOSX1 webar_reg ( .D(n223), .CLK(clk), .Q(webar) );
  DFFPOSX1 reset_out_reg ( .D(n155), .CLK(clk), .Q(reset_out) );
  DFFPOSX1 cke_reg ( .D(n154), .CLK(clk), .Q(cke) );
  DFFPOSX1 a_reg_10_ ( .D(n153), .CLK(clk), .Q(a[10]) );
  DFFPOSX1 a_reg_8_ ( .D(n226), .CLK(clk), .Q(a[8]) );
  DFFPOSX1 a_reg_4_ ( .D(n181), .CLK(clk), .Q(a[4]) );
  DFFPOSX1 ba_reg_1_ ( .D(n150), .CLK(clk), .Q(ba[1]) );
  DFFPOSX1 ba_reg_0_ ( .D(n229), .CLK(clk), .Q(ba[0]) );
  NAND3X1 U18 ( .A(n365), .B(n332), .C(n4), .Y(n2) );
  OAI21X1 U20 ( .A(n395), .B(n7), .C(n295), .Y(n150) );
  INVX1 U22 ( .A(n28), .Y(n7) );
  AOI21X1 U23 ( .A(n383), .B(n380), .C(n5), .Y(n28) );
  INVX1 U24 ( .A(n332), .Y(n5) );
  NAND3X1 U25 ( .A(n205), .B(n356), .C(n316), .Y(n151) );
  NAND3X1 U27 ( .A(n4), .B(n326), .C(n35), .Y(n31) );
  INVX1 U28 ( .A(n374), .Y(n35) );
  NAND3X1 U31 ( .A(n4), .B(n326), .C(n38), .Y(n32) );
  OAI21X1 U32 ( .A(n395), .B(n39), .C(n292), .Y(n153) );
  OAI21X1 U34 ( .A(n42), .B(n38), .C(n43), .Y(n39) );
  INVX1 U35 ( .A(n344), .Y(n43) );
  AOI21X1 U36 ( .A(n44), .B(n42), .C(n326), .Y(n41) );
  OAI21X1 U37 ( .A(n45), .B(n395), .C(n290), .Y(n154) );
  NAND3X1 U40 ( .A(n49), .B(n377), .C(n313), .Y(n48) );
  OAI21X1 U42 ( .A(n54), .B(n395), .C(n289), .Y(n155) );
  NAND3X1 U45 ( .A(n57), .B(n58), .C(n59), .Y(n56) );
  NOR3X1 U46 ( .A(n325), .B(n392), .C(n341), .Y(n59) );
  NAND3X1 U48 ( .A(counter[14]), .B(n63), .C(counter[16]), .Y(n60) );
  NOR3X1 U49 ( .A(counter[18]), .B(counter[5]), .C(counter[1]), .Y(n58) );
  NOR3X1 U50 ( .A(n371), .B(counter[17]), .C(counter[10]), .Y(n57) );
  OAI21X1 U51 ( .A(n65), .B(n395), .C(n288), .Y(n156) );
  NAND3X1 U54 ( .A(counter[1]), .B(counter[10]), .C(n68), .Y(n67) );
  AND2X1 U55 ( .A(n44), .B(n69), .Y(n68) );
  NAND3X1 U57 ( .A(n335), .B(n72), .C(n4), .Y(n71) );
  INVX1 U63 ( .A(n335), .Y(n73) );
  NAND3X1 U64 ( .A(n335), .B(n77), .C(n4), .Y(n74) );
  OAI21X1 U65 ( .A(n179), .B(n78), .C(n286), .Y(n160) );
  INVX1 U67 ( .A(counter[17]), .Y(n78) );
  OAI21X1 U68 ( .A(n179), .B(n81), .C(n283), .Y(n161) );
  OAI21X1 U70 ( .A(n179), .B(n83), .C(n280), .Y(n162) );
  INVX1 U72 ( .A(counter[15]), .Y(n83) );
  OAI21X1 U73 ( .A(n179), .B(n85), .C(n277), .Y(n163) );
  OAI21X1 U75 ( .A(n179), .B(n87), .C(n274), .Y(n164) );
  INVX1 U77 ( .A(counter[13]), .Y(n87) );
  OAI21X1 U78 ( .A(n179), .B(n89), .C(n271), .Y(n165) );
  OAI21X1 U80 ( .A(n179), .B(n91), .C(n268), .Y(n166) );
  INVX1 U82 ( .A(counter[11]), .Y(n91) );
  OAI21X1 U83 ( .A(n179), .B(n93), .C(n265), .Y(n167) );
  OAI21X1 U85 ( .A(n179), .B(n95), .C(n262), .Y(n168) );
  OAI21X1 U87 ( .A(n179), .B(n97), .C(n259), .Y(n169) );
  OAI21X1 U89 ( .A(n179), .B(n99), .C(n256), .Y(n170) );
  OAI21X1 U91 ( .A(n179), .B(n101), .C(n253), .Y(n171) );
  OAI21X1 U93 ( .A(n179), .B(n103), .C(n250), .Y(n172) );
  OAI21X1 U95 ( .A(n179), .B(n105), .C(n247), .Y(n173) );
  OAI21X1 U97 ( .A(n179), .B(n107), .C(n244), .Y(n174) );
  OAI21X1 U99 ( .A(n179), .B(n109), .C(n241), .Y(n175) );
  OAI21X1 U101 ( .A(n179), .B(n111), .C(n238), .Y(n176) );
  OAI21X1 U103 ( .A(n179), .B(n113), .C(n235), .Y(n177) );
  OAI21X1 U105 ( .A(n179), .B(n115), .C(n232), .Y(n178) );
  AND2X1 U107 ( .A(n179), .B(n359), .Y(n80) );
  INVX1 U108 ( .A(counter[18]), .Y(n115) );
  OAI21X1 U109 ( .A(RESET), .B(n359), .C(n395), .Y(n179) );
  INVX1 U111 ( .A(flag), .Y(n118) );
  OAI21X1 U112 ( .A(n119), .B(n392), .C(n47), .Y(n335) );
  NOR3X1 U113 ( .A(n330), .B(n77), .C(n365), .Y(n119) );
  OR2X1 U115 ( .A(n72), .B(n42), .Y(n77) );
  INVX1 U116 ( .A(n121), .Y(n42) );
  NAND3X1 U117 ( .A(n93), .B(n111), .C(n69), .Y(n121) );
  OAI21X1 U118 ( .A(n211), .B(n111), .C(n199), .Y(n72) );
  AOI21X1 U119 ( .A(n124), .B(counter[2]), .C(n125), .Y(n123) );
  NOR3X1 U120 ( .A(n322), .B(n386), .C(n105), .Y(n125) );
  NAND3X1 U121 ( .A(n111), .B(n109), .C(counter[3]), .Y(n126) );
  INVX1 U122 ( .A(n128), .Y(n124) );
  OAI21X1 U123 ( .A(n214), .B(n130), .C(n111), .Y(n128) );
  AOI21X1 U124 ( .A(n208), .B(n132), .C(n353), .Y(n129) );
  NAND3X1 U125 ( .A(counter[4]), .B(counter[6]), .C(n133), .Y(n53) );
  NOR3X1 U126 ( .A(n103), .B(counter[8]), .C(n99), .Y(n133) );
  INVX1 U127 ( .A(n377), .Y(n132) );
  NAND3X1 U128 ( .A(counter[3]), .B(n95), .C(n134), .Y(n131) );
  INVX1 U129 ( .A(counter[9]), .Y(n95) );
  AOI21X1 U130 ( .A(n135), .B(n62), .C(n69), .Y(n122) );
  AND2X1 U131 ( .A(n136), .B(n137), .Y(n69) );
  NOR3X1 U132 ( .A(n319), .B(counter[2]), .C(counter[11]), .Y(n137) );
  NAND3X1 U133 ( .A(n105), .B(n101), .C(n107), .Y(n138) );
  NOR3X1 U134 ( .A(n334), .B(n368), .C(n103), .Y(n136) );
  NOR3X1 U136 ( .A(counter[8]), .B(counter[9]), .C(counter[7]), .Y(n63) );
  OAI21X1 U138 ( .A(n392), .B(n383), .C(n389), .Y(n332) );
  NAND3X1 U139 ( .A(counter[2]), .B(counter[4]), .C(n142), .Y(n29) );
  NOR3X1 U140 ( .A(n386), .B(counter[3]), .C(n111), .Y(n142) );
  INVX1 U141 ( .A(n389), .Y(n326) );
  AOI21X1 U142 ( .A(n44), .B(n38), .C(n327), .Y(n34) );
  OR2X1 U143 ( .A(RESET), .B(n202), .Y(n327) );
  AOI21X1 U144 ( .A(n374), .B(n380), .C(n392), .Y(n143) );
  NAND3X1 U145 ( .A(n62), .B(n111), .C(n135), .Y(n30) );
  INVX1 U146 ( .A(n386), .Y(n135) );
  NAND3X1 U147 ( .A(counter[6]), .B(counter[5]), .C(n144), .Y(n127) );
  NOR3X1 U148 ( .A(n97), .B(counter[7]), .C(n362), .Y(n144) );
  INVX1 U149 ( .A(counter[1]), .Y(n111) );
  NOR3X1 U150 ( .A(counter[2]), .B(counter[4]), .C(n107), .Y(n62) );
  INVX1 U151 ( .A(counter[3]), .Y(n107) );
  NAND3X1 U152 ( .A(n49), .B(n105), .C(n130), .Y(n36) );
  INVX1 U153 ( .A(counter[4]), .Y(n105) );
  INVX1 U154 ( .A(n347), .Y(n38) );
  NAND3X1 U155 ( .A(n130), .B(n49), .C(counter[4]), .Y(n141) );
  AND2X1 U156 ( .A(counter[1]), .B(n109), .Y(n49) );
  INVX1 U157 ( .A(counter[2]), .Y(n109) );
  NOR3X1 U158 ( .A(n97), .B(n99), .C(n338), .Y(n130) );
  NAND3X1 U159 ( .A(n377), .B(n101), .C(n103), .Y(n146) );
  INVX1 U160 ( .A(counter[5]), .Y(n103) );
  INVX1 U161 ( .A(counter[6]), .Y(n101) );
  NOR3X1 U164 ( .A(n368), .B(n371), .C(n93), .Y(n134) );
  INVX1 U165 ( .A(counter[10]), .Y(n93) );
  INVX1 U167 ( .A(counter[12]), .Y(n89) );
  NAND3X1 U168 ( .A(counter[18]), .B(counter[17]), .C(n147), .Y(n140) );
  AND2X1 U169 ( .A(n81), .B(n85), .Y(n147) );
  INVX1 U170 ( .A(counter[14]), .Y(n85) );
  INVX1 U171 ( .A(counter[16]), .Y(n81) );
  INVX1 U172 ( .A(counter[7]), .Y(n99) );
  INVX1 U173 ( .A(counter[8]), .Y(n97) );
  INVX1 U174 ( .A(n392), .Y(n44) );
  NAND3X1 U175 ( .A(n4), .B(counter[15]), .C(n148), .Y(n52) );
  AND2X1 U176 ( .A(n113), .B(counter[13]), .Y(n148) );
  INVX1 U177 ( .A(counter[0]), .Y(n113) );
  INVX1 U178 ( .A(n395), .Y(n4) );
  INVX1 U180 ( .A(RESET), .Y(n47) );
  ddr3_init_engine_DW01_inc_0 add_88 ( .A(counter), .SUM({n27, n26, n25, n24, 
        n23, n22, n21, n20, n19, n18, n17, n16, n15, n14, n13, n12, n11, n10, 
        n9}) );
  INVX1 U17 ( .A(n182), .Y(n180) );
  INVX1 U19 ( .A(n180), .Y(n181) );
  BUFX2 U21 ( .A(n151), .Y(n182) );
  INVX1 U26 ( .A(n185), .Y(n183) );
  INVX1 U29 ( .A(n183), .Y(n184) );
  BUFX2 U30 ( .A(n71), .Y(n185) );
  INVX1 U33 ( .A(n188), .Y(n186) );
  INVX1 U38 ( .A(n186), .Y(n187) );
  BUFX2 U39 ( .A(n67), .Y(n188) );
  INVX1 U41 ( .A(n191), .Y(n189) );
  INVX1 U43 ( .A(n189), .Y(n190) );
  BUFX2 U44 ( .A(n56), .Y(n191) );
  INVX1 U47 ( .A(n194), .Y(n192) );
  INVX1 U52 ( .A(n192), .Y(n193) );
  BUFX2 U53 ( .A(n48), .Y(n194) );
  INVX1 U56 ( .A(n197), .Y(n195) );
  INVX1 U58 ( .A(n195), .Y(n196) );
  BUFX2 U59 ( .A(n2), .Y(n197) );
  INVX1 U60 ( .A(n200), .Y(n198) );
  INVX1 U61 ( .A(n198), .Y(n199) );
  BUFX2 U62 ( .A(n123), .Y(n200) );
  INVX1 U66 ( .A(n203), .Y(n201) );
  INVX1 U69 ( .A(n201), .Y(n202) );
  BUFX2 U71 ( .A(n143), .Y(n203) );
  INVX1 U74 ( .A(n206), .Y(n204) );
  INVX1 U76 ( .A(n204), .Y(n205) );
  BUFX2 U79 ( .A(n31), .Y(n206) );
  INVX1 U81 ( .A(n209), .Y(n207) );
  INVX1 U84 ( .A(n207), .Y(n208) );
  BUFX2 U86 ( .A(n131), .Y(n209) );
  INVX1 U88 ( .A(n212), .Y(n210) );
  INVX1 U90 ( .A(n210), .Y(n211) );
  BUFX2 U92 ( .A(n122), .Y(n212) );
  INVX1 U94 ( .A(n215), .Y(n213) );
  INVX1 U96 ( .A(n213), .Y(n214) );
  BUFX2 U98 ( .A(n129), .Y(n215) );
  INVX1 U100 ( .A(n218), .Y(n216) );
  INVX1 U102 ( .A(n216), .Y(n217) );
  AND2X1 U104 ( .A(n350), .B(n298), .Y(n159) );
  INVX1 U106 ( .A(n159), .Y(n218) );
  INVX1 U110 ( .A(n221), .Y(n219) );
  INVX1 U114 ( .A(n219), .Y(n220) );
  AND2X1 U135 ( .A(n350), .B(n301), .Y(n158) );
  INVX1 U137 ( .A(n158), .Y(n221) );
  INVX1 U162 ( .A(n224), .Y(n222) );
  INVX1 U163 ( .A(n222), .Y(n223) );
  AND2X2 U166 ( .A(n307), .B(n184), .Y(n157) );
  INVX1 U179 ( .A(n157), .Y(n224) );
  INVX1 U181 ( .A(n227), .Y(n225) );
  INVX1 U182 ( .A(n225), .Y(n226) );
  AND2X1 U183 ( .A(n356), .B(n304), .Y(n152) );
  INVX1 U184 ( .A(n152), .Y(n227) );
  INVX1 U185 ( .A(n230), .Y(n228) );
  INVX1 U186 ( .A(n228), .Y(n229) );
  AND2X2 U187 ( .A(n310), .B(n196), .Y(n149) );
  INVX1 U188 ( .A(n149), .Y(n230) );
  INVX1 U189 ( .A(n233), .Y(n231) );
  INVX1 U190 ( .A(n231), .Y(n232) );
  AND2X1 U191 ( .A(n27), .B(n80), .Y(n116) );
  INVX1 U192 ( .A(n116), .Y(n233) );
  INVX1 U193 ( .A(n236), .Y(n234) );
  INVX1 U194 ( .A(n234), .Y(n235) );
  AND2X1 U195 ( .A(n9), .B(n80), .Y(n114) );
  INVX1 U196 ( .A(n114), .Y(n236) );
  INVX1 U197 ( .A(n239), .Y(n237) );
  INVX1 U198 ( .A(n237), .Y(n238) );
  AND2X1 U199 ( .A(n10), .B(n80), .Y(n112) );
  INVX1 U200 ( .A(n112), .Y(n239) );
  INVX1 U201 ( .A(n242), .Y(n240) );
  INVX1 U202 ( .A(n240), .Y(n241) );
  AND2X1 U203 ( .A(n11), .B(n80), .Y(n110) );
  INVX1 U204 ( .A(n110), .Y(n242) );
  INVX1 U205 ( .A(n245), .Y(n243) );
  INVX1 U206 ( .A(n243), .Y(n244) );
  AND2X1 U207 ( .A(n12), .B(n80), .Y(n108) );
  INVX1 U208 ( .A(n108), .Y(n245) );
  INVX1 U209 ( .A(n248), .Y(n246) );
  INVX1 U210 ( .A(n246), .Y(n247) );
  AND2X1 U211 ( .A(n13), .B(n80), .Y(n106) );
  INVX1 U212 ( .A(n106), .Y(n248) );
  INVX1 U213 ( .A(n251), .Y(n249) );
  INVX1 U214 ( .A(n249), .Y(n250) );
  AND2X1 U215 ( .A(n14), .B(n80), .Y(n104) );
  INVX1 U216 ( .A(n104), .Y(n251) );
  INVX1 U217 ( .A(n254), .Y(n252) );
  INVX1 U218 ( .A(n252), .Y(n253) );
  AND2X1 U219 ( .A(n15), .B(n80), .Y(n102) );
  INVX1 U220 ( .A(n102), .Y(n254) );
  INVX1 U221 ( .A(n257), .Y(n255) );
  INVX1 U222 ( .A(n255), .Y(n256) );
  AND2X1 U223 ( .A(n16), .B(n80), .Y(n100) );
  INVX1 U224 ( .A(n100), .Y(n257) );
  INVX1 U225 ( .A(n260), .Y(n258) );
  INVX1 U226 ( .A(n258), .Y(n259) );
  AND2X1 U227 ( .A(n17), .B(n80), .Y(n98) );
  INVX1 U228 ( .A(n98), .Y(n260) );
  INVX1 U229 ( .A(n263), .Y(n261) );
  INVX1 U230 ( .A(n261), .Y(n262) );
  AND2X1 U231 ( .A(n18), .B(n80), .Y(n96) );
  INVX1 U232 ( .A(n96), .Y(n263) );
  INVX1 U233 ( .A(n266), .Y(n264) );
  INVX1 U234 ( .A(n264), .Y(n265) );
  AND2X1 U235 ( .A(n19), .B(n80), .Y(n94) );
  INVX1 U236 ( .A(n94), .Y(n266) );
  INVX1 U237 ( .A(n269), .Y(n267) );
  INVX1 U238 ( .A(n267), .Y(n268) );
  AND2X1 U239 ( .A(n20), .B(n80), .Y(n92) );
  INVX1 U240 ( .A(n92), .Y(n269) );
  INVX1 U241 ( .A(n272), .Y(n270) );
  INVX1 U242 ( .A(n270), .Y(n271) );
  AND2X1 U243 ( .A(n21), .B(n80), .Y(n90) );
  INVX1 U244 ( .A(n90), .Y(n272) );
  INVX1 U245 ( .A(n275), .Y(n273) );
  INVX1 U246 ( .A(n273), .Y(n274) );
  AND2X1 U247 ( .A(n22), .B(n80), .Y(n88) );
  INVX1 U248 ( .A(n88), .Y(n275) );
  INVX1 U249 ( .A(n278), .Y(n276) );
  INVX1 U250 ( .A(n276), .Y(n277) );
  AND2X1 U251 ( .A(n23), .B(n80), .Y(n86) );
  INVX1 U252 ( .A(n86), .Y(n278) );
  INVX1 U253 ( .A(n281), .Y(n279) );
  INVX1 U254 ( .A(n279), .Y(n280) );
  AND2X1 U255 ( .A(n24), .B(n80), .Y(n84) );
  INVX1 U256 ( .A(n84), .Y(n281) );
  INVX1 U257 ( .A(n284), .Y(n282) );
  INVX1 U258 ( .A(n282), .Y(n283) );
  AND2X1 U259 ( .A(n25), .B(n80), .Y(n82) );
  INVX1 U260 ( .A(n82), .Y(n284) );
  INVX1 U261 ( .A(n287), .Y(n285) );
  INVX1 U262 ( .A(n285), .Y(n286) );
  AND2X1 U263 ( .A(n26), .B(n80), .Y(n79) );
  INVX1 U264 ( .A(n79), .Y(n287) );
  AND2X2 U265 ( .A(ready), .B(n65), .Y(n66) );
  INVX1 U266 ( .A(n66), .Y(n288) );
  AND2X2 U267 ( .A(n47), .B(n187), .Y(n65) );
  AND2X1 U268 ( .A(reset_out), .B(n54), .Y(n55) );
  INVX1 U269 ( .A(n55), .Y(n289) );
  AND2X2 U270 ( .A(n47), .B(n190), .Y(n54) );
  AND2X1 U271 ( .A(cke), .B(n45), .Y(n46) );
  INVX1 U272 ( .A(n46), .Y(n290) );
  AND2X2 U273 ( .A(n47), .B(n193), .Y(n45) );
  INVX1 U274 ( .A(n293), .Y(n291) );
  INVX1 U275 ( .A(n291), .Y(n292) );
  AND2X1 U276 ( .A(a[10]), .B(n344), .Y(n40) );
  INVX1 U277 ( .A(n40), .Y(n293) );
  INVX1 U278 ( .A(n296), .Y(n294) );
  INVX1 U279 ( .A(n294), .Y(n295) );
  AND2X1 U280 ( .A(ba[1]), .B(n5), .Y(n8) );
  INVX1 U281 ( .A(n8), .Y(n296) );
  INVX1 U282 ( .A(n299), .Y(n297) );
  INVX1 U283 ( .A(n297), .Y(n298) );
  AND2X1 U284 ( .A(casbar), .B(n73), .Y(n76) );
  INVX1 U285 ( .A(n76), .Y(n299) );
  INVX1 U286 ( .A(n302), .Y(n300) );
  INVX1 U287 ( .A(n300), .Y(n301) );
  AND2X1 U288 ( .A(rasbar), .B(n73), .Y(n75) );
  INVX1 U289 ( .A(n75), .Y(n302) );
  INVX1 U290 ( .A(n305), .Y(n303) );
  INVX1 U291 ( .A(n303), .Y(n304) );
  AND2X1 U292 ( .A(a[8]), .B(n389), .Y(n37) );
  INVX1 U293 ( .A(n37), .Y(n305) );
  INVX1 U294 ( .A(n308), .Y(n306) );
  INVX1 U295 ( .A(n306), .Y(n307) );
  AND2X1 U296 ( .A(webar), .B(n73), .Y(n70) );
  INVX1 U297 ( .A(n70), .Y(n308) );
  INVX1 U298 ( .A(n311), .Y(n309) );
  INVX1 U299 ( .A(n309), .Y(n310) );
  AND2X1 U300 ( .A(ba[0]), .B(n5), .Y(n1) );
  INVX1 U301 ( .A(n1), .Y(n311) );
  INVX1 U302 ( .A(n314), .Y(n312) );
  INVX1 U303 ( .A(n312), .Y(n313) );
  OR2X1 U304 ( .A(n392), .B(n353), .Y(n51) );
  INVX1 U305 ( .A(n51), .Y(n314) );
  INVX1 U306 ( .A(n317), .Y(n315) );
  INVX1 U307 ( .A(n315), .Y(n316) );
  AND2X1 U308 ( .A(a[4]), .B(n389), .Y(n33) );
  INVX1 U309 ( .A(n33), .Y(n317) );
  INVX1 U310 ( .A(n320), .Y(n318) );
  INVX1 U311 ( .A(n318), .Y(n319) );
  BUFX2 U312 ( .A(n138), .Y(n320) );
  INVX1 U313 ( .A(n323), .Y(n321) );
  INVX1 U314 ( .A(n321), .Y(n322) );
  BUFX2 U315 ( .A(n126), .Y(n323) );
  INVX1 U316 ( .A(n328), .Y(n324) );
  INVX1 U317 ( .A(n324), .Y(n325) );
  BUFX2 U318 ( .A(n60), .Y(n328) );
  INVX1 U319 ( .A(n331), .Y(n329) );
  INVX1 U320 ( .A(n329), .Y(n330) );
  AND2X1 U321 ( .A(n347), .B(n380), .Y(n120) );
  INVX1 U322 ( .A(n120), .Y(n331) );
  INVX1 U323 ( .A(n336), .Y(n333) );
  INVX1 U324 ( .A(n333), .Y(n334) );
  AND2X1 U325 ( .A(counter[12]), .B(n63), .Y(n139) );
  INVX1 U326 ( .A(n139), .Y(n336) );
  INVX1 U327 ( .A(n339), .Y(n337) );
  INVX1 U328 ( .A(n337), .Y(n338) );
  BUFX2 U329 ( .A(n146), .Y(n339) );
  INVX1 U330 ( .A(n342), .Y(n340) );
  INVX1 U331 ( .A(n340), .Y(n341) );
  AND2X1 U332 ( .A(n62), .B(counter[6]), .Y(n61) );
  INVX1 U333 ( .A(n61), .Y(n342) );
  INVX1 U334 ( .A(n345), .Y(n343) );
  INVX1 U335 ( .A(n343), .Y(n344) );
  BUFX2 U336 ( .A(n41), .Y(n345) );
  INVX1 U337 ( .A(n348), .Y(n346) );
  INVX1 U338 ( .A(n346), .Y(n347) );
  BUFX2 U339 ( .A(n141), .Y(n348) );
  INVX1 U340 ( .A(n351), .Y(n349) );
  INVX1 U341 ( .A(n349), .Y(n350) );
  BUFX2 U342 ( .A(n74), .Y(n351) );
  INVX1 U343 ( .A(n354), .Y(n352) );
  INVX1 U344 ( .A(n352), .Y(n353) );
  BUFX2 U345 ( .A(n53), .Y(n354) );
  INVX1 U346 ( .A(n357), .Y(n355) );
  INVX1 U347 ( .A(n355), .Y(n356) );
  BUFX2 U348 ( .A(n32), .Y(n357) );
  INVX1 U349 ( .A(n360), .Y(n358) );
  INVX1 U350 ( .A(n358), .Y(n359) );
  AND2X1 U351 ( .A(INIT), .B(n118), .Y(n117) );
  INVX1 U352 ( .A(n117), .Y(n360) );
  INVX1 U353 ( .A(n363), .Y(n361) );
  INVX1 U354 ( .A(n361), .Y(n362) );
  AND2X1 U355 ( .A(counter[9]), .B(n134), .Y(n145) );
  INVX1 U356 ( .A(n145), .Y(n363) );
  INVX1 U357 ( .A(n366), .Y(n364) );
  INVX1 U358 ( .A(n364), .Y(n365) );
  AND2X1 U359 ( .A(n374), .B(n383), .Y(n3) );
  INVX1 U360 ( .A(n3), .Y(n366) );
  INVX1 U361 ( .A(n369), .Y(n367) );
  INVX1 U362 ( .A(n367), .Y(n368) );
  BUFX2 U363 ( .A(n140), .Y(n369) );
  INVX1 U364 ( .A(n372), .Y(n370) );
  INVX1 U365 ( .A(n370), .Y(n371) );
  AND2X1 U366 ( .A(counter[11]), .B(n89), .Y(n64) );
  INVX1 U367 ( .A(n64), .Y(n372) );
  INVX1 U368 ( .A(n375), .Y(n373) );
  INVX1 U369 ( .A(n373), .Y(n374) );
  BUFX2 U370 ( .A(n36), .Y(n375) );
  INVX1 U371 ( .A(n378), .Y(n376) );
  INVX1 U372 ( .A(n376), .Y(n377) );
  OR2X2 U373 ( .A(n362), .B(counter[3]), .Y(n50) );
  INVX1 U374 ( .A(n50), .Y(n378) );
  INVX1 U375 ( .A(n381), .Y(n379) );
  INVX1 U376 ( .A(n379), .Y(n380) );
  BUFX2 U377 ( .A(n30), .Y(n381) );
  INVX1 U378 ( .A(n384), .Y(n382) );
  INVX1 U379 ( .A(n382), .Y(n383) );
  BUFX2 U380 ( .A(n29), .Y(n384) );
  INVX1 U381 ( .A(n387), .Y(n385) );
  INVX1 U382 ( .A(n385), .Y(n386) );
  BUFX2 U383 ( .A(n127), .Y(n387) );
  INVX1 U384 ( .A(n390), .Y(n388) );
  INVX1 U385 ( .A(n388), .Y(n389) );
  BUFX2 U386 ( .A(n34), .Y(n390) );
  INVX1 U387 ( .A(n393), .Y(n391) );
  INVX1 U388 ( .A(n391), .Y(n392) );
  BUFX2 U389 ( .A(n52), .Y(n393) );
  INVX1 U390 ( .A(n396), .Y(n394) );
  INVX1 U391 ( .A(n394), .Y(n395) );
  AND2X1 U392 ( .A(flag), .B(n47), .Y(n6) );
  INVX1 U393 ( .A(n6), .Y(n396) );
endmodule


module ddr3_ring_buffer8 ( dout, listen, strobe, readPtr, din, reset );
  output [15:0] dout;
  input [2:0] readPtr;
  input [15:0] din;
  input listen, strobe, reset;
  wire   dStrobe0, dStrobe1, dStrobe2, dStrobe3, dStrobe, count_0_, F0,
         fStrobe, n43, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n125, n142, n241, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745;
  wire   [15:0] r0;
  wire   [15:0] r2;
  wire   [15:0] r4;
  wire   [15:0] r6;
  wire   [15:0] r1;
  wire   [15:0] r3;
  wire   [15:0] r5;
  wire   [15:0] r7;

  CLKBUF2 DELAY0 ( .A(strobe), .Y(dStrobe0) );
  CLKBUF2 DELAY1 ( .A(dStrobe0), .Y(dStrobe1) );
  CLKBUF2 DELAY2 ( .A(dStrobe1), .Y(dStrobe2) );
  CLKBUF2 DELAY3 ( .A(dStrobe2), .Y(dStrobe3) );
  CLKBUF2 DELAY4 ( .A(dStrobe3), .Y(dStrobe) );
  DFFSR F0_reg ( .D(n732), .CLK(n43), .R(n242), .S(n91), .Q(F0) );
  DFFSR count_reg_0_ ( .D(n465), .CLK(n43), .R(n242), .S(1'b1), .Q(count_0_)
         );
  DFFPOSX1 r2_reg_15_ ( .D(n464), .CLK(n734), .Q(r2[15]) );
  DFFPOSX1 r2_reg_14_ ( .D(n463), .CLK(n734), .Q(r2[14]) );
  DFFPOSX1 r2_reg_13_ ( .D(n462), .CLK(n734), .Q(r2[13]) );
  DFFPOSX1 r2_reg_12_ ( .D(n461), .CLK(n734), .Q(r2[12]) );
  DFFPOSX1 r2_reg_11_ ( .D(n460), .CLK(n734), .Q(r2[11]) );
  DFFPOSX1 r2_reg_10_ ( .D(n459), .CLK(n734), .Q(r2[10]) );
  DFFPOSX1 r2_reg_9_ ( .D(n458), .CLK(n735), .Q(r2[9]) );
  DFFPOSX1 r2_reg_8_ ( .D(n457), .CLK(n735), .Q(r2[8]) );
  DFFPOSX1 r2_reg_7_ ( .D(n456), .CLK(n734), .Q(r2[7]) );
  DFFPOSX1 r2_reg_6_ ( .D(n455), .CLK(n736), .Q(r2[6]) );
  DFFPOSX1 r2_reg_5_ ( .D(n454), .CLK(n736), .Q(r2[5]) );
  DFFPOSX1 r2_reg_4_ ( .D(n453), .CLK(n735), .Q(r2[4]) );
  DFFPOSX1 r2_reg_3_ ( .D(n452), .CLK(n736), .Q(r2[3]) );
  DFFPOSX1 r2_reg_2_ ( .D(n451), .CLK(n736), .Q(r2[2]) );
  DFFPOSX1 r2_reg_1_ ( .D(n450), .CLK(n735), .Q(r2[1]) );
  DFFPOSX1 r2_reg_0_ ( .D(n449), .CLK(n737), .Q(r2[0]) );
  DFFPOSX1 r4_reg_15_ ( .D(n448), .CLK(n737), .Q(r4[15]) );
  DFFPOSX1 r4_reg_14_ ( .D(n447), .CLK(n735), .Q(r4[14]) );
  DFFPOSX1 r4_reg_13_ ( .D(n446), .CLK(n737), .Q(r4[13]) );
  DFFPOSX1 r4_reg_12_ ( .D(n445), .CLK(n737), .Q(r4[12]) );
  DFFPOSX1 r4_reg_11_ ( .D(n444), .CLK(n736), .Q(r4[11]) );
  DFFPOSX1 r4_reg_10_ ( .D(n443), .CLK(n737), .Q(r4[10]) );
  DFFPOSX1 r4_reg_9_ ( .D(n442), .CLK(n737), .Q(r4[9]) );
  DFFPOSX1 r4_reg_8_ ( .D(n441), .CLK(n736), .Q(r4[8]) );
  DFFPOSX1 r4_reg_7_ ( .D(n440), .CLK(n737), .Q(r4[7]) );
  DFFPOSX1 r4_reg_6_ ( .D(n439), .CLK(n737), .Q(r4[6]) );
  DFFPOSX1 r4_reg_5_ ( .D(n438), .CLK(n736), .Q(r4[5]) );
  DFFPOSX1 r4_reg_4_ ( .D(n437), .CLK(n737), .Q(r4[4]) );
  DFFPOSX1 r4_reg_3_ ( .D(n436), .CLK(n735), .Q(r4[3]) );
  DFFPOSX1 r4_reg_2_ ( .D(n435), .CLK(n736), .Q(r4[2]) );
  DFFPOSX1 r4_reg_1_ ( .D(n434), .CLK(n738), .Q(r4[1]) );
  DFFPOSX1 r4_reg_0_ ( .D(n433), .CLK(n738), .Q(r4[0]) );
  DFFPOSX1 r6_reg_15_ ( .D(n432), .CLK(n736), .Q(r6[15]) );
  DFFPOSX1 r6_reg_14_ ( .D(n431), .CLK(n738), .Q(r6[14]) );
  DFFPOSX1 r6_reg_13_ ( .D(n430), .CLK(n738), .Q(r6[13]) );
  DFFPOSX1 r6_reg_12_ ( .D(n429), .CLK(n736), .Q(r6[12]) );
  DFFPOSX1 r6_reg_11_ ( .D(n428), .CLK(n738), .Q(r6[11]) );
  DFFPOSX1 r6_reg_10_ ( .D(n427), .CLK(n738), .Q(r6[10]) );
  DFFPOSX1 r6_reg_9_ ( .D(n426), .CLK(n737), .Q(r6[9]) );
  DFFPOSX1 r6_reg_8_ ( .D(n425), .CLK(n738), .Q(r6[8]) );
  DFFPOSX1 r6_reg_7_ ( .D(n424), .CLK(n738), .Q(r6[7]) );
  DFFPOSX1 r6_reg_6_ ( .D(n423), .CLK(n737), .Q(r6[6]) );
  DFFPOSX1 r6_reg_5_ ( .D(n422), .CLK(n738), .Q(r6[5]) );
  DFFPOSX1 r6_reg_4_ ( .D(n421), .CLK(n738), .Q(r6[4]) );
  DFFPOSX1 r6_reg_3_ ( .D(n420), .CLK(n737), .Q(r6[3]) );
  DFFPOSX1 r6_reg_2_ ( .D(n419), .CLK(n738), .Q(r6[2]) );
  DFFPOSX1 r6_reg_1_ ( .D(n418), .CLK(n738), .Q(r6[1]) );
  DFFPOSX1 r6_reg_0_ ( .D(n417), .CLK(n734), .Q(r6[0]) );
  DFFPOSX1 r0_reg_15_ ( .D(n416), .CLK(n734), .Q(r0[15]) );
  DFFPOSX1 r0_reg_14_ ( .D(n415), .CLK(n734), .Q(r0[14]) );
  DFFPOSX1 r0_reg_13_ ( .D(n414), .CLK(n734), .Q(r0[13]) );
  DFFPOSX1 r0_reg_12_ ( .D(n413), .CLK(n734), .Q(r0[12]) );
  DFFPOSX1 r0_reg_11_ ( .D(n412), .CLK(n735), .Q(r0[11]) );
  DFFPOSX1 r0_reg_10_ ( .D(n411), .CLK(n735), .Q(r0[10]) );
  DFFPOSX1 r0_reg_9_ ( .D(n410), .CLK(n734), .Q(r0[9]) );
  DFFPOSX1 r0_reg_8_ ( .D(n409), .CLK(n735), .Q(r0[8]) );
  DFFPOSX1 r0_reg_7_ ( .D(n408), .CLK(n735), .Q(r0[7]) );
  DFFPOSX1 r0_reg_6_ ( .D(n407), .CLK(n735), .Q(r0[6]) );
  DFFPOSX1 r0_reg_5_ ( .D(n406), .CLK(n736), .Q(r0[5]) );
  DFFPOSX1 r0_reg_4_ ( .D(n405), .CLK(n736), .Q(r0[4]) );
  DFFPOSX1 r0_reg_3_ ( .D(n404), .CLK(n735), .Q(r0[3]) );
  DFFPOSX1 r0_reg_2_ ( .D(n403), .CLK(n736), .Q(r0[2]) );
  DFFPOSX1 r0_reg_1_ ( .D(n402), .CLK(n737), .Q(r0[1]) );
  DFFPOSX1 r0_reg_0_ ( .D(n401), .CLK(n735), .Q(r0[0]) );
  DFFNEGX1 r3_reg_15_ ( .D(n400), .CLK(n742), .Q(r3[15]) );
  DFFNEGX1 r3_reg_14_ ( .D(n399), .CLK(n742), .Q(r3[14]) );
  DFFNEGX1 r3_reg_13_ ( .D(n398), .CLK(n742), .Q(r3[13]) );
  DFFNEGX1 r3_reg_12_ ( .D(n397), .CLK(n742), .Q(r3[12]) );
  DFFNEGX1 r3_reg_11_ ( .D(n396), .CLK(n742), .Q(r3[11]) );
  DFFNEGX1 r3_reg_10_ ( .D(n395), .CLK(n742), .Q(r3[10]) );
  DFFNEGX1 r3_reg_9_ ( .D(n394), .CLK(n742), .Q(r3[9]) );
  DFFNEGX1 r3_reg_8_ ( .D(n393), .CLK(n742), .Q(r3[8]) );
  DFFNEGX1 r3_reg_7_ ( .D(n392), .CLK(n741), .Q(r3[7]) );
  DFFNEGX1 r3_reg_6_ ( .D(n391), .CLK(n741), .Q(r3[6]) );
  DFFNEGX1 r3_reg_5_ ( .D(n390), .CLK(n741), .Q(r3[5]) );
  DFFNEGX1 r3_reg_4_ ( .D(n389), .CLK(n741), .Q(r3[4]) );
  DFFNEGX1 r3_reg_3_ ( .D(n388), .CLK(n741), .Q(r3[3]) );
  DFFNEGX1 r3_reg_2_ ( .D(n387), .CLK(n741), .Q(r3[2]) );
  DFFNEGX1 r3_reg_1_ ( .D(n386), .CLK(n741), .Q(r3[1]) );
  DFFNEGX1 r3_reg_0_ ( .D(n385), .CLK(n741), .Q(r3[0]) );
  DFFNEGX1 r5_reg_15_ ( .D(n384), .CLK(n740), .Q(r5[15]) );
  DFFNEGX1 r5_reg_14_ ( .D(n383), .CLK(n740), .Q(r5[14]) );
  DFFNEGX1 r5_reg_13_ ( .D(n382), .CLK(n740), .Q(r5[13]) );
  DFFNEGX1 r5_reg_12_ ( .D(n381), .CLK(n740), .Q(r5[12]) );
  DFFNEGX1 r5_reg_11_ ( .D(n380), .CLK(n740), .Q(r5[11]) );
  DFFNEGX1 r5_reg_10_ ( .D(n379), .CLK(n740), .Q(r5[10]) );
  DFFNEGX1 r5_reg_9_ ( .D(n378), .CLK(n739), .Q(r5[9]) );
  DFFNEGX1 r5_reg_8_ ( .D(n377), .CLK(n739), .Q(r5[8]) );
  DFFNEGX1 r5_reg_7_ ( .D(n376), .CLK(n739), .Q(r5[7]) );
  DFFNEGX1 r5_reg_6_ ( .D(n375), .CLK(n740), .Q(r5[6]) );
  DFFNEGX1 r5_reg_5_ ( .D(n374), .CLK(n740), .Q(r5[5]) );
  DFFNEGX1 r5_reg_4_ ( .D(n373), .CLK(n739), .Q(r5[4]) );
  DFFNEGX1 r5_reg_3_ ( .D(n372), .CLK(n739), .Q(r5[3]) );
  DFFNEGX1 r5_reg_2_ ( .D(n371), .CLK(n739), .Q(r5[2]) );
  DFFNEGX1 r5_reg_1_ ( .D(n370), .CLK(n739), .Q(r5[1]) );
  DFFNEGX1 r5_reg_0_ ( .D(n369), .CLK(n740), .Q(r5[0]) );
  DFFNEGX1 r7_reg_15_ ( .D(n368), .CLK(n740), .Q(r7[15]) );
  DFFNEGX1 r7_reg_14_ ( .D(n367), .CLK(n739), .Q(r7[14]) );
  DFFNEGX1 r7_reg_13_ ( .D(n366), .CLK(n739), .Q(r7[13]) );
  DFFNEGX1 r7_reg_12_ ( .D(n365), .CLK(n739), .Q(r7[12]) );
  DFFNEGX1 r7_reg_11_ ( .D(n364), .CLK(n739), .Q(r7[11]) );
  DFFNEGX1 r7_reg_10_ ( .D(n363), .CLK(n740), .Q(r7[10]) );
  DFFNEGX1 r7_reg_9_ ( .D(n362), .CLK(n740), .Q(r7[9]) );
  DFFNEGX1 r7_reg_8_ ( .D(n361), .CLK(n739), .Q(r7[8]) );
  DFFNEGX1 r7_reg_7_ ( .D(n360), .CLK(n739), .Q(r7[7]) );
  DFFNEGX1 r7_reg_6_ ( .D(n359), .CLK(n739), .Q(r7[6]) );
  DFFNEGX1 r7_reg_5_ ( .D(n358), .CLK(n739), .Q(r7[5]) );
  DFFNEGX1 r7_reg_4_ ( .D(n357), .CLK(n740), .Q(r7[4]) );
  DFFNEGX1 r7_reg_3_ ( .D(n356), .CLK(n740), .Q(r7[3]) );
  DFFNEGX1 r7_reg_2_ ( .D(n355), .CLK(n739), .Q(r7[2]) );
  DFFNEGX1 r7_reg_1_ ( .D(n354), .CLK(n738), .Q(r7[1]) );
  DFFNEGX1 r7_reg_0_ ( .D(n353), .CLK(n740), .Q(r7[0]) );
  DFFNEGX1 r1_reg_15_ ( .D(n352), .CLK(n740), .Q(r1[15]) );
  DFFNEGX1 r1_reg_14_ ( .D(n351), .CLK(n742), .Q(r1[14]) );
  DFFNEGX1 r1_reg_13_ ( .D(n350), .CLK(n742), .Q(r1[13]) );
  DFFNEGX1 r1_reg_12_ ( .D(n349), .CLK(n742), .Q(r1[12]) );
  DFFNEGX1 r1_reg_11_ ( .D(n348), .CLK(n742), .Q(r1[11]) );
  DFFNEGX1 r1_reg_10_ ( .D(n347), .CLK(n742), .Q(r1[10]) );
  DFFNEGX1 r1_reg_9_ ( .D(n346), .CLK(n742), .Q(r1[9]) );
  DFFNEGX1 r1_reg_8_ ( .D(n345), .CLK(n742), .Q(r1[8]) );
  DFFNEGX1 r1_reg_7_ ( .D(n344), .CLK(n741), .Q(r1[7]) );
  DFFNEGX1 r1_reg_6_ ( .D(n343), .CLK(n741), .Q(r1[6]) );
  DFFNEGX1 r1_reg_5_ ( .D(n342), .CLK(n741), .Q(r1[5]) );
  DFFNEGX1 r1_reg_4_ ( .D(n341), .CLK(n741), .Q(r1[4]) );
  DFFNEGX1 r1_reg_3_ ( .D(n340), .CLK(n741), .Q(r1[3]) );
  DFFNEGX1 r1_reg_2_ ( .D(n339), .CLK(n741), .Q(r1[2]) );
  DFFNEGX1 r1_reg_1_ ( .D(n338), .CLK(n741), .Q(r1[1]) );
  DFFNEGX1 r1_reg_0_ ( .D(n337), .CLK(n741), .Q(r1[0]) );
  INVX1 U8 ( .A(listen), .Y(n91) );
  OAI21X1 U9 ( .A(n92), .B(n93), .C(n662), .Y(n337) );
  OAI21X1 U11 ( .A(n92), .B(n95), .C(n659), .Y(n338) );
  OAI21X1 U13 ( .A(n92), .B(n97), .C(n656), .Y(n339) );
  OAI21X1 U15 ( .A(n92), .B(n99), .C(n653), .Y(n340) );
  OAI21X1 U17 ( .A(n92), .B(n101), .C(n650), .Y(n341) );
  OAI21X1 U19 ( .A(n92), .B(n103), .C(n647), .Y(n342) );
  OAI21X1 U21 ( .A(n92), .B(n105), .C(n644), .Y(n343) );
  OAI21X1 U23 ( .A(n92), .B(n107), .C(n641), .Y(n344) );
  OAI21X1 U25 ( .A(n92), .B(n109), .C(n638), .Y(n345) );
  OAI21X1 U27 ( .A(n92), .B(n111), .C(n635), .Y(n346) );
  OAI21X1 U29 ( .A(n92), .B(n113), .C(n632), .Y(n347) );
  OAI21X1 U31 ( .A(n92), .B(n115), .C(n629), .Y(n348) );
  OAI21X1 U33 ( .A(n92), .B(n117), .C(n626), .Y(n349) );
  OAI21X1 U35 ( .A(n92), .B(n119), .C(n623), .Y(n350) );
  OAI21X1 U37 ( .A(n92), .B(n121), .C(n620), .Y(n351) );
  OAI21X1 U39 ( .A(n92), .B(n123), .C(n617), .Y(n352) );
  OAI21X1 U105 ( .A(n93), .B(n159), .C(n614), .Y(n385) );
  OAI21X1 U107 ( .A(n95), .B(n159), .C(n611), .Y(n386) );
  OAI21X1 U109 ( .A(n97), .B(n159), .C(n608), .Y(n387) );
  OAI21X1 U111 ( .A(n99), .B(n159), .C(n605), .Y(n388) );
  OAI21X1 U113 ( .A(n101), .B(n159), .C(n602), .Y(n389) );
  OAI21X1 U115 ( .A(n103), .B(n159), .C(n599), .Y(n390) );
  OAI21X1 U117 ( .A(n105), .B(n159), .C(n596), .Y(n391) );
  OAI21X1 U119 ( .A(n107), .B(n159), .C(n593), .Y(n392) );
  OAI21X1 U121 ( .A(n109), .B(n159), .C(n590), .Y(n393) );
  OAI21X1 U123 ( .A(n111), .B(n159), .C(n587), .Y(n394) );
  OAI21X1 U125 ( .A(n113), .B(n159), .C(n584), .Y(n395) );
  OAI21X1 U127 ( .A(n115), .B(n159), .C(n581), .Y(n396) );
  OAI21X1 U129 ( .A(n117), .B(n159), .C(n578), .Y(n397) );
  OAI21X1 U131 ( .A(n119), .B(n159), .C(n575), .Y(n398) );
  OAI21X1 U133 ( .A(n121), .B(n159), .C(n572), .Y(n399) );
  OAI21X1 U135 ( .A(n123), .B(n159), .C(n569), .Y(n400) );
  OAI21X1 U137 ( .A(n92), .B(n93), .C(n566), .Y(n401) );
  OAI21X1 U139 ( .A(n92), .B(n95), .C(n563), .Y(n402) );
  OAI21X1 U141 ( .A(n92), .B(n97), .C(n560), .Y(n403) );
  OAI21X1 U143 ( .A(n92), .B(n99), .C(n557), .Y(n404) );
  OAI21X1 U145 ( .A(n92), .B(n101), .C(n554), .Y(n405) );
  OAI21X1 U147 ( .A(n92), .B(n103), .C(n551), .Y(n406) );
  OAI21X1 U149 ( .A(n92), .B(n105), .C(n548), .Y(n407) );
  OAI21X1 U151 ( .A(n92), .B(n107), .C(n545), .Y(n408) );
  OAI21X1 U153 ( .A(n92), .B(n109), .C(n542), .Y(n409) );
  OAI21X1 U155 ( .A(n92), .B(n111), .C(n539), .Y(n410) );
  OAI21X1 U157 ( .A(n92), .B(n113), .C(n536), .Y(n411) );
  OAI21X1 U159 ( .A(n92), .B(n115), .C(n533), .Y(n412) );
  OAI21X1 U161 ( .A(n92), .B(n117), .C(n530), .Y(n413) );
  OAI21X1 U163 ( .A(n92), .B(n119), .C(n527), .Y(n414) );
  OAI21X1 U165 ( .A(n92), .B(n121), .C(n524), .Y(n415) );
  OAI21X1 U167 ( .A(n92), .B(n123), .C(n521), .Y(n416) );
  OAI21X1 U233 ( .A(n93), .B(n159), .C(n518), .Y(n449) );
  INVX1 U235 ( .A(din[0]), .Y(n93) );
  OAI21X1 U236 ( .A(n95), .B(n159), .C(n515), .Y(n450) );
  INVX1 U238 ( .A(din[1]), .Y(n95) );
  OAI21X1 U239 ( .A(n97), .B(n159), .C(n512), .Y(n451) );
  INVX1 U241 ( .A(din[2]), .Y(n97) );
  OAI21X1 U242 ( .A(n99), .B(n159), .C(n509), .Y(n452) );
  INVX1 U244 ( .A(din[3]), .Y(n99) );
  OAI21X1 U245 ( .A(n101), .B(n159), .C(n506), .Y(n453) );
  INVX1 U247 ( .A(din[4]), .Y(n101) );
  OAI21X1 U248 ( .A(n103), .B(n159), .C(n503), .Y(n454) );
  INVX1 U250 ( .A(din[5]), .Y(n103) );
  OAI21X1 U251 ( .A(n105), .B(n159), .C(n500), .Y(n455) );
  INVX1 U253 ( .A(din[6]), .Y(n105) );
  OAI21X1 U254 ( .A(n107), .B(n159), .C(n497), .Y(n456) );
  INVX1 U256 ( .A(din[7]), .Y(n107) );
  OAI21X1 U257 ( .A(n109), .B(n159), .C(n494), .Y(n457) );
  INVX1 U259 ( .A(din[8]), .Y(n109) );
  OAI21X1 U260 ( .A(n111), .B(n159), .C(n491), .Y(n458) );
  INVX1 U262 ( .A(din[9]), .Y(n111) );
  OAI21X1 U263 ( .A(n113), .B(n159), .C(n488), .Y(n459) );
  INVX1 U265 ( .A(din[10]), .Y(n113) );
  OAI21X1 U266 ( .A(n115), .B(n159), .C(n485), .Y(n460) );
  INVX1 U268 ( .A(din[11]), .Y(n115) );
  OAI21X1 U269 ( .A(n117), .B(n159), .C(n482), .Y(n461) );
  INVX1 U271 ( .A(din[12]), .Y(n117) );
  OAI21X1 U272 ( .A(n119), .B(n159), .C(n479), .Y(n462) );
  INVX1 U274 ( .A(din[13]), .Y(n119) );
  OAI21X1 U275 ( .A(n121), .B(n159), .C(n476), .Y(n463) );
  INVX1 U277 ( .A(din[14]), .Y(n121) );
  OAI21X1 U278 ( .A(n123), .B(n159), .C(n473), .Y(n464) );
  INVX1 U281 ( .A(din[15]), .Y(n123) );
  OAI21X1 U282 ( .A(n466), .B(n92), .C(n224), .Y(n465) );
  INVX1 U284 ( .A(n729), .Y(n224) );
  AND2X1 U286 ( .A(n242), .B(listen), .Y(n466) );
  INVX1 U287 ( .A(reset), .Y(n242) );
  INVX1 U288 ( .A(n43), .Y(fStrobe) );
  OAI21X1 U289 ( .A(listen), .B(n732), .C(dStrobe), .Y(n43) );
  NAND3X1 U290 ( .A(n470), .B(n726), .C(n245), .Y(dout[9]) );
  AOI22X1 U292 ( .A(n248), .B(r7[9]), .C(n249), .D(r6[9]), .Y(n247) );
  AOI22X1 U293 ( .A(n250), .B(r5[9]), .C(n251), .D(r4[9]), .Y(n246) );
  AOI22X1 U294 ( .A(n252), .B(r3[9]), .C(n253), .D(r2[9]), .Y(n244) );
  AOI22X1 U295 ( .A(n254), .B(r1[9]), .C(n255), .D(r0[9]), .Y(n243) );
  NAND3X1 U296 ( .A(n467), .B(n723), .C(n258), .Y(dout[8]) );
  AOI22X1 U298 ( .A(n248), .B(r7[8]), .C(n249), .D(r6[8]), .Y(n260) );
  AOI22X1 U299 ( .A(n250), .B(r5[8]), .C(n251), .D(r4[8]), .Y(n259) );
  AOI22X1 U300 ( .A(n252), .B(r3[8]), .C(n253), .D(r2[8]), .Y(n257) );
  AOI22X1 U301 ( .A(n254), .B(r1[8]), .C(n255), .D(r0[8]), .Y(n256) );
  NAND3X1 U302 ( .A(n125), .B(n720), .C(n263), .Y(dout[7]) );
  AOI22X1 U304 ( .A(n248), .B(r7[7]), .C(n249), .D(r6[7]), .Y(n265) );
  AOI22X1 U305 ( .A(n250), .B(r5[7]), .C(n251), .D(r4[7]), .Y(n264) );
  AOI22X1 U306 ( .A(n252), .B(r3[7]), .C(n253), .D(r2[7]), .Y(n262) );
  AOI22X1 U307 ( .A(n254), .B(r1[7]), .C(n255), .D(r0[7]), .Y(n261) );
  NAND3X1 U308 ( .A(n87), .B(n717), .C(n268), .Y(dout[6]) );
  AOI22X1 U310 ( .A(n248), .B(r7[6]), .C(n249), .D(r6[6]), .Y(n270) );
  AOI22X1 U311 ( .A(n250), .B(r5[6]), .C(n251), .D(r4[6]), .Y(n269) );
  AOI22X1 U312 ( .A(n252), .B(r3[6]), .C(n253), .D(r2[6]), .Y(n267) );
  AOI22X1 U313 ( .A(n254), .B(r1[6]), .C(n255), .D(r0[6]), .Y(n266) );
  NAND3X1 U314 ( .A(n84), .B(n714), .C(n273), .Y(dout[5]) );
  AOI22X1 U316 ( .A(n248), .B(r7[5]), .C(n249), .D(r6[5]), .Y(n275) );
  AOI22X1 U317 ( .A(n250), .B(r5[5]), .C(n251), .D(r4[5]), .Y(n274) );
  AOI22X1 U318 ( .A(n252), .B(r3[5]), .C(n253), .D(r2[5]), .Y(n272) );
  AOI22X1 U319 ( .A(n254), .B(r1[5]), .C(n255), .D(r0[5]), .Y(n271) );
  NAND3X1 U320 ( .A(n81), .B(n711), .C(n278), .Y(dout[4]) );
  AOI22X1 U322 ( .A(n248), .B(r7[4]), .C(n249), .D(r6[4]), .Y(n280) );
  AOI22X1 U323 ( .A(n250), .B(r5[4]), .C(n251), .D(r4[4]), .Y(n279) );
  AOI22X1 U324 ( .A(n252), .B(r3[4]), .C(n253), .D(r2[4]), .Y(n277) );
  AOI22X1 U325 ( .A(n254), .B(r1[4]), .C(n255), .D(r0[4]), .Y(n276) );
  NAND3X1 U326 ( .A(n78), .B(n708), .C(n283), .Y(dout[3]) );
  AOI22X1 U328 ( .A(n248), .B(r7[3]), .C(n249), .D(r6[3]), .Y(n285) );
  AOI22X1 U329 ( .A(n250), .B(r5[3]), .C(n251), .D(r4[3]), .Y(n284) );
  AOI22X1 U330 ( .A(n252), .B(r3[3]), .C(n253), .D(r2[3]), .Y(n282) );
  AOI22X1 U331 ( .A(n254), .B(r1[3]), .C(n255), .D(r0[3]), .Y(n281) );
  NAND3X1 U332 ( .A(n75), .B(n705), .C(n288), .Y(dout[2]) );
  AOI22X1 U334 ( .A(n248), .B(r7[2]), .C(n249), .D(r6[2]), .Y(n290) );
  AOI22X1 U335 ( .A(n250), .B(r5[2]), .C(n251), .D(r4[2]), .Y(n289) );
  AOI22X1 U336 ( .A(n252), .B(r3[2]), .C(n253), .D(r2[2]), .Y(n287) );
  AOI22X1 U337 ( .A(n254), .B(r1[2]), .C(n255), .D(r0[2]), .Y(n286) );
  NAND3X1 U338 ( .A(n72), .B(n702), .C(n293), .Y(dout[1]) );
  AOI22X1 U340 ( .A(n248), .B(r7[1]), .C(n249), .D(r6[1]), .Y(n295) );
  AOI22X1 U341 ( .A(n250), .B(r5[1]), .C(n251), .D(r4[1]), .Y(n294) );
  AOI22X1 U342 ( .A(n252), .B(r3[1]), .C(n253), .D(r2[1]), .Y(n292) );
  AOI22X1 U343 ( .A(n254), .B(r1[1]), .C(n255), .D(r0[1]), .Y(n291) );
  NAND3X1 U344 ( .A(n69), .B(n699), .C(n298), .Y(dout[15]) );
  AOI22X1 U346 ( .A(n248), .B(r7[15]), .C(n249), .D(r6[15]), .Y(n300) );
  AOI22X1 U347 ( .A(n250), .B(r5[15]), .C(n251), .D(r4[15]), .Y(n299) );
  AOI22X1 U348 ( .A(n252), .B(r3[15]), .C(n253), .D(r2[15]), .Y(n297) );
  AOI22X1 U349 ( .A(n254), .B(r1[15]), .C(n255), .D(r0[15]), .Y(n296) );
  NAND3X1 U350 ( .A(n66), .B(n696), .C(n303), .Y(dout[14]) );
  AOI22X1 U352 ( .A(n248), .B(r7[14]), .C(n249), .D(r6[14]), .Y(n305) );
  AOI22X1 U353 ( .A(n250), .B(r5[14]), .C(n251), .D(r4[14]), .Y(n304) );
  AOI22X1 U354 ( .A(n252), .B(r3[14]), .C(n253), .D(r2[14]), .Y(n302) );
  AOI22X1 U355 ( .A(n254), .B(r1[14]), .C(n255), .D(r0[14]), .Y(n301) );
  NAND3X1 U356 ( .A(n63), .B(n693), .C(n308), .Y(dout[13]) );
  AOI22X1 U358 ( .A(n248), .B(r7[13]), .C(n249), .D(r6[13]), .Y(n310) );
  AOI22X1 U359 ( .A(n250), .B(r5[13]), .C(n251), .D(r4[13]), .Y(n309) );
  AOI22X1 U360 ( .A(n252), .B(r3[13]), .C(n253), .D(r2[13]), .Y(n307) );
  AOI22X1 U361 ( .A(n254), .B(r1[13]), .C(n255), .D(r0[13]), .Y(n306) );
  NAND3X1 U362 ( .A(n60), .B(n690), .C(n313), .Y(dout[12]) );
  AOI22X1 U364 ( .A(n248), .B(r7[12]), .C(n249), .D(r6[12]), .Y(n315) );
  AOI22X1 U365 ( .A(n250), .B(r5[12]), .C(n251), .D(r4[12]), .Y(n314) );
  AOI22X1 U366 ( .A(n252), .B(r3[12]), .C(n253), .D(r2[12]), .Y(n312) );
  AOI22X1 U367 ( .A(n254), .B(r1[12]), .C(n255), .D(r0[12]), .Y(n311) );
  NAND3X1 U368 ( .A(n57), .B(n687), .C(n318), .Y(dout[11]) );
  AOI22X1 U370 ( .A(n248), .B(r7[11]), .C(n249), .D(r6[11]), .Y(n320) );
  AOI22X1 U371 ( .A(n250), .B(r5[11]), .C(n251), .D(r4[11]), .Y(n319) );
  AOI22X1 U372 ( .A(n252), .B(r3[11]), .C(n253), .D(r2[11]), .Y(n317) );
  AOI22X1 U373 ( .A(n254), .B(r1[11]), .C(n255), .D(r0[11]), .Y(n316) );
  NAND3X1 U374 ( .A(n54), .B(n684), .C(n323), .Y(dout[10]) );
  AOI22X1 U376 ( .A(n248), .B(r7[10]), .C(n249), .D(r6[10]), .Y(n325) );
  AOI22X1 U377 ( .A(n250), .B(r5[10]), .C(n251), .D(r4[10]), .Y(n324) );
  AOI22X1 U378 ( .A(n252), .B(r3[10]), .C(n253), .D(r2[10]), .Y(n322) );
  AOI22X1 U379 ( .A(n254), .B(r1[10]), .C(n255), .D(r0[10]), .Y(n321) );
  NAND3X1 U380 ( .A(n51), .B(n681), .C(n328), .Y(dout[0]) );
  AOI22X1 U382 ( .A(n248), .B(r7[0]), .C(n249), .D(r6[0]), .Y(n330) );
  INVX1 U383 ( .A(n331), .Y(n249) );
  NAND3X1 U384 ( .A(readPtr[1]), .B(n332), .C(readPtr[2]), .Y(n331) );
  INVX1 U385 ( .A(n333), .Y(n248) );
  NAND3X1 U386 ( .A(readPtr[1]), .B(readPtr[0]), .C(readPtr[2]), .Y(n333) );
  AOI22X1 U387 ( .A(n250), .B(r5[0]), .C(n251), .D(r4[0]), .Y(n329) );
  INVX1 U388 ( .A(n334), .Y(n251) );
  NAND3X1 U389 ( .A(n332), .B(n335), .C(readPtr[2]), .Y(n334) );
  INVX1 U390 ( .A(n336), .Y(n250) );
  NAND3X1 U391 ( .A(readPtr[0]), .B(n335), .C(readPtr[2]), .Y(n336) );
  AOI22X1 U392 ( .A(n252), .B(r3[0]), .C(n253), .D(r2[0]), .Y(n327) );
  NOR3X1 U393 ( .A(readPtr[0]), .B(readPtr[2]), .C(n335), .Y(n253) );
  NOR3X1 U394 ( .A(n332), .B(readPtr[2]), .C(n335), .Y(n252) );
  INVX1 U395 ( .A(readPtr[1]), .Y(n335) );
  AOI22X1 U396 ( .A(n254), .B(r1[0]), .C(n255), .D(r0[0]), .Y(n326) );
  NOR3X1 U397 ( .A(readPtr[1]), .B(readPtr[2]), .C(readPtr[0]), .Y(n255) );
  NOR3X1 U398 ( .A(readPtr[1]), .B(readPtr[2]), .C(n332), .Y(n254) );
  INVX1 U399 ( .A(readPtr[0]), .Y(n332) );
  INVX1 U4 ( .A(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
  BUFX2 U6 ( .A(n329), .Y(n3) );
  INVX1 U7 ( .A(n6), .Y(n4) );
  INVX1 U10 ( .A(n4), .Y(n5) );
  BUFX2 U12 ( .A(n324), .Y(n6) );
  INVX1 U14 ( .A(n9), .Y(n7) );
  INVX1 U16 ( .A(n7), .Y(n8) );
  BUFX2 U18 ( .A(n319), .Y(n9) );
  INVX1 U20 ( .A(n12), .Y(n10) );
  INVX1 U22 ( .A(n10), .Y(n11) );
  BUFX2 U24 ( .A(n314), .Y(n12) );
  INVX1 U26 ( .A(n15), .Y(n13) );
  INVX1 U28 ( .A(n13), .Y(n14) );
  BUFX2 U30 ( .A(n309), .Y(n15) );
  INVX1 U32 ( .A(n18), .Y(n16) );
  INVX1 U34 ( .A(n16), .Y(n17) );
  BUFX2 U36 ( .A(n304), .Y(n18) );
  INVX1 U38 ( .A(n21), .Y(n19) );
  INVX1 U40 ( .A(n19), .Y(n20) );
  BUFX2 U41 ( .A(n299), .Y(n21) );
  INVX1 U42 ( .A(n24), .Y(n22) );
  INVX1 U43 ( .A(n22), .Y(n23) );
  BUFX2 U44 ( .A(n294), .Y(n24) );
  INVX1 U45 ( .A(n27), .Y(n25) );
  INVX1 U46 ( .A(n25), .Y(n26) );
  BUFX2 U47 ( .A(n289), .Y(n27) );
  INVX1 U48 ( .A(n30), .Y(n28) );
  INVX1 U49 ( .A(n28), .Y(n29) );
  BUFX2 U50 ( .A(n284), .Y(n30) );
  INVX1 U51 ( .A(n33), .Y(n31) );
  INVX1 U52 ( .A(n31), .Y(n32) );
  BUFX2 U53 ( .A(n279), .Y(n33) );
  INVX1 U54 ( .A(n36), .Y(n34) );
  INVX1 U55 ( .A(n34), .Y(n35) );
  BUFX2 U56 ( .A(n274), .Y(n36) );
  INVX1 U57 ( .A(n39), .Y(n37) );
  INVX1 U58 ( .A(n37), .Y(n38) );
  BUFX2 U59 ( .A(n269), .Y(n39) );
  INVX1 U60 ( .A(n42), .Y(n40) );
  INVX1 U61 ( .A(n40), .Y(n41) );
  BUFX2 U62 ( .A(n264), .Y(n42) );
  INVX1 U63 ( .A(n46), .Y(n44) );
  INVX1 U64 ( .A(n44), .Y(n45) );
  BUFX2 U65 ( .A(n259), .Y(n46) );
  INVX1 U66 ( .A(n49), .Y(n47) );
  INVX1 U67 ( .A(n47), .Y(n48) );
  BUFX2 U68 ( .A(n246), .Y(n49) );
  INVX1 U69 ( .A(n52), .Y(n50) );
  INVX1 U70 ( .A(n50), .Y(n51) );
  BUFX2 U71 ( .A(n326), .Y(n52) );
  INVX1 U72 ( .A(n55), .Y(n53) );
  INVX1 U73 ( .A(n53), .Y(n54) );
  BUFX2 U74 ( .A(n321), .Y(n55) );
  INVX1 U75 ( .A(n58), .Y(n56) );
  INVX1 U76 ( .A(n56), .Y(n57) );
  BUFX2 U77 ( .A(n316), .Y(n58) );
  INVX1 U78 ( .A(n61), .Y(n59) );
  INVX1 U79 ( .A(n59), .Y(n60) );
  BUFX2 U80 ( .A(n311), .Y(n61) );
  INVX1 U81 ( .A(n64), .Y(n62) );
  INVX1 U82 ( .A(n62), .Y(n63) );
  BUFX2 U83 ( .A(n306), .Y(n64) );
  INVX1 U84 ( .A(n67), .Y(n65) );
  INVX1 U85 ( .A(n65), .Y(n66) );
  BUFX2 U86 ( .A(n301), .Y(n67) );
  INVX1 U87 ( .A(n70), .Y(n68) );
  INVX1 U88 ( .A(n68), .Y(n69) );
  BUFX2 U89 ( .A(n296), .Y(n70) );
  INVX1 U90 ( .A(n73), .Y(n71) );
  INVX1 U91 ( .A(n71), .Y(n72) );
  BUFX2 U92 ( .A(n291), .Y(n73) );
  INVX1 U93 ( .A(n76), .Y(n74) );
  INVX1 U94 ( .A(n74), .Y(n75) );
  BUFX2 U95 ( .A(n286), .Y(n76) );
  INVX1 U96 ( .A(n79), .Y(n77) );
  INVX1 U97 ( .A(n77), .Y(n78) );
  BUFX2 U98 ( .A(n281), .Y(n79) );
  INVX1 U99 ( .A(n82), .Y(n80) );
  INVX1 U100 ( .A(n80), .Y(n81) );
  BUFX2 U101 ( .A(n276), .Y(n82) );
  INVX1 U102 ( .A(n85), .Y(n83) );
  INVX1 U103 ( .A(n83), .Y(n84) );
  BUFX2 U104 ( .A(n271), .Y(n85) );
  INVX1 U106 ( .A(n88), .Y(n86) );
  INVX1 U108 ( .A(n86), .Y(n87) );
  BUFX2 U110 ( .A(n266), .Y(n88) );
  INVX1 U112 ( .A(n142), .Y(n89) );
  INVX1 U114 ( .A(n89), .Y(n125) );
  BUFX2 U116 ( .A(n261), .Y(n142) );
  INVX1 U118 ( .A(n468), .Y(n241) );
  INVX1 U120 ( .A(n241), .Y(n467) );
  BUFX2 U122 ( .A(n256), .Y(n468) );
  INVX1 U124 ( .A(n471), .Y(n469) );
  INVX1 U126 ( .A(n469), .Y(n470) );
  BUFX2 U128 ( .A(n243), .Y(n471) );
  INVX1 U130 ( .A(n474), .Y(n472) );
  INVX1 U132 ( .A(n472), .Y(n473) );
  AND2X1 U134 ( .A(r2[15]), .B(n159), .Y(n240) );
  INVX1 U136 ( .A(n240), .Y(n474) );
  INVX1 U138 ( .A(n477), .Y(n475) );
  INVX1 U140 ( .A(n475), .Y(n476) );
  AND2X1 U142 ( .A(r2[14]), .B(n159), .Y(n239) );
  INVX1 U144 ( .A(n239), .Y(n477) );
  INVX1 U146 ( .A(n480), .Y(n478) );
  INVX1 U148 ( .A(n478), .Y(n479) );
  AND2X1 U150 ( .A(r2[13]), .B(n159), .Y(n238) );
  INVX1 U152 ( .A(n238), .Y(n480) );
  INVX1 U154 ( .A(n483), .Y(n481) );
  INVX1 U156 ( .A(n481), .Y(n482) );
  AND2X1 U158 ( .A(r2[12]), .B(n159), .Y(n237) );
  INVX1 U160 ( .A(n237), .Y(n483) );
  INVX1 U162 ( .A(n486), .Y(n484) );
  INVX1 U164 ( .A(n484), .Y(n485) );
  AND2X1 U166 ( .A(r2[11]), .B(n159), .Y(n236) );
  INVX1 U168 ( .A(n236), .Y(n486) );
  INVX1 U169 ( .A(n489), .Y(n487) );
  INVX1 U170 ( .A(n487), .Y(n488) );
  AND2X1 U171 ( .A(r2[10]), .B(n159), .Y(n235) );
  INVX1 U172 ( .A(n235), .Y(n489) );
  INVX1 U173 ( .A(n492), .Y(n490) );
  INVX1 U174 ( .A(n490), .Y(n491) );
  AND2X1 U175 ( .A(r2[9]), .B(n159), .Y(n234) );
  INVX1 U176 ( .A(n234), .Y(n492) );
  INVX1 U177 ( .A(n495), .Y(n493) );
  INVX1 U178 ( .A(n493), .Y(n494) );
  AND2X1 U179 ( .A(r2[8]), .B(n159), .Y(n233) );
  INVX1 U180 ( .A(n233), .Y(n495) );
  INVX1 U181 ( .A(n498), .Y(n496) );
  INVX1 U182 ( .A(n496), .Y(n497) );
  AND2X1 U183 ( .A(r2[7]), .B(n159), .Y(n232) );
  INVX1 U184 ( .A(n232), .Y(n498) );
  INVX1 U185 ( .A(n501), .Y(n499) );
  INVX1 U186 ( .A(n499), .Y(n500) );
  AND2X1 U187 ( .A(r2[6]), .B(n159), .Y(n231) );
  INVX1 U188 ( .A(n231), .Y(n501) );
  INVX1 U189 ( .A(n504), .Y(n502) );
  INVX1 U190 ( .A(n502), .Y(n503) );
  AND2X1 U191 ( .A(r2[5]), .B(n159), .Y(n230) );
  INVX1 U192 ( .A(n230), .Y(n504) );
  INVX1 U193 ( .A(n507), .Y(n505) );
  INVX1 U194 ( .A(n505), .Y(n506) );
  AND2X1 U195 ( .A(r2[4]), .B(n159), .Y(n229) );
  INVX1 U196 ( .A(n229), .Y(n507) );
  INVX1 U197 ( .A(n510), .Y(n508) );
  INVX1 U198 ( .A(n508), .Y(n509) );
  AND2X1 U199 ( .A(r2[3]), .B(n159), .Y(n228) );
  INVX1 U200 ( .A(n228), .Y(n510) );
  INVX1 U201 ( .A(n513), .Y(n511) );
  INVX1 U202 ( .A(n511), .Y(n512) );
  AND2X1 U203 ( .A(r2[2]), .B(n159), .Y(n227) );
  INVX1 U204 ( .A(n227), .Y(n513) );
  INVX1 U205 ( .A(n516), .Y(n514) );
  INVX1 U206 ( .A(n514), .Y(n515) );
  AND2X1 U207 ( .A(r2[1]), .B(n159), .Y(n226) );
  INVX1 U208 ( .A(n226), .Y(n516) );
  INVX1 U209 ( .A(n519), .Y(n517) );
  INVX1 U210 ( .A(n517), .Y(n518) );
  AND2X1 U211 ( .A(r2[0]), .B(n159), .Y(n225) );
  INVX1 U212 ( .A(n225), .Y(n519) );
  INVX1 U213 ( .A(n522), .Y(n520) );
  INVX1 U214 ( .A(n520), .Y(n521) );
  AND2X1 U215 ( .A(r0[15]), .B(n92), .Y(n191) );
  INVX1 U216 ( .A(n191), .Y(n522) );
  INVX1 U217 ( .A(n525), .Y(n523) );
  INVX1 U218 ( .A(n523), .Y(n524) );
  AND2X1 U219 ( .A(r0[14]), .B(n92), .Y(n190) );
  INVX1 U220 ( .A(n190), .Y(n525) );
  INVX1 U221 ( .A(n528), .Y(n526) );
  INVX1 U222 ( .A(n526), .Y(n527) );
  AND2X1 U223 ( .A(r0[13]), .B(n92), .Y(n189) );
  INVX1 U224 ( .A(n189), .Y(n528) );
  INVX1 U225 ( .A(n531), .Y(n529) );
  INVX1 U226 ( .A(n529), .Y(n530) );
  AND2X1 U227 ( .A(r0[12]), .B(n92), .Y(n188) );
  INVX1 U228 ( .A(n188), .Y(n531) );
  INVX1 U229 ( .A(n534), .Y(n532) );
  INVX1 U230 ( .A(n532), .Y(n533) );
  AND2X1 U231 ( .A(r0[11]), .B(n92), .Y(n187) );
  INVX1 U232 ( .A(n187), .Y(n534) );
  INVX1 U234 ( .A(n537), .Y(n535) );
  INVX1 U237 ( .A(n535), .Y(n536) );
  AND2X1 U240 ( .A(r0[10]), .B(n92), .Y(n186) );
  INVX1 U243 ( .A(n186), .Y(n537) );
  INVX1 U246 ( .A(n540), .Y(n538) );
  INVX1 U249 ( .A(n538), .Y(n539) );
  AND2X1 U252 ( .A(r0[9]), .B(n92), .Y(n185) );
  INVX1 U255 ( .A(n185), .Y(n540) );
  INVX1 U258 ( .A(n543), .Y(n541) );
  INVX1 U261 ( .A(n541), .Y(n542) );
  AND2X1 U264 ( .A(r0[8]), .B(n92), .Y(n184) );
  INVX1 U267 ( .A(n184), .Y(n543) );
  INVX1 U270 ( .A(n546), .Y(n544) );
  INVX1 U273 ( .A(n544), .Y(n545) );
  AND2X1 U276 ( .A(r0[7]), .B(n92), .Y(n183) );
  INVX1 U279 ( .A(n183), .Y(n546) );
  INVX1 U280 ( .A(n549), .Y(n547) );
  INVX1 U283 ( .A(n547), .Y(n548) );
  AND2X1 U285 ( .A(r0[6]), .B(n92), .Y(n182) );
  INVX1 U291 ( .A(n182), .Y(n549) );
  INVX1 U297 ( .A(n552), .Y(n550) );
  INVX1 U303 ( .A(n550), .Y(n551) );
  AND2X1 U309 ( .A(r0[5]), .B(n92), .Y(n181) );
  INVX1 U315 ( .A(n181), .Y(n552) );
  INVX1 U321 ( .A(n555), .Y(n553) );
  INVX1 U327 ( .A(n553), .Y(n554) );
  AND2X1 U333 ( .A(r0[4]), .B(n92), .Y(n180) );
  INVX1 U339 ( .A(n180), .Y(n555) );
  INVX1 U345 ( .A(n558), .Y(n556) );
  INVX1 U351 ( .A(n556), .Y(n557) );
  AND2X1 U357 ( .A(r0[3]), .B(n92), .Y(n179) );
  INVX1 U363 ( .A(n179), .Y(n558) );
  INVX1 U369 ( .A(n561), .Y(n559) );
  INVX1 U375 ( .A(n559), .Y(n560) );
  AND2X1 U381 ( .A(r0[2]), .B(n92), .Y(n178) );
  INVX1 U400 ( .A(n178), .Y(n561) );
  INVX1 U401 ( .A(n564), .Y(n562) );
  INVX1 U402 ( .A(n562), .Y(n563) );
  AND2X1 U403 ( .A(r0[1]), .B(n92), .Y(n177) );
  INVX1 U404 ( .A(n177), .Y(n564) );
  INVX1 U405 ( .A(n567), .Y(n565) );
  INVX1 U406 ( .A(n565), .Y(n566) );
  AND2X1 U407 ( .A(r0[0]), .B(n92), .Y(n176) );
  INVX1 U408 ( .A(n176), .Y(n567) );
  INVX1 U409 ( .A(n570), .Y(n568) );
  INVX1 U410 ( .A(n568), .Y(n569) );
  AND2X1 U411 ( .A(r3[15]), .B(n159), .Y(n175) );
  INVX1 U412 ( .A(n175), .Y(n570) );
  INVX1 U413 ( .A(n573), .Y(n571) );
  INVX1 U414 ( .A(n571), .Y(n572) );
  AND2X1 U415 ( .A(r3[14]), .B(n159), .Y(n174) );
  INVX1 U416 ( .A(n174), .Y(n573) );
  INVX1 U417 ( .A(n576), .Y(n574) );
  INVX1 U418 ( .A(n574), .Y(n575) );
  AND2X1 U419 ( .A(r3[13]), .B(n159), .Y(n173) );
  INVX1 U420 ( .A(n173), .Y(n576) );
  INVX1 U421 ( .A(n579), .Y(n577) );
  INVX1 U422 ( .A(n577), .Y(n578) );
  AND2X1 U423 ( .A(r3[12]), .B(n159), .Y(n172) );
  INVX1 U424 ( .A(n172), .Y(n579) );
  INVX1 U425 ( .A(n582), .Y(n580) );
  INVX1 U426 ( .A(n580), .Y(n581) );
  AND2X1 U427 ( .A(r3[11]), .B(n159), .Y(n171) );
  INVX1 U428 ( .A(n171), .Y(n582) );
  INVX1 U429 ( .A(n585), .Y(n583) );
  INVX1 U430 ( .A(n583), .Y(n584) );
  AND2X1 U431 ( .A(r3[10]), .B(n159), .Y(n170) );
  INVX1 U432 ( .A(n170), .Y(n585) );
  INVX1 U433 ( .A(n588), .Y(n586) );
  INVX1 U434 ( .A(n586), .Y(n587) );
  AND2X1 U435 ( .A(r3[9]), .B(n159), .Y(n169) );
  INVX1 U436 ( .A(n169), .Y(n588) );
  INVX1 U437 ( .A(n591), .Y(n589) );
  INVX1 U438 ( .A(n589), .Y(n590) );
  AND2X1 U439 ( .A(r3[8]), .B(n159), .Y(n168) );
  INVX1 U440 ( .A(n168), .Y(n591) );
  INVX1 U441 ( .A(n594), .Y(n592) );
  INVX1 U442 ( .A(n592), .Y(n593) );
  AND2X1 U443 ( .A(r3[7]), .B(n159), .Y(n167) );
  INVX1 U444 ( .A(n167), .Y(n594) );
  INVX1 U445 ( .A(n597), .Y(n595) );
  INVX1 U446 ( .A(n595), .Y(n596) );
  AND2X1 U447 ( .A(r3[6]), .B(n159), .Y(n166) );
  INVX1 U448 ( .A(n166), .Y(n597) );
  INVX1 U449 ( .A(n600), .Y(n598) );
  INVX1 U450 ( .A(n598), .Y(n599) );
  AND2X1 U451 ( .A(r3[5]), .B(n159), .Y(n165) );
  INVX1 U452 ( .A(n165), .Y(n600) );
  INVX1 U453 ( .A(n603), .Y(n601) );
  INVX1 U454 ( .A(n601), .Y(n602) );
  AND2X1 U455 ( .A(r3[4]), .B(n159), .Y(n164) );
  INVX1 U456 ( .A(n164), .Y(n603) );
  INVX1 U457 ( .A(n606), .Y(n604) );
  INVX1 U458 ( .A(n604), .Y(n605) );
  AND2X1 U459 ( .A(r3[3]), .B(n159), .Y(n163) );
  INVX1 U460 ( .A(n163), .Y(n606) );
  INVX1 U461 ( .A(n609), .Y(n607) );
  INVX1 U462 ( .A(n607), .Y(n608) );
  AND2X1 U463 ( .A(r3[2]), .B(n159), .Y(n162) );
  INVX1 U464 ( .A(n162), .Y(n609) );
  INVX1 U465 ( .A(n612), .Y(n610) );
  INVX1 U466 ( .A(n610), .Y(n611) );
  AND2X1 U467 ( .A(r3[1]), .B(n159), .Y(n161) );
  INVX1 U468 ( .A(n161), .Y(n612) );
  INVX1 U469 ( .A(n615), .Y(n613) );
  INVX1 U470 ( .A(n613), .Y(n614) );
  AND2X1 U471 ( .A(r3[0]), .B(n159), .Y(n160) );
  INVX1 U472 ( .A(n160), .Y(n615) );
  INVX1 U473 ( .A(n618), .Y(n616) );
  INVX1 U474 ( .A(n616), .Y(n617) );
  AND2X1 U475 ( .A(r1[15]), .B(n92), .Y(n124) );
  INVX1 U476 ( .A(n124), .Y(n618) );
  INVX1 U477 ( .A(n621), .Y(n619) );
  INVX1 U478 ( .A(n619), .Y(n620) );
  AND2X1 U479 ( .A(r1[14]), .B(n92), .Y(n122) );
  INVX1 U480 ( .A(n122), .Y(n621) );
  INVX1 U481 ( .A(n624), .Y(n622) );
  INVX1 U482 ( .A(n622), .Y(n623) );
  AND2X1 U483 ( .A(r1[13]), .B(n92), .Y(n120) );
  INVX1 U484 ( .A(n120), .Y(n624) );
  INVX1 U485 ( .A(n627), .Y(n625) );
  INVX1 U486 ( .A(n625), .Y(n626) );
  AND2X1 U487 ( .A(r1[12]), .B(n92), .Y(n118) );
  INVX1 U488 ( .A(n118), .Y(n627) );
  INVX1 U489 ( .A(n630), .Y(n628) );
  INVX1 U490 ( .A(n628), .Y(n629) );
  AND2X1 U491 ( .A(r1[11]), .B(n92), .Y(n116) );
  INVX1 U492 ( .A(n116), .Y(n630) );
  INVX1 U493 ( .A(n633), .Y(n631) );
  INVX1 U494 ( .A(n631), .Y(n632) );
  AND2X1 U495 ( .A(r1[10]), .B(n92), .Y(n114) );
  INVX1 U496 ( .A(n114), .Y(n633) );
  INVX1 U497 ( .A(n636), .Y(n634) );
  INVX1 U498 ( .A(n634), .Y(n635) );
  AND2X1 U499 ( .A(r1[9]), .B(n92), .Y(n112) );
  INVX1 U500 ( .A(n112), .Y(n636) );
  INVX1 U501 ( .A(n639), .Y(n637) );
  INVX1 U502 ( .A(n637), .Y(n638) );
  AND2X1 U503 ( .A(r1[8]), .B(n92), .Y(n110) );
  INVX1 U504 ( .A(n110), .Y(n639) );
  INVX1 U505 ( .A(n642), .Y(n640) );
  INVX1 U506 ( .A(n640), .Y(n641) );
  AND2X1 U507 ( .A(r1[7]), .B(n92), .Y(n108) );
  INVX1 U508 ( .A(n108), .Y(n642) );
  INVX1 U509 ( .A(n645), .Y(n643) );
  INVX1 U510 ( .A(n643), .Y(n644) );
  AND2X1 U511 ( .A(r1[6]), .B(n92), .Y(n106) );
  INVX1 U512 ( .A(n106), .Y(n645) );
  INVX1 U513 ( .A(n648), .Y(n646) );
  INVX1 U514 ( .A(n646), .Y(n647) );
  AND2X1 U515 ( .A(r1[5]), .B(n92), .Y(n104) );
  INVX1 U516 ( .A(n104), .Y(n648) );
  INVX1 U517 ( .A(n651), .Y(n649) );
  INVX1 U518 ( .A(n649), .Y(n650) );
  AND2X1 U519 ( .A(r1[4]), .B(n92), .Y(n102) );
  INVX1 U520 ( .A(n102), .Y(n651) );
  INVX1 U521 ( .A(n654), .Y(n652) );
  INVX1 U522 ( .A(n652), .Y(n653) );
  AND2X1 U523 ( .A(r1[3]), .B(n92), .Y(n100) );
  INVX1 U524 ( .A(n100), .Y(n654) );
  INVX1 U525 ( .A(n657), .Y(n655) );
  INVX1 U526 ( .A(n655), .Y(n656) );
  AND2X1 U527 ( .A(r1[2]), .B(n92), .Y(n98) );
  INVX1 U528 ( .A(n98), .Y(n657) );
  INVX1 U529 ( .A(n660), .Y(n658) );
  INVX1 U530 ( .A(n658), .Y(n659) );
  AND2X1 U531 ( .A(r1[1]), .B(n92), .Y(n96) );
  INVX1 U532 ( .A(n96), .Y(n660) );
  INVX1 U533 ( .A(n663), .Y(n661) );
  INVX1 U534 ( .A(n661), .Y(n662) );
  AND2X1 U535 ( .A(r1[0]), .B(n92), .Y(n94) );
  INVX1 U536 ( .A(n94), .Y(n663) );
  BUFX2 U537 ( .A(n330), .Y(n664) );
  AND2X2 U538 ( .A(n2), .B(n664), .Y(n328) );
  BUFX2 U539 ( .A(n325), .Y(n665) );
  AND2X2 U540 ( .A(n5), .B(n665), .Y(n323) );
  BUFX2 U541 ( .A(n320), .Y(n666) );
  AND2X2 U542 ( .A(n8), .B(n666), .Y(n318) );
  BUFX2 U543 ( .A(n315), .Y(n667) );
  AND2X2 U544 ( .A(n11), .B(n667), .Y(n313) );
  BUFX2 U545 ( .A(n310), .Y(n668) );
  AND2X2 U546 ( .A(n14), .B(n668), .Y(n308) );
  BUFX2 U547 ( .A(n305), .Y(n669) );
  AND2X2 U548 ( .A(n17), .B(n669), .Y(n303) );
  BUFX2 U549 ( .A(n300), .Y(n670) );
  AND2X2 U550 ( .A(n20), .B(n670), .Y(n298) );
  BUFX2 U551 ( .A(n295), .Y(n671) );
  AND2X2 U552 ( .A(n23), .B(n671), .Y(n293) );
  BUFX2 U553 ( .A(n290), .Y(n672) );
  AND2X2 U554 ( .A(n26), .B(n672), .Y(n288) );
  BUFX2 U555 ( .A(n285), .Y(n673) );
  AND2X2 U556 ( .A(n29), .B(n673), .Y(n283) );
  BUFX2 U557 ( .A(n280), .Y(n674) );
  AND2X2 U558 ( .A(n32), .B(n674), .Y(n278) );
  BUFX2 U559 ( .A(n275), .Y(n675) );
  AND2X2 U560 ( .A(n35), .B(n675), .Y(n273) );
  BUFX2 U561 ( .A(n270), .Y(n676) );
  AND2X2 U562 ( .A(n38), .B(n676), .Y(n268) );
  BUFX2 U563 ( .A(n265), .Y(n677) );
  AND2X2 U564 ( .A(n41), .B(n677), .Y(n263) );
  BUFX2 U565 ( .A(n260), .Y(n678) );
  AND2X2 U566 ( .A(n45), .B(n678), .Y(n258) );
  BUFX2 U567 ( .A(n247), .Y(n679) );
  AND2X2 U568 ( .A(n48), .B(n679), .Y(n245) );
  INVX1 U569 ( .A(n682), .Y(n680) );
  INVX1 U570 ( .A(n680), .Y(n681) );
  BUFX2 U571 ( .A(n327), .Y(n682) );
  INVX1 U572 ( .A(n685), .Y(n683) );
  INVX1 U573 ( .A(n683), .Y(n684) );
  BUFX2 U574 ( .A(n322), .Y(n685) );
  INVX1 U575 ( .A(n688), .Y(n686) );
  INVX1 U576 ( .A(n686), .Y(n687) );
  BUFX2 U577 ( .A(n317), .Y(n688) );
  INVX1 U578 ( .A(n691), .Y(n689) );
  INVX1 U579 ( .A(n689), .Y(n690) );
  BUFX2 U580 ( .A(n312), .Y(n691) );
  INVX1 U581 ( .A(n694), .Y(n692) );
  INVX1 U582 ( .A(n692), .Y(n693) );
  BUFX2 U583 ( .A(n307), .Y(n694) );
  INVX1 U584 ( .A(n697), .Y(n695) );
  INVX1 U585 ( .A(n695), .Y(n696) );
  BUFX2 U586 ( .A(n302), .Y(n697) );
  INVX1 U587 ( .A(n700), .Y(n698) );
  INVX1 U588 ( .A(n698), .Y(n699) );
  BUFX2 U589 ( .A(n297), .Y(n700) );
  INVX1 U590 ( .A(n703), .Y(n701) );
  INVX1 U591 ( .A(n701), .Y(n702) );
  BUFX2 U592 ( .A(n292), .Y(n703) );
  INVX1 U593 ( .A(n706), .Y(n704) );
  INVX1 U594 ( .A(n704), .Y(n705) );
  BUFX2 U595 ( .A(n287), .Y(n706) );
  INVX1 U596 ( .A(n709), .Y(n707) );
  INVX1 U597 ( .A(n707), .Y(n708) );
  BUFX2 U598 ( .A(n282), .Y(n709) );
  INVX1 U599 ( .A(n712), .Y(n710) );
  INVX1 U600 ( .A(n710), .Y(n711) );
  BUFX2 U601 ( .A(n277), .Y(n712) );
  INVX1 U602 ( .A(n715), .Y(n713) );
  INVX1 U603 ( .A(n713), .Y(n714) );
  BUFX2 U604 ( .A(n272), .Y(n715) );
  INVX1 U605 ( .A(n718), .Y(n716) );
  INVX1 U606 ( .A(n716), .Y(n717) );
  BUFX2 U607 ( .A(n267), .Y(n718) );
  INVX1 U608 ( .A(n721), .Y(n719) );
  INVX1 U609 ( .A(n719), .Y(n720) );
  BUFX2 U610 ( .A(n262), .Y(n721) );
  INVX1 U611 ( .A(n724), .Y(n722) );
  INVX1 U612 ( .A(n722), .Y(n723) );
  BUFX2 U613 ( .A(n257), .Y(n724) );
  INVX1 U614 ( .A(n727), .Y(n725) );
  INVX1 U615 ( .A(n725), .Y(n726) );
  BUFX2 U616 ( .A(n244), .Y(n727) );
  INVX1 U617 ( .A(n730), .Y(n728) );
  INVX1 U618 ( .A(n728), .Y(n729) );
  BUFX2 U619 ( .A(count_0_), .Y(n730) );
  INVX1 U620 ( .A(n733), .Y(n731) );
  INVX1 U621 ( .A(n731), .Y(n732) );
  BUFX2 U622 ( .A(F0), .Y(n733) );
  INVX8 U623 ( .A(n745), .Y(n734) );
  INVX8 U624 ( .A(n745), .Y(n735) );
  INVX8 U625 ( .A(n745), .Y(n736) );
  INVX8 U626 ( .A(n744), .Y(n737) );
  INVX8 U627 ( .A(n744), .Y(n738) );
  INVX8 U628 ( .A(n744), .Y(n739) );
  INVX8 U629 ( .A(n743), .Y(n740) );
  INVX8 U630 ( .A(n743), .Y(n741) );
  INVX8 U631 ( .A(n743), .Y(n742) );
  INVX8 U632 ( .A(fStrobe), .Y(n743) );
  INVX8 U633 ( .A(fStrobe), .Y(n744) );
  INVX8 U634 ( .A(fStrobe), .Y(n745) );
  INVX2 U635 ( .A(n729), .Y(n159) );
  INVX2 U636 ( .A(n224), .Y(n92) );
  INVX2 U637 ( .A(n143), .Y(n369) );
  INVX2 U638 ( .A(r5[0]), .Y(n143) );
  INVX2 U639 ( .A(n144), .Y(n370) );
  INVX2 U640 ( .A(r5[1]), .Y(n144) );
  INVX2 U641 ( .A(n145), .Y(n371) );
  INVX2 U642 ( .A(r5[2]), .Y(n145) );
  INVX2 U643 ( .A(n146), .Y(n372) );
  INVX2 U644 ( .A(r5[3]), .Y(n146) );
  INVX2 U645 ( .A(n147), .Y(n373) );
  INVX2 U646 ( .A(r5[4]), .Y(n147) );
  INVX2 U647 ( .A(n148), .Y(n374) );
  INVX2 U648 ( .A(r5[5]), .Y(n148) );
  INVX2 U649 ( .A(n149), .Y(n375) );
  INVX2 U650 ( .A(r5[6]), .Y(n149) );
  INVX2 U651 ( .A(n150), .Y(n376) );
  INVX2 U652 ( .A(r5[7]), .Y(n150) );
  INVX2 U653 ( .A(n151), .Y(n377) );
  INVX2 U654 ( .A(r5[8]), .Y(n151) );
  INVX2 U655 ( .A(n152), .Y(n378) );
  INVX2 U656 ( .A(r5[9]), .Y(n152) );
  INVX2 U657 ( .A(n153), .Y(n379) );
  INVX2 U658 ( .A(r5[10]), .Y(n153) );
  INVX2 U659 ( .A(n154), .Y(n380) );
  INVX2 U660 ( .A(r5[11]), .Y(n154) );
  INVX2 U661 ( .A(n155), .Y(n381) );
  INVX2 U662 ( .A(r5[12]), .Y(n155) );
  INVX2 U663 ( .A(n156), .Y(n382) );
  INVX2 U664 ( .A(r5[13]), .Y(n156) );
  INVX2 U665 ( .A(n157), .Y(n383) );
  INVX2 U666 ( .A(r5[14]), .Y(n157) );
  INVX2 U667 ( .A(n158), .Y(n384) );
  INVX2 U668 ( .A(r5[15]), .Y(n158) );
  INVX2 U669 ( .A(n208), .Y(n433) );
  INVX2 U670 ( .A(r4[0]), .Y(n208) );
  INVX2 U671 ( .A(n209), .Y(n434) );
  INVX2 U672 ( .A(r4[1]), .Y(n209) );
  INVX2 U673 ( .A(n210), .Y(n435) );
  INVX2 U674 ( .A(r4[2]), .Y(n210) );
  INVX2 U675 ( .A(n211), .Y(n436) );
  INVX2 U676 ( .A(r4[3]), .Y(n211) );
  INVX2 U677 ( .A(n212), .Y(n437) );
  INVX2 U678 ( .A(r4[4]), .Y(n212) );
  INVX2 U679 ( .A(n213), .Y(n438) );
  INVX2 U680 ( .A(r4[5]), .Y(n213) );
  INVX2 U681 ( .A(n214), .Y(n439) );
  INVX2 U682 ( .A(r4[6]), .Y(n214) );
  INVX2 U683 ( .A(n215), .Y(n440) );
  INVX2 U684 ( .A(r4[7]), .Y(n215) );
  INVX2 U685 ( .A(n216), .Y(n441) );
  INVX2 U686 ( .A(r4[8]), .Y(n216) );
  INVX2 U687 ( .A(n217), .Y(n442) );
  INVX2 U688 ( .A(r4[9]), .Y(n217) );
  INVX2 U689 ( .A(n218), .Y(n443) );
  INVX2 U690 ( .A(r4[10]), .Y(n218) );
  INVX2 U691 ( .A(n219), .Y(n444) );
  INVX2 U692 ( .A(r4[11]), .Y(n219) );
  INVX2 U693 ( .A(n220), .Y(n445) );
  INVX2 U694 ( .A(r4[12]), .Y(n220) );
  INVX2 U695 ( .A(n221), .Y(n446) );
  INVX2 U696 ( .A(r4[13]), .Y(n221) );
  INVX2 U697 ( .A(n222), .Y(n447) );
  INVX2 U698 ( .A(r4[14]), .Y(n222) );
  INVX2 U699 ( .A(n223), .Y(n448) );
  INVX2 U700 ( .A(r4[15]), .Y(n223) );
  INVX2 U701 ( .A(n126), .Y(n353) );
  INVX2 U702 ( .A(r7[0]), .Y(n126) );
  INVX2 U703 ( .A(n127), .Y(n354) );
  INVX2 U704 ( .A(r7[1]), .Y(n127) );
  INVX2 U705 ( .A(n128), .Y(n355) );
  INVX2 U706 ( .A(r7[2]), .Y(n128) );
  INVX2 U707 ( .A(n129), .Y(n356) );
  INVX2 U708 ( .A(r7[3]), .Y(n129) );
  INVX2 U709 ( .A(n130), .Y(n357) );
  INVX2 U710 ( .A(r7[4]), .Y(n130) );
  INVX2 U711 ( .A(n131), .Y(n358) );
  INVX2 U712 ( .A(r7[5]), .Y(n131) );
  INVX2 U713 ( .A(n132), .Y(n359) );
  INVX2 U714 ( .A(r7[6]), .Y(n132) );
  INVX2 U715 ( .A(n133), .Y(n360) );
  INVX2 U716 ( .A(r7[7]), .Y(n133) );
  INVX2 U717 ( .A(n134), .Y(n361) );
  INVX2 U718 ( .A(r7[8]), .Y(n134) );
  INVX2 U719 ( .A(n135), .Y(n362) );
  INVX2 U720 ( .A(r7[9]), .Y(n135) );
  INVX2 U721 ( .A(n136), .Y(n363) );
  INVX2 U722 ( .A(r7[10]), .Y(n136) );
  INVX2 U723 ( .A(n137), .Y(n364) );
  INVX2 U724 ( .A(r7[11]), .Y(n137) );
  INVX2 U725 ( .A(n138), .Y(n365) );
  INVX2 U726 ( .A(r7[12]), .Y(n138) );
  INVX2 U727 ( .A(n139), .Y(n366) );
  INVX2 U728 ( .A(r7[13]), .Y(n139) );
  INVX2 U729 ( .A(n140), .Y(n367) );
  INVX2 U730 ( .A(r7[14]), .Y(n140) );
  INVX2 U731 ( .A(n141), .Y(n368) );
  INVX2 U732 ( .A(r7[15]), .Y(n141) );
  INVX2 U733 ( .A(n192), .Y(n417) );
  INVX2 U734 ( .A(r6[0]), .Y(n192) );
  INVX2 U735 ( .A(n193), .Y(n418) );
  INVX2 U736 ( .A(r6[1]), .Y(n193) );
  INVX2 U737 ( .A(n194), .Y(n419) );
  INVX2 U738 ( .A(r6[2]), .Y(n194) );
  INVX2 U739 ( .A(n195), .Y(n420) );
  INVX2 U740 ( .A(r6[3]), .Y(n195) );
  INVX2 U741 ( .A(n196), .Y(n421) );
  INVX2 U742 ( .A(r6[4]), .Y(n196) );
  INVX2 U743 ( .A(n197), .Y(n422) );
  INVX2 U744 ( .A(r6[5]), .Y(n197) );
  INVX2 U745 ( .A(n198), .Y(n423) );
  INVX2 U746 ( .A(r6[6]), .Y(n198) );
  INVX2 U747 ( .A(n199), .Y(n424) );
  INVX2 U748 ( .A(r6[7]), .Y(n199) );
  INVX2 U749 ( .A(n200), .Y(n425) );
  INVX2 U750 ( .A(r6[8]), .Y(n200) );
  INVX2 U751 ( .A(n201), .Y(n426) );
  INVX2 U752 ( .A(r6[9]), .Y(n201) );
  INVX2 U753 ( .A(n202), .Y(n427) );
  INVX2 U754 ( .A(r6[10]), .Y(n202) );
  INVX2 U755 ( .A(n203), .Y(n428) );
  INVX2 U756 ( .A(r6[11]), .Y(n203) );
  INVX2 U757 ( .A(n204), .Y(n429) );
  INVX2 U758 ( .A(r6[12]), .Y(n204) );
  INVX2 U759 ( .A(n205), .Y(n430) );
  INVX2 U760 ( .A(r6[13]), .Y(n205) );
  INVX2 U761 ( .A(n206), .Y(n431) );
  INVX2 U762 ( .A(r6[14]), .Y(n206) );
  INVX2 U763 ( .A(n207), .Y(n432) );
  INVX2 U764 ( .A(r6[15]), .Y(n207) );
endmodule


module Processing_logic_DW01_inc_0 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;

  wire   [31:2] carry;

  HAX1 U1_1_30 ( .A(A[30]), .B(carry[30]), .YC(carry[31]), .YS(SUM[30]) );
  HAX1 U1_1_29 ( .A(A[29]), .B(carry[29]), .YC(carry[30]), .YS(SUM[29]) );
  HAX1 U1_1_28 ( .A(A[28]), .B(carry[28]), .YC(carry[29]), .YS(SUM[28]) );
  HAX1 U1_1_27 ( .A(A[27]), .B(carry[27]), .YC(carry[28]), .YS(SUM[27]) );
  HAX1 U1_1_26 ( .A(A[26]), .B(carry[26]), .YC(carry[27]), .YS(SUM[26]) );
  HAX1 U1_1_25 ( .A(A[25]), .B(carry[25]), .YC(carry[26]), .YS(SUM[25]) );
  HAX1 U1_1_24 ( .A(A[24]), .B(carry[24]), .YC(carry[25]), .YS(SUM[24]) );
  HAX1 U1_1_23 ( .A(A[23]), .B(carry[23]), .YC(carry[24]), .YS(SUM[23]) );
  HAX1 U1_1_22 ( .A(A[22]), .B(carry[22]), .YC(carry[23]), .YS(SUM[22]) );
  HAX1 U1_1_21 ( .A(A[21]), .B(carry[21]), .YC(carry[22]), .YS(SUM[21]) );
  HAX1 U1_1_20 ( .A(A[20]), .B(carry[20]), .YC(carry[21]), .YS(SUM[20]) );
  HAX1 U1_1_19 ( .A(A[19]), .B(carry[19]), .YC(carry[20]), .YS(SUM[19]) );
  HAX1 U1_1_18 ( .A(A[18]), .B(carry[18]), .YC(carry[19]), .YS(SUM[18]) );
  HAX1 U1_1_17 ( .A(A[17]), .B(carry[17]), .YC(carry[18]), .YS(SUM[17]) );
  HAX1 U1_1_16 ( .A(A[16]), .B(carry[16]), .YC(carry[17]), .YS(SUM[16]) );
  HAX1 U1_1_15 ( .A(A[15]), .B(carry[15]), .YC(carry[16]), .YS(SUM[15]) );
  HAX1 U1_1_14 ( .A(A[14]), .B(carry[14]), .YC(carry[15]), .YS(SUM[14]) );
  HAX1 U1_1_13 ( .A(A[13]), .B(carry[13]), .YC(carry[14]), .YS(SUM[13]) );
  HAX1 U1_1_12 ( .A(A[12]), .B(carry[12]), .YC(carry[13]), .YS(SUM[12]) );
  HAX1 U1_1_11 ( .A(A[11]), .B(carry[11]), .YC(carry[12]), .YS(SUM[11]) );
  HAX1 U1_1_10 ( .A(A[10]), .B(carry[10]), .YC(carry[11]), .YS(SUM[10]) );
  HAX1 U1_1_9 ( .A(A[9]), .B(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  HAX1 U1_1_8 ( .A(A[8]), .B(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  HAX1 U1_1_7 ( .A(A[7]), .B(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  HAX1 U1_1_6 ( .A(A[6]), .B(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  HAX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry[2]), .YS(SUM[1]) );
  XOR2X1 U1 ( .A(carry[31]), .B(A[31]), .Y(SUM[31]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module Processing_logic_DW01_inc_1 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;
  wire   n1;
  wire   [31:2] carry;

  HAX1 U1_1_30 ( .A(A[30]), .B(carry[30]), .YC(carry[31]), .YS(SUM[30]) );
  HAX1 U1_1_29 ( .A(A[29]), .B(carry[29]), .YC(carry[30]), .YS(SUM[29]) );
  HAX1 U1_1_28 ( .A(A[28]), .B(carry[28]), .YC(carry[29]), .YS(SUM[28]) );
  HAX1 U1_1_27 ( .A(A[27]), .B(carry[27]), .YC(carry[28]), .YS(SUM[27]) );
  HAX1 U1_1_26 ( .A(A[26]), .B(carry[26]), .YC(carry[27]), .YS(SUM[26]) );
  HAX1 U1_1_25 ( .A(A[25]), .B(carry[25]), .YC(carry[26]), .YS(SUM[25]) );
  HAX1 U1_1_24 ( .A(A[24]), .B(carry[24]), .YC(carry[25]), .YS(SUM[24]) );
  HAX1 U1_1_23 ( .A(A[23]), .B(carry[23]), .YC(carry[24]), .YS(SUM[23]) );
  HAX1 U1_1_22 ( .A(A[22]), .B(carry[22]), .YC(carry[23]), .YS(SUM[22]) );
  HAX1 U1_1_21 ( .A(A[21]), .B(carry[21]), .YC(carry[22]), .YS(SUM[21]) );
  HAX1 U1_1_20 ( .A(A[20]), .B(carry[20]), .YC(carry[21]), .YS(SUM[20]) );
  HAX1 U1_1_19 ( .A(A[19]), .B(carry[19]), .YC(carry[20]), .YS(SUM[19]) );
  HAX1 U1_1_18 ( .A(A[18]), .B(carry[18]), .YC(carry[19]), .YS(SUM[18]) );
  HAX1 U1_1_17 ( .A(A[17]), .B(carry[17]), .YC(carry[18]), .YS(SUM[17]) );
  HAX1 U1_1_16 ( .A(A[16]), .B(carry[16]), .YC(carry[17]), .YS(SUM[16]) );
  HAX1 U1_1_15 ( .A(A[15]), .B(carry[15]), .YC(carry[16]), .YS(SUM[15]) );
  HAX1 U1_1_14 ( .A(A[14]), .B(carry[14]), .YC(carry[15]), .YS(SUM[14]) );
  HAX1 U1_1_13 ( .A(A[13]), .B(carry[13]), .YC(carry[14]), .YS(SUM[13]) );
  HAX1 U1_1_12 ( .A(A[12]), .B(carry[12]), .YC(carry[13]), .YS(SUM[12]) );
  HAX1 U1_1_11 ( .A(A[11]), .B(carry[11]), .YC(carry[12]), .YS(SUM[11]) );
  HAX1 U1_1_10 ( .A(A[10]), .B(carry[10]), .YC(carry[11]), .YS(SUM[10]) );
  HAX1 U1_1_9 ( .A(A[9]), .B(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  HAX1 U1_1_8 ( .A(A[8]), .B(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  HAX1 U1_1_7 ( .A(A[7]), .B(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  HAX1 U1_1_6 ( .A(A[6]), .B(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  HAX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(n1), .YC(carry[2]), .YS(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  INVX8 U2 ( .A(SUM[0]), .Y(n1) );
  XOR2X1 U3 ( .A(carry[31]), .B(A[31]), .Y(SUM[31]) );
endmodule


module Processing_logic_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   carry_31_, carry_29_, carry_27_, carry_24_, carry_22_, carry_21_,
         carry_19_, carry_17_, carry_16_, carry_14_, carry_13_, carry_11_, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39;

  OR2X2 U1 ( .A(A[10]), .B(n27), .Y(n28) );
  INVX1 U2 ( .A(n28), .Y(n1) );
  OR2X2 U3 ( .A(A[12]), .B(n17), .Y(n29) );
  INVX1 U4 ( .A(n29), .Y(n2) );
  OR2X2 U5 ( .A(A[13]), .B(carry_13_), .Y(n30) );
  INVX1 U6 ( .A(n30), .Y(n3) );
  OR2X2 U7 ( .A(A[15]), .B(n18), .Y(n31) );
  INVX1 U8 ( .A(n31), .Y(n4) );
  OR2X2 U9 ( .A(A[16]), .B(carry_16_), .Y(n32) );
  INVX1 U10 ( .A(n32), .Y(n5) );
  OR2X2 U11 ( .A(A[18]), .B(n19), .Y(n33) );
  INVX1 U12 ( .A(n33), .Y(n6) );
  OR2X2 U13 ( .A(A[20]), .B(n20), .Y(n34) );
  INVX1 U14 ( .A(n34), .Y(n7) );
  OR2X2 U15 ( .A(A[21]), .B(carry_21_), .Y(n35) );
  INVX1 U16 ( .A(n35), .Y(n8) );
  OR2X2 U17 ( .A(A[23]), .B(n21), .Y(n36) );
  INVX1 U18 ( .A(n36), .Y(n9) );
  OR2X2 U19 ( .A(A[26]), .B(n22), .Y(n37) );
  INVX1 U20 ( .A(n37), .Y(n10) );
  OR2X2 U21 ( .A(A[28]), .B(n23), .Y(n38) );
  INVX1 U22 ( .A(n38), .Y(n11) );
  OR2X2 U23 ( .A(A[30]), .B(n14), .Y(n39) );
  INVX1 U24 ( .A(n39), .Y(n12) );
  OR2X1 U25 ( .A(A[24]), .B(carry_24_), .Y(n13) );
  OR2X1 U26 ( .A(A[29]), .B(carry_29_), .Y(n14) );
  OR2X1 U27 ( .A(A[5]), .B(n24), .Y(n15) );
  OR2X2 U28 ( .A(A[6]), .B(n15), .Y(n16) );
  INVX1 U29 ( .A(n1), .Y(carry_11_) );
  OR2X2 U30 ( .A(A[11]), .B(carry_11_), .Y(n17) );
  INVX1 U31 ( .A(n3), .Y(carry_14_) );
  INVX1 U32 ( .A(n2), .Y(carry_13_) );
  OR2X2 U33 ( .A(A[14]), .B(carry_14_), .Y(n18) );
  INVX1 U34 ( .A(n5), .Y(carry_17_) );
  INVX1 U35 ( .A(n4), .Y(carry_16_) );
  OR2X2 U36 ( .A(A[17]), .B(carry_17_), .Y(n19) );
  INVX1 U37 ( .A(n6), .Y(carry_19_) );
  OR2X2 U38 ( .A(A[19]), .B(carry_19_), .Y(n20) );
  INVX1 U39 ( .A(n8), .Y(carry_22_) );
  INVX1 U40 ( .A(n7), .Y(carry_21_) );
  OR2X2 U41 ( .A(A[22]), .B(carry_22_), .Y(n21) );
  INVX1 U42 ( .A(n9), .Y(carry_24_) );
  OR2X2 U43 ( .A(A[25]), .B(n13), .Y(n22) );
  INVX1 U44 ( .A(n10), .Y(carry_27_) );
  OR2X2 U45 ( .A(A[27]), .B(carry_27_), .Y(n23) );
  INVX1 U46 ( .A(n11), .Y(carry_29_) );
  OR2X2 U47 ( .A(A[4]), .B(A[3]), .Y(n24) );
  OR2X2 U48 ( .A(A[7]), .B(n16), .Y(n25) );
  OR2X2 U49 ( .A(A[8]), .B(n25), .Y(n26) );
  OR2X2 U50 ( .A(A[9]), .B(n26), .Y(n27) );
  INVX1 U51 ( .A(n12), .Y(carry_31_) );
  XNOR2X1 U52 ( .A(n27), .B(A[10]), .Y(DIFF[10]) );
  XNOR2X1 U53 ( .A(carry_11_), .B(A[11]), .Y(DIFF[11]) );
  XNOR2X1 U54 ( .A(n17), .B(A[12]), .Y(DIFF[12]) );
  XNOR2X1 U55 ( .A(carry_13_), .B(A[13]), .Y(DIFF[13]) );
  XNOR2X1 U56 ( .A(carry_14_), .B(A[14]), .Y(DIFF[14]) );
  XNOR2X1 U57 ( .A(n18), .B(A[15]), .Y(DIFF[15]) );
  XNOR2X1 U58 ( .A(carry_16_), .B(A[16]), .Y(DIFF[16]) );
  XNOR2X1 U59 ( .A(carry_17_), .B(A[17]), .Y(DIFF[17]) );
  XNOR2X1 U60 ( .A(n19), .B(A[18]), .Y(DIFF[18]) );
  XNOR2X1 U61 ( .A(carry_19_), .B(A[19]), .Y(DIFF[19]) );
  XNOR2X1 U62 ( .A(n20), .B(A[20]), .Y(DIFF[20]) );
  XNOR2X1 U63 ( .A(carry_21_), .B(A[21]), .Y(DIFF[21]) );
  XNOR2X1 U64 ( .A(carry_22_), .B(A[22]), .Y(DIFF[22]) );
  XNOR2X1 U65 ( .A(n21), .B(A[23]), .Y(DIFF[23]) );
  XNOR2X1 U66 ( .A(carry_24_), .B(A[24]), .Y(DIFF[24]) );
  XNOR2X1 U67 ( .A(n13), .B(A[25]), .Y(DIFF[25]) );
  XNOR2X1 U68 ( .A(n22), .B(A[26]), .Y(DIFF[26]) );
  XNOR2X1 U69 ( .A(carry_27_), .B(A[27]), .Y(DIFF[27]) );
  XNOR2X1 U70 ( .A(n23), .B(A[28]), .Y(DIFF[28]) );
  XNOR2X1 U71 ( .A(carry_29_), .B(A[29]), .Y(DIFF[29]) );
  XNOR2X1 U72 ( .A(n14), .B(A[30]), .Y(DIFF[30]) );
  XNOR2X1 U73 ( .A(A[31]), .B(carry_31_), .Y(DIFF[31]) );
  XNOR2X1 U74 ( .A(A[3]), .B(A[4]), .Y(DIFF[4]) );
  XNOR2X1 U75 ( .A(n24), .B(A[5]), .Y(DIFF[5]) );
  XNOR2X1 U76 ( .A(n15), .B(A[6]), .Y(DIFF[6]) );
  XNOR2X1 U77 ( .A(n16), .B(A[7]), .Y(DIFF[7]) );
  XNOR2X1 U78 ( .A(n25), .B(A[8]), .Y(DIFF[8]) );
  XNOR2X1 U79 ( .A(n26), .B(A[9]), .Y(DIFF[9]) );
  INVX2 U80 ( .A(A[3]), .Y(DIFF[3]) );
endmodule


module Processing_logic_DW01_cmp6_1 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330;

  NOR3X1 U1 ( .A(n4), .B(n2), .C(n3), .Y(n1) );
  INVX8 U2 ( .A(n194), .Y(n2) );
  INVX8 U3 ( .A(n191), .Y(n3) );
  INVX1 U4 ( .A(n269), .Y(n4) );
  NOR3X1 U5 ( .A(n7), .B(n6), .C(n155), .Y(n5) );
  INVX8 U6 ( .A(n295), .Y(n6) );
  INVX1 U7 ( .A(n296), .Y(n7) );
  NOR3X1 U8 ( .A(n9), .B(n10), .C(n11), .Y(n8) );
  INVX2 U9 ( .A(n8), .Y(n320) );
  INVX8 U10 ( .A(n253), .Y(n9) );
  INVX8 U11 ( .A(n256), .Y(n10) );
  INVX1 U12 ( .A(n321), .Y(n11) );
  NOR3X1 U13 ( .A(n13), .B(n112), .C(n14), .Y(n12) );
  INVX1 U14 ( .A(n12), .Y(n211) );
  INVX8 U15 ( .A(n216), .Y(n13) );
  INVX1 U16 ( .A(n214), .Y(n14) );
  NOR3X1 U17 ( .A(n16), .B(n143), .C(n17), .Y(n15) );
  INVX8 U18 ( .A(n242), .Y(n16) );
  INVX1 U19 ( .A(n240), .Y(n17) );
  INVX1 U20 ( .A(n48), .Y(n195) );
  NOR3X1 U21 ( .A(n19), .B(n97), .C(n45), .Y(n18) );
  INVX2 U22 ( .A(n18), .Y(n184) );
  INVX8 U23 ( .A(n188), .Y(n19) );
  INVX1 U24 ( .A(n25), .Y(n203) );
  INVX1 U25 ( .A(n20), .Y(n262) );
  INVX1 U26 ( .A(n27), .Y(n82) );
  NOR3X1 U27 ( .A(n91), .B(n94), .C(n21), .Y(n20) );
  INVX1 U28 ( .A(n264), .Y(n21) );
  NOR3X1 U29 ( .A(n23), .B(n109), .C(n24), .Y(n22) );
  INVX8 U30 ( .A(n210), .Y(n23) );
  INVX1 U31 ( .A(n208), .Y(n24) );
  NOR3X1 U32 ( .A(n26), .B(n161), .C(n22), .Y(n25) );
  INVX8 U33 ( .A(n207), .Y(n26) );
  NOR3X1 U34 ( .A(n30), .B(n28), .C(n29), .Y(n27) );
  INVX8 U35 ( .A(n239), .Y(n28) );
  INVX8 U36 ( .A(n237), .Y(n29) );
  INVX1 U37 ( .A(n306), .Y(n30) );
  INVX1 U38 ( .A(A[1]), .Y(n176) );
  INVX1 U39 ( .A(n31), .Y(n265) );
  NOR3X1 U40 ( .A(n32), .B(n33), .C(n1), .Y(n31) );
  INVX8 U41 ( .A(n174), .Y(n32) );
  INVX8 U42 ( .A(n268), .Y(n33) );
  INVX1 U43 ( .A(n43), .Y(n235) );
  NOR3X1 U44 ( .A(n35), .B(n164), .C(n36), .Y(n34) );
  INVX8 U45 ( .A(n202), .Y(n35) );
  INVX1 U46 ( .A(n200), .Y(n36) );
  NOR3X1 U47 ( .A(n39), .B(n38), .C(n5), .Y(n37) );
  INVX8 U48 ( .A(n222), .Y(n38) );
  INVX8 U49 ( .A(n219), .Y(n39) );
  INVX1 U50 ( .A(A[0]), .Y(n177) );
  INVX1 U51 ( .A(n40), .Y(n289) );
  NOR3X1 U52 ( .A(n41), .B(n42), .C(n37), .Y(n40) );
  INVX8 U53 ( .A(n159), .Y(n41) );
  INVX8 U54 ( .A(n292), .Y(n42) );
  NOR3X1 U55 ( .A(n44), .B(n124), .C(n15), .Y(n43) );
  INVX8 U56 ( .A(n239), .Y(n44) );
  NOR3X1 U57 ( .A(n47), .B(n170), .C(n46), .Y(n45) );
  INVX8 U58 ( .A(n191), .Y(n46) );
  INVX1 U59 ( .A(n189), .Y(n47) );
  NOR3X1 U60 ( .A(n49), .B(n103), .C(n34), .Y(n48) );
  INVX8 U61 ( .A(n199), .Y(n49) );
  AND2X2 U62 ( .A(n319), .B(n131), .Y(n253) );
  AND2X2 U63 ( .A(n180), .B(n95), .Y(n179) );
  OR2X2 U64 ( .A(n323), .B(A[5]), .Y(n256) );
  AND2X2 U65 ( .A(A[5]), .B(n323), .Y(n252) );
  OR2X2 U66 ( .A(n327), .B(B[4]), .Y(n324) );
  OR2X2 U67 ( .A(n76), .B(n77), .Y(n79) );
  AND2X2 U68 ( .A(B[4]), .B(n327), .Y(n255) );
  AND2X2 U69 ( .A(n324), .B(n133), .Y(n259) );
  OR2X2 U70 ( .A(n78), .B(n79), .Y(n75) );
  AND2X2 U71 ( .A(n177), .B(n176), .Y(n330) );
  INVX1 U72 ( .A(n330), .Y(n50) );
  BUFX2 U73 ( .A(n183), .Y(n51) );
  BUFX2 U74 ( .A(n192), .Y(n52) );
  BUFX2 U75 ( .A(n217), .Y(n53) );
  BUFX2 U76 ( .A(n220), .Y(n54) );
  BUFX2 U77 ( .A(n223), .Y(n55) );
  BUFX2 U78 ( .A(n226), .Y(n56) );
  BUFX2 U79 ( .A(n229), .Y(n57) );
  BUFX2 U80 ( .A(n232), .Y(n58) );
  BUFX2 U81 ( .A(n243), .Y(n59) );
  BUFX2 U82 ( .A(n246), .Y(n60) );
  BUFX2 U83 ( .A(n249), .Y(n61) );
  BUFX2 U84 ( .A(n274), .Y(n62) );
  BUFX2 U85 ( .A(n279), .Y(n63) );
  BUFX2 U86 ( .A(n284), .Y(n64) );
  BUFX2 U87 ( .A(n297), .Y(n65) );
  BUFX2 U88 ( .A(n302), .Y(n66) );
  BUFX2 U89 ( .A(n311), .Y(n67) );
  BUFX2 U90 ( .A(n316), .Y(n68) );
  BUFX2 U91 ( .A(n326), .Y(n69) );
  BUFX2 U92 ( .A(n273), .Y(n70) );
  BUFX2 U93 ( .A(n278), .Y(n71) );
  BUFX2 U94 ( .A(n283), .Y(n72) );
  BUFX2 U95 ( .A(n288), .Y(n73) );
  INVX1 U96 ( .A(n179), .Y(n74) );
  INVX1 U97 ( .A(n256), .Y(n76) );
  INVX1 U98 ( .A(n133), .Y(n77) );
  INVX1 U99 ( .A(n254), .Y(n78) );
  INVX1 U100 ( .A(n301), .Y(n80) );
  INVX1 U101 ( .A(n80), .Y(n81) );
  INVX1 U102 ( .A(n310), .Y(n83) );
  INVX1 U103 ( .A(n83), .Y(n84) );
  INVX1 U104 ( .A(n315), .Y(n85) );
  INVX1 U105 ( .A(n85), .Y(n86) );
  BUFX2 U106 ( .A(n325), .Y(n87) );
  INVX1 U107 ( .A(n90), .Y(n88) );
  INVX1 U108 ( .A(n88), .Y(n89) );
  AND2X2 U109 ( .A(n50), .B(n261), .Y(n329) );
  INVX1 U110 ( .A(n329), .Y(n90) );
  INVX1 U111 ( .A(n93), .Y(n91) );
  INVX1 U112 ( .A(n91), .Y(n92) );
  AND2X1 U113 ( .A(A[30]), .B(n182), .Y(n263) );
  INVX1 U114 ( .A(n263), .Y(n93) );
  INVX1 U115 ( .A(n96), .Y(n94) );
  INVX1 U116 ( .A(n94), .Y(n95) );
  AND2X1 U117 ( .A(B[31]), .B(n178), .Y(n181) );
  INVX1 U118 ( .A(n181), .Y(n96) );
  INVX1 U119 ( .A(n99), .Y(n97) );
  INVX1 U120 ( .A(n97), .Y(n98) );
  AND2X1 U121 ( .A(B[28]), .B(n270), .Y(n187) );
  INVX1 U122 ( .A(n187), .Y(n99) );
  INVX1 U123 ( .A(n102), .Y(n100) );
  INVX1 U124 ( .A(n100), .Y(n101) );
  AND2X1 U125 ( .A(B[26]), .B(n275), .Y(n193) );
  INVX1 U126 ( .A(n193), .Y(n102) );
  INVX1 U127 ( .A(n105), .Y(n103) );
  INVX1 U128 ( .A(n103), .Y(n104) );
  AND2X1 U129 ( .A(B[24]), .B(n280), .Y(n198) );
  INVX1 U130 ( .A(n198), .Y(n105) );
  INVX1 U131 ( .A(n108), .Y(n106) );
  INVX1 U132 ( .A(n106), .Y(n107) );
  AND2X1 U133 ( .A(B[22]), .B(n285), .Y(n204) );
  INVX1 U134 ( .A(n204), .Y(n108) );
  INVX1 U135 ( .A(n111), .Y(n109) );
  INVX1 U136 ( .A(n109), .Y(n110) );
  AND2X1 U137 ( .A(B[20]), .B(n290), .Y(n209) );
  INVX1 U138 ( .A(n209), .Y(n111) );
  INVX1 U139 ( .A(n114), .Y(n112) );
  INVX1 U140 ( .A(n112), .Y(n113) );
  AND2X1 U141 ( .A(B[18]), .B(n293), .Y(n215) );
  INVX1 U142 ( .A(n215), .Y(n114) );
  INVX1 U143 ( .A(n117), .Y(n115) );
  INVX1 U144 ( .A(n115), .Y(n116) );
  AND2X1 U145 ( .A(B[16]), .B(n298), .Y(n221) );
  INVX1 U146 ( .A(n221), .Y(n117) );
  INVX1 U147 ( .A(n120), .Y(n118) );
  INVX1 U148 ( .A(n118), .Y(n119) );
  AND2X1 U149 ( .A(B[14]), .B(n303), .Y(n227) );
  INVX1 U150 ( .A(n227), .Y(n120) );
  INVX1 U151 ( .A(n123), .Y(n121) );
  INVX1 U152 ( .A(n121), .Y(n122) );
  AND2X1 U153 ( .A(B[12]), .B(n307), .Y(n233) );
  INVX1 U154 ( .A(n233), .Y(n123) );
  INVX1 U155 ( .A(n126), .Y(n124) );
  INVX1 U156 ( .A(n124), .Y(n125) );
  AND2X1 U157 ( .A(B[10]), .B(n312), .Y(n238) );
  INVX1 U158 ( .A(n238), .Y(n126) );
  INVX1 U159 ( .A(n129), .Y(n127) );
  INVX1 U160 ( .A(n127), .Y(n128) );
  AND2X1 U161 ( .A(B[8]), .B(n317), .Y(n244) );
  INVX1 U162 ( .A(n244), .Y(n129) );
  INVX1 U163 ( .A(n132), .Y(n130) );
  INVX1 U164 ( .A(n130), .Y(n131) );
  AND2X1 U165 ( .A(B[6]), .B(n322), .Y(n250) );
  INVX1 U166 ( .A(n250), .Y(n132) );
  INVX1 U167 ( .A(n255), .Y(n133) );
  INVX1 U168 ( .A(n136), .Y(n134) );
  INVX1 U169 ( .A(n134), .Y(n135) );
  AND2X1 U170 ( .A(A[3]), .B(n328), .Y(n258) );
  INVX1 U171 ( .A(n258), .Y(n136) );
  INVX1 U172 ( .A(n139), .Y(n137) );
  INVX1 U173 ( .A(n137), .Y(n138) );
  INVX1 U174 ( .A(n252), .Y(n139) );
  INVX1 U175 ( .A(n142), .Y(n140) );
  INVX1 U176 ( .A(n140), .Y(n141) );
  AND2X1 U177 ( .A(A[7]), .B(n318), .Y(n247) );
  INVX1 U178 ( .A(n247), .Y(n142) );
  INVX1 U179 ( .A(n145), .Y(n143) );
  INVX1 U180 ( .A(n143), .Y(n144) );
  AND2X1 U181 ( .A(A[9]), .B(n313), .Y(n241) );
  INVX1 U182 ( .A(n241), .Y(n145) );
  INVX1 U183 ( .A(n148), .Y(n146) );
  INVX1 U184 ( .A(n146), .Y(n147) );
  AND2X1 U185 ( .A(A[11]), .B(n308), .Y(n236) );
  INVX1 U186 ( .A(n236), .Y(n148) );
  INVX1 U187 ( .A(n151), .Y(n149) );
  INVX1 U188 ( .A(n149), .Y(n150) );
  AND2X1 U189 ( .A(A[13]), .B(n304), .Y(n230) );
  INVX1 U190 ( .A(n230), .Y(n151) );
  INVX1 U191 ( .A(n154), .Y(n152) );
  INVX1 U192 ( .A(n152), .Y(n153) );
  AND2X1 U193 ( .A(A[15]), .B(n299), .Y(n224) );
  INVX1 U194 ( .A(n224), .Y(n154) );
  INVX1 U195 ( .A(n157), .Y(n155) );
  INVX1 U196 ( .A(n155), .Y(n156) );
  AND2X1 U197 ( .A(A[17]), .B(n294), .Y(n218) );
  INVX1 U198 ( .A(n218), .Y(n157) );
  INVX1 U199 ( .A(n160), .Y(n158) );
  INVX1 U200 ( .A(n158), .Y(n159) );
  AND2X1 U201 ( .A(A[19]), .B(n291), .Y(n212) );
  INVX1 U202 ( .A(n212), .Y(n160) );
  INVX1 U203 ( .A(n163), .Y(n161) );
  INVX1 U204 ( .A(n161), .Y(n162) );
  AND2X1 U205 ( .A(A[21]), .B(n286), .Y(n206) );
  INVX1 U206 ( .A(n206), .Y(n163) );
  INVX1 U207 ( .A(n166), .Y(n164) );
  INVX1 U208 ( .A(n164), .Y(n165) );
  AND2X1 U209 ( .A(A[23]), .B(n281), .Y(n201) );
  INVX1 U210 ( .A(n201), .Y(n166) );
  INVX1 U211 ( .A(n169), .Y(n167) );
  INVX1 U212 ( .A(n167), .Y(n168) );
  AND2X1 U213 ( .A(A[25]), .B(n276), .Y(n196) );
  INVX1 U214 ( .A(n196), .Y(n169) );
  INVX1 U215 ( .A(n172), .Y(n170) );
  INVX1 U216 ( .A(n170), .Y(n171) );
  AND2X1 U217 ( .A(A[27]), .B(n271), .Y(n190) );
  INVX1 U218 ( .A(n190), .Y(n172) );
  INVX1 U219 ( .A(n175), .Y(n173) );
  INVX1 U220 ( .A(n173), .Y(n174) );
  AND2X1 U221 ( .A(A[29]), .B(n267), .Y(n185) );
  INVX1 U222 ( .A(n185), .Y(n175) );
  INVX2 U223 ( .A(n260), .Y(n257) );
  OAI21X1 U224 ( .A(B[31]), .B(n178), .C(n74), .Y(LT) );
  OAI21X1 U225 ( .A(A[30]), .B(n182), .C(n51), .Y(n180) );
  NAND3X1 U226 ( .A(n186), .B(n174), .C(n184), .Y(n183) );
  NAND3X1 U227 ( .A(n194), .B(n101), .C(n52), .Y(n189) );
  NAND3X1 U228 ( .A(n195), .B(n168), .C(n197), .Y(n192) );
  NAND3X1 U229 ( .A(n205), .B(n107), .C(n203), .Y(n200) );
  NAND3X1 U230 ( .A(n213), .B(n159), .C(n211), .Y(n208) );
  NAND3X1 U231 ( .A(n219), .B(n156), .C(n53), .Y(n214) );
  NAND3X1 U232 ( .A(n222), .B(n116), .C(n54), .Y(n217) );
  NAND3X1 U233 ( .A(n225), .B(n153), .C(n55), .Y(n220) );
  NAND3X1 U234 ( .A(n228), .B(n119), .C(n56), .Y(n223) );
  NAND3X1 U235 ( .A(n57), .B(n150), .C(n231), .Y(n226) );
  NAND3X1 U236 ( .A(n234), .B(n122), .C(n58), .Y(n229) );
  NAND3X1 U237 ( .A(n237), .B(n147), .C(n235), .Y(n232) );
  NAND3X1 U238 ( .A(n245), .B(n128), .C(n59), .Y(n240) );
  NAND3X1 U239 ( .A(n60), .B(n141), .C(n248), .Y(n243) );
  NAND3X1 U240 ( .A(n61), .B(n131), .C(n251), .Y(n246) );
  NAND3X1 U241 ( .A(n138), .B(n253), .C(n75), .Y(n249) );
  NAND3X1 U242 ( .A(n257), .B(n135), .C(n259), .Y(n254) );
  OAI21X1 U243 ( .A(B[31]), .B(n178), .C(n262), .Y(LE) );
  NAND3X1 U244 ( .A(n265), .B(n188), .C(n186), .Y(n264) );
  INVX1 U245 ( .A(n266), .Y(n186) );
  OAI21X1 U246 ( .A(A[30]), .B(n182), .C(n92), .Y(n266) );
  OR2X1 U247 ( .A(n267), .B(A[29]), .Y(n188) );
  AND2X1 U248 ( .A(n268), .B(n98), .Y(n191) );
  OR2X1 U249 ( .A(n271), .B(A[27]), .Y(n194) );
  NAND3X1 U250 ( .A(n171), .B(n272), .C(n70), .Y(n269) );
  NAND3X1 U251 ( .A(n62), .B(n199), .C(n197), .Y(n273) );
  AND2X1 U252 ( .A(n272), .B(n101), .Y(n197) );
  OR2X1 U253 ( .A(n276), .B(A[25]), .Y(n199) );
  NAND3X1 U254 ( .A(n168), .B(n277), .C(n71), .Y(n274) );
  NAND3X1 U255 ( .A(n63), .B(n205), .C(n202), .Y(n278) );
  AND2X1 U256 ( .A(n277), .B(n104), .Y(n202) );
  OR2X1 U257 ( .A(n281), .B(A[23]), .Y(n205) );
  NAND3X1 U258 ( .A(n165), .B(n282), .C(n72), .Y(n279) );
  NAND3X1 U259 ( .A(n64), .B(n210), .C(n207), .Y(n283) );
  AND2X1 U260 ( .A(n282), .B(n107), .Y(n207) );
  OR2X1 U261 ( .A(n286), .B(A[21]), .Y(n210) );
  NAND3X1 U262 ( .A(n162), .B(n287), .C(n73), .Y(n284) );
  NAND3X1 U263 ( .A(n289), .B(n216), .C(n213), .Y(n288) );
  AND2X1 U264 ( .A(n287), .B(n110), .Y(n213) );
  OR2X1 U265 ( .A(n291), .B(A[19]), .Y(n216) );
  AND2X1 U266 ( .A(n292), .B(n113), .Y(n219) );
  OR2X1 U267 ( .A(n294), .B(A[17]), .Y(n222) );
  NAND3X1 U268 ( .A(n65), .B(n228), .C(n225), .Y(n296) );
  AND2X1 U269 ( .A(n295), .B(n116), .Y(n225) );
  OR2X1 U270 ( .A(n299), .B(A[15]), .Y(n228) );
  NAND3X1 U271 ( .A(n153), .B(n300), .C(n81), .Y(n297) );
  NAND3X1 U272 ( .A(n231), .B(n234), .C(n66), .Y(n301) );
  AND2X1 U273 ( .A(n300), .B(n119), .Y(n231) );
  OR2X1 U274 ( .A(n304), .B(A[13]), .Y(n234) );
  NAND3X1 U275 ( .A(n150), .B(n305), .C(n82), .Y(n302) );
  AND2X1 U276 ( .A(n305), .B(n122), .Y(n237) );
  OR2X1 U277 ( .A(n308), .B(A[11]), .Y(n239) );
  NAND3X1 U278 ( .A(n147), .B(n309), .C(n84), .Y(n306) );
  NAND3X1 U279 ( .A(n67), .B(n245), .C(n242), .Y(n310) );
  AND2X1 U280 ( .A(n309), .B(n125), .Y(n242) );
  OR2X1 U281 ( .A(n313), .B(A[9]), .Y(n245) );
  NAND3X1 U282 ( .A(n144), .B(n314), .C(n86), .Y(n311) );
  NAND3X1 U283 ( .A(n248), .B(n251), .C(n68), .Y(n315) );
  AND2X1 U284 ( .A(n314), .B(n128), .Y(n248) );
  OR2X1 U285 ( .A(n318), .B(A[7]), .Y(n251) );
  NAND3X1 U286 ( .A(n141), .B(n319), .C(n320), .Y(n316) );
  NAND3X1 U287 ( .A(n138), .B(n324), .C(n87), .Y(n321) );
  NAND3X1 U288 ( .A(n69), .B(n260), .C(n259), .Y(n325) );
  OR2X1 U289 ( .A(n328), .B(A[3]), .Y(n260) );
  NAND3X1 U290 ( .A(n135), .B(n261), .C(n89), .Y(n326) );
  INVX1 U291 ( .A(A[2]), .Y(n261) );
  INVX1 U292 ( .A(B[3]), .Y(n328) );
  INVX1 U293 ( .A(A[4]), .Y(n327) );
  INVX1 U294 ( .A(B[5]), .Y(n323) );
  OR2X1 U295 ( .A(n322), .B(B[6]), .Y(n319) );
  INVX1 U296 ( .A(A[6]), .Y(n322) );
  INVX1 U297 ( .A(B[7]), .Y(n318) );
  OR2X1 U298 ( .A(n317), .B(B[8]), .Y(n314) );
  INVX1 U299 ( .A(A[8]), .Y(n317) );
  INVX1 U300 ( .A(B[9]), .Y(n313) );
  OR2X1 U301 ( .A(n312), .B(B[10]), .Y(n309) );
  INVX1 U302 ( .A(A[10]), .Y(n312) );
  INVX1 U303 ( .A(B[11]), .Y(n308) );
  OR2X1 U304 ( .A(n307), .B(B[12]), .Y(n305) );
  INVX1 U305 ( .A(A[12]), .Y(n307) );
  INVX1 U306 ( .A(B[13]), .Y(n304) );
  OR2X1 U307 ( .A(n303), .B(B[14]), .Y(n300) );
  INVX1 U308 ( .A(A[14]), .Y(n303) );
  INVX1 U309 ( .A(B[15]), .Y(n299) );
  OR2X1 U310 ( .A(n298), .B(B[16]), .Y(n295) );
  INVX1 U311 ( .A(A[16]), .Y(n298) );
  INVX1 U312 ( .A(B[17]), .Y(n294) );
  OR2X1 U313 ( .A(n293), .B(B[18]), .Y(n292) );
  INVX1 U314 ( .A(A[18]), .Y(n293) );
  INVX1 U315 ( .A(B[19]), .Y(n291) );
  OR2X1 U316 ( .A(n290), .B(B[20]), .Y(n287) );
  INVX1 U317 ( .A(A[20]), .Y(n290) );
  INVX1 U318 ( .A(B[21]), .Y(n286) );
  OR2X1 U319 ( .A(n285), .B(B[22]), .Y(n282) );
  INVX1 U320 ( .A(A[22]), .Y(n285) );
  INVX1 U321 ( .A(B[23]), .Y(n281) );
  OR2X1 U322 ( .A(n280), .B(B[24]), .Y(n277) );
  INVX1 U323 ( .A(A[24]), .Y(n280) );
  INVX1 U324 ( .A(B[25]), .Y(n276) );
  OR2X1 U325 ( .A(n275), .B(B[26]), .Y(n272) );
  INVX1 U326 ( .A(A[26]), .Y(n275) );
  INVX1 U327 ( .A(B[27]), .Y(n271) );
  OR2X1 U328 ( .A(n270), .B(B[28]), .Y(n268) );
  INVX1 U329 ( .A(A[28]), .Y(n270) );
  INVX1 U330 ( .A(B[29]), .Y(n267) );
  INVX1 U331 ( .A(B[30]), .Y(n182) );
  INVX1 U332 ( .A(A[31]), .Y(n178) );
endmodule


module Processing_logic_DW01_dec_0 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138;

  XOR2X1 U1 ( .A(n71), .B(n4), .Y(SUM[30]) );
  AND2X2 U2 ( .A(n2), .B(n3), .Y(n39) );
  INVX1 U3 ( .A(n72), .Y(n1) );
  AND2X1 U4 ( .A(n83), .B(n79), .Y(n2) );
  AND2X1 U5 ( .A(n138), .B(n76), .Y(n3) );
  INVX8 U6 ( .A(A[30]), .Y(n4) );
  AND2X2 U7 ( .A(n97), .B(n7), .Y(n5) );
  AND2X1 U8 ( .A(n97), .B(n8), .Y(n6) );
  INVX1 U9 ( .A(A[27]), .Y(n8) );
  AND2X2 U10 ( .A(n101), .B(n8), .Y(n7) );
  OR2X2 U11 ( .A(n15), .B(A[11]), .Y(n68) );
  OR2X2 U12 ( .A(A[29]), .B(n27), .Y(n71) );
  OR2X2 U13 ( .A(A[16]), .B(n54), .Y(n72) );
  INVX1 U14 ( .A(n72), .Y(n9) );
  OR2X2 U15 ( .A(n14), .B(A[18]), .Y(n73) );
  AND2X2 U16 ( .A(n66), .B(n119), .Y(n118) );
  AND2X2 U17 ( .A(n129), .B(n128), .Y(n127) );
  AND2X2 U18 ( .A(n32), .B(n130), .Y(n129) );
  AND2X2 U19 ( .A(n64), .B(n133), .Y(n132) );
  AND2X2 U20 ( .A(n76), .B(n80), .Y(n77) );
  INVX1 U21 ( .A(n77), .Y(n10) );
  AND2X2 U22 ( .A(n79), .B(n83), .Y(n80) );
  AND2X2 U23 ( .A(n82), .B(n86), .Y(n83) );
  INVX1 U24 ( .A(n83), .Y(n11) );
  AND2X2 U25 ( .A(n85), .B(n84), .Y(n86) );
  INVX1 U26 ( .A(n86), .Y(n12) );
  AND2X2 U27 ( .A(n87), .B(n22), .Y(n88) );
  INVX1 U28 ( .A(n88), .Y(n13) );
  INVX1 U29 ( .A(n38), .Y(n14) );
  INVX1 U30 ( .A(n39), .Y(n15) );
  OR2X2 U31 ( .A(n26), .B(A[25]), .Y(n70) );
  INVX1 U32 ( .A(n70), .Y(n16) );
  INVX1 U33 ( .A(n70), .Y(n17) );
  OR2X2 U34 ( .A(n30), .B(A[23]), .Y(n74) );
  INVX1 U35 ( .A(n74), .Y(n18) );
  INVX1 U36 ( .A(n74), .Y(n19) );
  OR2X2 U37 ( .A(n24), .B(A[21]), .Y(n75) );
  INVX1 U38 ( .A(n75), .Y(n20) );
  INVX1 U39 ( .A(n75), .Y(n21) );
  OR2X2 U40 ( .A(n92), .B(A[4]), .Y(n69) );
  INVX1 U41 ( .A(n69), .Y(n22) );
  INVX1 U42 ( .A(n69), .Y(n23) );
  AND2X2 U43 ( .A(n118), .B(n117), .Y(n116) );
  INVX1 U44 ( .A(n116), .Y(n24) );
  INVX1 U45 ( .A(n116), .Y(n25) );
  AND2X2 U46 ( .A(n107), .B(n18), .Y(n106) );
  INVX1 U47 ( .A(n106), .Y(n26) );
  AND2X2 U48 ( .A(n101), .B(n6), .Y(n96) );
  INVX1 U49 ( .A(n96), .Y(n27) );
  INVX1 U50 ( .A(n5), .Y(n28) );
  AND2X2 U51 ( .A(n102), .B(n16), .Y(n101) );
  INVX1 U52 ( .A(n101), .Y(n29) );
  AND2X2 U53 ( .A(n112), .B(n20), .Y(n111) );
  INVX1 U54 ( .A(n111), .Y(n30) );
  INVX1 U55 ( .A(n111), .Y(n31) );
  AND2X2 U56 ( .A(n131), .B(n132), .Y(n32) );
  BUFX2 U57 ( .A(n132), .Y(n33) );
  AND2X2 U58 ( .A(n123), .B(n1), .Y(n38) );
  INVX1 U59 ( .A(n38), .Y(n34) );
  INVX1 U60 ( .A(n39), .Y(n35) );
  INVX1 U61 ( .A(n12), .Y(n81) );
  INVX1 U62 ( .A(n118), .Y(n36) );
  INVX1 U63 ( .A(n137), .Y(n37) );
  INVX1 U64 ( .A(n129), .Y(n40) );
  INVX1 U65 ( .A(n32), .Y(n41) );
  INVX1 U66 ( .A(n33), .Y(n42) );
  INVX1 U67 ( .A(n80), .Y(n43) );
  INVX1 U68 ( .A(n78), .Y(n44) );
  INVX1 U69 ( .A(n11), .Y(n78) );
  INVX1 U70 ( .A(n81), .Y(n45) );
  INVX1 U71 ( .A(n84), .Y(n46) );
  INVX1 U72 ( .A(n13), .Y(n84) );
  INVX1 U73 ( .A(n104), .Y(n47) );
  BUFX2 U74 ( .A(n25), .Y(n48) );
  BUFX2 U75 ( .A(n34), .Y(n49) );
  BUFX2 U76 ( .A(n35), .Y(n50) );
  INVX1 U77 ( .A(n10), .Y(n137) );
  INVX1 U78 ( .A(n94), .Y(n51) );
  INVX1 U79 ( .A(n99), .Y(n52) );
  INVX1 U80 ( .A(n109), .Y(n53) );
  INVX1 U81 ( .A(n127), .Y(n54) );
  INVX1 U82 ( .A(n127), .Y(n55) );
  BUFX2 U83 ( .A(n23), .Y(n56) );
  INVX1 U84 ( .A(n103), .Y(n57) );
  INVX1 U85 ( .A(n98), .Y(n58) );
  INVX1 U86 ( .A(n9), .Y(n59) );
  INVX1 U87 ( .A(n59), .Y(n60) );
  INVX1 U88 ( .A(n108), .Y(n61) );
  INVX1 U89 ( .A(n21), .Y(n62) );
  INVX1 U90 ( .A(n62), .Y(n63) );
  INVX1 U91 ( .A(n68), .Y(n64) );
  INVX1 U92 ( .A(n68), .Y(n65) );
  INVX1 U93 ( .A(n73), .Y(n66) );
  INVX1 U94 ( .A(n73), .Y(n67) );
  INVX1 U95 ( .A(n65), .Y(n134) );
  INVX1 U96 ( .A(n50), .Y(n135) );
  INVX1 U97 ( .A(n56), .Y(n91) );
  INVX1 U98 ( .A(n17), .Y(n103) );
  INVX1 U99 ( .A(n26), .Y(n104) );
  INVX1 U100 ( .A(n7), .Y(n98) );
  INVX1 U101 ( .A(n29), .Y(n99) );
  INVX1 U102 ( .A(n28), .Y(n94) );
  INVX1 U103 ( .A(n60), .Y(n124) );
  INVX1 U104 ( .A(n55), .Y(n125) );
  INVX1 U105 ( .A(n67), .Y(n120) );
  INVX1 U106 ( .A(n49), .Y(n121) );
  INVX1 U107 ( .A(n19), .Y(n108) );
  INVX1 U108 ( .A(n31), .Y(n109) );
  INVX1 U109 ( .A(n63), .Y(n113) );
  INVX1 U110 ( .A(n48), .Y(n114) );
  INVX8 U111 ( .A(A[3]), .Y(SUM[3]) );
  INVX1 U112 ( .A(SUM[3]), .Y(n92) );
  OR2X2 U113 ( .A(n71), .B(A[30]), .Y(n93) );
  OAI21X1 U114 ( .A(n80), .B(n76), .C(n37), .Y(SUM[9]) );
  OAI21X1 U115 ( .A(n78), .B(n79), .C(n43), .Y(SUM[8]) );
  OAI21X1 U116 ( .A(n81), .B(n82), .C(n44), .Y(SUM[7]) );
  OAI21X1 U117 ( .A(n84), .B(n85), .C(n45), .Y(SUM[6]) );
  OAI21X1 U118 ( .A(n56), .B(n87), .C(n46), .Y(SUM[5]) );
  OAI21X1 U119 ( .A(n89), .B(n90), .C(n91), .Y(SUM[4]) );
  XNOR2X1 U120 ( .A(A[31]), .B(n93), .Y(SUM[31]) );
  OAI21X1 U121 ( .A(n94), .B(n95), .C(n71), .Y(SUM[29]) );
  INVX1 U122 ( .A(A[29]), .Y(n95) );
  OAI21X1 U123 ( .A(n58), .B(n97), .C(n51), .Y(SUM[28]) );
  INVX1 U124 ( .A(A[28]), .Y(n97) );
  OAI21X1 U125 ( .A(n99), .B(n100), .C(n98), .Y(SUM[27]) );
  INVX1 U126 ( .A(A[27]), .Y(n100) );
  OAI21X1 U127 ( .A(n57), .B(n102), .C(n52), .Y(SUM[26]) );
  INVX1 U128 ( .A(A[26]), .Y(n102) );
  OAI21X1 U129 ( .A(n104), .B(n105), .C(n103), .Y(SUM[25]) );
  INVX1 U130 ( .A(A[25]), .Y(n105) );
  OAI21X1 U131 ( .A(n61), .B(n107), .C(n47), .Y(SUM[24]) );
  INVX1 U132 ( .A(A[24]), .Y(n107) );
  OAI21X1 U133 ( .A(n109), .B(n110), .C(n108), .Y(SUM[23]) );
  INVX1 U134 ( .A(A[23]), .Y(n110) );
  OAI21X1 U135 ( .A(n63), .B(n112), .C(n53), .Y(SUM[22]) );
  INVX1 U136 ( .A(A[22]), .Y(n112) );
  OAI21X1 U137 ( .A(n114), .B(n115), .C(n113), .Y(SUM[21]) );
  INVX1 U138 ( .A(A[21]), .Y(n115) );
  OAI21X1 U139 ( .A(n118), .B(n117), .C(n48), .Y(SUM[20]) );
  INVX1 U140 ( .A(A[20]), .Y(n117) );
  OAI21X1 U141 ( .A(n67), .B(n119), .C(n36), .Y(SUM[19]) );
  INVX1 U142 ( .A(A[19]), .Y(n119) );
  OAI21X1 U143 ( .A(n121), .B(n122), .C(n120), .Y(SUM[18]) );
  INVX1 U144 ( .A(A[18]), .Y(n122) );
  OAI21X1 U145 ( .A(n60), .B(n123), .C(n49), .Y(SUM[17]) );
  INVX1 U146 ( .A(A[17]), .Y(n123) );
  OAI21X1 U147 ( .A(n125), .B(n126), .C(n124), .Y(SUM[16]) );
  INVX1 U148 ( .A(A[16]), .Y(n126) );
  OAI21X1 U149 ( .A(n129), .B(n128), .C(n55), .Y(SUM[15]) );
  INVX1 U150 ( .A(A[15]), .Y(n128) );
  OAI21X1 U151 ( .A(n32), .B(n130), .C(n40), .Y(SUM[14]) );
  INVX1 U152 ( .A(A[14]), .Y(n130) );
  OAI21X1 U153 ( .A(n33), .B(n131), .C(n41), .Y(SUM[13]) );
  INVX1 U154 ( .A(A[13]), .Y(n131) );
  OAI21X1 U155 ( .A(n65), .B(n133), .C(n42), .Y(SUM[12]) );
  INVX1 U156 ( .A(A[12]), .Y(n133) );
  OAI21X1 U157 ( .A(n135), .B(n136), .C(n134), .Y(SUM[11]) );
  INVX1 U158 ( .A(A[11]), .Y(n136) );
  OAI21X1 U159 ( .A(n137), .B(n138), .C(n50), .Y(SUM[10]) );
  INVX1 U160 ( .A(A[10]), .Y(n138) );
  INVX1 U161 ( .A(A[9]), .Y(n76) );
  INVX1 U162 ( .A(A[8]), .Y(n79) );
  INVX1 U163 ( .A(A[7]), .Y(n82) );
  INVX1 U164 ( .A(A[6]), .Y(n85) );
  INVX1 U165 ( .A(A[5]), .Y(n87) );
  INVX1 U166 ( .A(A[4]), .Y(n90) );
  INVX1 U167 ( .A(n92), .Y(n89) );
endmodule


module Processing_logic_DW01_inc_2 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;

  wire   [31:2] carry;

  HAX1 U1_1_30 ( .A(A[30]), .B(carry[30]), .YC(carry[31]), .YS(SUM[30]) );
  HAX1 U1_1_29 ( .A(A[29]), .B(carry[29]), .YC(carry[30]), .YS(SUM[29]) );
  HAX1 U1_1_28 ( .A(A[28]), .B(carry[28]), .YC(carry[29]), .YS(SUM[28]) );
  HAX1 U1_1_27 ( .A(A[27]), .B(carry[27]), .YC(carry[28]), .YS(SUM[27]) );
  HAX1 U1_1_26 ( .A(A[26]), .B(carry[26]), .YC(carry[27]), .YS(SUM[26]) );
  HAX1 U1_1_25 ( .A(A[25]), .B(carry[25]), .YC(carry[26]), .YS(SUM[25]) );
  HAX1 U1_1_24 ( .A(A[24]), .B(carry[24]), .YC(carry[25]), .YS(SUM[24]) );
  HAX1 U1_1_23 ( .A(A[23]), .B(carry[23]), .YC(carry[24]), .YS(SUM[23]) );
  HAX1 U1_1_22 ( .A(A[22]), .B(carry[22]), .YC(carry[23]), .YS(SUM[22]) );
  HAX1 U1_1_21 ( .A(A[21]), .B(carry[21]), .YC(carry[22]), .YS(SUM[21]) );
  HAX1 U1_1_20 ( .A(A[20]), .B(carry[20]), .YC(carry[21]), .YS(SUM[20]) );
  HAX1 U1_1_19 ( .A(A[19]), .B(carry[19]), .YC(carry[20]), .YS(SUM[19]) );
  HAX1 U1_1_18 ( .A(A[18]), .B(carry[18]), .YC(carry[19]), .YS(SUM[18]) );
  HAX1 U1_1_17 ( .A(A[17]), .B(carry[17]), .YC(carry[18]), .YS(SUM[17]) );
  HAX1 U1_1_16 ( .A(A[16]), .B(carry[16]), .YC(carry[17]), .YS(SUM[16]) );
  HAX1 U1_1_15 ( .A(A[15]), .B(carry[15]), .YC(carry[16]), .YS(SUM[15]) );
  HAX1 U1_1_14 ( .A(A[14]), .B(carry[14]), .YC(carry[15]), .YS(SUM[14]) );
  HAX1 U1_1_13 ( .A(A[13]), .B(carry[13]), .YC(carry[14]), .YS(SUM[13]) );
  HAX1 U1_1_12 ( .A(A[12]), .B(carry[12]), .YC(carry[13]), .YS(SUM[12]) );
  HAX1 U1_1_11 ( .A(A[11]), .B(carry[11]), .YC(carry[12]), .YS(SUM[11]) );
  HAX1 U1_1_10 ( .A(A[10]), .B(carry[10]), .YC(carry[11]), .YS(SUM[10]) );
  HAX1 U1_1_9 ( .A(A[9]), .B(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  HAX1 U1_1_8 ( .A(A[8]), .B(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  HAX1 U1_1_7 ( .A(A[7]), .B(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  HAX1 U1_1_6 ( .A(A[6]), .B(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  HAX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry[2]), .YS(SUM[1]) );
  XOR2X1 U1 ( .A(carry[31]), .B(A[31]), .Y(SUM[31]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module Processing_logic_DW_cmp_8 ( A, B, TC, GE_LT, GE_GT_EQ, GE_LT_GT_LE, 
        EQ_NE );
  input [31:0] A;
  input [31:0] B;
  input TC, GE_LT, GE_GT_EQ;
  output GE_LT_GT_LE, EQ_NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n11, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493;

  OAI21X1 U1 ( .A(n436), .B(n234), .C(n264), .Y(GE_LT_GT_LE) );
  AOI21X1 U3 ( .A(n2), .B(n244), .C(n7), .Y(n5) );
  OAI21X1 U5 ( .A(n248), .B(n442), .C(n262), .Y(n7) );
  AOI21X1 U7 ( .A(n15), .B(n491), .C(n11), .Y(n9) );
  OAI21X1 U13 ( .A(n233), .B(n246), .C(n271), .Y(n15) );
  AOI21X1 U19 ( .A(n29), .B(n242), .C(n23), .Y(n21) );
  OAI21X1 U21 ( .A(n282), .B(n250), .C(n269), .Y(n23) );
  OAI21X1 U27 ( .A(n280), .B(n288), .C(n266), .Y(n29) );
  OAI21X1 U33 ( .A(n286), .B(n439), .C(n260), .Y(n2) );
  AOI21X1 U35 ( .A(n43), .B(n457), .C(n37), .Y(n35) );
  OAI21X1 U37 ( .A(n289), .B(n427), .C(n339), .Y(n37) );
  OAI21X1 U43 ( .A(n424), .B(n489), .C(n336), .Y(n43) );
  AOI21X1 U49 ( .A(n57), .B(n454), .C(n51), .Y(n49) );
  OAI21X1 U51 ( .A(n421), .B(n486), .C(n333), .Y(n51) );
  OAI21X1 U57 ( .A(n418), .B(n483), .C(n330), .Y(n57) );
  AOI21X1 U62 ( .A(n92), .B(n388), .C(n63), .Y(n1) );
  OAI21X1 U64 ( .A(n459), .B(n433), .C(n257), .Y(n63) );
  AOI21X1 U66 ( .A(n73), .B(n445), .C(n67), .Y(n65) );
  OAI21X1 U68 ( .A(n415), .B(n480), .C(n327), .Y(n67) );
  OAI21X1 U74 ( .A(n412), .B(n477), .C(n324), .Y(n73) );
  AOI21X1 U80 ( .A(n87), .B(n451), .C(n81), .Y(n79) );
  OAI21X1 U82 ( .A(n409), .B(n474), .C(n321), .Y(n81) );
  OAI21X1 U88 ( .A(n406), .B(n471), .C(n318), .Y(n87) );
  OAI21X1 U93 ( .A(n403), .B(n430), .C(n254), .Y(n92) );
  AOI21X1 U95 ( .A(n102), .B(n448), .C(n96), .Y(n94) );
  OAI21X1 U97 ( .A(n400), .B(n468), .C(n315), .Y(n96) );
  OAI21X1 U103 ( .A(n397), .B(n465), .C(n312), .Y(n102) );
  AOI21X1 U108 ( .A(n391), .B(n385), .C(n109), .Y(n107) );
  OAI21X1 U110 ( .A(n394), .B(n462), .C(n309), .Y(n109) );
  INVX1 U119 ( .A(A[30]), .Y(n145) );
  INVX1 U120 ( .A(A[29]), .Y(n144) );
  INVX1 U121 ( .A(A[28]), .Y(n143) );
  INVX1 U122 ( .A(A[27]), .Y(n142) );
  INVX1 U123 ( .A(A[26]), .Y(n141) );
  INVX1 U124 ( .A(A[25]), .Y(n140) );
  INVX1 U125 ( .A(A[24]), .Y(n139) );
  INVX1 U126 ( .A(A[23]), .Y(n138) );
  INVX1 U127 ( .A(A[22]), .Y(n137) );
  INVX1 U128 ( .A(A[21]), .Y(n136) );
  INVX1 U129 ( .A(A[20]), .Y(n135) );
  INVX1 U130 ( .A(A[19]), .Y(n134) );
  INVX1 U131 ( .A(A[18]), .Y(n133) );
  INVX1 U132 ( .A(A[17]), .Y(n132) );
  INVX1 U133 ( .A(A[16]), .Y(n131) );
  INVX1 U134 ( .A(A[15]), .Y(n130) );
  INVX1 U135 ( .A(A[14]), .Y(n129) );
  INVX1 U136 ( .A(A[13]), .Y(n128) );
  INVX1 U137 ( .A(A[12]), .Y(n127) );
  INVX1 U138 ( .A(A[11]), .Y(n126) );
  INVX1 U139 ( .A(A[10]), .Y(n125) );
  INVX1 U140 ( .A(A[9]), .Y(n124) );
  INVX1 U141 ( .A(A[8]), .Y(n123) );
  INVX1 U142 ( .A(A[7]), .Y(n122) );
  INVX1 U143 ( .A(A[6]), .Y(n121) );
  INVX1 U144 ( .A(A[5]), .Y(n120) );
  INVX1 U145 ( .A(A[4]), .Y(n119) );
  INVX1 U146 ( .A(A[3]), .Y(n118) );
  BUFX2 U152 ( .A(B[30]), .Y(n221) );
  INVX1 U153 ( .A(n245), .Y(n222) );
  OR2X1 U154 ( .A(B[30]), .B(n145), .Y(n16) );
  INVX1 U155 ( .A(n249), .Y(n223) );
  OR2X1 U156 ( .A(B[28]), .B(n143), .Y(n24) );
  OR2X1 U157 ( .A(B[29]), .B(n144), .Y(n18) );
  INVX1 U158 ( .A(A[0]), .Y(n493) );
  INVX1 U159 ( .A(A[1]), .Y(n492) );
  OR2X2 U160 ( .A(n138), .B(B[23]), .Y(n40) );
  INVX1 U161 ( .A(n40), .Y(n224) );
  AND2X2 U162 ( .A(B[25]), .B(n140), .Y(n33) );
  INVX1 U163 ( .A(n33), .Y(n225) );
  OR2X2 U164 ( .A(n140), .B(B[25]), .Y(n32) );
  INVX1 U165 ( .A(n32), .Y(n226) );
  AND2X2 U166 ( .A(B[27]), .B(n142), .Y(n27) );
  INVX1 U167 ( .A(n27), .Y(n227) );
  OR2X2 U168 ( .A(n142), .B(B[27]), .Y(n26) );
  INVX1 U169 ( .A(n26), .Y(n228) );
  AND2X2 U170 ( .A(B[28]), .B(n143), .Y(n25) );
  INVX1 U171 ( .A(n25), .Y(n229) );
  AND2X2 U172 ( .A(n221), .B(n145), .Y(n17) );
  INVX1 U173 ( .A(n17), .Y(n230) );
  OR2X2 U174 ( .A(n245), .B(n278), .Y(n14) );
  INVX1 U175 ( .A(n14), .Y(n231) );
  AND2X2 U176 ( .A(A[31]), .B(n146), .Y(n13) );
  INVX1 U177 ( .A(n13), .Y(n232) );
  AND2X2 U178 ( .A(n144), .B(B[29]), .Y(n19) );
  INVX1 U179 ( .A(n19), .Y(n233) );
  AND2X2 U180 ( .A(n243), .B(n343), .Y(n4) );
  INVX1 U181 ( .A(n4), .Y(n234) );
  AND2X2 U182 ( .A(n341), .B(n284), .Y(n34) );
  INVX1 U183 ( .A(n34), .Y(n235) );
  INVX1 U184 ( .A(n34), .Y(n236) );
  OR2X2 U185 ( .A(n141), .B(B[26]), .Y(n30) );
  INVX1 U186 ( .A(n30), .Y(n237) );
  INVX1 U187 ( .A(n30), .Y(n238) );
  OR2X2 U188 ( .A(n139), .B(B[24]), .Y(n38) );
  INVX1 U189 ( .A(n38), .Y(n239) );
  INVX1 U190 ( .A(n38), .Y(n240) );
  OR2X2 U191 ( .A(n249), .B(n275), .Y(n22) );
  INVX1 U192 ( .A(n22), .Y(n241) );
  INVX1 U193 ( .A(n22), .Y(n242) );
  OR2X2 U194 ( .A(n247), .B(n364), .Y(n6) );
  INVX1 U195 ( .A(n6), .Y(n243) );
  INVX1 U196 ( .A(n6), .Y(n244) );
  INVX1 U197 ( .A(n16), .Y(n245) );
  INVX1 U198 ( .A(n222), .Y(n246) );
  AND2X2 U199 ( .A(n490), .B(n231), .Y(n8) );
  INVX1 U200 ( .A(n8), .Y(n247) );
  INVX1 U201 ( .A(n8), .Y(n248) );
  INVX1 U202 ( .A(n24), .Y(n249) );
  INVX1 U203 ( .A(n223), .Y(n250) );
  OR2X2 U204 ( .A(n137), .B(B[22]), .Y(n44) );
  INVX1 U205 ( .A(n44), .Y(n251) );
  OR2X2 U206 ( .A(n273), .B(n239), .Y(n36) );
  INVX1 U207 ( .A(n36), .Y(n252) );
  INVX1 U208 ( .A(B[31]), .Y(n146) );
  INVX1 U209 ( .A(n255), .Y(n253) );
  INVX1 U210 ( .A(n253), .Y(n254) );
  BUFX2 U211 ( .A(n94), .Y(n255) );
  INVX1 U212 ( .A(n258), .Y(n256) );
  INVX1 U213 ( .A(n256), .Y(n257) );
  BUFX2 U214 ( .A(n65), .Y(n258) );
  INVX1 U215 ( .A(n35), .Y(n259) );
  INVX1 U216 ( .A(n259), .Y(n260) );
  INVX1 U217 ( .A(n9), .Y(n261) );
  INVX1 U218 ( .A(n261), .Y(n262) );
  INVX1 U219 ( .A(n5), .Y(n263) );
  INVX1 U220 ( .A(n263), .Y(n264) );
  INVX1 U221 ( .A(n267), .Y(n265) );
  INVX1 U222 ( .A(n265), .Y(n266) );
  AND2X2 U223 ( .A(B[26]), .B(n141), .Y(n31) );
  INVX1 U224 ( .A(n31), .Y(n267) );
  INVX1 U225 ( .A(n229), .Y(n268) );
  INVX1 U226 ( .A(n268), .Y(n269) );
  INVX1 U227 ( .A(n230), .Y(n270) );
  INVX1 U228 ( .A(n270), .Y(n271) );
  INVX1 U229 ( .A(n224), .Y(n272) );
  INVX1 U230 ( .A(n272), .Y(n273) );
  INVX1 U231 ( .A(n228), .Y(n274) );
  INVX1 U232 ( .A(n274), .Y(n275) );
  INVX1 U233 ( .A(n226), .Y(n276) );
  INVX1 U234 ( .A(n276), .Y(n277) );
  INVX1 U235 ( .A(n18), .Y(n278) );
  INVX1 U236 ( .A(n232), .Y(n11) );
  INVX1 U237 ( .A(n225), .Y(n279) );
  INVX1 U238 ( .A(n279), .Y(n280) );
  INVX1 U239 ( .A(n227), .Y(n281) );
  INVX1 U240 ( .A(n281), .Y(n282) );
  INVX1 U241 ( .A(n252), .Y(n283) );
  INVX1 U242 ( .A(n283), .Y(n284) );
  INVX1 U243 ( .A(n235), .Y(n285) );
  INVX1 U244 ( .A(n285), .Y(n286) );
  INVX1 U245 ( .A(n237), .Y(n287) );
  INVX1 U246 ( .A(n287), .Y(n288) );
  BUFX2 U247 ( .A(n240), .Y(n289) );
  INVX1 U248 ( .A(n292), .Y(n290) );
  INVX1 U249 ( .A(n290), .Y(n291) );
  OR2X1 U250 ( .A(n492), .B(n493), .Y(n115) );
  INVX1 U251 ( .A(n115), .Y(n292) );
  INVX1 U252 ( .A(n295), .Y(n293) );
  INVX1 U253 ( .A(n293), .Y(n294) );
  OR2X1 U254 ( .A(n346), .B(n465), .Y(n101) );
  INVX1 U255 ( .A(n101), .Y(n295) );
  INVX1 U256 ( .A(n298), .Y(n296) );
  INVX1 U257 ( .A(n296), .Y(n297) );
  OR2X1 U258 ( .A(n349), .B(n471), .Y(n86) );
  INVX1 U259 ( .A(n86), .Y(n298) );
  INVX1 U260 ( .A(n301), .Y(n299) );
  INVX1 U261 ( .A(n299), .Y(n300) );
  OR2X1 U262 ( .A(n352), .B(n477), .Y(n72) );
  INVX1 U263 ( .A(n72), .Y(n301) );
  INVX1 U264 ( .A(n304), .Y(n302) );
  INVX1 U265 ( .A(n302), .Y(n303) );
  OR2X1 U266 ( .A(n355), .B(n483), .Y(n56) );
  INVX1 U267 ( .A(n56), .Y(n304) );
  INVX1 U268 ( .A(n307), .Y(n305) );
  INVX1 U269 ( .A(n305), .Y(n306) );
  OR2X2 U270 ( .A(n238), .B(n277), .Y(n28) );
  INVX1 U271 ( .A(n28), .Y(n307) );
  INVX1 U272 ( .A(n310), .Y(n308) );
  INVX1 U273 ( .A(n308), .Y(n309) );
  AND2X1 U274 ( .A(B[4]), .B(n119), .Y(n111) );
  INVX1 U275 ( .A(n111), .Y(n310) );
  INVX1 U276 ( .A(n313), .Y(n311) );
  INVX1 U277 ( .A(n311), .Y(n312) );
  AND2X1 U278 ( .A(B[6]), .B(n121), .Y(n104) );
  INVX1 U279 ( .A(n104), .Y(n313) );
  INVX1 U280 ( .A(n316), .Y(n314) );
  INVX1 U281 ( .A(n314), .Y(n315) );
  AND2X1 U282 ( .A(B[8]), .B(n123), .Y(n98) );
  INVX1 U283 ( .A(n98), .Y(n316) );
  INVX1 U284 ( .A(n319), .Y(n317) );
  INVX1 U285 ( .A(n317), .Y(n318) );
  AND2X1 U286 ( .A(B[10]), .B(n125), .Y(n89) );
  INVX1 U287 ( .A(n89), .Y(n319) );
  INVX1 U288 ( .A(n322), .Y(n320) );
  INVX1 U289 ( .A(n320), .Y(n321) );
  AND2X1 U290 ( .A(B[12]), .B(n127), .Y(n83) );
  INVX1 U291 ( .A(n83), .Y(n322) );
  INVX1 U292 ( .A(n325), .Y(n323) );
  INVX1 U293 ( .A(n323), .Y(n324) );
  AND2X1 U294 ( .A(B[14]), .B(n129), .Y(n75) );
  INVX1 U295 ( .A(n75), .Y(n325) );
  INVX1 U296 ( .A(n328), .Y(n326) );
  INVX1 U297 ( .A(n326), .Y(n327) );
  AND2X1 U298 ( .A(B[16]), .B(n131), .Y(n69) );
  INVX1 U299 ( .A(n69), .Y(n328) );
  INVX1 U300 ( .A(n331), .Y(n329) );
  INVX1 U301 ( .A(n329), .Y(n330) );
  AND2X1 U302 ( .A(B[18]), .B(n133), .Y(n59) );
  INVX1 U303 ( .A(n59), .Y(n331) );
  INVX1 U304 ( .A(n334), .Y(n332) );
  INVX1 U305 ( .A(n332), .Y(n333) );
  AND2X1 U306 ( .A(B[20]), .B(n135), .Y(n53) );
  INVX1 U307 ( .A(n53), .Y(n334) );
  INVX1 U308 ( .A(n337), .Y(n335) );
  INVX1 U309 ( .A(n335), .Y(n336) );
  AND2X1 U310 ( .A(B[22]), .B(n137), .Y(n45) );
  INVX1 U311 ( .A(n45), .Y(n337) );
  INVX1 U312 ( .A(n340), .Y(n338) );
  INVX1 U313 ( .A(n338), .Y(n339) );
  AND2X2 U314 ( .A(B[24]), .B(n139), .Y(n39) );
  INVX1 U315 ( .A(n39), .Y(n340) );
  OR2X2 U316 ( .A(n361), .B(n489), .Y(n42) );
  INVX1 U317 ( .A(n42), .Y(n341) );
  INVX1 U318 ( .A(n344), .Y(n342) );
  INVX1 U319 ( .A(n342), .Y(n343) );
  OR2X2 U320 ( .A(n236), .B(n358), .Y(n3) );
  INVX1 U321 ( .A(n3), .Y(n344) );
  INVX1 U322 ( .A(n347), .Y(n345) );
  INVX1 U323 ( .A(n345), .Y(n346) );
  OR2X1 U324 ( .A(n120), .B(B[5]), .Y(n105) );
  INVX1 U325 ( .A(n105), .Y(n347) );
  INVX1 U326 ( .A(n350), .Y(n348) );
  INVX1 U327 ( .A(n348), .Y(n349) );
  OR2X1 U328 ( .A(n124), .B(B[9]), .Y(n90) );
  INVX1 U329 ( .A(n90), .Y(n350) );
  INVX1 U330 ( .A(n353), .Y(n351) );
  INVX1 U331 ( .A(n351), .Y(n352) );
  OR2X1 U332 ( .A(n128), .B(B[13]), .Y(n76) );
  INVX1 U333 ( .A(n76), .Y(n353) );
  INVX1 U334 ( .A(n356), .Y(n354) );
  INVX1 U335 ( .A(n354), .Y(n355) );
  OR2X1 U336 ( .A(n132), .B(B[17]), .Y(n60) );
  INVX1 U337 ( .A(n60), .Y(n356) );
  INVX1 U338 ( .A(n359), .Y(n357) );
  INVX1 U339 ( .A(n357), .Y(n358) );
  AND2X2 U340 ( .A(n454), .B(n303), .Y(n48) );
  INVX1 U341 ( .A(n48), .Y(n359) );
  INVX1 U342 ( .A(n362), .Y(n360) );
  INVX1 U343 ( .A(n360), .Y(n361) );
  OR2X2 U344 ( .A(n136), .B(B[21]), .Y(n46) );
  INVX1 U345 ( .A(n46), .Y(n362) );
  INVX1 U346 ( .A(n365), .Y(n363) );
  INVX1 U347 ( .A(n363), .Y(n364) );
  AND2X2 U348 ( .A(n241), .B(n306), .Y(n20) );
  INVX1 U349 ( .A(n20), .Y(n365) );
  INVX1 U350 ( .A(n368), .Y(n366) );
  INVX1 U351 ( .A(n366), .Y(n367) );
  OR2X2 U352 ( .A(n118), .B(B[3]), .Y(n112) );
  INVX1 U353 ( .A(n112), .Y(n368) );
  INVX1 U354 ( .A(n371), .Y(n369) );
  INVX1 U355 ( .A(n369), .Y(n370) );
  OR2X1 U356 ( .A(n122), .B(B[7]), .Y(n99) );
  INVX1 U357 ( .A(n99), .Y(n371) );
  INVX1 U358 ( .A(n374), .Y(n372) );
  INVX1 U359 ( .A(n372), .Y(n373) );
  OR2X1 U360 ( .A(n126), .B(B[11]), .Y(n84) );
  INVX1 U361 ( .A(n84), .Y(n374) );
  INVX1 U362 ( .A(n377), .Y(n375) );
  INVX1 U363 ( .A(n375), .Y(n376) );
  AND2X2 U364 ( .A(n451), .B(n297), .Y(n78) );
  INVX1 U365 ( .A(n78), .Y(n377) );
  INVX1 U366 ( .A(n380), .Y(n378) );
  INVX1 U367 ( .A(n378), .Y(n379) );
  OR2X1 U368 ( .A(n130), .B(B[15]), .Y(n70) );
  INVX1 U369 ( .A(n70), .Y(n380) );
  INVX1 U370 ( .A(n383), .Y(n381) );
  INVX1 U371 ( .A(n381), .Y(n382) );
  OR2X1 U372 ( .A(n134), .B(B[19]), .Y(n54) );
  INVX1 U373 ( .A(n54), .Y(n383) );
  INVX1 U374 ( .A(n386), .Y(n384) );
  INVX1 U375 ( .A(n384), .Y(n385) );
  AND2X2 U376 ( .A(A[2]), .B(n291), .Y(n114) );
  INVX1 U377 ( .A(n114), .Y(n386) );
  INVX1 U378 ( .A(n389), .Y(n387) );
  INVX1 U379 ( .A(n387), .Y(n388) );
  OR2X2 U380 ( .A(n376), .B(n459), .Y(n62) );
  INVX1 U381 ( .A(n62), .Y(n389) );
  INVX1 U382 ( .A(n392), .Y(n390) );
  INVX1 U383 ( .A(n390), .Y(n391) );
  OR2X2 U384 ( .A(n367), .B(n462), .Y(n108) );
  INVX1 U385 ( .A(n108), .Y(n392) );
  INVX1 U386 ( .A(n395), .Y(n393) );
  INVX1 U387 ( .A(n393), .Y(n394) );
  AND2X2 U388 ( .A(B[3]), .B(n118), .Y(n113) );
  INVX1 U389 ( .A(n113), .Y(n395) );
  INVX1 U390 ( .A(n398), .Y(n396) );
  INVX1 U391 ( .A(n396), .Y(n397) );
  AND2X1 U392 ( .A(B[5]), .B(n120), .Y(n106) );
  INVX1 U393 ( .A(n106), .Y(n398) );
  INVX1 U394 ( .A(n401), .Y(n399) );
  INVX1 U395 ( .A(n399), .Y(n400) );
  AND2X1 U396 ( .A(B[7]), .B(n122), .Y(n100) );
  INVX1 U397 ( .A(n100), .Y(n401) );
  INVX1 U398 ( .A(n404), .Y(n402) );
  INVX1 U399 ( .A(n402), .Y(n403) );
  AND2X2 U400 ( .A(n448), .B(n294), .Y(n93) );
  INVX1 U401 ( .A(n93), .Y(n404) );
  INVX1 U402 ( .A(n407), .Y(n405) );
  INVX1 U403 ( .A(n405), .Y(n406) );
  AND2X1 U404 ( .A(B[9]), .B(n124), .Y(n91) );
  INVX1 U405 ( .A(n91), .Y(n407) );
  INVX1 U406 ( .A(n410), .Y(n408) );
  INVX1 U407 ( .A(n408), .Y(n409) );
  AND2X1 U408 ( .A(B[11]), .B(n126), .Y(n85) );
  INVX1 U409 ( .A(n85), .Y(n410) );
  INVX1 U410 ( .A(n413), .Y(n411) );
  INVX1 U411 ( .A(n411), .Y(n412) );
  AND2X1 U412 ( .A(B[13]), .B(n128), .Y(n77) );
  INVX1 U413 ( .A(n77), .Y(n413) );
  INVX1 U414 ( .A(n416), .Y(n414) );
  INVX1 U415 ( .A(n414), .Y(n415) );
  AND2X1 U416 ( .A(B[15]), .B(n130), .Y(n71) );
  INVX1 U417 ( .A(n71), .Y(n416) );
  INVX1 U418 ( .A(n419), .Y(n417) );
  INVX1 U419 ( .A(n417), .Y(n418) );
  AND2X1 U420 ( .A(B[17]), .B(n132), .Y(n61) );
  INVX1 U421 ( .A(n61), .Y(n419) );
  INVX1 U422 ( .A(n422), .Y(n420) );
  INVX1 U423 ( .A(n420), .Y(n421) );
  AND2X1 U424 ( .A(B[19]), .B(n134), .Y(n55) );
  INVX1 U425 ( .A(n55), .Y(n422) );
  INVX1 U426 ( .A(n425), .Y(n423) );
  INVX1 U427 ( .A(n423), .Y(n424) );
  AND2X1 U428 ( .A(B[21]), .B(n136), .Y(n47) );
  INVX1 U429 ( .A(n47), .Y(n425) );
  INVX1 U430 ( .A(n428), .Y(n426) );
  INVX1 U431 ( .A(n426), .Y(n427) );
  AND2X1 U432 ( .A(B[23]), .B(n138), .Y(n41) );
  INVX1 U433 ( .A(n41), .Y(n428) );
  INVX1 U434 ( .A(n431), .Y(n429) );
  INVX1 U435 ( .A(n429), .Y(n430) );
  BUFX2 U436 ( .A(n107), .Y(n431) );
  INVX1 U437 ( .A(n434), .Y(n432) );
  INVX1 U438 ( .A(n432), .Y(n433) );
  BUFX2 U439 ( .A(n79), .Y(n434) );
  INVX1 U440 ( .A(n437), .Y(n435) );
  INVX1 U441 ( .A(n435), .Y(n436) );
  BUFX2 U442 ( .A(n1), .Y(n437) );
  INVX1 U443 ( .A(n440), .Y(n438) );
  INVX1 U444 ( .A(n438), .Y(n439) );
  BUFX2 U445 ( .A(n49), .Y(n440) );
  INVX1 U446 ( .A(n443), .Y(n441) );
  INVX1 U447 ( .A(n441), .Y(n442) );
  BUFX2 U448 ( .A(n21), .Y(n443) );
  INVX1 U449 ( .A(n446), .Y(n444) );
  INVX1 U450 ( .A(n444), .Y(n445) );
  OR2X2 U451 ( .A(n379), .B(n480), .Y(n66) );
  INVX1 U452 ( .A(n66), .Y(n446) );
  INVX1 U453 ( .A(n449), .Y(n447) );
  INVX1 U454 ( .A(n447), .Y(n448) );
  OR2X2 U455 ( .A(n370), .B(n468), .Y(n95) );
  INVX1 U456 ( .A(n95), .Y(n449) );
  INVX1 U457 ( .A(n452), .Y(n450) );
  INVX1 U458 ( .A(n450), .Y(n451) );
  OR2X2 U459 ( .A(n373), .B(n474), .Y(n80) );
  INVX1 U460 ( .A(n80), .Y(n452) );
  INVX1 U461 ( .A(n455), .Y(n453) );
  INVX1 U462 ( .A(n453), .Y(n454) );
  OR2X2 U463 ( .A(n382), .B(n486), .Y(n50) );
  INVX1 U464 ( .A(n50), .Y(n455) );
  INVX1 U465 ( .A(n284), .Y(n456) );
  INVX1 U466 ( .A(n456), .Y(n457) );
  INVX1 U467 ( .A(n460), .Y(n458) );
  INVX1 U468 ( .A(n458), .Y(n459) );
  AND2X2 U469 ( .A(n445), .B(n300), .Y(n64) );
  INVX1 U470 ( .A(n64), .Y(n460) );
  INVX1 U471 ( .A(n463), .Y(n461) );
  INVX1 U472 ( .A(n461), .Y(n462) );
  OR2X1 U473 ( .A(n119), .B(B[4]), .Y(n110) );
  INVX1 U474 ( .A(n110), .Y(n463) );
  INVX1 U475 ( .A(n466), .Y(n464) );
  INVX1 U476 ( .A(n464), .Y(n465) );
  OR2X1 U477 ( .A(n121), .B(B[6]), .Y(n103) );
  INVX1 U478 ( .A(n103), .Y(n466) );
  INVX1 U479 ( .A(n469), .Y(n467) );
  INVX1 U480 ( .A(n467), .Y(n468) );
  OR2X1 U481 ( .A(n123), .B(B[8]), .Y(n97) );
  INVX1 U482 ( .A(n97), .Y(n469) );
  INVX1 U483 ( .A(n472), .Y(n470) );
  INVX1 U484 ( .A(n470), .Y(n471) );
  OR2X1 U485 ( .A(n125), .B(B[10]), .Y(n88) );
  INVX1 U486 ( .A(n88), .Y(n472) );
  INVX1 U487 ( .A(n475), .Y(n473) );
  INVX1 U488 ( .A(n473), .Y(n474) );
  OR2X1 U489 ( .A(n127), .B(B[12]), .Y(n82) );
  INVX1 U490 ( .A(n82), .Y(n475) );
  INVX1 U491 ( .A(n478), .Y(n476) );
  INVX1 U492 ( .A(n476), .Y(n477) );
  OR2X1 U493 ( .A(n129), .B(B[14]), .Y(n74) );
  INVX1 U494 ( .A(n74), .Y(n478) );
  INVX1 U495 ( .A(n481), .Y(n479) );
  INVX1 U496 ( .A(n479), .Y(n480) );
  OR2X1 U497 ( .A(n131), .B(B[16]), .Y(n68) );
  INVX1 U498 ( .A(n68), .Y(n481) );
  INVX1 U499 ( .A(n484), .Y(n482) );
  INVX1 U500 ( .A(n482), .Y(n483) );
  OR2X1 U501 ( .A(n133), .B(B[18]), .Y(n58) );
  INVX1 U502 ( .A(n58), .Y(n484) );
  INVX1 U503 ( .A(n487), .Y(n485) );
  INVX1 U504 ( .A(n485), .Y(n486) );
  OR2X1 U505 ( .A(n135), .B(B[20]), .Y(n52) );
  INVX1 U506 ( .A(n52), .Y(n487) );
  INVX1 U507 ( .A(n251), .Y(n488) );
  INVX1 U508 ( .A(n488), .Y(n489) );
  OR2X2 U509 ( .A(n146), .B(A[31]), .Y(n490) );
  OR2X2 U510 ( .A(n146), .B(A[31]), .Y(n491) );
endmodule


module Processing_logic ( clk, ck, reset, ready, DATA_data_out, DATA_get, 
        CMD_empty, CMD_data_out, CMD_get, RETURN_full, RETURN_put, 
        RETURN_address, RETURN_data, DQ_in, DQS_in, DQS_bar_in, cs_bar, 
        ras_bar, cas_bar, we_bar, DQ_out, DQS_out, DQS_bar_out, BA, A, DM, 
        ts_con, ri_o );
  input [15:0] DATA_data_out;
  input [33:0] CMD_data_out;
  output [25:0] RETURN_address;
  output [15:0] RETURN_data;
  input [15:0] DQ_in;
  input [1:0] DQS_in;
  input [1:0] DQS_bar_in;
  output [15:0] DQ_out;
  output [1:0] DQS_out;
  output [1:0] DQS_bar_out;
  output [2:0] BA;
  output [12:0] A;
  output [1:0] DM;
  input clk, ck, reset, ready, CMD_empty, RETURN_full;
  output DATA_get, CMD_get, RETURN_put, cs_bar, ras_bar, cas_bar, we_bar,
         ts_con, ri_o;
  wire   n229, n230, n231, n232, listen, flag_bl_write, flag_bl_read, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, flag_at_read, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n1752, n1753, n1754, n1755, n1756,
         n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
         n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
         n1777, n1778, n1779, n1780, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n2077, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2442, n2509, n3036,
         n3073, n3079, n3126, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n669, n703, n737, n805,
         n839, n873, n907, n942, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n2439, n2546, n2547, n2548, n2551, n2553, n2555, n2557,
         n2559, n2561, n2563, n2565, n2567, n2569, n2571, n2573, n2575, n2577,
         n2579, n2581, n2583, n2585, n2587, n2589, n2591, n2593, n2595, n2597,
         n2599, n2601, n2603, n2605, n2607, n2609, n2611, n2613, n2615, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2647, n2648, n2649,
         n2650, n2651, n2653, n2654, n2656, n2657, n2658, n2659, n2660, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2707, n2708, n2709, n2710, n2711, n2713, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2724, n2725, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2749,
         n2750, n2752, n2753, n2754, n2756, n2757, n2758, n2760, n2761, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2771, n2772, n2773, n2774,
         n2775, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2796,
         n2798, n2799, n2801, n2802, n2803, n2804, n2806, n2807, n2808, n2810,
         n2811, n2814, n2815, n2816, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2828, n2829, n2830, n2831, n2832, n2834, n2835,
         n2836, n2837, n2838, n2839, n2841, n2842, n2843, n2847, n2849, n2850,
         n2851, n2852, n2854, n2855, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2874, n2876, n2877, n2879, n2880, n2881, n2882, n2883, n2885, n2887,
         n2888, n2889, n2900, n2901, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2923, n2924, n2926, n2927, n2928, n2934, n2936, n2937,
         n2938, n2939, n2940, n2941, n2942, n2946, n2947, n2948, n2949, n2950,
         n2952, n2953, n2954, n2957, n2959, n2961, n2962, n2963, n2964, n2966,
         n2968, n2969, n2970, n2971, n2972, n2973, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2998, n2999, n3000,
         n3001, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3021, n3022,
         n3023, n3024, n3025, n3027, n3028, n3029, n3031, n3032, n3034, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3063, n3064, n3065, n3066, n3067, n3069, n3070,
         n3071, n3072, n3075, n3076, n3077, n3078, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3104,
         n3106, n3107, n3108, n3110, n3111, n3112, n3113, n3115, n3117, n3118,
         n3121, n3122, n3123, n3124, n3128, n3129, n3130, n3131, n3132, n3134,
         n3135, n3136, n3137, n3138, n3140, n3142, n3144, n3146, n3148, n3150,
         n3152, n3154, n3156, n3158, n3160, n3162, n3164, n3166, n3168, n3170,
         n3172, n3174, n3176, n3178, n3180, n3182, n3184, n3186, n3188, n3190,
         n3192, n3194, n3196, n3198, n3200, n3202, n3204, n3206, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3223, n3225, n3227, n3229, n3231, n3233, n3235, n3237,
         n3239, n3241, n3243, n3245, n3247, n3249, n3251, n3253, n3255, n3257,
         n3259, n3261, n3263, n3265, n3267, n3269, n3271, n3273, n3275, n3277,
         n3279, n3281, n3283, n3285, n3287, n3289, n3291, n3293, n3295, n3297,
         n3299, n3301, n3303, n3305, n3307, n3309, n3311, n3313, n3315, n3317,
         n3319, n3321, n3323, n3325, n3327, n3329, n3331, n3333, n3335, n3337,
         n3339, n3341, n3343, n3345, n3347, n3349, n3351, n3353, n3355, n3357,
         n3359, n3361, n3363, n3365, n3367, n3369, n3371, n3373, n3375, n3377,
         n3379, n3381, n3383, n3385, n3387, n3389, n3391, n3393, n3395, n3397,
         n3399, n3401, n3403, n3405, n3407, n3409, n3411, n3413, n3415, n3417,
         n3419, n3421, n3427, net67203, net67172, net67122, net67120, net66975,
         net66974, net66962, net66953, net66834, net66714, net66503, net66499,
         net66482, net66423, net66385, net66383, net66381, net66380, net66378,
         net66376, net66374, net66372, net66370, net66368, net66352, net66350,
         net66348, net66346, net66344, net66342, net66339, net66338, net66336,
         net66330, net66328, net66325, net66319, net66290, net66289, net66283,
         net66168, net66166, net66160, net66151, net66149, net66140, net66116,
         net66114, net66112, net66110, net66108, net66106, net66104, net66102,
         net66100, net66098, net66096, net66094, net66092, net66090, net66088,
         net66086, net66084, net66082, net66080, net66078, net66076, net66073,
         net66063, net66062, net66061, net66060, net66046, net66042, net66031,
         net66007, net65999, net65992, net65987, net65981, r577_net62534,
         r577_GE_LT_GT_LE, r576_net62635, r576_net62636, add_576_carry_7_,
         add_576_carry_8_, add_576_carry_9_, add_576_carry_10_,
         add_576_carry_11_, add_576_carry_12_, C25909_net2920, C25909_net2767,
         C25909_net2740, C25909_net2624, net79422, net79420, net79416,
         net79414, net79412, net79410, net79408, net79402, net79400, net79398,
         net79440, net79436, net79434, net79432, net79430, net79428, net79482,
         net79510, net79514, net79518, net79534, net79533, net79538, net79541,
         net79593, net79605, net79794, net80322, net80376, net80382, net80435,
         net80464, net80463, net80519, net80518, net80561, net80598, net80596,
         net80595, net80661, net80682, net80709, net80708, net80723, net80736,
         net80747, net80760, net80775, net80781, net80783, net80791, net80839,
         net80862, net80872, net80914, net80718, net80717, net66539, net66327,
         net82094, net82125, net82138, net82191, net82209, net82215, net82336,
         net82349, net82348, net82428, net82427, net82435, net82472, net82506,
         net82538, net82567, net82576, net82455, net82454, net66558, net66329,
         net84792, net66956, net66955, r576_net62631, r576_net62630,
         r576_net62619, r576_GE_LT_GT_LE, net89555, net89705, net89562,
         net89554, net66954, net92619, net92789, net92764, net92761, net92751,
         net92748, net92746, net92732, net92731, net92836, net92856, net92867,
         net92933, net93022, net93057, net93072, net93077, net92773, net92735,
         net89563, net89561, net89543, net80232, net66970, net92747, net92757,
         net92738, net92651, net79438, net66441, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n249, n250, n251, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n628, n629, n630, n631, n632, n633, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1751, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2078, n2079, n2080, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2376, n2377, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2440,
         n2441, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2549, n2629, n2646, n2652, n2655, n2661, n2671,
         n2706, n2712, n2714, n2723, n2726, n2748, n2751, n2755, n2759, n2762,
         n2770, n2776, n2795, n2797, n2800, n2805, n2809, n2812, n2813, n2817,
         n2827, n2833, n2840, n2844, n2845, n2846, n2848, n2853, n2856, n2873,
         n2875, n2878, n2884, n2886, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2902, n2903, n2922, n2925, n2929, n2930,
         n2931, n2932, n2933, n2935, n2943, n2944, n2945, n2951, n2955, n2956,
         n2958, n2960, n2965, n2967, n2974, n2983, n2997, n3002, n3020, n3026,
         n3030, n3033, n3035, n3052, n3062, n3068, n3074, n3103, n3105, n3109,
         n3114, n3116, n3119, n3120, n3125, n3127, n3133, n3423, n3424, n3425,
         n3426, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
         n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877,
         n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887,
         n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897,
         n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
         n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
         n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987,
         n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997,
         n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007,
         n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017,
         n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
         n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037,
         n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047,
         n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057,
         n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067,
         n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077,
         n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087,
         n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097,
         n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107,
         n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117,
         n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
         n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
         n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
         n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
         n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
         n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
         n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
         n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
         n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
         n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
         n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
         n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257,
         n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267,
         n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
         n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6;
  wire   [2:0] ring_ptr;
  wire   [31:0] clkcount;
  wire   [4:0] state;
  wire   [31:0] i;
  wire   [31:5] j;
  wire   [31:0] blk_cnt;
  wire   [2:0] buff_bank_addr;
  wire   [9:0] buff_col_addr;
  wire   [511:0] buff_data;
  assign RETURN_address[25] = CMD_data_out[25];
  assign RETURN_address[24] = CMD_data_out[24];
  assign RETURN_address[23] = CMD_data_out[23];
  assign RETURN_address[22] = CMD_data_out[22];
  assign RETURN_address[21] = CMD_data_out[21];
  assign RETURN_address[20] = CMD_data_out[20];
  assign RETURN_address[19] = CMD_data_out[19];
  assign RETURN_address[18] = CMD_data_out[18];
  assign RETURN_address[17] = CMD_data_out[17];
  assign RETURN_address[16] = CMD_data_out[16];
  assign RETURN_address[15] = CMD_data_out[15];
  assign RETURN_address[14] = CMD_data_out[14];
  assign RETURN_address[13] = CMD_data_out[13];
  assign RETURN_address[12] = CMD_data_out[12];
  assign RETURN_address[11] = CMD_data_out[11];
  assign RETURN_address[10] = CMD_data_out[10];
  assign RETURN_address[9] = CMD_data_out[9];
  assign RETURN_address[8] = CMD_data_out[8];
  assign RETURN_address[7] = CMD_data_out[7];
  assign RETURN_address[6] = CMD_data_out[6];
  assign RETURN_address[5] = CMD_data_out[5];
  assign RETURN_address[4] = CMD_data_out[4];
  assign RETURN_address[3] = CMD_data_out[3];
  assign RETURN_address[2] = CMD_data_out[2];
  assign RETURN_address[1] = CMD_data_out[1];
  assign RETURN_address[0] = CMD_data_out[0];
  assign cs_bar = 1'b0;
  assign DM[1] = 1'b0;
  assign DM[0] = 1'b0;

  ddr3_ring_buffer8 ring_buffer ( .dout(RETURN_data), .listen(listen), 
        .strobe(DQS_in[0]), .readPtr(ring_ptr), .din(DQ_in), .reset(reset) );
  DFFNEGX1 buff_bank_addr_reg_2_ ( .D(n3208), .CLK(clk), .Q(buff_bank_addr[2])
         );
  DFFNEGX1 buff_bank_addr_reg_1_ ( .D(n3209), .CLK(clk), .Q(buff_bank_addr[1])
         );
  DFFNEGX1 buff_bank_addr_reg_0_ ( .D(n3210), .CLK(clk), .Q(buff_bank_addr[0])
         );
  DFFNEGX1 buff_col_addr_reg_9_ ( .D(n3211), .CLK(clk), .Q(buff_col_addr[9])
         );
  DFFNEGX1 buff_col_addr_reg_8_ ( .D(n3212), .CLK(clk), .Q(buff_col_addr[8])
         );
  DFFNEGX1 buff_col_addr_reg_7_ ( .D(n3213), .CLK(clk), .Q(buff_col_addr[7])
         );
  DFFNEGX1 buff_col_addr_reg_6_ ( .D(n3214), .CLK(clk), .Q(buff_col_addr[6])
         );
  DFFNEGX1 buff_col_addr_reg_5_ ( .D(n3215), .CLK(clk), .Q(buff_col_addr[5])
         );
  DFFNEGX1 buff_col_addr_reg_4_ ( .D(n3216), .CLK(clk), .Q(buff_col_addr[4])
         );
  DFFNEGX1 buff_col_addr_reg_3_ ( .D(n3217), .CLK(clk), .Q(buff_col_addr[3])
         );
  DFFNEGX1 buff_col_addr_reg_2_ ( .D(n3218), .CLK(clk), .Q(buff_col_addr[2])
         );
  DFFNEGX1 buff_col_addr_reg_1_ ( .D(n3219), .CLK(clk), .Q(buff_col_addr[1])
         );
  DFFNEGX1 buff_col_addr_reg_0_ ( .D(n3220), .CLK(clk), .Q(buff_col_addr[0])
         );
  DFFNEGX1 buff_data_reg_1__1_ ( .D(n2633), .CLK(clk), .Q(buff_data[481]) );
  DFFNEGX1 buff_data_reg_1__0_ ( .D(n2634), .CLK(clk), .Q(buff_data[480]) );
  DFFNEGX1 buff_data_reg_1__15_ ( .D(n2635), .CLK(clk), .Q(buff_data[495]) );
  DFFNEGX1 buff_data_reg_1__14_ ( .D(n2636), .CLK(clk), .Q(buff_data[494]) );
  DFFNEGX1 buff_data_reg_1__13_ ( .D(n2637), .CLK(clk), .Q(buff_data[493]) );
  DFFNEGX1 buff_data_reg_1__12_ ( .D(n2638), .CLK(clk), .Q(buff_data[492]) );
  DFFNEGX1 buff_data_reg_1__11_ ( .D(n2639), .CLK(clk), .Q(buff_data[491]) );
  DFFNEGX1 buff_data_reg_1__10_ ( .D(n2640), .CLK(clk), .Q(buff_data[490]) );
  DFFNEGX1 buff_data_reg_1__9_ ( .D(n2641), .CLK(clk), .Q(buff_data[489]) );
  DFFNEGX1 buff_data_reg_1__8_ ( .D(n2642), .CLK(clk), .Q(buff_data[488]) );
  DFFNEGX1 buff_data_reg_1__7_ ( .D(n2643), .CLK(clk), .Q(buff_data[487]) );
  DFFNEGX1 buff_data_reg_1__6_ ( .D(n2644), .CLK(clk), .Q(buff_data[486]) );
  DFFNEGX1 buff_data_reg_1__5_ ( .D(n2645), .CLK(clk), .Q(buff_data[485]) );
  DFFNEGX1 buff_data_reg_1__4_ ( .D(n2120), .CLK(clk), .Q(buff_data[484]) );
  DFFNEGX1 buff_data_reg_1__3_ ( .D(n2647), .CLK(clk), .Q(buff_data[483]) );
  DFFNEGX1 buff_data_reg_1__2_ ( .D(n2648), .CLK(clk), .Q(buff_data[482]) );
  DFFNEGX1 buff_data_reg_8__14_ ( .D(n2745), .CLK(clk), .Q(buff_data[382]) );
  DFFNEGX1 buff_data_reg_8__13_ ( .D(n2746), .CLK(clk), .Q(buff_data[381]) );
  DFFNEGX1 buff_data_reg_8__12_ ( .D(n2747), .CLK(clk), .Q(buff_data[380]) );
  DFFNEGX1 buff_data_reg_8__11_ ( .D(n1976), .CLK(clk), .Q(buff_data[379]) );
  DFFNEGX1 buff_data_reg_8__10_ ( .D(n2749), .CLK(clk), .Q(buff_data[378]) );
  DFFNEGX1 buff_data_reg_8__9_ ( .D(n2750), .CLK(clk), .Q(buff_data[377]) );
  DFFNEGX1 buff_data_reg_8__8_ ( .D(n2006), .CLK(clk), .Q(buff_data[376]) );
  DFFNEGX1 buff_data_reg_8__7_ ( .D(n2752), .CLK(clk), .Q(buff_data[375]) );
  DFFNEGX1 buff_data_reg_8__6_ ( .D(n2753), .CLK(clk), .Q(buff_data[374]) );
  DFFNEGX1 buff_data_reg_8__5_ ( .D(n2754), .CLK(clk), .Q(buff_data[373]) );
  DFFNEGX1 buff_data_reg_8__4_ ( .D(n1993), .CLK(clk), .Q(buff_data[372]) );
  DFFNEGX1 buff_data_reg_8__3_ ( .D(n2756), .CLK(clk), .Q(buff_data[371]) );
  DFFNEGX1 buff_data_reg_8__2_ ( .D(n2757), .CLK(clk), .Q(buff_data[370]) );
  DFFNEGX1 buff_data_reg_8__1_ ( .D(n2758), .CLK(clk), .Q(buff_data[369]) );
  DFFNEGX1 buff_data_reg_8__0_ ( .D(n2130), .CLK(clk), .Q(buff_data[368]) );
  DFFNEGX1 buff_data_reg_8__15_ ( .D(n2760), .CLK(clk), .Q(buff_data[383]) );
  DFFNEGX1 buff_data_reg_14__11_ ( .D(n2841), .CLK(clk), .Q(buff_data[283]) );
  DFFNEGX1 buff_data_reg_14__10_ ( .D(n2842), .CLK(clk), .Q(buff_data[282]) );
  DFFNEGX1 buff_data_reg_14__9_ ( .D(n2843), .CLK(clk), .Q(buff_data[281]) );
  DFFNEGX1 buff_data_reg_14__8_ ( .D(n1974), .CLK(clk), .Q(buff_data[280]) );
  DFFNEGX1 buff_data_reg_14__7_ ( .D(n1981), .CLK(clk), .Q(buff_data[279]) );
  DFFNEGX1 buff_data_reg_14__6_ ( .D(n1961), .CLK(clk), .Q(buff_data[278]) );
  DFFNEGX1 buff_data_reg_14__5_ ( .D(n2847), .CLK(clk), .Q(buff_data[277]) );
  DFFNEGX1 buff_data_reg_14__4_ ( .D(n1838), .CLK(clk), .Q(buff_data[276]) );
  DFFNEGX1 buff_data_reg_14__3_ ( .D(n2849), .CLK(clk), .Q(buff_data[275]) );
  DFFNEGX1 buff_data_reg_14__2_ ( .D(n2850), .CLK(clk), .Q(buff_data[274]) );
  DFFNEGX1 buff_data_reg_14__1_ ( .D(n2851), .CLK(clk), .Q(buff_data[273]) );
  DFFNEGX1 buff_data_reg_14__0_ ( .D(n2852), .CLK(clk), .Q(buff_data[272]) );
  DFFNEGX1 buff_data_reg_14__15_ ( .D(n1963), .CLK(clk), .Q(buff_data[287]) );
  DFFNEGX1 buff_data_reg_14__14_ ( .D(n2854), .CLK(clk), .Q(buff_data[286]) );
  DFFNEGX1 buff_data_reg_14__13_ ( .D(n2855), .CLK(clk), .Q(buff_data[285]) );
  DFFNEGX1 buff_data_reg_14__12_ ( .D(n2140), .CLK(clk), .Q(buff_data[284]) );
  DFFNEGX1 buff_data_reg_20__8_ ( .D(n2937), .CLK(clk), .Q(buff_data[184]) );
  DFFNEGX1 buff_data_reg_20__7_ ( .D(n2938), .CLK(clk), .Q(buff_data[183]) );
  DFFNEGX1 buff_data_reg_20__6_ ( .D(n2939), .CLK(clk), .Q(buff_data[182]) );
  DFFNEGX1 buff_data_reg_20__5_ ( .D(n2940), .CLK(clk), .Q(buff_data[181]) );
  DFFNEGX1 buff_data_reg_20__4_ ( .D(n2941), .CLK(clk), .Q(buff_data[180]) );
  DFFNEGX1 buff_data_reg_20__3_ ( .D(n2942), .CLK(clk), .Q(buff_data[179]) );
  DFFNEGX1 buff_data_reg_20__2_ ( .D(n1967), .CLK(clk), .Q(buff_data[178]) );
  DFFNEGX1 buff_data_reg_20__1_ ( .D(n1969), .CLK(clk), .Q(buff_data[177]) );
  DFFNEGX1 buff_data_reg_20__0_ ( .D(n1951), .CLK(clk), .Q(buff_data[176]) );
  DFFNEGX1 buff_data_reg_20__15_ ( .D(n2946), .CLK(clk), .Q(buff_data[191]) );
  DFFNEGX1 buff_data_reg_20__14_ ( .D(n2947), .CLK(clk), .Q(buff_data[190]) );
  DFFNEGX1 buff_data_reg_20__13_ ( .D(n2948), .CLK(clk), .Q(buff_data[189]) );
  DFFNEGX1 buff_data_reg_20__12_ ( .D(n2949), .CLK(clk), .Q(buff_data[188]) );
  DFFNEGX1 buff_data_reg_20__11_ ( .D(n2950), .CLK(clk), .Q(buff_data[187]) );
  DFFNEGX1 buff_data_reg_20__10_ ( .D(n2145), .CLK(clk), .Q(buff_data[186]) );
  DFFNEGX1 buff_data_reg_20__9_ ( .D(n2952), .CLK(clk), .Q(buff_data[185]) );
  DFFNEGX1 buff_data_reg_26__5_ ( .D(n2171), .CLK(clk), .Q(buff_data[85]) );
  DFFNEGX1 buff_data_reg_26__4_ ( .D(n3037), .CLK(clk), .Q(buff_data[84]) );
  DFFNEGX1 buff_data_reg_26__3_ ( .D(n3038), .CLK(clk), .Q(buff_data[83]) );
  DFFNEGX1 buff_data_reg_26__2_ ( .D(n3039), .CLK(clk), .Q(buff_data[82]) );
  DFFNEGX1 buff_data_reg_26__1_ ( .D(n3040), .CLK(clk), .Q(buff_data[81]) );
  DFFNEGX1 buff_data_reg_26__0_ ( .D(n3041), .CLK(clk), .Q(buff_data[80]) );
  DFFNEGX1 buff_data_reg_26__15_ ( .D(n3042), .CLK(clk), .Q(buff_data[95]) );
  DFFNEGX1 buff_data_reg_26__14_ ( .D(n3043), .CLK(clk), .Q(buff_data[94]) );
  DFFNEGX1 buff_data_reg_26__13_ ( .D(n3044), .CLK(clk), .Q(buff_data[93]) );
  DFFNEGX1 buff_data_reg_26__12_ ( .D(n3045), .CLK(clk), .Q(buff_data[92]) );
  DFFNEGX1 buff_data_reg_26__11_ ( .D(n3046), .CLK(clk), .Q(buff_data[91]) );
  DFFNEGX1 buff_data_reg_26__10_ ( .D(n3047), .CLK(clk), .Q(buff_data[90]) );
  DFFNEGX1 buff_data_reg_26__9_ ( .D(n3048), .CLK(clk), .Q(buff_data[89]) );
  DFFNEGX1 buff_data_reg_26__8_ ( .D(n3049), .CLK(clk), .Q(buff_data[88]) );
  DFFNEGX1 buff_data_reg_26__7_ ( .D(n3050), .CLK(clk), .Q(buff_data[87]) );
  DFFNEGX1 buff_data_reg_26__6_ ( .D(n3051), .CLK(clk), .Q(buff_data[86]) );
  DFFNEGX1 buff_data_reg_0__15_ ( .D(n2617), .CLK(clk), .Q(buff_data[511]) );
  DFFNEGX1 buff_data_reg_0__14_ ( .D(n2618), .CLK(clk), .Q(buff_data[510]) );
  DFFNEGX1 buff_data_reg_0__13_ ( .D(n2619), .CLK(clk), .Q(buff_data[509]) );
  DFFNEGX1 buff_data_reg_0__12_ ( .D(n2620), .CLK(clk), .Q(buff_data[508]) );
  DFFNEGX1 buff_data_reg_0__11_ ( .D(n2621), .CLK(clk), .Q(buff_data[507]) );
  DFFNEGX1 buff_data_reg_0__10_ ( .D(n2622), .CLK(clk), .Q(buff_data[506]) );
  DFFNEGX1 buff_data_reg_0__9_ ( .D(n2623), .CLK(clk), .Q(buff_data[505]) );
  DFFNEGX1 buff_data_reg_0__8_ ( .D(n2624), .CLK(clk), .Q(buff_data[504]) );
  DFFNEGX1 buff_data_reg_0__7_ ( .D(n2625), .CLK(clk), .Q(buff_data[503]) );
  DFFNEGX1 buff_data_reg_0__6_ ( .D(n2626), .CLK(clk), .Q(buff_data[502]) );
  DFFNEGX1 buff_data_reg_0__5_ ( .D(n2627), .CLK(clk), .Q(buff_data[501]) );
  DFFNEGX1 buff_data_reg_0__4_ ( .D(n2628), .CLK(clk), .Q(buff_data[500]) );
  DFFNEGX1 buff_data_reg_0__3_ ( .D(n2118), .CLK(clk), .Q(buff_data[499]) );
  DFFNEGX1 buff_data_reg_0__2_ ( .D(n2630), .CLK(clk), .Q(buff_data[498]) );
  DFFNEGX1 buff_data_reg_0__1_ ( .D(n2631), .CLK(clk), .Q(buff_data[497]) );
  DFFNEGX1 buff_data_reg_0__0_ ( .D(n2632), .CLK(clk), .Q(buff_data[496]) );
  DFFNEGX1 buff_data_reg_2__15_ ( .D(n2649), .CLK(clk), .Q(buff_data[479]) );
  DFFNEGX1 buff_data_reg_2__14_ ( .D(n2650), .CLK(clk), .Q(buff_data[478]) );
  DFFNEGX1 buff_data_reg_2__13_ ( .D(n2651), .CLK(clk), .Q(buff_data[477]) );
  DFFNEGX1 buff_data_reg_2__12_ ( .D(n1900), .CLK(clk), .Q(buff_data[476]) );
  DFFNEGX1 buff_data_reg_2__11_ ( .D(n2653), .CLK(clk), .Q(buff_data[475]) );
  DFFNEGX1 buff_data_reg_2__10_ ( .D(n2654), .CLK(clk), .Q(buff_data[474]) );
  DFFNEGX1 buff_data_reg_2__9_ ( .D(n1955), .CLK(clk), .Q(buff_data[473]) );
  DFFNEGX1 buff_data_reg_2__8_ ( .D(n2656), .CLK(clk), .Q(buff_data[472]) );
  DFFNEGX1 buff_data_reg_2__7_ ( .D(n2657), .CLK(clk), .Q(buff_data[471]) );
  DFFNEGX1 buff_data_reg_2__6_ ( .D(n2658), .CLK(clk), .Q(buff_data[470]) );
  DFFNEGX1 buff_data_reg_2__5_ ( .D(n2659), .CLK(clk), .Q(buff_data[469]) );
  DFFNEGX1 buff_data_reg_2__4_ ( .D(n2660), .CLK(clk), .Q(buff_data[468]) );
  DFFNEGX1 buff_data_reg_2__3_ ( .D(n2122), .CLK(clk), .Q(buff_data[467]) );
  DFFNEGX1 buff_data_reg_2__2_ ( .D(n2662), .CLK(clk), .Q(buff_data[466]) );
  DFFNEGX1 buff_data_reg_2__1_ ( .D(n2663), .CLK(clk), .Q(buff_data[465]) );
  DFFNEGX1 buff_data_reg_2__0_ ( .D(n2664), .CLK(clk), .Q(buff_data[464]) );
  DFFNEGX1 buff_data_reg_3__15_ ( .D(n2665), .CLK(clk), .Q(buff_data[463]) );
  DFFNEGX1 buff_data_reg_3__14_ ( .D(n2666), .CLK(clk), .Q(buff_data[462]) );
  DFFNEGX1 buff_data_reg_3__13_ ( .D(n2667), .CLK(clk), .Q(buff_data[461]) );
  DFFNEGX1 buff_data_reg_3__12_ ( .D(n2668), .CLK(clk), .Q(buff_data[460]) );
  DFFNEGX1 buff_data_reg_3__11_ ( .D(n2669), .CLK(clk), .Q(buff_data[459]) );
  DFFNEGX1 buff_data_reg_3__10_ ( .D(n2670), .CLK(clk), .Q(buff_data[458]) );
  DFFNEGX1 buff_data_reg_3__9_ ( .D(n1989), .CLK(clk), .Q(buff_data[457]) );
  DFFNEGX1 buff_data_reg_3__8_ ( .D(n2672), .CLK(clk), .Q(buff_data[456]) );
  DFFNEGX1 buff_data_reg_3__7_ ( .D(n2673), .CLK(clk), .Q(buff_data[455]) );
  DFFNEGX1 buff_data_reg_3__6_ ( .D(n2674), .CLK(clk), .Q(buff_data[454]) );
  DFFNEGX1 buff_data_reg_3__5_ ( .D(n2675), .CLK(clk), .Q(buff_data[453]) );
  DFFNEGX1 buff_data_reg_3__4_ ( .D(n2676), .CLK(clk), .Q(buff_data[452]) );
  DFFNEGX1 buff_data_reg_3__3_ ( .D(n2677), .CLK(clk), .Q(buff_data[451]) );
  DFFNEGX1 buff_data_reg_3__2_ ( .D(n2678), .CLK(clk), .Q(buff_data[450]) );
  DFFNEGX1 buff_data_reg_3__1_ ( .D(n2679), .CLK(clk), .Q(buff_data[449]) );
  DFFNEGX1 buff_data_reg_3__0_ ( .D(n2680), .CLK(clk), .Q(buff_data[448]) );
  DFFNEGX1 buff_data_reg_4__15_ ( .D(n2681), .CLK(clk), .Q(buff_data[447]) );
  DFFNEGX1 buff_data_reg_4__14_ ( .D(n2682), .CLK(clk), .Q(buff_data[446]) );
  DFFNEGX1 buff_data_reg_4__13_ ( .D(n2683), .CLK(clk), .Q(buff_data[445]) );
  DFFNEGX1 buff_data_reg_4__12_ ( .D(n2684), .CLK(clk), .Q(buff_data[444]) );
  DFFNEGX1 buff_data_reg_4__11_ ( .D(n2685), .CLK(clk), .Q(buff_data[443]) );
  DFFNEGX1 buff_data_reg_4__10_ ( .D(n2686), .CLK(clk), .Q(buff_data[442]) );
  DFFNEGX1 buff_data_reg_4__9_ ( .D(n2687), .CLK(clk), .Q(buff_data[441]) );
  DFFNEGX1 buff_data_reg_4__8_ ( .D(n2688), .CLK(clk), .Q(buff_data[440]) );
  DFFNEGX1 buff_data_reg_4__7_ ( .D(n2689), .CLK(clk), .Q(buff_data[439]) );
  DFFNEGX1 buff_data_reg_4__6_ ( .D(n2690), .CLK(clk), .Q(buff_data[438]) );
  DFFNEGX1 buff_data_reg_4__5_ ( .D(n2691), .CLK(clk), .Q(buff_data[437]) );
  DFFNEGX1 buff_data_reg_4__4_ ( .D(n2692), .CLK(clk), .Q(buff_data[436]) );
  DFFNEGX1 buff_data_reg_4__3_ ( .D(n2693), .CLK(clk), .Q(buff_data[435]) );
  DFFNEGX1 buff_data_reg_4__2_ ( .D(n2694), .CLK(clk), .Q(buff_data[434]) );
  DFFNEGX1 buff_data_reg_4__1_ ( .D(n2695), .CLK(clk), .Q(buff_data[433]) );
  DFFNEGX1 buff_data_reg_4__0_ ( .D(n2696), .CLK(clk), .Q(buff_data[432]) );
  DFFNEGX1 buff_data_reg_5__15_ ( .D(n2697), .CLK(clk), .Q(buff_data[431]) );
  DFFNEGX1 buff_data_reg_5__14_ ( .D(n2698), .CLK(clk), .Q(buff_data[430]) );
  DFFNEGX1 buff_data_reg_5__13_ ( .D(n2699), .CLK(clk), .Q(buff_data[429]) );
  DFFNEGX1 buff_data_reg_5__12_ ( .D(n2700), .CLK(clk), .Q(buff_data[428]) );
  DFFNEGX1 buff_data_reg_5__11_ ( .D(n2701), .CLK(clk), .Q(buff_data[427]) );
  DFFNEGX1 buff_data_reg_5__10_ ( .D(n2702), .CLK(clk), .Q(buff_data[426]) );
  DFFNEGX1 buff_data_reg_5__9_ ( .D(n2703), .CLK(clk), .Q(buff_data[425]) );
  DFFNEGX1 buff_data_reg_5__8_ ( .D(n2704), .CLK(clk), .Q(buff_data[424]) );
  DFFNEGX1 buff_data_reg_5__7_ ( .D(n2705), .CLK(clk), .Q(buff_data[423]) );
  DFFNEGX1 buff_data_reg_5__6_ ( .D(n2058), .CLK(clk), .Q(buff_data[422]) );
  DFFNEGX1 buff_data_reg_5__5_ ( .D(n2707), .CLK(clk), .Q(buff_data[421]) );
  DFFNEGX1 buff_data_reg_5__4_ ( .D(n2708), .CLK(clk), .Q(buff_data[420]) );
  DFFNEGX1 buff_data_reg_5__3_ ( .D(n2709), .CLK(clk), .Q(buff_data[419]) );
  DFFNEGX1 buff_data_reg_5__2_ ( .D(n2710), .CLK(clk), .Q(buff_data[418]) );
  DFFNEGX1 buff_data_reg_5__1_ ( .D(n2711), .CLK(clk), .Q(buff_data[417]) );
  DFFNEGX1 buff_data_reg_5__0_ ( .D(n1979), .CLK(clk), .Q(buff_data[416]) );
  DFFNEGX1 buff_data_reg_6__15_ ( .D(n2713), .CLK(clk), .Q(buff_data[415]) );
  DFFNEGX1 buff_data_reg_6__14_ ( .D(n1954), .CLK(clk), .Q(buff_data[414]) );
  DFFNEGX1 buff_data_reg_6__13_ ( .D(n2715), .CLK(clk), .Q(buff_data[413]) );
  DFFNEGX1 buff_data_reg_6__12_ ( .D(n2716), .CLK(clk), .Q(buff_data[412]) );
  DFFNEGX1 buff_data_reg_6__11_ ( .D(n2717), .CLK(clk), .Q(buff_data[411]) );
  DFFNEGX1 buff_data_reg_6__10_ ( .D(n2718), .CLK(clk), .Q(buff_data[410]) );
  DFFNEGX1 buff_data_reg_6__9_ ( .D(n2719), .CLK(clk), .Q(buff_data[409]) );
  DFFNEGX1 buff_data_reg_6__8_ ( .D(n2720), .CLK(clk), .Q(buff_data[408]) );
  DFFNEGX1 buff_data_reg_6__7_ ( .D(n2721), .CLK(clk), .Q(buff_data[407]) );
  DFFNEGX1 buff_data_reg_6__6_ ( .D(n2722), .CLK(clk), .Q(buff_data[406]) );
  DFFNEGX1 buff_data_reg_6__5_ ( .D(n1905), .CLK(clk), .Q(buff_data[405]) );
  DFFNEGX1 buff_data_reg_6__4_ ( .D(n2724), .CLK(clk), .Q(buff_data[404]) );
  DFFNEGX1 buff_data_reg_6__3_ ( .D(n2725), .CLK(clk), .Q(buff_data[403]) );
  DFFNEGX1 buff_data_reg_6__2_ ( .D(n2124), .CLK(clk), .Q(buff_data[402]) );
  DFFNEGX1 buff_data_reg_6__1_ ( .D(n2727), .CLK(clk), .Q(buff_data[401]) );
  DFFNEGX1 buff_data_reg_6__0_ ( .D(n2728), .CLK(clk), .Q(buff_data[400]) );
  DFFNEGX1 buff_data_reg_7__15_ ( .D(n2729), .CLK(clk), .Q(buff_data[399]) );
  DFFNEGX1 buff_data_reg_7__14_ ( .D(n2730), .CLK(clk), .Q(buff_data[398]) );
  DFFNEGX1 buff_data_reg_7__13_ ( .D(n2731), .CLK(clk), .Q(buff_data[397]) );
  DFFNEGX1 buff_data_reg_7__12_ ( .D(n2732), .CLK(clk), .Q(buff_data[396]) );
  DFFNEGX1 buff_data_reg_7__11_ ( .D(n2733), .CLK(clk), .Q(buff_data[395]) );
  DFFNEGX1 buff_data_reg_7__10_ ( .D(n2734), .CLK(clk), .Q(buff_data[394]) );
  DFFNEGX1 buff_data_reg_7__9_ ( .D(n2735), .CLK(clk), .Q(buff_data[393]) );
  DFFNEGX1 buff_data_reg_7__8_ ( .D(n2736), .CLK(clk), .Q(buff_data[392]) );
  DFFNEGX1 buff_data_reg_7__7_ ( .D(n2737), .CLK(clk), .Q(buff_data[391]) );
  DFFNEGX1 buff_data_reg_7__6_ ( .D(n2738), .CLK(clk), .Q(buff_data[390]) );
  DFFNEGX1 buff_data_reg_7__5_ ( .D(n2739), .CLK(clk), .Q(buff_data[389]) );
  DFFNEGX1 buff_data_reg_7__4_ ( .D(n2740), .CLK(clk), .Q(buff_data[388]) );
  DFFNEGX1 buff_data_reg_7__3_ ( .D(n2741), .CLK(clk), .Q(buff_data[387]) );
  DFFNEGX1 buff_data_reg_7__2_ ( .D(n2742), .CLK(clk), .Q(buff_data[386]) );
  DFFNEGX1 buff_data_reg_7__1_ ( .D(n2743), .CLK(clk), .Q(buff_data[385]) );
  DFFNEGX1 buff_data_reg_7__0_ ( .D(n2744), .CLK(clk), .Q(buff_data[384]) );
  DFFNEGX1 buff_data_reg_9__15_ ( .D(n2761), .CLK(clk), .Q(buff_data[367]) );
  DFFNEGX1 buff_data_reg_9__14_ ( .D(n1902), .CLK(clk), .Q(buff_data[366]) );
  DFFNEGX1 buff_data_reg_9__13_ ( .D(n2763), .CLK(clk), .Q(buff_data[365]) );
  DFFNEGX1 buff_data_reg_9__12_ ( .D(n2764), .CLK(clk), .Q(buff_data[364]) );
  DFFNEGX1 buff_data_reg_9__11_ ( .D(n2765), .CLK(clk), .Q(buff_data[363]) );
  DFFNEGX1 buff_data_reg_9__10_ ( .D(n2766), .CLK(clk), .Q(buff_data[362]) );
  DFFNEGX1 buff_data_reg_9__9_ ( .D(n2767), .CLK(clk), .Q(buff_data[361]) );
  DFFNEGX1 buff_data_reg_9__8_ ( .D(n2768), .CLK(clk), .Q(buff_data[360]) );
  DFFNEGX1 buff_data_reg_9__7_ ( .D(n2769), .CLK(clk), .Q(buff_data[359]) );
  DFFNEGX1 buff_data_reg_9__6_ ( .D(n2023), .CLK(clk), .Q(buff_data[358]) );
  DFFNEGX1 buff_data_reg_9__5_ ( .D(n2771), .CLK(clk), .Q(buff_data[357]) );
  DFFNEGX1 buff_data_reg_9__4_ ( .D(n2772), .CLK(clk), .Q(buff_data[356]) );
  DFFNEGX1 buff_data_reg_9__3_ ( .D(n2773), .CLK(clk), .Q(buff_data[355]) );
  DFFNEGX1 buff_data_reg_9__2_ ( .D(n2774), .CLK(clk), .Q(buff_data[354]) );
  DFFNEGX1 buff_data_reg_9__1_ ( .D(n2775), .CLK(clk), .Q(buff_data[353]) );
  DFFNEGX1 buff_data_reg_9__0_ ( .D(n2137), .CLK(clk), .Q(buff_data[352]) );
  DFFNEGX1 buff_data_reg_10__15_ ( .D(n2777), .CLK(clk), .Q(buff_data[351]) );
  DFFNEGX1 buff_data_reg_10__14_ ( .D(n2778), .CLK(clk), .Q(buff_data[350]) );
  DFFNEGX1 buff_data_reg_10__13_ ( .D(n2779), .CLK(clk), .Q(buff_data[349]) );
  DFFNEGX1 buff_data_reg_10__12_ ( .D(n2780), .CLK(clk), .Q(buff_data[348]) );
  DFFNEGX1 buff_data_reg_10__11_ ( .D(n2781), .CLK(clk), .Q(buff_data[347]) );
  DFFNEGX1 buff_data_reg_10__10_ ( .D(n2782), .CLK(clk), .Q(buff_data[346]) );
  DFFNEGX1 buff_data_reg_10__9_ ( .D(n2783), .CLK(clk), .Q(buff_data[345]) );
  DFFNEGX1 buff_data_reg_10__8_ ( .D(n2784), .CLK(clk), .Q(buff_data[344]) );
  DFFNEGX1 buff_data_reg_10__7_ ( .D(n2785), .CLK(clk), .Q(buff_data[343]) );
  DFFNEGX1 buff_data_reg_10__6_ ( .D(n2786), .CLK(clk), .Q(buff_data[342]) );
  DFFNEGX1 buff_data_reg_10__5_ ( .D(n2787), .CLK(clk), .Q(buff_data[341]) );
  DFFNEGX1 buff_data_reg_10__4_ ( .D(n2788), .CLK(clk), .Q(buff_data[340]) );
  DFFNEGX1 buff_data_reg_10__3_ ( .D(n2789), .CLK(clk), .Q(buff_data[339]) );
  DFFNEGX1 buff_data_reg_10__2_ ( .D(n2790), .CLK(clk), .Q(buff_data[338]) );
  DFFNEGX1 buff_data_reg_10__1_ ( .D(n2791), .CLK(clk), .Q(buff_data[337]) );
  DFFNEGX1 buff_data_reg_10__0_ ( .D(n2792), .CLK(clk), .Q(buff_data[336]) );
  DFFNEGX1 buff_data_reg_11__15_ ( .D(n2793), .CLK(clk), .Q(buff_data[335]) );
  DFFNEGX1 buff_data_reg_11__14_ ( .D(n2794), .CLK(clk), .Q(buff_data[334]) );
  DFFNEGX1 buff_data_reg_11__13_ ( .D(n1984), .CLK(clk), .Q(buff_data[333]) );
  DFFNEGX1 buff_data_reg_11__12_ ( .D(n2796), .CLK(clk), .Q(buff_data[332]) );
  DFFNEGX1 buff_data_reg_11__11_ ( .D(n1907), .CLK(clk), .Q(buff_data[331]) );
  DFFNEGX1 buff_data_reg_11__10_ ( .D(n2798), .CLK(clk), .Q(buff_data[330]) );
  DFFNEGX1 buff_data_reg_11__9_ ( .D(n2799), .CLK(clk), .Q(buff_data[329]) );
  DFFNEGX1 buff_data_reg_11__8_ ( .D(n2008), .CLK(clk), .Q(buff_data[328]) );
  DFFNEGX1 buff_data_reg_11__7_ ( .D(n2801), .CLK(clk), .Q(buff_data[327]) );
  DFFNEGX1 buff_data_reg_11__6_ ( .D(n2802), .CLK(clk), .Q(buff_data[326]) );
  DFFNEGX1 buff_data_reg_11__5_ ( .D(n2803), .CLK(clk), .Q(buff_data[325]) );
  DFFNEGX1 buff_data_reg_11__4_ ( .D(n2804), .CLK(clk), .Q(buff_data[324]) );
  DFFNEGX1 buff_data_reg_11__3_ ( .D(n2133), .CLK(clk), .Q(buff_data[323]) );
  DFFNEGX1 buff_data_reg_11__2_ ( .D(n2806), .CLK(clk), .Q(buff_data[322]) );
  DFFNEGX1 buff_data_reg_11__1_ ( .D(n2807), .CLK(clk), .Q(buff_data[321]) );
  DFFNEGX1 buff_data_reg_11__0_ ( .D(n2808), .CLK(clk), .Q(buff_data[320]) );
  DFFNEGX1 buff_data_reg_12__15_ ( .D(n2175), .CLK(clk), .Q(buff_data[319]) );
  DFFNEGX1 buff_data_reg_12__14_ ( .D(n2810), .CLK(clk), .Q(buff_data[318]) );
  DFFNEGX1 buff_data_reg_12__13_ ( .D(n2811), .CLK(clk), .Q(buff_data[317]) );
  DFFNEGX1 buff_data_reg_12__12_ ( .D(n2003), .CLK(clk), .Q(buff_data[316]) );
  DFFNEGX1 buff_data_reg_12__11_ ( .D(n2017), .CLK(clk), .Q(buff_data[315]) );
  DFFNEGX1 buff_data_reg_12__10_ ( .D(n2814), .CLK(clk), .Q(buff_data[314]) );
  DFFNEGX1 buff_data_reg_12__9_ ( .D(n2815), .CLK(clk), .Q(buff_data[313]) );
  DFFNEGX1 buff_data_reg_12__8_ ( .D(n2816), .CLK(clk), .Q(buff_data[312]) );
  DFFNEGX1 buff_data_reg_12__7_ ( .D(n2019), .CLK(clk), .Q(buff_data[311]) );
  DFFNEGX1 buff_data_reg_12__6_ ( .D(n2818), .CLK(clk), .Q(buff_data[310]) );
  DFFNEGX1 buff_data_reg_12__5_ ( .D(n2819), .CLK(clk), .Q(buff_data[309]) );
  DFFNEGX1 buff_data_reg_12__4_ ( .D(n2820), .CLK(clk), .Q(buff_data[308]) );
  DFFNEGX1 buff_data_reg_12__3_ ( .D(n2821), .CLK(clk), .Q(buff_data[307]) );
  DFFNEGX1 buff_data_reg_12__2_ ( .D(n2822), .CLK(clk), .Q(buff_data[306]) );
  DFFNEGX1 buff_data_reg_12__1_ ( .D(n2823), .CLK(clk), .Q(buff_data[305]) );
  DFFNEGX1 buff_data_reg_12__0_ ( .D(n2824), .CLK(clk), .Q(buff_data[304]) );
  DFFNEGX1 buff_data_reg_13__15_ ( .D(n2825), .CLK(clk), .Q(buff_data[303]) );
  DFFNEGX1 buff_data_reg_13__14_ ( .D(n2826), .CLK(clk), .Q(buff_data[302]) );
  DFFNEGX1 buff_data_reg_13__13_ ( .D(n1986), .CLK(clk), .Q(buff_data[301]) );
  DFFNEGX1 buff_data_reg_13__12_ ( .D(n2828), .CLK(clk), .Q(buff_data[300]) );
  DFFNEGX1 buff_data_reg_13__11_ ( .D(n2829), .CLK(clk), .Q(buff_data[299]) );
  DFFNEGX1 buff_data_reg_13__10_ ( .D(n2830), .CLK(clk), .Q(buff_data[298]) );
  DFFNEGX1 buff_data_reg_13__9_ ( .D(n2831), .CLK(clk), .Q(buff_data[297]) );
  DFFNEGX1 buff_data_reg_13__8_ ( .D(n2832), .CLK(clk), .Q(buff_data[296]) );
  DFFNEGX1 buff_data_reg_13__7_ ( .D(n2010), .CLK(clk), .Q(buff_data[295]) );
  DFFNEGX1 buff_data_reg_13__6_ ( .D(n2834), .CLK(clk), .Q(buff_data[294]) );
  DFFNEGX1 buff_data_reg_13__5_ ( .D(n2835), .CLK(clk), .Q(buff_data[293]) );
  DFFNEGX1 buff_data_reg_13__4_ ( .D(n2836), .CLK(clk), .Q(buff_data[292]) );
  DFFNEGX1 buff_data_reg_13__3_ ( .D(n2837), .CLK(clk), .Q(buff_data[291]) );
  DFFNEGX1 buff_data_reg_13__2_ ( .D(n2838), .CLK(clk), .Q(buff_data[290]) );
  DFFNEGX1 buff_data_reg_13__1_ ( .D(n2839), .CLK(clk), .Q(buff_data[289]) );
  DFFNEGX1 buff_data_reg_13__0_ ( .D(n2135), .CLK(clk), .Q(buff_data[288]) );
  DFFNEGX1 buff_data_reg_15__15_ ( .D(n2857), .CLK(clk), .Q(buff_data[271]) );
  DFFNEGX1 buff_data_reg_15__14_ ( .D(n2858), .CLK(clk), .Q(buff_data[270]) );
  DFFNEGX1 buff_data_reg_15__13_ ( .D(n2859), .CLK(clk), .Q(buff_data[269]) );
  DFFNEGX1 buff_data_reg_15__12_ ( .D(n2860), .CLK(clk), .Q(buff_data[268]) );
  DFFNEGX1 buff_data_reg_15__11_ ( .D(n2861), .CLK(clk), .Q(buff_data[267]) );
  DFFNEGX1 buff_data_reg_15__10_ ( .D(n2862), .CLK(clk), .Q(buff_data[266]) );
  DFFNEGX1 buff_data_reg_15__9_ ( .D(n2863), .CLK(clk), .Q(buff_data[265]) );
  DFFNEGX1 buff_data_reg_15__8_ ( .D(n2864), .CLK(clk), .Q(buff_data[264]) );
  DFFNEGX1 buff_data_reg_15__7_ ( .D(n2865), .CLK(clk), .Q(buff_data[263]) );
  DFFNEGX1 buff_data_reg_15__6_ ( .D(n2866), .CLK(clk), .Q(buff_data[262]) );
  DFFNEGX1 buff_data_reg_15__5_ ( .D(n2867), .CLK(clk), .Q(buff_data[261]) );
  DFFNEGX1 buff_data_reg_15__4_ ( .D(n2868), .CLK(clk), .Q(buff_data[260]) );
  DFFNEGX1 buff_data_reg_15__3_ ( .D(n2869), .CLK(clk), .Q(buff_data[259]) );
  DFFNEGX1 buff_data_reg_15__2_ ( .D(n2870), .CLK(clk), .Q(buff_data[258]) );
  DFFNEGX1 buff_data_reg_15__1_ ( .D(n2871), .CLK(clk), .Q(buff_data[257]) );
  DFFNEGX1 buff_data_reg_15__0_ ( .D(n2872), .CLK(clk), .Q(buff_data[256]) );
  DFFNEGX1 buff_data_reg_16__15_ ( .D(n1919), .CLK(clk), .Q(buff_data[255]) );
  DFFNEGX1 buff_data_reg_16__14_ ( .D(n2874), .CLK(clk), .Q(buff_data[254]) );
  DFFNEGX1 buff_data_reg_16__13_ ( .D(net80914), .CLK(clk), .Q(buff_data[253])
         );
  DFFNEGX1 buff_data_reg_16__12_ ( .D(n2876), .CLK(clk), .Q(buff_data[252]) );
  DFFNEGX1 buff_data_reg_16__11_ ( .D(n2877), .CLK(clk), .Q(buff_data[251]) );
  DFFNEGX1 buff_data_reg_16__10_ ( .D(n1958), .CLK(clk), .Q(buff_data[250]) );
  DFFNEGX1 buff_data_reg_16__9_ ( .D(n2879), .CLK(clk), .Q(buff_data[249]) );
  DFFNEGX1 buff_data_reg_16__8_ ( .D(n2880), .CLK(clk), .Q(buff_data[248]) );
  DFFNEGX1 buff_data_reg_16__7_ ( .D(n2881), .CLK(clk), .Q(buff_data[247]) );
  DFFNEGX1 buff_data_reg_16__6_ ( .D(n2882), .CLK(clk), .Q(buff_data[246]) );
  DFFNEGX1 buff_data_reg_16__5_ ( .D(n2883), .CLK(clk), .Q(buff_data[245]) );
  DFFNEGX1 buff_data_reg_16__4_ ( .D(n1913), .CLK(clk), .Q(buff_data[244]) );
  DFFNEGX1 buff_data_reg_16__3_ ( .D(n2885), .CLK(clk), .Q(buff_data[243]) );
  DFFNEGX1 buff_data_reg_16__2_ ( .D(n2147), .CLK(clk), .Q(buff_data[242]) );
  DFFNEGX1 buff_data_reg_16__1_ ( .D(n2887), .CLK(clk), .Q(buff_data[241]) );
  DFFNEGX1 buff_data_reg_16__0_ ( .D(n2888), .CLK(clk), .Q(buff_data[240]) );
  DFFNEGX1 buff_data_reg_17__15_ ( .D(n2889), .CLK(clk), .Q(buff_data[239]) );
  DFFNEGX1 buff_data_reg_17__14_ ( .D(n1949), .CLK(clk), .Q(buff_data[238]) );
  DFFNEGX1 buff_data_reg_17__13_ ( .D(n2031), .CLK(clk), .Q(buff_data[237]) );
  DFFNEGX1 buff_data_reg_17__12_ ( .D(n2042), .CLK(clk), .Q(buff_data[236]) );
  DFFNEGX1 buff_data_reg_17__11_ ( .D(n2065), .CLK(clk), .Q(buff_data[235]) );
  DFFNEGX1 buff_data_reg_17__10_ ( .D(n1932), .CLK(clk), .Q(buff_data[234]) );
  DFFNEGX1 buff_data_reg_17__9_ ( .D(n1934), .CLK(clk), .Q(buff_data[233]) );
  DFFNEGX1 buff_data_reg_17__8_ ( .D(n2033), .CLK(clk), .Q(buff_data[232]) );
  DFFNEGX1 buff_data_reg_17__7_ ( .D(n2045), .CLK(clk), .Q(buff_data[231]) );
  DFFNEGX1 buff_data_reg_17__6_ ( .D(n2054), .CLK(clk), .Q(buff_data[230]) );
  DFFNEGX1 buff_data_reg_17__5_ ( .D(n2061), .CLK(clk), .Q(buff_data[229]) );
  DFFNEGX1 buff_data_reg_17__4_ ( .D(n2900), .CLK(clk), .Q(buff_data[228]) );
  DFFNEGX1 buff_data_reg_17__3_ ( .D(n2901), .CLK(clk), .Q(buff_data[227]) );
  DFFNEGX1 buff_data_reg_17__2_ ( .D(n2152), .CLK(clk), .Q(buff_data[226]) );
  DFFNEGX1 buff_data_reg_17__1_ ( .D(n1943), .CLK(clk), .Q(buff_data[225]) );
  DFFNEGX1 buff_data_reg_17__0_ ( .D(n2904), .CLK(clk), .Q(buff_data[224]) );
  DFFNEGX1 buff_data_reg_18__15_ ( .D(n2905), .CLK(clk), .Q(buff_data[223]) );
  DFFNEGX1 buff_data_reg_18__14_ ( .D(n2906), .CLK(clk), .Q(buff_data[222]) );
  DFFNEGX1 buff_data_reg_18__13_ ( .D(n2907), .CLK(clk), .Q(buff_data[221]) );
  DFFNEGX1 buff_data_reg_18__12_ ( .D(n2908), .CLK(clk), .Q(buff_data[220]) );
  DFFNEGX1 buff_data_reg_18__11_ ( .D(n2909), .CLK(clk), .Q(buff_data[219]) );
  DFFNEGX1 buff_data_reg_18__10_ ( .D(n2910), .CLK(clk), .Q(buff_data[218]) );
  DFFNEGX1 buff_data_reg_18__9_ ( .D(n2911), .CLK(clk), .Q(buff_data[217]) );
  DFFNEGX1 buff_data_reg_18__8_ ( .D(n2912), .CLK(clk), .Q(buff_data[216]) );
  DFFNEGX1 buff_data_reg_18__7_ ( .D(n2913), .CLK(clk), .Q(buff_data[215]) );
  DFFNEGX1 buff_data_reg_18__6_ ( .D(n2914), .CLK(clk), .Q(buff_data[214]) );
  DFFNEGX1 buff_data_reg_18__5_ ( .D(n2915), .CLK(clk), .Q(buff_data[213]) );
  DFFNEGX1 buff_data_reg_18__4_ ( .D(n2916), .CLK(clk), .Q(buff_data[212]) );
  DFFNEGX1 buff_data_reg_18__3_ ( .D(n2917), .CLK(clk), .Q(buff_data[211]) );
  DFFNEGX1 buff_data_reg_18__2_ ( .D(n2918), .CLK(clk), .Q(buff_data[210]) );
  DFFNEGX1 buff_data_reg_18__1_ ( .D(n2919), .CLK(clk), .Q(buff_data[209]) );
  DFFNEGX1 buff_data_reg_18__0_ ( .D(n2920), .CLK(clk), .Q(buff_data[208]) );
  DFFNEGX1 buff_data_reg_19__15_ ( .D(n2921), .CLK(clk), .Q(buff_data[207]) );
  DFFNEGX1 buff_data_reg_19__14_ ( .D(n1948), .CLK(clk), .Q(buff_data[206]) );
  DFFNEGX1 buff_data_reg_19__13_ ( .D(n2923), .CLK(clk), .Q(buff_data[205]) );
  DFFNEGX1 buff_data_reg_19__12_ ( .D(n2924), .CLK(clk), .Q(buff_data[204]) );
  DFFNEGX1 buff_data_reg_19__11_ ( .D(n2067), .CLK(clk), .Q(buff_data[203]) );
  DFFNEGX1 buff_data_reg_19__10_ ( .D(n2926), .CLK(clk), .Q(buff_data[202]) );
  DFFNEGX1 buff_data_reg_19__9_ ( .D(n2927), .CLK(clk), .Q(buff_data[201]) );
  DFFNEGX1 buff_data_reg_19__8_ ( .D(n2928), .CLK(clk), .Q(buff_data[200]) );
  DFFNEGX1 buff_data_reg_19__7_ ( .D(n1923), .CLK(clk), .Q(buff_data[199]) );
  DFFNEGX1 buff_data_reg_19__6_ ( .D(n2050), .CLK(clk), .Q(buff_data[198]) );
  DFFNEGX1 buff_data_reg_19__5_ ( .D(n2063), .CLK(clk), .Q(buff_data[197]) );
  DFFNEGX1 buff_data_reg_19__4_ ( .D(n2056), .CLK(clk), .Q(buff_data[196]) );
  DFFNEGX1 buff_data_reg_19__3_ ( .D(n1926), .CLK(clk), .Q(buff_data[195]) );
  DFFNEGX1 buff_data_reg_19__2_ ( .D(n2934), .CLK(clk), .Q(buff_data[194]) );
  DFFNEGX1 buff_data_reg_19__1_ ( .D(n2154), .CLK(clk), .Q(buff_data[193]) );
  DFFNEGX1 buff_data_reg_19__0_ ( .D(n2936), .CLK(clk), .Q(buff_data[192]) );
  DFFNEGX1 buff_data_reg_21__15_ ( .D(n2953), .CLK(clk), .Q(buff_data[175]) );
  DFFNEGX1 buff_data_reg_21__14_ ( .D(n2954), .CLK(clk), .Q(buff_data[174]) );
  DFFNEGX1 buff_data_reg_21__13_ ( .D(n1915), .CLK(clk), .Q(buff_data[173]) );
  DFFNEGX1 buff_data_reg_21__12_ ( .D(n1946), .CLK(clk), .Q(buff_data[172]) );
  DFFNEGX1 buff_data_reg_21__11_ ( .D(n2957), .CLK(clk), .Q(buff_data[171]) );
  DFFNEGX1 buff_data_reg_21__10_ ( .D(n2069), .CLK(clk), .Q(buff_data[170]) );
  DFFNEGX1 buff_data_reg_21__9_ ( .D(n2959), .CLK(clk), .Q(buff_data[169]) );
  DFFNEGX1 buff_data_reg_21__8_ ( .D(n1917), .CLK(clk), .Q(buff_data[168]) );
  DFFNEGX1 buff_data_reg_21__7_ ( .D(n2961), .CLK(clk), .Q(buff_data[167]) );
  DFFNEGX1 buff_data_reg_21__6_ ( .D(n2962), .CLK(clk), .Q(buff_data[166]) );
  DFFNEGX1 buff_data_reg_21__5_ ( .D(n2963), .CLK(clk), .Q(buff_data[165]) );
  DFFNEGX1 buff_data_reg_21__4_ ( .D(n2964), .CLK(clk), .Q(buff_data[164]) );
  DFFNEGX1 buff_data_reg_21__3_ ( .D(n2025), .CLK(clk), .Q(buff_data[163]) );
  DFFNEGX1 buff_data_reg_21__2_ ( .D(n2966), .CLK(clk), .Q(buff_data[162]) );
  DFFNEGX1 buff_data_reg_21__1_ ( .D(n2157), .CLK(clk), .Q(buff_data[161]) );
  DFFNEGX1 buff_data_reg_21__0_ ( .D(n2968), .CLK(clk), .Q(buff_data[160]) );
  DFFNEGX1 buff_data_reg_22__15_ ( .D(n2969), .CLK(clk), .Q(buff_data[159]) );
  DFFNEGX1 buff_data_reg_22__14_ ( .D(n2970), .CLK(clk), .Q(buff_data[158]) );
  DFFNEGX1 buff_data_reg_22__13_ ( .D(n2971), .CLK(clk), .Q(buff_data[157]) );
  DFFNEGX1 buff_data_reg_22__12_ ( .D(n2972), .CLK(clk), .Q(buff_data[156]) );
  DFFNEGX1 buff_data_reg_22__11_ ( .D(n2973), .CLK(clk), .Q(buff_data[155]) );
  DFFNEGX1 buff_data_reg_22__10_ ( .D(n2071), .CLK(clk), .Q(buff_data[154]) );
  DFFNEGX1 buff_data_reg_22__9_ ( .D(n2975), .CLK(clk), .Q(buff_data[153]) );
  DFFNEGX1 buff_data_reg_22__8_ ( .D(n2976), .CLK(clk), .Q(buff_data[152]) );
  DFFNEGX1 buff_data_reg_22__7_ ( .D(n2977), .CLK(clk), .Q(buff_data[151]) );
  DFFNEGX1 buff_data_reg_22__6_ ( .D(n2978), .CLK(clk), .Q(buff_data[150]) );
  DFFNEGX1 buff_data_reg_22__5_ ( .D(n2979), .CLK(clk), .Q(buff_data[149]) );
  DFFNEGX1 buff_data_reg_22__4_ ( .D(n2980), .CLK(clk), .Q(buff_data[148]) );
  DFFNEGX1 buff_data_reg_22__3_ ( .D(n2981), .CLK(clk), .Q(buff_data[147]) );
  DFFNEGX1 buff_data_reg_22__2_ ( .D(n2982), .CLK(clk), .Q(buff_data[146]) );
  DFFNEGX1 buff_data_reg_22__1_ ( .D(n2149), .CLK(clk), .Q(buff_data[145]) );
  DFFNEGX1 buff_data_reg_22__0_ ( .D(n2984), .CLK(clk), .Q(buff_data[144]) );
  DFFNEGX1 buff_data_reg_23__15_ ( .D(n2985), .CLK(clk), .Q(buff_data[143]) );
  DFFNEGX1 buff_data_reg_23__14_ ( .D(n2986), .CLK(clk), .Q(buff_data[142]) );
  DFFNEGX1 buff_data_reg_23__13_ ( .D(n2987), .CLK(clk), .Q(buff_data[141]) );
  DFFNEGX1 buff_data_reg_23__12_ ( .D(n2988), .CLK(clk), .Q(buff_data[140]) );
  DFFNEGX1 buff_data_reg_23__11_ ( .D(n2989), .CLK(clk), .Q(buff_data[139]) );
  DFFNEGX1 buff_data_reg_23__10_ ( .D(n2990), .CLK(clk), .Q(buff_data[138]) );
  DFFNEGX1 buff_data_reg_23__9_ ( .D(n2991), .CLK(clk), .Q(buff_data[137]) );
  DFFNEGX1 buff_data_reg_23__8_ ( .D(n2992), .CLK(clk), .Q(buff_data[136]) );
  DFFNEGX1 buff_data_reg_23__7_ ( .D(n2993), .CLK(clk), .Q(buff_data[135]) );
  DFFNEGX1 buff_data_reg_23__6_ ( .D(n2994), .CLK(clk), .Q(buff_data[134]) );
  DFFNEGX1 buff_data_reg_23__5_ ( .D(n2995), .CLK(clk), .Q(buff_data[133]) );
  DFFNEGX1 buff_data_reg_23__4_ ( .D(n2996), .CLK(clk), .Q(buff_data[132]) );
  DFFNEGX1 buff_data_reg_23__3_ ( .D(n2998), .CLK(clk), .Q(buff_data[131]) );
  DFFNEGX1 buff_data_reg_23__2_ ( .D(n2999), .CLK(clk), .Q(buff_data[130]) );
  DFFNEGX1 buff_data_reg_23__1_ ( .D(n3000), .CLK(clk), .Q(buff_data[129]) );
  DFFNEGX1 buff_data_reg_23__0_ ( .D(n3001), .CLK(clk), .Q(buff_data[128]) );
  DFFNEGX1 buff_data_reg_24__15_ ( .D(n2166), .CLK(clk), .Q(buff_data[127]) );
  DFFNEGX1 buff_data_reg_24__14_ ( .D(n3003), .CLK(clk), .Q(buff_data[126]) );
  DFFNEGX1 buff_data_reg_24__13_ ( .D(n3004), .CLK(clk), .Q(buff_data[125]) );
  DFFNEGX1 buff_data_reg_24__12_ ( .D(n3005), .CLK(clk), .Q(buff_data[124]) );
  DFFNEGX1 buff_data_reg_24__11_ ( .D(n3006), .CLK(clk), .Q(buff_data[123]) );
  DFFNEGX1 buff_data_reg_24__10_ ( .D(n3007), .CLK(clk), .Q(buff_data[122]) );
  DFFNEGX1 buff_data_reg_24__9_ ( .D(n3008), .CLK(clk), .Q(buff_data[121]) );
  DFFNEGX1 buff_data_reg_24__8_ ( .D(n3009), .CLK(clk), .Q(buff_data[120]) );
  DFFNEGX1 buff_data_reg_24__7_ ( .D(n3010), .CLK(clk), .Q(buff_data[119]) );
  DFFNEGX1 buff_data_reg_24__6_ ( .D(n3011), .CLK(clk), .Q(buff_data[118]) );
  DFFNEGX1 buff_data_reg_24__5_ ( .D(n3012), .CLK(clk), .Q(buff_data[117]) );
  DFFNEGX1 buff_data_reg_24__4_ ( .D(n3013), .CLK(clk), .Q(buff_data[116]) );
  DFFNEGX1 buff_data_reg_24__3_ ( .D(n3014), .CLK(clk), .Q(buff_data[115]) );
  DFFNEGX1 buff_data_reg_24__2_ ( .D(n3015), .CLK(clk), .Q(buff_data[114]) );
  DFFNEGX1 buff_data_reg_24__1_ ( .D(n3016), .CLK(clk), .Q(buff_data[113]) );
  DFFNEGX1 buff_data_reg_24__0_ ( .D(n3017), .CLK(clk), .Q(buff_data[112]) );
  DFFNEGX1 buff_data_reg_25__15_ ( .D(n3018), .CLK(clk), .Q(buff_data[111]) );
  DFFNEGX1 buff_data_reg_25__14_ ( .D(n3019), .CLK(clk), .Q(buff_data[110]) );
  DFFNEGX1 buff_data_reg_25__13_ ( .D(n1821), .CLK(clk), .Q(buff_data[109]) );
  DFFNEGX1 buff_data_reg_25__12_ ( .D(n3021), .CLK(clk), .Q(buff_data[108]) );
  DFFNEGX1 buff_data_reg_25__11_ ( .D(n3022), .CLK(clk), .Q(buff_data[107]) );
  DFFNEGX1 buff_data_reg_25__10_ ( .D(n3023), .CLK(clk), .Q(buff_data[106]) );
  DFFNEGX1 buff_data_reg_25__9_ ( .D(n3024), .CLK(clk), .Q(buff_data[105]) );
  DFFNEGX1 buff_data_reg_25__8_ ( .D(n3025), .CLK(clk), .Q(buff_data[104]) );
  DFFNEGX1 buff_data_reg_25__7_ ( .D(n1826), .CLK(clk), .Q(buff_data[103]) );
  DFFNEGX1 buff_data_reg_25__6_ ( .D(n3027), .CLK(clk), .Q(buff_data[102]) );
  DFFNEGX1 buff_data_reg_25__5_ ( .D(n3028), .CLK(clk), .Q(buff_data[101]) );
  DFFNEGX1 buff_data_reg_25__4_ ( .D(n3029), .CLK(clk), .Q(buff_data[100]) );
  DFFNEGX1 buff_data_reg_25__3_ ( .D(n3031), .CLK(clk), .Q(buff_data[99]) );
  DFFNEGX1 buff_data_reg_25__2_ ( .D(n3032), .CLK(clk), .Q(buff_data[98]) );
  DFFNEGX1 buff_data_reg_25__1_ ( .D(n1830), .CLK(clk), .Q(buff_data[97]) );
  DFFNEGX1 buff_data_reg_25__0_ ( .D(n3034), .CLK(clk), .Q(buff_data[96]) );
  DFFNEGX1 buff_data_reg_27__15_ ( .D(n2165), .CLK(clk), .Q(buff_data[79]) );
  DFFNEGX1 buff_data_reg_27__14_ ( .D(n3053), .CLK(clk), .Q(buff_data[78]) );
  DFFNEGX1 buff_data_reg_27__13_ ( .D(n3054), .CLK(clk), .Q(buff_data[77]) );
  DFFNEGX1 buff_data_reg_27__12_ ( .D(n3055), .CLK(clk), .Q(buff_data[76]) );
  DFFNEGX1 buff_data_reg_27__11_ ( .D(n3056), .CLK(clk), .Q(buff_data[75]) );
  DFFNEGX1 buff_data_reg_27__10_ ( .D(n3057), .CLK(clk), .Q(buff_data[74]) );
  DFFNEGX1 buff_data_reg_27__9_ ( .D(n3058), .CLK(clk), .Q(buff_data[73]) );
  DFFNEGX1 buff_data_reg_27__8_ ( .D(n3059), .CLK(clk), .Q(buff_data[72]) );
  DFFNEGX1 buff_data_reg_27__7_ ( .D(n3060), .CLK(clk), .Q(buff_data[71]) );
  DFFNEGX1 buff_data_reg_27__6_ ( .D(n3061), .CLK(clk), .Q(buff_data[70]) );
  DFFNEGX1 buff_data_reg_27__5_ ( .D(n1964), .CLK(clk), .Q(buff_data[69]) );
  DFFNEGX1 buff_data_reg_27__4_ ( .D(n3063), .CLK(clk), .Q(buff_data[68]) );
  DFFNEGX1 buff_data_reg_27__3_ ( .D(n3064), .CLK(clk), .Q(buff_data[67]) );
  DFFNEGX1 buff_data_reg_27__2_ ( .D(n3065), .CLK(clk), .Q(buff_data[66]) );
  DFFNEGX1 buff_data_reg_27__1_ ( .D(n3066), .CLK(clk), .Q(buff_data[65]) );
  DFFNEGX1 buff_data_reg_27__0_ ( .D(n3067), .CLK(clk), .Q(buff_data[64]) );
  DFFNEGX1 buff_data_reg_28__15_ ( .D(n2168), .CLK(clk), .Q(buff_data[63]) );
  DFFNEGX1 buff_data_reg_28__14_ ( .D(n3069), .CLK(clk), .Q(buff_data[62]) );
  DFFNEGX1 buff_data_reg_28__13_ ( .D(n3070), .CLK(clk), .Q(buff_data[61]) );
  DFFNEGX1 buff_data_reg_28__12_ ( .D(n3071), .CLK(clk), .Q(buff_data[60]) );
  DFFNEGX1 buff_data_reg_28__11_ ( .D(n3072), .CLK(clk), .Q(buff_data[59]) );
  DFFNEGX1 buff_data_reg_28__10_ ( .D(n3075), .CLK(clk), .Q(buff_data[58]) );
  DFFNEGX1 buff_data_reg_28__9_ ( .D(n3076), .CLK(clk), .Q(buff_data[57]) );
  DFFNEGX1 buff_data_reg_28__8_ ( .D(n3077), .CLK(clk), .Q(buff_data[56]) );
  DFFNEGX1 buff_data_reg_28__7_ ( .D(n3078), .CLK(clk), .Q(buff_data[55]) );
  DFFNEGX1 buff_data_reg_28__6_ ( .D(n3080), .CLK(clk), .Q(buff_data[54]) );
  DFFNEGX1 buff_data_reg_28__5_ ( .D(n3081), .CLK(clk), .Q(buff_data[53]) );
  DFFNEGX1 buff_data_reg_28__4_ ( .D(n3082), .CLK(clk), .Q(buff_data[52]) );
  DFFNEGX1 buff_data_reg_28__3_ ( .D(n3083), .CLK(clk), .Q(buff_data[51]) );
  DFFNEGX1 buff_data_reg_28__2_ ( .D(n3084), .CLK(clk), .Q(buff_data[50]) );
  DFFNEGX1 buff_data_reg_28__1_ ( .D(n3085), .CLK(clk), .Q(buff_data[49]) );
  DFFNEGX1 buff_data_reg_28__0_ ( .D(n3086), .CLK(clk), .Q(buff_data[48]) );
  DFFNEGX1 buff_data_reg_29__15_ ( .D(n3087), .CLK(clk), .Q(buff_data[47]) );
  DFFNEGX1 buff_data_reg_29__14_ ( .D(n3088), .CLK(clk), .Q(buff_data[46]) );
  DFFNEGX1 buff_data_reg_29__13_ ( .D(n3089), .CLK(clk), .Q(buff_data[45]) );
  DFFNEGX1 buff_data_reg_29__12_ ( .D(n3090), .CLK(clk), .Q(buff_data[44]) );
  DFFNEGX1 buff_data_reg_29__11_ ( .D(n3091), .CLK(clk), .Q(buff_data[43]) );
  DFFNEGX1 buff_data_reg_29__10_ ( .D(n3092), .CLK(clk), .Q(buff_data[42]) );
  DFFNEGX1 buff_data_reg_29__9_ ( .D(n3093), .CLK(clk), .Q(buff_data[41]) );
  DFFNEGX1 buff_data_reg_29__8_ ( .D(n3094), .CLK(clk), .Q(buff_data[40]) );
  DFFNEGX1 buff_data_reg_29__7_ ( .D(n3095), .CLK(clk), .Q(buff_data[39]) );
  DFFNEGX1 buff_data_reg_29__6_ ( .D(n3096), .CLK(clk), .Q(buff_data[38]) );
  DFFNEGX1 buff_data_reg_29__5_ ( .D(n3097), .CLK(clk), .Q(buff_data[37]) );
  DFFNEGX1 buff_data_reg_29__4_ ( .D(n3098), .CLK(clk), .Q(buff_data[36]) );
  DFFNEGX1 buff_data_reg_29__3_ ( .D(n3099), .CLK(clk), .Q(buff_data[35]) );
  DFFNEGX1 buff_data_reg_29__2_ ( .D(n3100), .CLK(clk), .Q(buff_data[34]) );
  DFFNEGX1 buff_data_reg_29__1_ ( .D(n3101), .CLK(clk), .Q(buff_data[33]) );
  DFFNEGX1 buff_data_reg_29__0_ ( .D(n3102), .CLK(clk), .Q(buff_data[32]) );
  DFFNEGX1 buff_data_reg_30__15_ ( .D(n2142), .CLK(clk), .Q(buff_data[31]) );
  DFFNEGX1 buff_data_reg_30__14_ ( .D(n3104), .CLK(clk), .Q(buff_data[30]) );
  DFFNEGX1 buff_data_reg_30__13_ ( .D(n1936), .CLK(clk), .Q(buff_data[29]) );
  DFFNEGX1 buff_data_reg_30__12_ ( .D(n3106), .CLK(clk), .Q(buff_data[28]) );
  DFFNEGX1 buff_data_reg_30__11_ ( .D(n3107), .CLK(clk), .Q(buff_data[27]) );
  DFFNEGX1 buff_data_reg_30__10_ ( .D(n3108), .CLK(clk), .Q(buff_data[26]) );
  DFFNEGX1 buff_data_reg_30__9_ ( .D(n1940), .CLK(clk), .Q(buff_data[25]) );
  DFFNEGX1 buff_data_reg_30__8_ ( .D(n3110), .CLK(clk), .Q(buff_data[24]) );
  DFFNEGX1 buff_data_reg_30__7_ ( .D(n3111), .CLK(clk), .Q(buff_data[23]) );
  DFFNEGX1 buff_data_reg_30__6_ ( .D(n3112), .CLK(clk), .Q(buff_data[22]) );
  DFFNEGX1 buff_data_reg_30__5_ ( .D(n3113), .CLK(clk), .Q(buff_data[21]) );
  DFFNEGX1 buff_data_reg_30__4_ ( .D(n2079), .CLK(clk), .Q(buff_data[20]) );
  DFFNEGX1 buff_data_reg_30__3_ ( .D(n3115), .CLK(clk), .Q(buff_data[19]) );
  DFFNEGX1 buff_data_reg_30__2_ ( .D(n1929), .CLK(clk), .Q(buff_data[18]) );
  DFFNEGX1 buff_data_reg_30__1_ ( .D(n3117), .CLK(clk), .Q(buff_data[17]) );
  DFFNEGX1 buff_data_reg_30__0_ ( .D(n3118), .CLK(clk), .Q(buff_data[16]) );
  DFFNEGX1 buff_data_reg_31__15_ ( .D(n2173), .CLK(clk), .Q(buff_data[15]) );
  DFFNEGX1 buff_data_reg_31__14_ ( .D(n1938), .CLK(clk), .Q(buff_data[14]) );
  DFFNEGX1 buff_data_reg_31__13_ ( .D(n3121), .CLK(clk), .Q(buff_data[13]) );
  DFFNEGX1 buff_data_reg_31__12_ ( .D(n3122), .CLK(clk), .Q(buff_data[12]) );
  DFFNEGX1 buff_data_reg_31__11_ ( .D(n3123), .CLK(clk), .Q(buff_data[11]) );
  DFFNEGX1 buff_data_reg_31__10_ ( .D(n3124), .CLK(clk), .Q(buff_data[10]) );
  DFFNEGX1 buff_data_reg_31__9_ ( .D(n1960), .CLK(clk), .Q(buff_data[9]) );
  DFFNEGX1 buff_data_reg_31__8_ ( .D(n3128), .CLK(clk), .Q(buff_data[8]) );
  DFFNEGX1 buff_data_reg_31__7_ ( .D(n3129), .CLK(clk), .Q(buff_data[7]) );
  DFFNEGX1 buff_data_reg_31__6_ ( .D(n3130), .CLK(clk), .Q(buff_data[6]) );
  DFFNEGX1 buff_data_reg_31__5_ ( .D(n3131), .CLK(clk), .Q(buff_data[5]) );
  DFFNEGX1 buff_data_reg_31__4_ ( .D(n3132), .CLK(clk), .Q(buff_data[4]) );
  DFFNEGX1 buff_data_reg_31__3_ ( .D(n3134), .CLK(clk), .Q(buff_data[3]) );
  DFFNEGX1 buff_data_reg_31__2_ ( .D(n3135), .CLK(clk), .Q(buff_data[2]) );
  DFFNEGX1 buff_data_reg_31__1_ ( .D(n3136), .CLK(clk), .Q(buff_data[1]) );
  DFFNEGX1 buff_data_reg_31__0_ ( .D(n3137), .CLK(clk), .Q(buff_data[0]) );
  DFFPOSX1 DQS_out_reg_1_ ( .D(n2547), .CLK(clk), .Q(DQS_out[1]) );
  DFFPOSX1 DQS_out_reg_0_ ( .D(n2548), .CLK(clk), .Q(DQS_out[0]) );
  DFFPOSX1 ts_con_reg ( .D(n909), .CLK(clk), .Q(ts_con) );
  INVX1 U2060 ( .A(clk), .Y(n252) );
  Processing_logic_DW01_inc_0 add_199 ( .A(clkcount), .SUM({n284, n283, n282, 
        n281, n280, n279, n278, n277, n276, n275, n274, n273, n272, n271, n270, 
        n269, n268, n267, n266, n265, n264, n263, n262, n261, n260, n259, n258, 
        n257, n256, n255, n254, n253}) );
  Processing_logic_DW01_inc_1 r586 ( .A({j, n232, n231, n230, net79430, 
        net79400}), .SUM({n2112, n2111, n2110, n2109, n2108, n2107, n2106, 
        n2105, n2104, n2103, n2102, n2101, n2100, n2099, n2098, n2097, n2096, 
        n2095, n2094, n2093, n2092, n2091, n2090, n2089, n2088, n2087, n2086, 
        n2085, n2084, n2083, n2082, n2081}) );
  Processing_logic_DW01_sub_0 r582 ( .A({blk_cnt[31:3], 1'b0, 1'b0, 1'b0}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .DIFF({n1780, n1779, n1778, n1777, n1776, n1775, n1774, n1773, n1772, 
        n1771, n1770, n1769, n1768, n1767, n1766, n1765, n1764, n1763, n1762, 
        n1761, n1760, n1759, n1758, n1757, n1756, n1755, n1754, n1753, n1752, 
        SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3}), .CO() );
  Processing_logic_DW01_cmp6_1 r589 ( .A({j, n232, n231, n230, net79428, 
        net79398}), .B({blk_cnt[31:3], 1'b0, 1'b0, 1'b0}), .TC(1'b1), .LT(
        n2442), .GT(), .EQ(), .LE(n2509), .GE(), .NE() );
  Processing_logic_DW01_dec_0 sub_657 ( .A({blk_cnt[31:3], 1'b0, 1'b0, 1'b0}), 
        .SUM({n2406, n2405, n2404, n2403, n2402, n2401, n2400, n2399, n2398, 
        n2397, n2396, n2395, n2394, n2393, n2392, n2391, n2390, n2389, n2388, 
        n2387, n2386, n2385, n2384, n2383, n2382, n2381, n2380, n2379, n2378, 
        SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6}) );
  Processing_logic_DW01_inc_2 r575 ( .A(i), .SUM({n634, n635, n636, n637, n638, 
        n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n669, n703, 
        n737, n805, n839, n873, n907, n942, n976, n977, n978, n979, n980, n981, 
        n982, n983, n984}) );
  \**SEQGEN**  blk_cnt_reg_31_ ( .clear(reset), .preset(1'b0), .next_state(
        n3427), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        blk_cnt[31]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  state_reg_0_ ( .clear(reset), .preset(1'b0), .next_state(n3361), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(state[0]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  i_reg_31_ ( .clear(reset), .preset(1'b0), .next_state(n3365), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(i[31]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  flag_bl_write_reg ( .clear(reset), .preset(1'b0), .next_state(
        n3221), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        flag_bl_write), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  state_reg_4_ ( .clear(reset), .preset(1'b0), .next_state(n3353), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(state[4]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  i_reg_30_ ( .clear(reset), .preset(1'b0), .next_state(n3291), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(i[30]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  i_reg_29_ ( .clear(reset), .preset(1'b0), .next_state(n3293), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(i[29]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  i_reg_28_ ( .clear(reset), .preset(1'b0), .next_state(n3295), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(i[28]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  i_reg_27_ ( .clear(reset), .preset(1'b0), .next_state(n3297), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(i[27]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  i_reg_26_ ( .clear(reset), .preset(1'b0), .next_state(n3299), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(i[26]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  i_reg_25_ ( .clear(reset), .preset(1'b0), .next_state(n3301), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(i[25]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  i_reg_24_ ( .clear(reset), .preset(1'b0), .next_state(n3303), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(i[24]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  i_reg_23_ ( .clear(reset), .preset(1'b0), .next_state(n3305), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(i[23]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  i_reg_22_ ( .clear(reset), .preset(1'b0), .next_state(n3307), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(i[22]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  i_reg_21_ ( .clear(reset), .preset(1'b0), .next_state(n3309), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(i[21]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  i_reg_20_ ( .clear(reset), .preset(1'b0), .next_state(n3311), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(i[20]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  i_reg_19_ ( .clear(reset), .preset(1'b0), .next_state(n3313), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(i[19]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  i_reg_18_ ( .clear(reset), .preset(1'b0), .next_state(n3315), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(i[18]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  i_reg_17_ ( .clear(reset), .preset(1'b0), .next_state(n3317), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(i[17]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  i_reg_16_ ( .clear(reset), .preset(1'b0), .next_state(n3319), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(i[16]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  i_reg_15_ ( .clear(reset), .preset(1'b0), .next_state(n3321), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(i[15]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  i_reg_14_ ( .clear(reset), .preset(1'b0), .next_state(n3323), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(i[14]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  i_reg_13_ ( .clear(reset), .preset(1'b0), .next_state(n3325), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(i[13]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  i_reg_12_ ( .clear(reset), .preset(1'b0), .next_state(n3327), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(i[12]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  i_reg_11_ ( .clear(reset), .preset(1'b0), .next_state(n3329), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(i[11]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  i_reg_10_ ( .clear(reset), .preset(1'b0), .next_state(n3331), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(i[10]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  i_reg_9_ ( .clear(reset), .preset(1'b0), .next_state(n3333), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(i[9]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  i_reg_8_ ( .clear(reset), .preset(1'b0), .next_state(n3335), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(i[8]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  i_reg_7_ ( .clear(reset), .preset(1'b0), .next_state(n3337), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(i[7]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  i_reg_6_ ( .clear(reset), .preset(1'b0), .next_state(n3339), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(i[6]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  i_reg_5_ ( .clear(reset), .preset(1'b0), .next_state(n3341), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(i[5]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  i_reg_4_ ( .clear(reset), .preset(1'b0), .next_state(n3343), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(i[4]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  i_reg_3_ ( .clear(reset), .preset(1'b0), .next_state(n3345), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(i[3]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  i_reg_2_ ( .clear(reset), .preset(1'b0), .next_state(n3347), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(i[2]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  i_reg_1_ ( .clear(reset), .preset(1'b0), .next_state(n3349), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(i[1]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  i_reg_0_ ( .clear(reset), .preset(1'b0), .next_state(n3351), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(i[0]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  state_reg_1_ ( .clear(reset), .preset(1'b0), .next_state(n3359), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(state[1]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  state_reg_3_ ( .clear(reset), .preset(1'b0), .next_state(n3355), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(state[3]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  state_reg_2_ ( .clear(reset), .preset(1'b0), .next_state(n3357), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(state[2]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  listen_reg ( .clear(reset), .preset(1'b0), .next_state(n2439), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(listen), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  ring_ptr_reg_2_ ( .clear(reset), .preset(1'b0), .next_state(
        n3227), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        ring_ptr[2]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  ring_ptr_reg_0_ ( .clear(reset), .preset(1'b0), .next_state(
        n3225), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        ring_ptr[0]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  ring_ptr_reg_1_ ( .clear(reset), .preset(1'b0), .next_state(
        n3223), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        ring_ptr[1]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  flag_at_read_reg ( .clear(reset), .preset(1'b0), .next_state(
        n3206), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        flag_at_read), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  RETURN_put_reg ( .clear(reset), .preset(1'b0), .next_state(
        n3079), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        RETURN_put), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  clkcount_reg_30_ ( .clear(reset), .preset(1'b0), .next_state(
        n3229), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        clkcount[30]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  clkcount_reg_29_ ( .clear(reset), .preset(1'b0), .next_state(
        n3231), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        clkcount[29]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  clkcount_reg_28_ ( .clear(reset), .preset(1'b0), .next_state(
        n3233), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        clkcount[28]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  clkcount_reg_27_ ( .clear(reset), .preset(1'b0), .next_state(
        n3235), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        clkcount[27]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  clkcount_reg_26_ ( .clear(reset), .preset(1'b0), .next_state(
        n3237), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        clkcount[26]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  clkcount_reg_25_ ( .clear(reset), .preset(1'b0), .next_state(
        n3239), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        clkcount[25]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  clkcount_reg_24_ ( .clear(reset), .preset(1'b0), .next_state(
        n3241), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        clkcount[24]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  clkcount_reg_23_ ( .clear(reset), .preset(1'b0), .next_state(
        n3243), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        clkcount[23]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  clkcount_reg_22_ ( .clear(reset), .preset(1'b0), .next_state(
        n3245), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        clkcount[22]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  clkcount_reg_21_ ( .clear(reset), .preset(1'b0), .next_state(
        n3247), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        clkcount[21]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  clkcount_reg_20_ ( .clear(reset), .preset(1'b0), .next_state(
        n3249), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        clkcount[20]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  clkcount_reg_19_ ( .clear(reset), .preset(1'b0), .next_state(
        n3251), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        clkcount[19]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  clkcount_reg_18_ ( .clear(reset), .preset(1'b0), .next_state(
        n3253), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        clkcount[18]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  clkcount_reg_17_ ( .clear(reset), .preset(1'b0), .next_state(
        n3255), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        clkcount[17]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  clkcount_reg_16_ ( .clear(reset), .preset(1'b0), .next_state(
        n3257), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        clkcount[16]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  clkcount_reg_15_ ( .clear(reset), .preset(1'b0), .next_state(
        n3259), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        clkcount[15]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  clkcount_reg_14_ ( .clear(reset), .preset(1'b0), .next_state(
        n3261), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        clkcount[14]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  clkcount_reg_13_ ( .clear(reset), .preset(1'b0), .next_state(
        n3263), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        clkcount[13]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  clkcount_reg_12_ ( .clear(reset), .preset(1'b0), .next_state(
        n3265), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        clkcount[12]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  clkcount_reg_11_ ( .clear(reset), .preset(1'b0), .next_state(
        n3267), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        clkcount[11]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  clkcount_reg_10_ ( .clear(reset), .preset(1'b0), .next_state(
        n3269), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        clkcount[10]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  clkcount_reg_9_ ( .clear(reset), .preset(1'b0), .next_state(
        n3271), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        clkcount[9]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  clkcount_reg_8_ ( .clear(reset), .preset(1'b0), .next_state(
        n3273), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        clkcount[8]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  clkcount_reg_7_ ( .clear(reset), .preset(1'b0), .next_state(
        n3275), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        clkcount[7]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  clkcount_reg_6_ ( .clear(reset), .preset(1'b0), .next_state(
        n3277), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        clkcount[6]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  clkcount_reg_5_ ( .clear(reset), .preset(1'b0), .next_state(
        n3279), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        clkcount[5]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  clkcount_reg_4_ ( .clear(reset), .preset(1'b0), .next_state(
        n3281), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        clkcount[4]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  clkcount_reg_3_ ( .clear(reset), .preset(1'b0), .next_state(
        n3283), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        clkcount[3]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  clkcount_reg_2_ ( .clear(reset), .preset(1'b0), .next_state(
        n3285), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        clkcount[2]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  clkcount_reg_1_ ( .clear(reset), .preset(1'b0), .next_state(
        n3287), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        clkcount[1]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  clkcount_reg_0_ ( .clear(reset), .preset(1'b0), .next_state(
        n3289), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        clkcount[0]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  clkcount_reg_31_ ( .clear(reset), .preset(1'b0), .next_state(
        n3363), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        clkcount[31]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  blk_cnt_reg_30_ ( .clear(reset), .preset(1'b0), .next_state(
        n3367), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        blk_cnt[30]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  blk_cnt_reg_29_ ( .clear(reset), .preset(1'b0), .next_state(
        n3369), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        blk_cnt[29]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  blk_cnt_reg_28_ ( .clear(reset), .preset(1'b0), .next_state(
        n3371), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        blk_cnt[28]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  blk_cnt_reg_27_ ( .clear(reset), .preset(1'b0), .next_state(
        n3373), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        blk_cnt[27]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  blk_cnt_reg_26_ ( .clear(reset), .preset(1'b0), .next_state(
        n3375), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        blk_cnt[26]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  blk_cnt_reg_25_ ( .clear(reset), .preset(1'b0), .next_state(
        n3377), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        blk_cnt[25]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  blk_cnt_reg_24_ ( .clear(reset), .preset(1'b0), .next_state(
        n3379), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        blk_cnt[24]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  blk_cnt_reg_23_ ( .clear(reset), .preset(1'b0), .next_state(
        n3381), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        blk_cnt[23]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  blk_cnt_reg_22_ ( .clear(reset), .preset(1'b0), .next_state(
        n3383), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        blk_cnt[22]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  blk_cnt_reg_21_ ( .clear(reset), .preset(1'b0), .next_state(
        n3385), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        blk_cnt[21]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  blk_cnt_reg_20_ ( .clear(reset), .preset(1'b0), .next_state(
        n3387), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        blk_cnt[20]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  blk_cnt_reg_19_ ( .clear(reset), .preset(1'b0), .next_state(
        n3389), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        blk_cnt[19]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  blk_cnt_reg_18_ ( .clear(reset), .preset(1'b0), .next_state(
        n3391), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        blk_cnt[18]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  blk_cnt_reg_17_ ( .clear(reset), .preset(1'b0), .next_state(
        n3393), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        blk_cnt[17]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  blk_cnt_reg_16_ ( .clear(reset), .preset(1'b0), .next_state(
        n3395), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        blk_cnt[16]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  blk_cnt_reg_15_ ( .clear(reset), .preset(1'b0), .next_state(
        n3397), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        blk_cnt[15]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  blk_cnt_reg_14_ ( .clear(reset), .preset(1'b0), .next_state(
        n3399), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        blk_cnt[14]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  blk_cnt_reg_13_ ( .clear(reset), .preset(1'b0), .next_state(
        n3401), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        blk_cnt[13]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  blk_cnt_reg_12_ ( .clear(reset), .preset(1'b0), .next_state(
        n3403), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        blk_cnt[12]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  blk_cnt_reg_11_ ( .clear(reset), .preset(1'b0), .next_state(
        n3405), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        blk_cnt[11]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  blk_cnt_reg_10_ ( .clear(reset), .preset(1'b0), .next_state(
        n3407), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        blk_cnt[10]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  blk_cnt_reg_9_ ( .clear(reset), .preset(1'b0), .next_state(
        n3409), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        blk_cnt[9]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  blk_cnt_reg_8_ ( .clear(reset), .preset(1'b0), .next_state(
        n3411), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        blk_cnt[8]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  blk_cnt_reg_7_ ( .clear(reset), .preset(1'b0), .next_state(
        n3413), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        blk_cnt[7]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  blk_cnt_reg_6_ ( .clear(reset), .preset(1'b0), .next_state(
        n3415), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        blk_cnt[6]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  blk_cnt_reg_5_ ( .clear(reset), .preset(1'b0), .next_state(
        n3417), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        blk_cnt[5]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  blk_cnt_reg_4_ ( .clear(reset), .preset(1'b0), .next_state(
        n3419), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        blk_cnt[4]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  blk_cnt_reg_3_ ( .clear(reset), .preset(1'b0), .next_state(
        n3421), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        blk_cnt[3]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  j_reg_0_ ( .clear(reset), .preset(1'b0), .next_state(n3200), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(net79414), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  j_reg_1_ ( .clear(reset), .preset(1'b0), .next_state(n3198), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(n229), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  j_reg_2_ ( .clear(reset), .preset(1'b0), .next_state(n3196), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(n230), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  j_reg_3_ ( .clear(reset), .preset(1'b0), .next_state(n3194), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(n231), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  j_reg_4_ ( .clear(reset), .preset(1'b0), .next_state(n3192), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(n232), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  j_reg_5_ ( .clear(reset), .preset(1'b0), .next_state(n3190), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(j[5]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  j_reg_6_ ( .clear(reset), .preset(1'b0), .next_state(n3188), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(j[6]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  j_reg_7_ ( .clear(reset), .preset(1'b0), .next_state(n3186), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(j[7]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  j_reg_8_ ( .clear(reset), .preset(1'b0), .next_state(n3184), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(j[8]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  j_reg_9_ ( .clear(reset), .preset(1'b0), .next_state(n3182), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(j[9]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  j_reg_10_ ( .clear(reset), .preset(1'b0), .next_state(n3180), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(j[10]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  j_reg_11_ ( .clear(reset), .preset(1'b0), .next_state(n3178), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(j[11]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  j_reg_12_ ( .clear(reset), .preset(1'b0), .next_state(n3176), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(j[12]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  j_reg_13_ ( .clear(reset), .preset(1'b0), .next_state(n3174), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(j[13]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  j_reg_14_ ( .clear(reset), .preset(1'b0), .next_state(n3172), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(j[14]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  j_reg_15_ ( .clear(reset), .preset(1'b0), .next_state(n3170), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(j[15]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  j_reg_16_ ( .clear(reset), .preset(1'b0), .next_state(n3168), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(j[16]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  j_reg_17_ ( .clear(reset), .preset(1'b0), .next_state(n3166), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(j[17]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  j_reg_18_ ( .clear(reset), .preset(1'b0), .next_state(n3164), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(j[18]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  j_reg_19_ ( .clear(reset), .preset(1'b0), .next_state(n3162), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(j[19]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  j_reg_20_ ( .clear(reset), .preset(1'b0), .next_state(n3160), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(j[20]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  j_reg_21_ ( .clear(reset), .preset(1'b0), .next_state(n3158), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(j[21]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  j_reg_22_ ( .clear(reset), .preset(1'b0), .next_state(n3156), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(j[22]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  j_reg_23_ ( .clear(reset), .preset(1'b0), .next_state(n3154), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(j[23]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  j_reg_24_ ( .clear(reset), .preset(1'b0), .next_state(n3152), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(j[24]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  j_reg_25_ ( .clear(reset), .preset(1'b0), .next_state(n3150), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(j[25]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  j_reg_26_ ( .clear(reset), .preset(1'b0), .next_state(n3148), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(j[26]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  j_reg_27_ ( .clear(reset), .preset(1'b0), .next_state(n3146), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(j[27]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  j_reg_28_ ( .clear(reset), .preset(1'b0), .next_state(n3144), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(j[28]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  j_reg_29_ ( .clear(reset), .preset(1'b0), .next_state(n3142), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(j[29]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  j_reg_30_ ( .clear(reset), .preset(1'b0), .next_state(n3140), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(j[30]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  j_reg_31_ ( .clear(reset), .preset(1'b0), .next_state(n3138), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(j[31]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  CMD_get_reg ( .clear(reset), .preset(1'b0), .next_state(n3036), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(CMD_get), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  DATA_get_reg ( .clear(reset), .preset(1'b0), .next_state(n3036), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(DATA_get), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  ras_bar_reg ( .clear(1'b0), .preset(reset), .next_state(n3204), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(ras_bar), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  we_bar_reg ( .clear(1'b0), .preset(reset), .next_state(n3202), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(we_bar), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  DQ_out_reg_15_ ( .clear(reset), .preset(1'b0), .next_state(
        n2615), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        DQ_out[15]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DQ_out_reg_14_ ( .clear(reset), .preset(1'b0), .next_state(
        n2613), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        DQ_out[14]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DQ_out_reg_13_ ( .clear(reset), .preset(1'b0), .next_state(
        n2611), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        DQ_out[13]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DQ_out_reg_12_ ( .clear(reset), .preset(1'b0), .next_state(
        n2609), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        DQ_out[12]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DQ_out_reg_11_ ( .clear(reset), .preset(1'b0), .next_state(
        n2607), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        DQ_out[11]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DQ_out_reg_10_ ( .clear(reset), .preset(1'b0), .next_state(
        n2605), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        DQ_out[10]), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  DQ_out_reg_9_ ( .clear(reset), .preset(1'b0), .next_state(n2603), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(DQ_out[9]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  DQ_out_reg_8_ ( .clear(reset), .preset(1'b0), .next_state(n2601), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(DQ_out[8]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  DQ_out_reg_7_ ( .clear(reset), .preset(1'b0), .next_state(n2599), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(DQ_out[7]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  DQ_out_reg_6_ ( .clear(reset), .preset(1'b0), .next_state(n2597), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(DQ_out[6]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  DQ_out_reg_5_ ( .clear(reset), .preset(1'b0), .next_state(n2595), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(DQ_out[5]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  DQ_out_reg_4_ ( .clear(reset), .preset(1'b0), .next_state(n2593), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(DQ_out[4]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  DQ_out_reg_3_ ( .clear(reset), .preset(1'b0), .next_state(n2591), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(DQ_out[3]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  DQ_out_reg_2_ ( .clear(reset), .preset(1'b0), .next_state(n2589), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(DQ_out[2]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  DQ_out_reg_1_ ( .clear(reset), .preset(1'b0), .next_state(n2587), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(DQ_out[1]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  DQ_out_reg_0_ ( .clear(reset), .preset(1'b0), .next_state(n2585), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(DQ_out[0]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  flag_bl_read_reg ( .clear(reset), .preset(1'b0), .next_state(
        n2583), .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(
        flag_bl_read), .QN(), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  A_reg_12_ ( .clear(reset), .preset(1'b0), .next_state(n2551), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(A[12]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  A_reg_11_ ( .clear(reset), .preset(1'b0), .next_state(n2553), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(A[11]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  A_reg_10_ ( .clear(reset), .preset(1'b0), .next_state(n2555), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(A[10]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  A_reg_9_ ( .clear(reset), .preset(1'b0), .next_state(n2557), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(A[9]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  A_reg_8_ ( .clear(reset), .preset(1'b0), .next_state(n2559), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(A[8]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  A_reg_7_ ( .clear(reset), .preset(1'b0), .next_state(n2561), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(A[7]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  A_reg_6_ ( .clear(reset), .preset(1'b0), .next_state(n2563), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(A[6]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  A_reg_5_ ( .clear(reset), .preset(1'b0), .next_state(n2565), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(A[5]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  A_reg_4_ ( .clear(reset), .preset(1'b0), .next_state(n2567), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(A[4]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  A_reg_3_ ( .clear(reset), .preset(1'b0), .next_state(n2569), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(A[3]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  A_reg_2_ ( .clear(reset), .preset(1'b0), .next_state(n2571), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(A[2]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  A_reg_1_ ( .clear(reset), .preset(1'b0), .next_state(n2573), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(A[1]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  A_reg_0_ ( .clear(reset), .preset(1'b0), .next_state(n2575), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(A[0]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  BA_reg_2_ ( .clear(reset), .preset(1'b0), .next_state(n2577), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(BA[2]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  BA_reg_1_ ( .clear(reset), .preset(1'b0), .next_state(n2579), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(BA[1]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  BA_reg_0_ ( .clear(reset), .preset(1'b0), .next_state(n2581), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(BA[0]), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  ri_o_reg ( .clear(reset), .preset(1'b0), .next_state(n3073), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(ri_o), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  cas_bar_reg ( .clear(1'b0), .preset(reset), .next_state(n114), 
        .clocked_on(n252), .data_in(1'b0), .enable(1'b0), .Q(cas_bar), .QN(), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  Processing_logic_DW_cmp_8 lt_657 ( .A({j, n232, n231, n230, net79430, 
        net79402}), .B({n2406, n2405, n2404, n2403, n2402, n2401, n2400, n2399, 
        n2398, n2397, n2396, n2395, n2394, n2393, n2392, n2391, n2390, n2389, 
        n2388, n2387, n2386, n2385, n2384, n2383, n2382, n2381, n2380, n2379, 
        n2378, 1'b1, 1'b1, 1'b1}), .TC(1'b1), .GE_LT(1'b1), .GE_GT_EQ(1'b0), 
        .GE_LT_GT_LE(n2407), .EQ_NE() );
  INVX1 U6 ( .A(n438), .Y(n1) );
  INVX1 U7 ( .A(n438), .Y(n1607) );
  MUX2X1 U8 ( .B(n573), .A(buff_data[272]), .S(n99), .Y(n4183) );
  INVX1 U9 ( .A(net82538), .Y(n327) );
  INVX4 U10 ( .A(n2000), .Y(net80839) );
  INVX4 U11 ( .A(n11), .Y(net80464) );
  INVX1 U12 ( .A(n2074), .Y(n2) );
  INVX1 U13 ( .A(net82538), .Y(n3) );
  INVX1 U14 ( .A(n1801), .Y(n4) );
  INVX1 U15 ( .A(n1801), .Y(n5) );
  INVX1 U16 ( .A(n1801), .Y(n2053) );
  MUX2X1 U17 ( .B(n565), .A(buff_data[185]), .S(n537), .Y(n4112) );
  INVX2 U18 ( .A(n6), .Y(n537) );
  AND2X2 U19 ( .A(net89705), .B(n4011), .Y(n6) );
  INVX1 U20 ( .A(n6), .Y(n7) );
  INVX1 U21 ( .A(n6), .Y(n8) );
  INVX1 U22 ( .A(n428), .Y(n9) );
  INVX1 U23 ( .A(net92867), .Y(n10) );
  AND2X2 U24 ( .A(net80596), .B(net66441), .Y(n11) );
  INVX1 U25 ( .A(n3), .Y(n12) );
  MUX2X1 U26 ( .B(n575), .A(buff_data[207]), .S(n406), .Y(n4131) );
  INVX1 U27 ( .A(n30), .Y(n13) );
  INVX1 U28 ( .A(n29), .Y(n14) );
  MUX2X1 U29 ( .B(buff_data[468]), .A(n576), .S(n1850), .Y(n195) );
  INVX2 U30 ( .A(n149), .Y(n181) );
  INVX1 U31 ( .A(n561), .Y(n15) );
  INVX1 U32 ( .A(n15), .Y(n16) );
  INVX1 U33 ( .A(n2194), .Y(n17) );
  INVX1 U34 ( .A(n2194), .Y(n18) );
  INVX2 U35 ( .A(n1842), .Y(n19) );
  INVX1 U36 ( .A(n1842), .Y(n466) );
  INVX1 U37 ( .A(n325), .Y(n20) );
  INVX1 U38 ( .A(n326), .Y(n21) );
  INVX1 U39 ( .A(n210), .Y(n22) );
  MUX2X1 U40 ( .B(n573), .A(buff_data[400]), .S(n546), .Y(n4287) );
  INVX1 U41 ( .A(n1835), .Y(n23) );
  INVX1 U42 ( .A(n25), .Y(n24) );
  INVX1 U43 ( .A(n1966), .Y(n25) );
  INVX1 U44 ( .A(n19), .Y(n26) );
  INVX1 U45 ( .A(n179), .Y(n27) );
  MUX2X1 U46 ( .B(n567), .A(buff_data[414]), .S(n181), .Y(n28) );
  INVX8 U47 ( .A(n28), .Y(n1954) );
  INVX2 U48 ( .A(n1848), .Y(n29) );
  INVX2 U49 ( .A(n1848), .Y(n30) );
  INVX1 U50 ( .A(n1848), .Y(n563) );
  INVX1 U51 ( .A(n179), .Y(n31) );
  INVX4 U52 ( .A(n160), .Y(net93057) );
  INVX2 U53 ( .A(n1804), .Y(n160) );
  INVX2 U54 ( .A(n1843), .Y(n32) );
  INVX2 U55 ( .A(n1843), .Y(n2194) );
  INVX1 U56 ( .A(n187), .Y(n33) );
  INVX8 U57 ( .A(n562), .Y(n34) );
  INVX4 U58 ( .A(n1825), .Y(n562) );
  INVX1 U59 ( .A(n70), .Y(n35) );
  INVX1 U60 ( .A(n1912), .Y(n36) );
  INVX1 U61 ( .A(net80322), .Y(n37) );
  INVX1 U62 ( .A(n203), .Y(n38) );
  AND2X2 U63 ( .A(net82472), .B(n3963), .Y(n39) );
  MUX2X1 U64 ( .B(n41), .A(n572), .S(n14), .Y(n40) );
  INVX8 U65 ( .A(n40), .Y(n1900) );
  INVX8 U66 ( .A(n1901), .Y(n41) );
  INVX1 U67 ( .A(n559), .Y(n42) );
  INVX1 U68 ( .A(n559), .Y(n43) );
  INVX1 U69 ( .A(n175), .Y(n2198) );
  INVX1 U70 ( .A(n33), .Y(n44) );
  INVX1 U71 ( .A(n175), .Y(n45) );
  INVX8 U72 ( .A(n2194), .Y(n2195) );
  INVX1 U73 ( .A(n2116), .Y(n370) );
  INVX1 U74 ( .A(n558), .Y(n46) );
  INVX1 U75 ( .A(n416), .Y(n185) );
  MUX2X1 U76 ( .B(n48), .A(n565), .S(n1817), .Y(n47) );
  INVX8 U77 ( .A(n47), .Y(n1989) );
  INVX8 U78 ( .A(n1990), .Y(n48) );
  INVX4 U79 ( .A(n160), .Y(net79538) );
  INVX1 U80 ( .A(n210), .Y(n60) );
  INVX1 U81 ( .A(n218), .Y(n49) );
  INVX4 U82 ( .A(n218), .Y(n444) );
  INVX1 U83 ( .A(n72), .Y(n50) );
  INVX4 U84 ( .A(n72), .Y(n443) );
  INVX1 U85 ( .A(n407), .Y(n51) );
  INVX1 U86 ( .A(n381), .Y(n366) );
  INVX8 U87 ( .A(n462), .Y(net80783) );
  INVX1 U88 ( .A(n80), .Y(n52) );
  INVX1 U89 ( .A(n66), .Y(n53) );
  INVX2 U90 ( .A(n1911), .Y(n54) );
  INVX1 U91 ( .A(n1911), .Y(n55) );
  INVX1 U92 ( .A(n1911), .Y(n1815) );
  INVX1 U93 ( .A(net80791), .Y(n56) );
  AND2X2 U94 ( .A(net80872), .B(net66503), .Y(n57) );
  MUX2X1 U95 ( .B(n59), .A(n571), .S(n174), .Y(n58) );
  INVX8 U96 ( .A(n58), .Y(n2017) );
  INVX8 U97 ( .A(n2018), .Y(n59) );
  MUX2X1 U98 ( .B(n574), .A(buff_data[274]), .S(n415), .Y(n4185) );
  MUX2X1 U99 ( .B(n62), .A(n573), .S(net80783), .Y(n61) );
  INVX8 U100 ( .A(n61), .Y(n1979) );
  INVX8 U101 ( .A(n1980), .Y(n62) );
  MUX2X1 U102 ( .B(n565), .A(n64), .S(n328), .Y(n63) );
  INVX8 U103 ( .A(n63), .Y(n1934) );
  INVX8 U104 ( .A(n1935), .Y(n64) );
  MUX2X1 U105 ( .B(n575), .A(buff_data[79]), .S(n531), .Y(n65) );
  INVX8 U106 ( .A(n65), .Y(n2165) );
  INVX1 U107 ( .A(net80322), .Y(n66) );
  INVX1 U108 ( .A(n203), .Y(n67) );
  INVX1 U109 ( .A(n66), .Y(n68) );
  INVX1 U110 ( .A(n37), .Y(n336) );
  INVX1 U111 ( .A(net80322), .Y(n203) );
  MUX2X1 U112 ( .B(n575), .A(buff_data[287]), .S(n99), .Y(n69) );
  INVX8 U113 ( .A(n69), .Y(n1963) );
  INVX1 U114 ( .A(n580), .Y(n70) );
  INVX1 U115 ( .A(n468), .Y(n71) );
  OR2X2 U116 ( .A(n56), .B(n219), .Y(n72) );
  MUX2X1 U117 ( .B(n74), .A(n568), .S(net80781), .Y(n73) );
  INVX8 U118 ( .A(n73), .Y(n2118) );
  INVX8 U119 ( .A(n2119), .Y(n74) );
  INVX1 U120 ( .A(n103), .Y(n75) );
  INVX1 U121 ( .A(n103), .Y(n76) );
  MUX2X1 U122 ( .B(n571), .A(buff_data[331]), .S(n358), .Y(n77) );
  INVX8 U123 ( .A(n77), .Y(n1907) );
  MUX2X1 U124 ( .B(n79), .A(n573), .S(n107), .Y(n78) );
  INVX8 U125 ( .A(n78), .Y(n1951) );
  INVX8 U126 ( .A(n1952), .Y(n79) );
  INVX1 U127 ( .A(n1802), .Y(n80) );
  INVX1 U128 ( .A(n438), .Y(n81) );
  INVX1 U129 ( .A(net92856), .Y(n82) );
  INVX1 U130 ( .A(n536), .Y(n83) );
  INVX1 U131 ( .A(n8), .Y(n84) );
  MUX2X1 U132 ( .B(n312), .A(n574), .S(n107), .Y(n311) );
  INVX1 U133 ( .A(n9), .Y(n85) );
  INVX1 U134 ( .A(n1931), .Y(n86) );
  INVX1 U135 ( .A(n550), .Y(n87) );
  INVX1 U136 ( .A(n550), .Y(n88) );
  INVX1 U137 ( .A(n70), .Y(net79510) );
  INVX1 U138 ( .A(n580), .Y(n228) );
  INVX1 U139 ( .A(net82538), .Y(net79533) );
  MUX2X1 U140 ( .B(n567), .A(n90), .S(n1824), .Y(n89) );
  INVX8 U141 ( .A(n89), .Y(n1949) );
  INVX8 U142 ( .A(n1950), .Y(n90) );
  INVX1 U143 ( .A(n228), .Y(n91) );
  MUX2X1 U144 ( .B(n93), .A(n564), .S(n20), .Y(n92) );
  INVX8 U145 ( .A(n92), .Y(n2071) );
  INVX8 U146 ( .A(n2072), .Y(n93) );
  INVX1 U147 ( .A(n154), .Y(n94) );
  MUX2X1 U148 ( .B(n572), .A(n96), .S(n415), .Y(n95) );
  INVX8 U149 ( .A(n95), .Y(n2140) );
  INVX8 U150 ( .A(n2141), .Y(n96) );
  AND2X2 U151 ( .A(net66503), .B(net80598), .Y(n97) );
  INVX1 U152 ( .A(n1569), .Y(net66503) );
  AND2X2 U153 ( .A(n320), .B(net66423), .Y(n98) );
  INVX1 U154 ( .A(n1931), .Y(n99) );
  INVX1 U155 ( .A(n1931), .Y(n100) );
  MUX2X1 U156 ( .B(n568), .A(buff_data[195]), .S(n406), .Y(n101) );
  INVX8 U157 ( .A(n101), .Y(n1926) );
  MUX2X1 U162 ( .B(n567), .A(buff_data[206]), .S(n401), .Y(n102) );
  INVX8 U163 ( .A(n102), .Y(n1948) );
  INVX1 U164 ( .A(n11), .Y(n103) );
  MUX2X1 U165 ( .B(n571), .A(n105), .S(n51), .Y(n104) );
  INVX8 U166 ( .A(n104), .Y(n2065) );
  INVX8 U167 ( .A(n2066), .Y(n105) );
  INVX1 U168 ( .A(n2053), .Y(n106) );
  INVX1 U169 ( .A(n5), .Y(n107) );
  INVX1 U170 ( .A(n29), .Y(n108) );
  INVX1 U171 ( .A(n30), .Y(n109) );
  INVX1 U172 ( .A(n30), .Y(net80760) );
  INVX1 U173 ( .A(n30), .Y(n110) );
  INVX1 U174 ( .A(n30), .Y(n111) );
  INVX1 U175 ( .A(n29), .Y(n112) );
  INVX1 U176 ( .A(n181), .Y(n113) );
  MUX2X1 U177 ( .B(n860), .A(n115), .S(n1670), .Y(n114) );
  INVX8 U178 ( .A(cas_bar), .Y(n115) );
  MUX2X1 U179 ( .B(buff_data[452]), .A(n576), .S(n2030), .Y(n4332) );
  INVX8 U180 ( .A(n32), .Y(n2030) );
  AND2X2 U181 ( .A(net89543), .B(n117), .Y(n116) );
  INVX1 U182 ( .A(n116), .Y(net92773) );
  INVX8 U183 ( .A(n1230), .Y(n117) );
  INVX1 U184 ( .A(n179), .Y(n118) );
  INVX2 U185 ( .A(n1842), .Y(n179) );
  INVX1 U186 ( .A(n29), .Y(n119) );
  INVX1 U187 ( .A(n29), .Y(n120) );
  INVX1 U188 ( .A(n557), .Y(n121) );
  INVX1 U189 ( .A(n557), .Y(n122) );
  INVX1 U190 ( .A(n557), .Y(n2200) );
  MUX2X1 U191 ( .B(n564), .A(buff_data[506]), .S(n16), .Y(n4380) );
  INVX1 U192 ( .A(n207), .Y(n123) );
  INVX1 U193 ( .A(n123), .Y(n124) );
  INVX1 U194 ( .A(n1835), .Y(n125) );
  INVX1 U195 ( .A(n556), .Y(n126) );
  INVX1 U196 ( .A(n556), .Y(n127) );
  INVX1 U197 ( .A(n29), .Y(n128) );
  INVX1 U198 ( .A(n30), .Y(n129) );
  INVX1 U199 ( .A(n29), .Y(n130) );
  INVX1 U200 ( .A(n30), .Y(n131) );
  INVX1 U201 ( .A(n19), .Y(n132) );
  INVX1 U202 ( .A(n25), .Y(n133) );
  INVX1 U203 ( .A(n398), .Y(n134) );
  INVX1 U204 ( .A(n25), .Y(n135) );
  INVX1 U205 ( .A(n19), .Y(n136) );
  INVX1 U206 ( .A(n179), .Y(n137) );
  INVX1 U207 ( .A(n19), .Y(n138) );
  INVX1 U208 ( .A(n179), .Y(n2199) );
  INVX1 U209 ( .A(n557), .Y(n139) );
  INVX1 U210 ( .A(n557), .Y(n140) );
  INVX1 U211 ( .A(n163), .Y(n141) );
  INVX1 U212 ( .A(n19), .Y(n142) );
  INVX1 U213 ( .A(n1841), .Y(n143) );
  INVX1 U214 ( .A(n557), .Y(n144) );
  INVX1 U215 ( .A(n557), .Y(n145) );
  INVX1 U216 ( .A(n1841), .Y(n556) );
  INVX1 U217 ( .A(n326), .Y(n146) );
  INVX1 U218 ( .A(n556), .Y(n147) );
  INVX1 U219 ( .A(n1835), .Y(n148) );
  AND2X2 U220 ( .A(net92619), .B(net66423), .Y(n149) );
  MUX2X1 U221 ( .B(n151), .A(n568), .S(n120), .Y(n150) );
  INVX8 U222 ( .A(n150), .Y(n2122) );
  INVX8 U223 ( .A(n2123), .Y(n151) );
  INVX1 U224 ( .A(net79416), .Y(net79398) );
  INVX1 U225 ( .A(net79416), .Y(net79400) );
  INVX2 U226 ( .A(net79416), .Y(net79402) );
  MUX2X1 U227 ( .B(n153), .A(n576), .S(n118), .Y(n152) );
  INVX8 U228 ( .A(n152), .Y(n2120) );
  INVX8 U229 ( .A(n2121), .Y(n153) );
  INVX1 U230 ( .A(n398), .Y(n154) );
  INVX1 U231 ( .A(n203), .Y(n155) );
  INVX1 U232 ( .A(n37), .Y(n156) );
  INVX1 U233 ( .A(n37), .Y(n157) );
  INVX1 U234 ( .A(n66), .Y(n158) );
  INVX1 U235 ( .A(n179), .Y(n159) );
  INVX1 U236 ( .A(n325), .Y(n161) );
  INVX1 U237 ( .A(n325), .Y(n162) );
  INVX1 U238 ( .A(n326), .Y(n432) );
  INVX1 U239 ( .A(net66714), .Y(n163) );
  INVX1 U240 ( .A(n208), .Y(n164) );
  INVX1 U241 ( .A(n208), .Y(n165) );
  INVX1 U242 ( .A(n208), .Y(n344) );
  INVX2 U243 ( .A(n1841), .Y(n557) );
  BUFX2 U244 ( .A(n2407), .Y(n166) );
  INVX4 U245 ( .A(n143), .Y(n1928) );
  INVX2 U246 ( .A(n318), .Y(n866) );
  INVX1 U247 ( .A(n551), .Y(n167) );
  INVX1 U248 ( .A(n551), .Y(n168) );
  INVX1 U249 ( .A(n551), .Y(n2181) );
  INVX1 U250 ( .A(n551), .Y(n169) );
  INVX1 U251 ( .A(n551), .Y(n170) );
  INVX1 U252 ( .A(n417), .Y(n171) );
  INVX1 U253 ( .A(n163), .Y(n172) );
  AND2X2 U254 ( .A(net92619), .B(net66482), .Y(n1843) );
  INVX1 U255 ( .A(n52), .Y(n173) );
  INVX1 U256 ( .A(n337), .Y(n174) );
  INVX1 U257 ( .A(n187), .Y(n175) );
  INVX2 U258 ( .A(n2002), .Y(n349) );
  INVX1 U259 ( .A(n25), .Y(n176) );
  INVX1 U260 ( .A(n398), .Y(n177) );
  INVX1 U261 ( .A(n326), .Y(n2128) );
  INVX1 U262 ( .A(net80775), .Y(n178) );
  INVX1 U263 ( .A(n4056), .Y(n431) );
  INVX1 U264 ( .A(n431), .Y(n188) );
  INVX1 U265 ( .A(n1836), .Y(n440) );
  INVX1 U266 ( .A(n179), .Y(n180) );
  INVX1 U267 ( .A(n208), .Y(n182) );
  INVX1 U268 ( .A(n208), .Y(n183) );
  INVX1 U269 ( .A(n1992), .Y(n184) );
  INVX2 U270 ( .A(n1992), .Y(net79518) );
  AND2X2 U271 ( .A(net80519), .B(n4056), .Y(n186) );
  AND2X2 U272 ( .A(n548), .B(n188), .Y(n187) );
  INVX1 U273 ( .A(n187), .Y(n210) );
  INVX1 U274 ( .A(n551), .Y(n189) );
  INVX1 U275 ( .A(n551), .Y(n190) );
  INVX1 U276 ( .A(n551), .Y(n191) );
  INVX1 U277 ( .A(n551), .Y(n192) );
  INVX1 U278 ( .A(n558), .Y(n193) );
  INVX1 U279 ( .A(n203), .Y(n194) );
  INVX1 U280 ( .A(n429), .Y(n1927) );
  INVX8 U281 ( .A(n195), .Y(n2660) );
  INVX1 U282 ( .A(n208), .Y(n196) );
  INVX1 U283 ( .A(n208), .Y(n197) );
  INVX1 U284 ( .A(n208), .Y(n198) );
  INVX1 U285 ( .A(n559), .Y(n199) );
  INVX1 U286 ( .A(n1922), .Y(n406) );
  MUX2X1 U287 ( .B(n565), .A(buff_data[9]), .S(n2117), .Y(n200) );
  INVX8 U288 ( .A(n200), .Y(n1960) );
  MUX2X1 U289 ( .B(n566), .A(n202), .S(n51), .Y(n201) );
  INVX8 U290 ( .A(n201), .Y(n2033) );
  INVX8 U291 ( .A(n2034), .Y(n202) );
  INVX2 U292 ( .A(net80322), .Y(n558) );
  INVX1 U293 ( .A(n337), .Y(n204) );
  INVX1 U294 ( .A(n381), .Y(n2185) );
  INVX1 U295 ( .A(n228), .Y(n205) );
  INVX1 U296 ( .A(n228), .Y(n206) );
  INVX1 U297 ( .A(n70), .Y(n305) );
  INVX1 U298 ( .A(n429), .Y(n207) );
  INVX2 U299 ( .A(n1972), .Y(n208) );
  INVX2 U300 ( .A(n1972), .Y(n559) );
  INVX1 U301 ( .A(n1966), .Y(n398) );
  INVX4 U302 ( .A(n2052), .Y(n551) );
  INVX1 U303 ( .A(n468), .Y(n209) );
  INVX2 U304 ( .A(n2073), .Y(n553) );
  INVX1 U305 ( .A(n359), .Y(n211) );
  INVX1 U306 ( .A(n359), .Y(n212) );
  INVX1 U307 ( .A(n295), .Y(n2178) );
  INVX1 U308 ( .A(n361), .Y(n531) );
  MUX2X1 U309 ( .B(n574), .A(n214), .S(n181), .Y(n213) );
  INVX8 U310 ( .A(n213), .Y(n2124) );
  INVX8 U311 ( .A(n2125), .Y(n214) );
  INVX1 U312 ( .A(n429), .Y(n215) );
  INVX1 U313 ( .A(n4218), .Y(n216) );
  INVX2 U314 ( .A(n1804), .Y(n462) );
  INVX1 U315 ( .A(n544), .Y(n217) );
  OR2X2 U316 ( .A(n463), .B(n219), .Y(n218) );
  INVX8 U317 ( .A(n3963), .Y(n219) );
  MUX2X1 U318 ( .B(n572), .A(n221), .S(n3), .Y(n220) );
  INVX8 U319 ( .A(n220), .Y(n1946) );
  INVX8 U320 ( .A(n1947), .Y(n221) );
  INVX1 U321 ( .A(n553), .Y(n222) );
  INVX1 U322 ( .A(n553), .Y(n223) );
  INVX1 U323 ( .A(n359), .Y(n224) );
  INVX1 U324 ( .A(n359), .Y(n225) );
  INVX1 U325 ( .A(n359), .Y(n4043) );
  INVX1 U326 ( .A(n2029), .Y(n359) );
  MUX2X1 U327 ( .B(n227), .A(n564), .S(n173), .Y(n226) );
  INVX8 U328 ( .A(n226), .Y(n1932) );
  INVX8 U329 ( .A(n1933), .Y(n227) );
  INVX1 U330 ( .A(n580), .Y(n550) );
  MUX2X1 U331 ( .B(n570), .A(n250), .S(n2048), .Y(n249) );
  INVX8 U332 ( .A(n249), .Y(n1961) );
  INVX8 U333 ( .A(n1962), .Y(n250) );
  MUX2X1 U334 ( .B(n566), .A(n285), .S(n2048), .Y(n251) );
  INVX8 U335 ( .A(n251), .Y(n1974) );
  INVX8 U336 ( .A(n1975), .Y(n285) );
  INVX1 U337 ( .A(n433), .Y(n286) );
  INVX1 U338 ( .A(n433), .Y(n287) );
  INVX1 U339 ( .A(n307), .Y(n288) );
  INVX1 U340 ( .A(n307), .Y(n289) );
  INVX1 U341 ( .A(n433), .Y(n290) );
  INVX1 U342 ( .A(n295), .Y(n291) );
  INVX1 U343 ( .A(n429), .Y(n1953) );
  MUX2X1 U344 ( .B(n293), .A(n569), .S(n611), .Y(n292) );
  INVX8 U345 ( .A(n292), .Y(n1905) );
  INVX8 U346 ( .A(n1906), .Y(n293) );
  INVX1 U347 ( .A(n2184), .Y(n294) );
  INVX1 U348 ( .A(n361), .Y(n295) );
  MUX2X1 U349 ( .B(n297), .A(n573), .S(n367), .Y(n296) );
  INVX8 U350 ( .A(n296), .Y(n2135) );
  INVX8 U351 ( .A(n2136), .Y(n297) );
  INVX1 U352 ( .A(net80775), .Y(net80682) );
  INVX1 U353 ( .A(n467), .Y(n298) );
  INVX1 U354 ( .A(n560), .Y(n299) );
  INVX1 U355 ( .A(n468), .Y(n300) );
  MUX2X1 U356 ( .B(n568), .A(n302), .S(net80464), .Y(n301) );
  INVX8 U357 ( .A(n301), .Y(n2025) );
  INVX8 U358 ( .A(n2026), .Y(n302) );
  INVX1 U359 ( .A(n307), .Y(n303) );
  INVX1 U360 ( .A(n307), .Y(n304) );
  INVX1 U361 ( .A(n307), .Y(net79593) );
  INVX1 U362 ( .A(n1973), .Y(n307) );
  BUFX4 U363 ( .A(n2073), .Y(n306) );
  INVX1 U364 ( .A(n1973), .Y(n433) );
  INVX1 U365 ( .A(n337), .Y(n308) );
  MUX2X1 U366 ( .B(n575), .A(n310), .S(n54), .Y(n309) );
  INVX8 U367 ( .A(n309), .Y(n1919) );
  INVX8 U368 ( .A(n1920), .Y(n310) );
  INVX8 U369 ( .A(n311), .Y(n1967) );
  INVX8 U370 ( .A(n1968), .Y(n312) );
  MUX2X1 U371 ( .B(n569), .A(n314), .S(n553), .Y(n313) );
  INVX8 U372 ( .A(n313), .Y(n2171) );
  INVX8 U373 ( .A(n2172), .Y(n314) );
  INVX1 U374 ( .A(n2184), .Y(n2161) );
  MUX2X1 U375 ( .B(n566), .A(n316), .S(net80464), .Y(n315) );
  INVX8 U376 ( .A(n315), .Y(n1917) );
  INVX8 U377 ( .A(n1918), .Y(n316) );
  INVX1 U378 ( .A(net92751), .Y(n317) );
  NOR3X1 U379 ( .A(n319), .B(n1306), .C(n864), .Y(n318) );
  INVX8 U380 ( .A(n4524), .Y(n319) );
  INVX1 U381 ( .A(net92856), .Y(n320) );
  MUX2X1 U382 ( .B(n574), .A(n322), .S(n2075), .Y(n321) );
  INVX8 U383 ( .A(n321), .Y(n2152) );
  INVX8 U384 ( .A(n2153), .Y(n322) );
  MUX2X1 U385 ( .B(n569), .A(n324), .S(n2075), .Y(n323) );
  INVX8 U386 ( .A(n323), .Y(n2061) );
  INVX8 U387 ( .A(n2062), .Y(n324) );
  INVX1 U388 ( .A(n1966), .Y(n325) );
  INVX1 U389 ( .A(n1966), .Y(n326) );
  MUX2X1 U390 ( .B(buff_data[190]), .A(n567), .S(n1816), .Y(n4116) );
  OR2X2 U391 ( .A(net80595), .B(n1803), .Y(n328) );
  INVX1 U392 ( .A(n4056), .Y(n1803) );
  MUX2X1 U393 ( .B(n564), .A(n330), .S(net80464), .Y(n329) );
  INVX8 U394 ( .A(n329), .Y(n2069) );
  INVX8 U395 ( .A(n2070), .Y(n330) );
  INVX1 U396 ( .A(n1837), .Y(n331) );
  INVX1 U397 ( .A(n433), .Y(n332) );
  INVX1 U398 ( .A(n433), .Y(n333) );
  INVX1 U399 ( .A(n407), .Y(n334) );
  INVX1 U400 ( .A(n407), .Y(n335) );
  INVX1 U401 ( .A(n2074), .Y(n2075) );
  INVX1 U402 ( .A(n4205), .Y(n337) );
  INVX1 U403 ( .A(n403), .Y(n338) );
  MUX2X1 U404 ( .B(n564), .A(n340), .S(n537), .Y(n339) );
  INVX8 U405 ( .A(n339), .Y(n2145) );
  INVX8 U406 ( .A(n2146), .Y(n340) );
  INVX1 U407 ( .A(n317), .Y(n341) );
  INVX1 U408 ( .A(n536), .Y(n342) );
  INVX1 U409 ( .A(n8), .Y(n343) );
  MUX2X1 U410 ( .B(n578), .A(buff_data[71]), .S(n123), .Y(n4018) );
  MUX2X1 U411 ( .B(n573), .A(buff_data[64]), .S(n2076), .Y(n4012) );
  INVX1 U412 ( .A(n2053), .Y(n345) );
  INVX1 U413 ( .A(n4205), .Y(n2184) );
  MUX2X1 U414 ( .B(n347), .A(n570), .S(n2126), .Y(n346) );
  INVX8 U415 ( .A(n346), .Y(n2054) );
  INVX8 U416 ( .A(n2055), .Y(n347) );
  INVX1 U417 ( .A(n2074), .Y(n1824) );
  MUX2X1 U418 ( .B(n568), .A(buff_data[3]), .S(n370), .Y(n3953) );
  INVX1 U419 ( .A(n399), .Y(n348) );
  MUX2X1 U420 ( .B(n574), .A(buff_data[2]), .S(n370), .Y(n3952) );
  INVX4 U421 ( .A(n377), .Y(n2179) );
  INVX1 U422 ( .A(n2002), .Y(n350) );
  INVX1 U423 ( .A(n553), .Y(n351) );
  INVX1 U424 ( .A(n553), .Y(n379) );
  INVX1 U425 ( .A(n468), .Y(n352) );
  INVX1 U426 ( .A(n381), .Y(n353) );
  MUX2X1 U427 ( .B(n355), .A(n566), .S(n184), .Y(n354) );
  INVX8 U428 ( .A(n354), .Y(n2006) );
  INVX8 U429 ( .A(n2007), .Y(n355) );
  MUX2X1 U430 ( .B(n357), .A(n575), .S(n2162), .Y(n356) );
  INVX8 U431 ( .A(n356), .Y(n2173) );
  INVX8 U432 ( .A(n2174), .Y(n357) );
  INVX1 U433 ( .A(n2193), .Y(n358) );
  INVX2 U434 ( .A(n2029), .Y(n560) );
  INVX1 U435 ( .A(n429), .Y(n360) );
  INVX1 U436 ( .A(n429), .Y(n361) );
  MUX2X1 U437 ( .B(n363), .A(n567), .S(n2162), .Y(n362) );
  INVX8 U438 ( .A(n362), .Y(n1938) );
  INVX8 U439 ( .A(n1939), .Y(n363) );
  MUX2X1 U440 ( .B(n365), .A(n570), .S(n22), .Y(n364) );
  INVX8 U441 ( .A(n364), .Y(n2023) );
  INVX8 U442 ( .A(n2024), .Y(n365) );
  INVX1 U443 ( .A(n187), .Y(n2041) );
  INVX1 U444 ( .A(n416), .Y(n367) );
  INVX1 U445 ( .A(net79541), .Y(net80775) );
  MUX2X1 U446 ( .B(n568), .A(buff_data[67]), .S(n531), .Y(n4015) );
  INVX8 U447 ( .A(n560), .Y(n368) );
  INVX1 U448 ( .A(n551), .Y(n369) );
  INVX2 U449 ( .A(n2052), .Y(n552) );
  INVX1 U450 ( .A(n98), .Y(n371) );
  INVX1 U451 ( .A(n2035), .Y(n372) );
  INVX1 U452 ( .A(n2035), .Y(n2196) );
  INVX1 U453 ( .A(n538), .Y(n373) );
  MUX2X1 U454 ( .B(n569), .A(n375), .S(n2076), .Y(n374) );
  INVX8 U455 ( .A(n374), .Y(n1964) );
  INVX8 U456 ( .A(n1965), .Y(n375) );
  INVX1 U457 ( .A(n551), .Y(n2049) );
  AND2X1 U458 ( .A(n549), .B(n376), .Y(net80232) );
  AND2X1 U459 ( .A(net66007), .B(ready), .Y(n376) );
  BUFX2 U460 ( .A(n445), .Y(n377) );
  INVX4 U461 ( .A(n445), .Y(n2162) );
  INVX1 U462 ( .A(net79794), .Y(n378) );
  INVX1 U463 ( .A(RETURN_full), .Y(n380) );
  INVX2 U464 ( .A(n420), .Y(n423) );
  OR2X1 U465 ( .A(n2407), .B(n2442), .Y(net89543) );
  INVX1 U466 ( .A(n4205), .Y(n381) );
  INVX2 U467 ( .A(n428), .Y(n384) );
  INVX2 U468 ( .A(n428), .Y(n401) );
  MUX2X1 U469 ( .B(n383), .A(n574), .S(n170), .Y(n382) );
  INVX8 U470 ( .A(n382), .Y(n1929) );
  INVX8 U471 ( .A(n1930), .Y(n383) );
  MUX2X1 U472 ( .B(n573), .A(buff_data[0]), .S(n2117), .Y(n3950) );
  INVX1 U473 ( .A(n2116), .Y(n2117) );
  OR2X2 U474 ( .A(n380), .B(n555), .Y(n385) );
  INVX1 U475 ( .A(n554), .Y(net92764) );
  INVX1 U476 ( .A(n33), .Y(n2040) );
  INVX1 U477 ( .A(n4), .Y(n386) );
  INVX1 U478 ( .A(n425), .Y(n387) );
  MUX2X1 U479 ( .B(n571), .A(n389), .S(n401), .Y(n388) );
  INVX8 U480 ( .A(n388), .Y(n2067) );
  INVX8 U481 ( .A(n2068), .Y(n389) );
  MUX2X1 U482 ( .B(n570), .A(n391), .S(n401), .Y(n390) );
  INVX8 U483 ( .A(n390), .Y(n2050) );
  INVX8 U484 ( .A(n2051), .Y(n391) );
  MUX2X1 U485 ( .B(n569), .A(n393), .S(n401), .Y(n392) );
  INVX8 U486 ( .A(n392), .Y(n2063) );
  INVX8 U487 ( .A(n2064), .Y(n393) );
  MUX2X1 U488 ( .B(n574), .A(n395), .S(n55), .Y(n394) );
  INVX8 U489 ( .A(n394), .Y(n2147) );
  INVX8 U490 ( .A(n2148), .Y(n395) );
  MUX2X1 U491 ( .B(n564), .A(n397), .S(n54), .Y(n396) );
  INVX8 U492 ( .A(n396), .Y(n1958) );
  INVX8 U493 ( .A(n1959), .Y(n397) );
  INVX1 U494 ( .A(n544), .Y(n2127) );
  INVX1 U495 ( .A(n1922), .Y(n544) );
  INVX1 U496 ( .A(n1911), .Y(n399) );
  INVX1 U497 ( .A(n399), .Y(n400) );
  INVX1 U498 ( .A(n403), .Y(n402) );
  INVX1 U499 ( .A(n80), .Y(n403) );
  INVX1 U500 ( .A(net65981), .Y(net82094) );
  OR2X2 U501 ( .A(n387), .B(n405), .Y(n404) );
  INVX8 U502 ( .A(net66482), .Y(n405) );
  MUX2X1 U503 ( .B(n568), .A(buff_data[227]), .S(n328), .Y(n4150) );
  MUX2X1 U504 ( .B(n573), .A(buff_data[224]), .S(n328), .Y(n4149) );
  INVX1 U505 ( .A(n1802), .Y(n407) );
  INVX1 U506 ( .A(n72), .Y(n408) );
  INVX1 U507 ( .A(n218), .Y(n409) );
  MUX2X1 U508 ( .B(n411), .A(n568), .S(n2038), .Y(n410) );
  INVX8 U509 ( .A(n410), .Y(n2133) );
  INVX8 U510 ( .A(n2134), .Y(n411) );
  INVX1 U511 ( .A(n2193), .Y(n2036) );
  MUX2X1 U512 ( .B(n413), .A(n566), .S(n2039), .Y(n412) );
  INVX8 U513 ( .A(n412), .Y(n2008) );
  INVX8 U514 ( .A(n2009), .Y(n413) );
  INVX1 U515 ( .A(n1931), .Y(n414) );
  INVX1 U516 ( .A(n98), .Y(n415) );
  INVX1 U517 ( .A(n1931), .Y(n2048) );
  INVX1 U518 ( .A(n2161), .Y(n2160) );
  INVX1 U519 ( .A(net66714), .Y(n416) );
  INVX1 U520 ( .A(net66714), .Y(n417) );
  INVX1 U521 ( .A(net66714), .Y(net79541) );
  INVX1 U522 ( .A(n2161), .Y(n418) );
  INVX1 U523 ( .A(n294), .Y(n419) );
  INVX4 U524 ( .A(n1997), .Y(n426) );
  INVX1 U525 ( .A(n3565), .Y(n420) );
  INVX1 U526 ( .A(n420), .Y(n421) );
  INVX1 U527 ( .A(n420), .Y(n422) );
  INVX1 U528 ( .A(n1807), .Y(n424) );
  INVX1 U529 ( .A(n441), .Y(n425) );
  NOR3X1 U530 ( .A(net82094), .B(n1998), .C(n1494), .Y(n427) );
  INVX4 U531 ( .A(n427), .Y(n3565) );
  AND2X2 U532 ( .A(n425), .B(net66482), .Y(n428) );
  INVX1 U533 ( .A(net92746), .Y(n539) );
  INVX1 U534 ( .A(n232), .Y(net66329) );
  OR2X2 U535 ( .A(n539), .B(n430), .Y(n429) );
  INVX8 U536 ( .A(net66482), .Y(n430) );
  INVX1 U537 ( .A(n4440), .Y(n434) );
  INVX1 U538 ( .A(n468), .Y(n435) );
  INVX1 U539 ( .A(n468), .Y(n436) );
  INVX1 U540 ( .A(n468), .Y(n2078) );
  BUFX2 U541 ( .A(n4508), .Y(n437) );
  INVX1 U542 ( .A(RETURN_full), .Y(n1807) );
  INVX8 U543 ( .A(n229), .Y(net79440) );
  OR2X2 U544 ( .A(n441), .B(n439), .Y(n438) );
  INVX8 U545 ( .A(n3963), .Y(n439) );
  INVX1 U546 ( .A(n2192), .Y(n2193) );
  INVX1 U547 ( .A(n4218), .Y(n2192) );
  INVX1 U548 ( .A(n535), .Y(n441) );
  INVX1 U549 ( .A(n2000), .Y(n2002) );
  INVX1 U550 ( .A(n98), .Y(n2035) );
  INVX1 U551 ( .A(n116), .Y(n442) );
  OR2X2 U552 ( .A(n539), .B(n446), .Y(n445) );
  INVX8 U553 ( .A(n3963), .Y(n446) );
  INVX1 U554 ( .A(n325), .Y(n2197) );
  INVX2 U555 ( .A(n2073), .Y(n468) );
  INVX1 U556 ( .A(n535), .Y(net92867) );
  INVX2 U557 ( .A(n1973), .Y(n467) );
  INVX8 U558 ( .A(n467), .Y(net80376) );
  INVX8 U559 ( .A(n438), .Y(n2191) );
  INVX4 U560 ( .A(n3630), .Y(n3568) );
  AND2X2 U561 ( .A(CMD_data_out[30]), .B(n3571), .Y(n3578) );
  INVX2 U562 ( .A(n1740), .Y(n1741) );
  OR2X2 U563 ( .A(n780), .B(n529), .Y(n4440) );
  INVX1 U564 ( .A(n4440), .Y(n447) );
  OR2X1 U565 ( .A(n1033), .B(n1035), .Y(n4389) );
  INVX1 U566 ( .A(n4389), .Y(n448) );
  OR2X1 U567 ( .A(n1046), .B(n1049), .Y(n4394) );
  INVX1 U568 ( .A(n4394), .Y(n449) );
  OR2X1 U569 ( .A(n1059), .B(n1061), .Y(n4396) );
  INVX1 U570 ( .A(n4396), .Y(n450) );
  OR2X1 U571 ( .A(n1070), .B(n1073), .Y(n4398) );
  INVX1 U572 ( .A(n4398), .Y(n451) );
  OR2X1 U573 ( .A(n1084), .B(n1087), .Y(n4400) );
  INVX1 U574 ( .A(n4400), .Y(n452) );
  OR2X1 U575 ( .A(n1098), .B(n1101), .Y(n4402) );
  INVX1 U576 ( .A(n4402), .Y(n453) );
  OR2X1 U577 ( .A(n1112), .B(n1115), .Y(n4404) );
  INVX1 U578 ( .A(n4404), .Y(n454) );
  OR2X1 U579 ( .A(n1126), .B(n1129), .Y(n4406) );
  INVX1 U580 ( .A(n4406), .Y(n455) );
  OR2X1 U581 ( .A(n1139), .B(n1141), .Y(n4408) );
  INVX1 U582 ( .A(n4408), .Y(n456) );
  OR2X1 U583 ( .A(n1150), .B(n1153), .Y(n4410) );
  INVX1 U584 ( .A(n4410), .Y(n457) );
  OR2X1 U585 ( .A(n1164), .B(n1167), .Y(n4412) );
  INVX1 U586 ( .A(n4412), .Y(n458) );
  OR2X1 U587 ( .A(n1177), .B(n1179), .Y(n4414) );
  INVX1 U588 ( .A(n4414), .Y(n459) );
  OR2X1 U589 ( .A(n1188), .B(n1191), .Y(n4416) );
  INVX1 U590 ( .A(n4416), .Y(n460) );
  OR2X1 U591 ( .A(n1201), .B(n1203), .Y(n4420) );
  INVX1 U592 ( .A(n4420), .Y(n461) );
  AND2X2 U593 ( .A(net92619), .B(net66441), .Y(n1804) );
  AND2X2 U594 ( .A(n10), .B(net66441), .Y(net82538) );
  AND2X2 U595 ( .A(net92651), .B(net92761), .Y(net80791) );
  INVX1 U596 ( .A(net80791), .Y(n463) );
  AND2X2 U597 ( .A(n1810), .B(n1808), .Y(net89563) );
  INVX1 U598 ( .A(net89563), .Y(n464) );
  INVX1 U599 ( .A(net80232), .Y(n465) );
  AND2X2 U600 ( .A(n1847), .B(net92764), .Y(n1834) );
  AND2X2 U601 ( .A(net92619), .B(n4056), .Y(n1842) );
  AND2X2 U602 ( .A(n535), .B(net66423), .Y(n1966) );
  AND2X2 U603 ( .A(net66539), .B(net93077), .Y(n1973) );
  AND2X2 U604 ( .A(net66503), .B(n378), .Y(n2073) );
  AND2X2 U605 ( .A(n607), .B(CMD_data_out[3]), .Y(n3512) );
  INVX1 U606 ( .A(n3512), .Y(n469) );
  OR2X2 U607 ( .A(n866), .B(n1581), .Y(n4516) );
  INVX1 U608 ( .A(n4516), .Y(n470) );
  BUFX2 U609 ( .A(n3651), .Y(n471) );
  BUFX2 U610 ( .A(n3772), .Y(n472) );
  AND2X2 U611 ( .A(n424), .B(n1834), .Y(n1846) );
  INVX1 U612 ( .A(n1846), .Y(n473) );
  AND2X1 U613 ( .A(n1894), .B(n3914), .Y(n4513) );
  INVX1 U614 ( .A(n4513), .Y(n474) );
  BUFX2 U615 ( .A(n3570), .Y(n475) );
  BUFX2 U616 ( .A(n3574), .Y(n476) );
  BUFX2 U617 ( .A(n3577), .Y(n477) );
  BUFX2 U618 ( .A(n3916), .Y(n478) );
  AND2X2 U619 ( .A(n1780), .B(n3568), .Y(n3567) );
  INVX1 U620 ( .A(n3567), .Y(n479) );
  AND2X2 U621 ( .A(n634), .B(n3641), .Y(n3640) );
  INVX1 U622 ( .A(n3640), .Y(n480) );
  AND2X2 U623 ( .A(n284), .B(n1788), .Y(n3644) );
  INVX1 U624 ( .A(n3644), .Y(n481) );
  AND2X2 U625 ( .A(n984), .B(n3641), .Y(n3710) );
  INVX1 U626 ( .A(n3710), .Y(n482) );
  AND2X2 U627 ( .A(n983), .B(n3641), .Y(n3711) );
  INVX1 U628 ( .A(n3711), .Y(n483) );
  AND2X2 U629 ( .A(n982), .B(n3641), .Y(n3712) );
  INVX1 U630 ( .A(n3712), .Y(n484) );
  AND2X2 U631 ( .A(n981), .B(n3641), .Y(n3713) );
  INVX1 U632 ( .A(n3713), .Y(n485) );
  AND2X2 U633 ( .A(n980), .B(n3641), .Y(n3714) );
  INVX1 U634 ( .A(n3714), .Y(n486) );
  AND2X2 U635 ( .A(n979), .B(n3641), .Y(n3715) );
  INVX1 U636 ( .A(n3715), .Y(n487) );
  AND2X2 U637 ( .A(n978), .B(n3641), .Y(n3716) );
  INVX1 U638 ( .A(n3716), .Y(n488) );
  AND2X2 U639 ( .A(n977), .B(n3641), .Y(n3717) );
  INVX1 U640 ( .A(n3717), .Y(n489) );
  AND2X2 U641 ( .A(n976), .B(n3641), .Y(n3718) );
  INVX1 U642 ( .A(n3718), .Y(n490) );
  AND2X2 U643 ( .A(n942), .B(n3641), .Y(n3719) );
  INVX1 U644 ( .A(n3719), .Y(n491) );
  AND2X2 U645 ( .A(n907), .B(n3641), .Y(n3720) );
  INVX1 U646 ( .A(n3720), .Y(n492) );
  AND2X2 U647 ( .A(n873), .B(n3641), .Y(n3721) );
  INVX1 U648 ( .A(n3721), .Y(n493) );
  AND2X2 U649 ( .A(n839), .B(n3641), .Y(n3722) );
  INVX1 U650 ( .A(n3722), .Y(n494) );
  AND2X2 U651 ( .A(n805), .B(n3641), .Y(n3723) );
  INVX1 U652 ( .A(n3723), .Y(n495) );
  AND2X2 U653 ( .A(n737), .B(n3641), .Y(n3724) );
  INVX1 U654 ( .A(n3724), .Y(n496) );
  AND2X2 U655 ( .A(n703), .B(n3641), .Y(n3725) );
  INVX1 U656 ( .A(n3725), .Y(n497) );
  AND2X2 U657 ( .A(n669), .B(n3641), .Y(n3726) );
  INVX1 U658 ( .A(n3726), .Y(n498) );
  AND2X2 U659 ( .A(n648), .B(n3641), .Y(n3727) );
  INVX1 U660 ( .A(n3727), .Y(n499) );
  AND2X2 U661 ( .A(n647), .B(n3641), .Y(n3728) );
  INVX1 U662 ( .A(n3728), .Y(n500) );
  AND2X2 U663 ( .A(n646), .B(n3641), .Y(n3729) );
  INVX1 U664 ( .A(n3729), .Y(n501) );
  AND2X2 U665 ( .A(n645), .B(n3641), .Y(n3730) );
  INVX1 U666 ( .A(n3730), .Y(n502) );
  AND2X2 U667 ( .A(n644), .B(n3641), .Y(n3731) );
  INVX1 U668 ( .A(n3731), .Y(n503) );
  AND2X2 U669 ( .A(n643), .B(n3641), .Y(n3732) );
  INVX1 U670 ( .A(n3732), .Y(n504) );
  AND2X2 U671 ( .A(n642), .B(n3641), .Y(n3734) );
  INVX1 U672 ( .A(n3734), .Y(n505) );
  AND2X2 U673 ( .A(n641), .B(n3641), .Y(n3736) );
  INVX1 U674 ( .A(n3736), .Y(n506) );
  AND2X2 U675 ( .A(n640), .B(n3641), .Y(n3738) );
  INVX1 U676 ( .A(n3738), .Y(n507) );
  AND2X2 U677 ( .A(n639), .B(n3641), .Y(n3740) );
  INVX1 U678 ( .A(n3740), .Y(n508) );
  AND2X2 U679 ( .A(n638), .B(n3641), .Y(n3742) );
  INVX1 U680 ( .A(n3742), .Y(n509) );
  AND2X2 U681 ( .A(n637), .B(n3641), .Y(n3744) );
  INVX1 U682 ( .A(n3744), .Y(n510) );
  AND2X2 U683 ( .A(n636), .B(n3641), .Y(n3746) );
  INVX1 U684 ( .A(n3746), .Y(n511) );
  AND2X2 U685 ( .A(n283), .B(n1788), .Y(n3840) );
  INVX1 U686 ( .A(n3840), .Y(n512) );
  AND2X2 U687 ( .A(n2110), .B(n3925), .Y(net66380) );
  INVX1 U688 ( .A(net66380), .Y(n513) );
  AND2X2 U689 ( .A(n2111), .B(n3925), .Y(n3947) );
  INVX1 U690 ( .A(n3947), .Y(n514) );
  AND2X2 U691 ( .A(n2112), .B(n3925), .Y(n3948) );
  INVX1 U692 ( .A(n3948), .Y(n515) );
  BUFX2 U693 ( .A(n4438), .Y(n516) );
  BUFX2 U694 ( .A(n4443), .Y(n517) );
  BUFX2 U695 ( .A(n4445), .Y(n518) );
  AND2X2 U696 ( .A(CMD_data_out[13]), .B(n4451), .Y(n4455) );
  INVX1 U697 ( .A(n4455), .Y(n519) );
  AND2X2 U698 ( .A(CMD_data_out[14]), .B(n4451), .Y(n4461) );
  INVX1 U699 ( .A(n4461), .Y(n520) );
  AND2X2 U700 ( .A(CMD_data_out[15]), .B(n4451), .Y(n4467) );
  INVX1 U701 ( .A(n4467), .Y(n521) );
  AND2X2 U702 ( .A(CMD_data_out[16]), .B(n4451), .Y(n4472) );
  INVX1 U703 ( .A(n4472), .Y(n522) );
  AND2X2 U704 ( .A(CMD_data_out[17]), .B(n4451), .Y(n4477) );
  INVX1 U705 ( .A(n4477), .Y(n523) );
  AND2X2 U706 ( .A(CMD_data_out[18]), .B(n4451), .Y(n4482) );
  INVX1 U707 ( .A(n4482), .Y(n524) );
  AND2X2 U708 ( .A(CMD_data_out[19]), .B(n4451), .Y(n4487) );
  INVX1 U709 ( .A(n4487), .Y(n525) );
  AND2X2 U710 ( .A(CMD_data_out[20]), .B(n4451), .Y(n4492) );
  INVX1 U711 ( .A(n4492), .Y(n526) );
  AND2X2 U712 ( .A(CMD_data_out[21]), .B(n4451), .Y(n4497) );
  INVX1 U713 ( .A(n4497), .Y(n527) );
  AND2X2 U714 ( .A(CMD_data_out[22]), .B(n4451), .Y(n4502) );
  INVX1 U715 ( .A(n4502), .Y(n528) );
  BUFX2 U716 ( .A(n4507), .Y(n529) );
  BUFX2 U717 ( .A(n3895), .Y(n530) );
  AND2X2 U718 ( .A(n82), .B(net66423), .Y(n1931) );
  BUFX2 U719 ( .A(n3893), .Y(n532) );
  BUFX2 U720 ( .A(n3903), .Y(n533) );
  AND2X2 U721 ( .A(n770), .B(n474), .Y(n4505) );
  INVX1 U722 ( .A(n4505), .Y(n534) );
  BUFX2 U723 ( .A(net66558), .Y(n535) );
  AND2X2 U724 ( .A(net89705), .B(n4011), .Y(n1801) );
  INVX1 U725 ( .A(n6), .Y(n536) );
  OR2X2 U726 ( .A(net80595), .B(n1803), .Y(n1802) );
  AND2X2 U727 ( .A(net92747), .B(net92748), .Y(net92746) );
  INVX1 U728 ( .A(net92746), .Y(n538) );
  AND2X2 U729 ( .A(n471), .B(n1692), .Y(n3650) );
  INVX1 U730 ( .A(n3650), .Y(n540) );
  AND2X2 U731 ( .A(net82506), .B(n1808), .Y(net66168) );
  INVX1 U732 ( .A(net66168), .Y(n541) );
  INVX1 U733 ( .A(net66168), .Y(n542) );
  INVX1 U734 ( .A(n2129), .Y(n543) );
  AND2X2 U735 ( .A(net80598), .B(net66482), .Y(n1922) );
  BUFX2 U736 ( .A(n2188), .Y(n545) );
  AND2X2 U737 ( .A(net92619), .B(net66423), .Y(n611) );
  INVX1 U738 ( .A(n149), .Y(n546) );
  AND2X2 U739 ( .A(n1845), .B(n473), .Y(net92751) );
  INVX1 U740 ( .A(net92751), .Y(n547) );
  INVX1 U741 ( .A(net92751), .Y(n548) );
  BUFX2 U742 ( .A(CMD_empty), .Y(n549) );
  AND2X2 U743 ( .A(net66539), .B(n10), .Y(n1911) );
  AND2X2 U744 ( .A(net66423), .B(net80518), .Y(n2052) );
  AND2X2 U745 ( .A(n1224), .B(n1813), .Y(net92735) );
  INVX1 U746 ( .A(net92735), .Y(n554) );
  INVX1 U747 ( .A(net92735), .Y(n555) );
  AND2X2 U748 ( .A(net92619), .B(n4011), .Y(n1841) );
  AND2X2 U749 ( .A(net66441), .B(net80518), .Y(net80322) );
  AND2X2 U750 ( .A(net80518), .B(n4011), .Y(n1972) );
  AND2X2 U751 ( .A(n4056), .B(n1800), .Y(n2029) );
  AND2X2 U752 ( .A(net66539), .B(net92619), .Y(n1825) );
  INVX1 U753 ( .A(n1825), .Y(n561) );
  AND2X2 U754 ( .A(net92761), .B(n1227), .Y(n1848) );
  BUFX2 U755 ( .A(DATA_data_out[10]), .Y(n564) );
  BUFX2 U756 ( .A(DATA_data_out[9]), .Y(n565) );
  BUFX2 U757 ( .A(DATA_data_out[8]), .Y(n566) );
  BUFX2 U758 ( .A(DATA_data_out[14]), .Y(n567) );
  BUFX2 U759 ( .A(DATA_data_out[3]), .Y(n568) );
  BUFX2 U760 ( .A(DATA_data_out[5]), .Y(n569) );
  BUFX2 U761 ( .A(DATA_data_out[6]), .Y(n570) );
  BUFX2 U762 ( .A(DATA_data_out[11]), .Y(n571) );
  BUFX2 U763 ( .A(DATA_data_out[12]), .Y(n572) );
  BUFX2 U764 ( .A(DATA_data_out[0]), .Y(n573) );
  BUFX2 U765 ( .A(DATA_data_out[2]), .Y(n574) );
  BUFX2 U766 ( .A(DATA_data_out[15]), .Y(n575) );
  BUFX2 U767 ( .A(DATA_data_out[4]), .Y(n576) );
  BUFX2 U768 ( .A(DATA_data_out[1]), .Y(n577) );
  BUFX2 U769 ( .A(DATA_data_out[7]), .Y(n578) );
  BUFX2 U770 ( .A(DATA_data_out[13]), .Y(n579) );
  AND2X2 U771 ( .A(n3579), .B(n426), .Y(n3571) );
  AND2X2 U772 ( .A(net80596), .B(net66539), .Y(n580) );
  AND2X1 U773 ( .A(CMD_data_out[0]), .B(CMD_data_out[1]), .Y(n581) );
  AND2X2 U774 ( .A(n1755), .B(n3568), .Y(n3581) );
  INVX1 U775 ( .A(n3581), .Y(n582) );
  AND2X2 U776 ( .A(n1756), .B(n3568), .Y(n3583) );
  INVX1 U777 ( .A(n3583), .Y(n583) );
  AND2X2 U778 ( .A(n1757), .B(n3568), .Y(n3585) );
  INVX1 U779 ( .A(n3585), .Y(n584) );
  AND2X2 U780 ( .A(n1758), .B(n3568), .Y(n3587) );
  INVX1 U781 ( .A(n3587), .Y(n585) );
  AND2X2 U782 ( .A(n1759), .B(n3568), .Y(n3589) );
  INVX1 U783 ( .A(n3589), .Y(n586) );
  AND2X2 U784 ( .A(n1760), .B(n3568), .Y(n3591) );
  INVX1 U785 ( .A(n3591), .Y(n587) );
  AND2X2 U786 ( .A(n1761), .B(n3568), .Y(n3593) );
  INVX1 U787 ( .A(n3593), .Y(n588) );
  AND2X2 U788 ( .A(n1762), .B(n3568), .Y(n3595) );
  INVX1 U789 ( .A(n3595), .Y(n589) );
  AND2X2 U790 ( .A(n1763), .B(n3568), .Y(n3597) );
  INVX1 U791 ( .A(n3597), .Y(n590) );
  AND2X2 U792 ( .A(n1764), .B(n3568), .Y(n3599) );
  INVX1 U793 ( .A(n3599), .Y(n591) );
  AND2X2 U794 ( .A(n1765), .B(n3568), .Y(n3601) );
  INVX1 U795 ( .A(n3601), .Y(n592) );
  AND2X2 U796 ( .A(n1766), .B(n3568), .Y(n3603) );
  INVX1 U797 ( .A(n3603), .Y(n593) );
  AND2X2 U798 ( .A(n1767), .B(n3568), .Y(n3605) );
  INVX1 U799 ( .A(n3605), .Y(n594) );
  AND2X2 U800 ( .A(n1768), .B(n3568), .Y(n3607) );
  INVX1 U801 ( .A(n3607), .Y(n595) );
  AND2X2 U802 ( .A(n1769), .B(n3568), .Y(n3609) );
  INVX1 U803 ( .A(n3609), .Y(n596) );
  AND2X2 U804 ( .A(n1770), .B(n3568), .Y(n3611) );
  INVX1 U805 ( .A(n3611), .Y(n597) );
  AND2X2 U806 ( .A(n1771), .B(n3568), .Y(n3613) );
  INVX1 U807 ( .A(n3613), .Y(n598) );
  AND2X2 U808 ( .A(n1772), .B(n3568), .Y(n3615) );
  INVX1 U809 ( .A(n3615), .Y(n599) );
  AND2X2 U810 ( .A(n1773), .B(n3568), .Y(n3617) );
  INVX1 U811 ( .A(n3617), .Y(n600) );
  AND2X2 U812 ( .A(n1774), .B(n3568), .Y(n3619) );
  INVX1 U813 ( .A(n3619), .Y(n601) );
  AND2X2 U814 ( .A(n1775), .B(n3568), .Y(n3621) );
  INVX1 U815 ( .A(n3621), .Y(n602) );
  AND2X2 U816 ( .A(n1776), .B(n3568), .Y(n3623) );
  INVX1 U817 ( .A(n3623), .Y(n603) );
  AND2X2 U818 ( .A(n1777), .B(n3568), .Y(n3625) );
  INVX1 U819 ( .A(n3625), .Y(n604) );
  AND2X2 U820 ( .A(n1778), .B(n3568), .Y(n3627) );
  INVX1 U821 ( .A(n3627), .Y(n605) );
  AND2X2 U822 ( .A(n1779), .B(n3568), .Y(n3629) );
  INVX1 U823 ( .A(n3629), .Y(n606) );
  OR2X1 U824 ( .A(n231), .B(n232), .Y(net92738) );
  AND2X1 U825 ( .A(n581), .B(CMD_data_out[2]), .Y(n607) );
  BUFX2 U826 ( .A(add_576_carry_7_), .Y(n608) );
  INVX1 U827 ( .A(n469), .Y(add_576_carry_7_) );
  BUFX2 U828 ( .A(n549), .Y(n609) );
  INVX1 U829 ( .A(n149), .Y(n610) );
  INVX1 U830 ( .A(n4457), .Y(n612) );
  INVX1 U831 ( .A(n612), .Y(n613) );
  INVX1 U832 ( .A(n4463), .Y(n614) );
  INVX1 U833 ( .A(n614), .Y(n615) );
  INVX1 U834 ( .A(n4469), .Y(n616) );
  INVX1 U835 ( .A(n616), .Y(n617) );
  INVX1 U836 ( .A(n4474), .Y(n618) );
  INVX1 U837 ( .A(n618), .Y(n619) );
  INVX1 U838 ( .A(n4479), .Y(n620) );
  INVX1 U839 ( .A(n620), .Y(n621) );
  INVX1 U840 ( .A(n4484), .Y(n622) );
  INVX1 U841 ( .A(n622), .Y(n623) );
  INVX1 U842 ( .A(n4489), .Y(n628) );
  INVX1 U843 ( .A(n628), .Y(n629) );
  INVX1 U844 ( .A(n4494), .Y(n630) );
  INVX1 U845 ( .A(n630), .Y(n631) );
  INVX1 U846 ( .A(n4499), .Y(n632) );
  INVX1 U847 ( .A(n632), .Y(n633) );
  INVX1 U848 ( .A(n651), .Y(n649) );
  INVX1 U849 ( .A(n649), .Y(n650) );
  BUFX2 U850 ( .A(n3634), .Y(n651) );
  INVX1 U851 ( .A(n654), .Y(n652) );
  INVX1 U852 ( .A(n652), .Y(n653) );
  BUFX2 U853 ( .A(n3707), .Y(n654) );
  INVX1 U854 ( .A(n657), .Y(n655) );
  INVX1 U855 ( .A(n655), .Y(n656) );
  BUFX2 U856 ( .A(n4572), .Y(n657) );
  INVX1 U857 ( .A(n660), .Y(n658) );
  INVX1 U858 ( .A(n658), .Y(n659) );
  BUFX2 U859 ( .A(n4582), .Y(n660) );
  INVX1 U860 ( .A(n663), .Y(n661) );
  INVX1 U861 ( .A(n661), .Y(n662) );
  BUFX2 U862 ( .A(net66060), .Y(n663) );
  INVX1 U863 ( .A(n666), .Y(n664) );
  INVX1 U864 ( .A(n664), .Y(n665) );
  BUFX2 U865 ( .A(n4543), .Y(n666) );
  INVX1 U866 ( .A(n670), .Y(n667) );
  INVX1 U867 ( .A(n667), .Y(n668) );
  BUFX2 U868 ( .A(n3764), .Y(n670) );
  INVX1 U869 ( .A(n673), .Y(n671) );
  INVX1 U870 ( .A(n671), .Y(n672) );
  BUFX2 U871 ( .A(n4006), .Y(n673) );
  INVX1 U872 ( .A(n676), .Y(n674) );
  INVX1 U873 ( .A(n674), .Y(n675) );
  AND2X1 U874 ( .A(n253), .B(n1788), .Y(n3780) );
  INVX1 U875 ( .A(n3780), .Y(n676) );
  INVX1 U876 ( .A(n679), .Y(n677) );
  INVX1 U877 ( .A(n677), .Y(n678) );
  AND2X1 U878 ( .A(n255), .B(n1788), .Y(n3784) );
  INVX1 U879 ( .A(n3784), .Y(n679) );
  INVX1 U880 ( .A(n682), .Y(n680) );
  INVX1 U881 ( .A(n680), .Y(n681) );
  AND2X1 U882 ( .A(n256), .B(n1788), .Y(n3786) );
  INVX1 U883 ( .A(n3786), .Y(n682) );
  INVX1 U884 ( .A(n685), .Y(n683) );
  INVX1 U885 ( .A(n683), .Y(n684) );
  AND2X1 U886 ( .A(n257), .B(n1788), .Y(n3788) );
  INVX1 U887 ( .A(n3788), .Y(n685) );
  INVX1 U888 ( .A(n688), .Y(n686) );
  INVX1 U889 ( .A(n686), .Y(n687) );
  AND2X1 U890 ( .A(n258), .B(n1788), .Y(n3790) );
  INVX1 U891 ( .A(n3790), .Y(n688) );
  INVX1 U892 ( .A(n691), .Y(n689) );
  INVX1 U893 ( .A(n689), .Y(n690) );
  AND2X1 U894 ( .A(n259), .B(n1788), .Y(n3792) );
  INVX1 U895 ( .A(n3792), .Y(n691) );
  INVX1 U896 ( .A(n694), .Y(n692) );
  INVX1 U897 ( .A(n692), .Y(n693) );
  AND2X1 U898 ( .A(n260), .B(n1788), .Y(n3794) );
  INVX1 U899 ( .A(n3794), .Y(n694) );
  INVX1 U900 ( .A(n697), .Y(n695) );
  INVX1 U901 ( .A(n695), .Y(n696) );
  AND2X1 U902 ( .A(n261), .B(n1788), .Y(n3796) );
  INVX1 U903 ( .A(n3796), .Y(n697) );
  INVX1 U904 ( .A(n700), .Y(n698) );
  INVX1 U905 ( .A(n698), .Y(n699) );
  AND2X1 U906 ( .A(n262), .B(n1788), .Y(n3798) );
  INVX1 U907 ( .A(n3798), .Y(n700) );
  INVX1 U908 ( .A(n704), .Y(n701) );
  INVX1 U909 ( .A(n701), .Y(n702) );
  AND2X1 U910 ( .A(n263), .B(n1788), .Y(n3800) );
  INVX1 U911 ( .A(n3800), .Y(n704) );
  INVX1 U912 ( .A(n707), .Y(n705) );
  INVX1 U913 ( .A(n705), .Y(n706) );
  AND2X1 U914 ( .A(n264), .B(n1788), .Y(n3802) );
  INVX1 U915 ( .A(n3802), .Y(n707) );
  INVX1 U916 ( .A(n710), .Y(n708) );
  INVX1 U917 ( .A(n708), .Y(n709) );
  AND2X1 U918 ( .A(n265), .B(n1788), .Y(n3804) );
  INVX1 U919 ( .A(n3804), .Y(n710) );
  INVX1 U920 ( .A(n713), .Y(n711) );
  INVX1 U921 ( .A(n711), .Y(n712) );
  AND2X1 U922 ( .A(n266), .B(n1788), .Y(n3806) );
  INVX1 U923 ( .A(n3806), .Y(n713) );
  INVX1 U924 ( .A(n716), .Y(n714) );
  INVX1 U925 ( .A(n714), .Y(n715) );
  AND2X1 U926 ( .A(n267), .B(n1788), .Y(n3808) );
  INVX1 U927 ( .A(n3808), .Y(n716) );
  INVX1 U928 ( .A(n719), .Y(n717) );
  INVX1 U929 ( .A(n717), .Y(n718) );
  AND2X1 U930 ( .A(n268), .B(n1788), .Y(n3810) );
  INVX1 U931 ( .A(n3810), .Y(n719) );
  INVX1 U932 ( .A(n722), .Y(n720) );
  INVX1 U933 ( .A(n720), .Y(n721) );
  AND2X1 U934 ( .A(n269), .B(n1788), .Y(n3812) );
  INVX1 U935 ( .A(n3812), .Y(n722) );
  INVX1 U936 ( .A(n725), .Y(n723) );
  INVX1 U937 ( .A(n723), .Y(n724) );
  AND2X1 U938 ( .A(n270), .B(n1788), .Y(n3814) );
  INVX1 U939 ( .A(n3814), .Y(n725) );
  INVX1 U940 ( .A(n728), .Y(n726) );
  INVX1 U941 ( .A(n726), .Y(n727) );
  AND2X1 U942 ( .A(n271), .B(n1788), .Y(n3816) );
  INVX1 U943 ( .A(n3816), .Y(n728) );
  INVX1 U944 ( .A(n731), .Y(n729) );
  INVX1 U945 ( .A(n729), .Y(n730) );
  AND2X1 U946 ( .A(n272), .B(n1788), .Y(n3818) );
  INVX1 U947 ( .A(n3818), .Y(n731) );
  INVX1 U948 ( .A(n734), .Y(n732) );
  INVX1 U949 ( .A(n732), .Y(n733) );
  AND2X1 U950 ( .A(n273), .B(n1788), .Y(n3820) );
  INVX1 U951 ( .A(n3820), .Y(n734) );
  INVX1 U952 ( .A(n738), .Y(n735) );
  INVX1 U953 ( .A(n735), .Y(n736) );
  AND2X1 U954 ( .A(n274), .B(n1788), .Y(n3822) );
  INVX1 U955 ( .A(n3822), .Y(n738) );
  INVX1 U956 ( .A(n741), .Y(n739) );
  INVX1 U957 ( .A(n739), .Y(n740) );
  AND2X1 U958 ( .A(n275), .B(n1788), .Y(n3824) );
  INVX1 U959 ( .A(n3824), .Y(n741) );
  INVX1 U960 ( .A(n744), .Y(n742) );
  INVX1 U961 ( .A(n742), .Y(n743) );
  AND2X1 U962 ( .A(n276), .B(n1788), .Y(n3826) );
  INVX1 U963 ( .A(n3826), .Y(n744) );
  INVX1 U964 ( .A(n747), .Y(n745) );
  INVX1 U965 ( .A(n745), .Y(n746) );
  AND2X1 U966 ( .A(n277), .B(n1788), .Y(n3828) );
  INVX1 U967 ( .A(n3828), .Y(n747) );
  INVX1 U968 ( .A(n750), .Y(n748) );
  INVX1 U969 ( .A(n748), .Y(n749) );
  AND2X1 U970 ( .A(n278), .B(n1788), .Y(n3830) );
  INVX1 U971 ( .A(n3830), .Y(n750) );
  INVX1 U972 ( .A(n753), .Y(n751) );
  INVX1 U973 ( .A(n751), .Y(n752) );
  AND2X1 U974 ( .A(n279), .B(n1788), .Y(n3832) );
  INVX1 U975 ( .A(n3832), .Y(n753) );
  INVX1 U976 ( .A(n756), .Y(n754) );
  INVX1 U977 ( .A(n754), .Y(n755) );
  AND2X1 U978 ( .A(n280), .B(n1788), .Y(n3834) );
  INVX1 U979 ( .A(n3834), .Y(n756) );
  INVX1 U980 ( .A(n759), .Y(n757) );
  INVX1 U981 ( .A(n757), .Y(n758) );
  AND2X1 U982 ( .A(n281), .B(n1788), .Y(n3836) );
  INVX1 U983 ( .A(n3836), .Y(n759) );
  INVX1 U984 ( .A(n762), .Y(n760) );
  INVX1 U985 ( .A(n760), .Y(n761) );
  AND2X1 U986 ( .A(n282), .B(n1788), .Y(n3838) );
  INVX1 U987 ( .A(n3838), .Y(n762) );
  INVX1 U988 ( .A(n765), .Y(n763) );
  INVX1 U989 ( .A(n763), .Y(n764) );
  BUFX2 U990 ( .A(n4418), .Y(n765) );
  INVX1 U991 ( .A(n768), .Y(n766) );
  INVX1 U992 ( .A(n766), .Y(n767) );
  BUFX2 U993 ( .A(n4422), .Y(n768) );
  INVX1 U994 ( .A(n4512), .Y(n769) );
  INVX1 U995 ( .A(n769), .Y(n770) );
  INVX1 U996 ( .A(n450), .Y(n771) );
  INVX1 U997 ( .A(n771), .Y(n772) );
  INVX1 U998 ( .A(n456), .Y(n773) );
  INVX1 U999 ( .A(n773), .Y(n774) );
  INVX1 U1000 ( .A(n459), .Y(n775) );
  INVX1 U1001 ( .A(n775), .Y(n776) );
  INVX1 U1002 ( .A(n461), .Y(n777) );
  INVX1 U1003 ( .A(n777), .Y(n778) );
  INVX1 U1004 ( .A(n781), .Y(n779) );
  INVX1 U1005 ( .A(n779), .Y(n780) );
  BUFX2 U1006 ( .A(n4506), .Y(n781) );
  AND2X2 U1007 ( .A(n472), .B(n1627), .Y(n3760) );
  INVX1 U1008 ( .A(n784), .Y(n782) );
  INVX1 U1009 ( .A(n782), .Y(n783) );
  BUFX2 U1010 ( .A(n3888), .Y(n784) );
  INVX1 U1011 ( .A(n787), .Y(n785) );
  INVX1 U1012 ( .A(n785), .Y(n786) );
  BUFX2 U1013 ( .A(n3853), .Y(n787) );
  INVX1 U1014 ( .A(n790), .Y(n788) );
  INVX1 U1015 ( .A(n788), .Y(n789) );
  BUFX2 U1016 ( .A(n4557), .Y(n790) );
  INVX1 U1017 ( .A(n793), .Y(n791) );
  INVX1 U1018 ( .A(n791), .Y(n792) );
  BUFX2 U1019 ( .A(n4559), .Y(n793) );
  INVX1 U1020 ( .A(n796), .Y(n794) );
  INVX1 U1021 ( .A(n794), .Y(n795) );
  BUFX2 U1022 ( .A(n4585), .Y(n796) );
  INVX1 U1023 ( .A(n799), .Y(n797) );
  INVX1 U1024 ( .A(n797), .Y(n798) );
  BUFX2 U1025 ( .A(n4623), .Y(n799) );
  INVX1 U1026 ( .A(n802), .Y(n800) );
  INVX1 U1027 ( .A(n800), .Y(n801) );
  BUFX2 U1028 ( .A(n4615), .Y(n802) );
  INVX1 U1029 ( .A(n806), .Y(n803) );
  INVX1 U1030 ( .A(n803), .Y(n804) );
  BUFX2 U1031 ( .A(n3854), .Y(n806) );
  INVX1 U1032 ( .A(n809), .Y(n807) );
  INVX1 U1033 ( .A(n807), .Y(n808) );
  BUFX2 U1034 ( .A(n4558), .Y(n809) );
  INVX1 U1035 ( .A(n812), .Y(n810) );
  INVX1 U1036 ( .A(n810), .Y(n811) );
  BUFX2 U1037 ( .A(n4560), .Y(n812) );
  INVX1 U1038 ( .A(n815), .Y(n813) );
  INVX1 U1039 ( .A(n813), .Y(n814) );
  BUFX2 U1040 ( .A(n4586), .Y(n815) );
  INVX1 U1041 ( .A(n818), .Y(n816) );
  INVX1 U1042 ( .A(n816), .Y(n817) );
  BUFX2 U1043 ( .A(n4616), .Y(n818) );
  INVX1 U1044 ( .A(n821), .Y(n819) );
  INVX1 U1045 ( .A(n819), .Y(n820) );
  BUFX2 U1046 ( .A(n4624), .Y(n821) );
  INVX1 U1047 ( .A(n824), .Y(n822) );
  INVX1 U1048 ( .A(n822), .Y(n823) );
  BUFX2 U1049 ( .A(n4424), .Y(n824) );
  INVX1 U1050 ( .A(n827), .Y(n825) );
  INVX1 U1051 ( .A(n825), .Y(n826) );
  BUFX2 U1052 ( .A(n4437), .Y(n827) );
  INVX1 U1053 ( .A(n830), .Y(n828) );
  INVX1 U1054 ( .A(n828), .Y(n829) );
  BUFX2 U1055 ( .A(n4556), .Y(n830) );
  INVX1 U1056 ( .A(n833), .Y(n831) );
  INVX1 U1057 ( .A(n831), .Y(n832) );
  BUFX2 U1058 ( .A(n4555), .Y(n833) );
  INVX1 U1059 ( .A(n836), .Y(n834) );
  INVX1 U1060 ( .A(n834), .Y(n835) );
  BUFX2 U1061 ( .A(n3904), .Y(n836) );
  INVX1 U1062 ( .A(n840), .Y(n837) );
  INVX1 U1063 ( .A(n837), .Y(n838) );
  BUFX2 U1064 ( .A(n3550), .Y(n840) );
  INVX1 U1065 ( .A(n843), .Y(n841) );
  INVX1 U1066 ( .A(n841), .Y(n842) );
  BUFX2 U1067 ( .A(n3692), .Y(n843) );
  INVX1 U1068 ( .A(n470), .Y(n844) );
  INVX1 U1069 ( .A(n844), .Y(n845) );
  INVX1 U1070 ( .A(net66970), .Y(n1810) );
  AND2X1 U1071 ( .A(add_576_carry_7_), .B(CMD_data_out[4]), .Y(n3513) );
  INVX1 U1072 ( .A(n3513), .Y(n846) );
  INVX1 U1073 ( .A(n846), .Y(add_576_carry_8_) );
  AND2X1 U1074 ( .A(add_576_carry_8_), .B(CMD_data_out[5]), .Y(n3514) );
  INVX1 U1075 ( .A(n3514), .Y(n847) );
  INVX1 U1076 ( .A(n847), .Y(add_576_carry_9_) );
  INVX1 U1077 ( .A(n850), .Y(n848) );
  INVX1 U1078 ( .A(n848), .Y(n849) );
  BUFX2 U1079 ( .A(n4590), .Y(n850) );
  INVX1 U1080 ( .A(n853), .Y(n851) );
  INVX1 U1081 ( .A(n851), .Y(n852) );
  BUFX2 U1082 ( .A(n3750), .Y(n853) );
  INVX1 U1083 ( .A(n856), .Y(n854) );
  INVX1 U1084 ( .A(n854), .Y(n855) );
  BUFX2 U1085 ( .A(n4562), .Y(n856) );
  INVX1 U1086 ( .A(n859), .Y(n857) );
  INVX1 U1087 ( .A(n857), .Y(n858) );
  BUFX2 U1088 ( .A(n3898), .Y(n859) );
  INVX1 U1089 ( .A(n861), .Y(n860) );
  BUFX2 U1090 ( .A(n4515), .Y(n861) );
  INVX1 U1091 ( .A(n3910), .Y(n862) );
  INVX1 U1092 ( .A(n862), .Y(n863) );
  INVX1 U1093 ( .A(n4526), .Y(n864) );
  INVX1 U1094 ( .A(n437), .Y(n865) );
  AND2X1 U1095 ( .A(n1221), .B(net79414), .Y(net92757) );
  INVX1 U1096 ( .A(net92757), .Y(n867) );
  INVX1 U1097 ( .A(n867), .Y(net66441) );
  INVX2 U1098 ( .A(n3642), .Y(n3782) );
  INVX1 U1099 ( .A(net66385), .Y(n1855) );
  AND2X2 U1100 ( .A(net66499), .B(n3643), .Y(n4532) );
  AND2X2 U1101 ( .A(net66975), .B(net66974), .Y(n4547) );
  OR2X1 U1102 ( .A(n1320), .B(n1321), .Y(n1317) );
  INVX1 U1103 ( .A(n1317), .Y(n868) );
  OR2X1 U1104 ( .A(n1318), .B(n1319), .Y(n1322) );
  INVX1 U1105 ( .A(n1322), .Y(n869) );
  OR2X1 U1106 ( .A(n1329), .B(n1330), .Y(n1326) );
  INVX1 U1107 ( .A(n1326), .Y(n870) );
  OR2X1 U1108 ( .A(n1327), .B(n1328), .Y(n1331) );
  INVX1 U1109 ( .A(n1331), .Y(n871) );
  OR2X1 U1110 ( .A(n1338), .B(n1339), .Y(n1335) );
  INVX1 U1111 ( .A(n1335), .Y(n872) );
  OR2X1 U1112 ( .A(n1336), .B(n1337), .Y(n1340) );
  INVX1 U1113 ( .A(n1340), .Y(n874) );
  OR2X1 U1114 ( .A(n1412), .B(n1413), .Y(n1409) );
  INVX1 U1115 ( .A(n1409), .Y(n875) );
  OR2X1 U1116 ( .A(n1410), .B(n1411), .Y(n1414) );
  INVX1 U1117 ( .A(n1414), .Y(n876) );
  OR2X1 U1118 ( .A(n1595), .B(n1596), .Y(n1592) );
  INVX1 U1119 ( .A(n1592), .Y(n877) );
  OR2X1 U1120 ( .A(n1593), .B(n1594), .Y(n1597) );
  INVX1 U1121 ( .A(n1597), .Y(n878) );
  AND2X2 U1122 ( .A(CMD_data_out[32]), .B(n1718), .Y(n3659) );
  INVX1 U1123 ( .A(n3659), .Y(n879) );
  AND2X2 U1124 ( .A(n4546), .B(net66974), .Y(n1719) );
  INVX1 U1125 ( .A(n1719), .Y(n880) );
  OR2X1 U1126 ( .A(n1796), .B(n1797), .Y(n1793) );
  INVX1 U1127 ( .A(n1793), .Y(n881) );
  OR2X1 U1128 ( .A(n1794), .B(n1795), .Y(n1798) );
  INVX1 U1129 ( .A(n1798), .Y(n882) );
  AND2X1 U1130 ( .A(add_576_carry_10_), .B(CMD_data_out[7]), .Y(n3516) );
  INVX1 U1131 ( .A(n3516), .Y(n883) );
  OR2X1 U1132 ( .A(i[20]), .B(i[19]), .Y(n3526) );
  INVX1 U1133 ( .A(n3526), .Y(n884) );
  OR2X1 U1134 ( .A(i[22]), .B(i[21]), .Y(n3525) );
  INVX1 U1135 ( .A(n3525), .Y(n885) );
  OR2X1 U1136 ( .A(i[23]), .B(i[22]), .Y(n3553) );
  INVX1 U1137 ( .A(n3553), .Y(n886) );
  OR2X1 U1138 ( .A(i[25]), .B(i[24]), .Y(n3552) );
  INVX1 U1139 ( .A(n3552), .Y(n887) );
  AND2X1 U1140 ( .A(n3660), .B(n3661), .Y(n3673) );
  INVX1 U1141 ( .A(n3673), .Y(n888) );
  AND2X1 U1142 ( .A(n3756), .B(n1545), .Y(n3753) );
  INVX1 U1143 ( .A(n3753), .Y(n889) );
  AND2X1 U1144 ( .A(n4545), .B(n1717), .Y(n4504) );
  INVX1 U1145 ( .A(n4504), .Y(n890) );
  OR2X2 U1146 ( .A(net66975), .B(net66974), .Y(n4612) );
  INVX1 U1147 ( .A(n4612), .Y(n891) );
  INVX4 U1148 ( .A(CMD_data_out[31]), .Y(net66974) );
  INVX1 U1149 ( .A(n894), .Y(n892) );
  INVX1 U1150 ( .A(n892), .Y(n893) );
  OR2X1 U1151 ( .A(net79414), .B(n230), .Y(net92732) );
  INVX1 U1152 ( .A(net92732), .Y(n894) );
  INVX1 U1153 ( .A(n897), .Y(n895) );
  INVX1 U1154 ( .A(n895), .Y(n896) );
  OR2X1 U1155 ( .A(j[14]), .B(j[15]), .Y(n1863) );
  INVX1 U1156 ( .A(n1863), .Y(n897) );
  INVX1 U1157 ( .A(n900), .Y(n898) );
  INVX1 U1158 ( .A(n898), .Y(n899) );
  OR2X1 U1159 ( .A(j[12]), .B(j[13]), .Y(n1865) );
  INVX1 U1160 ( .A(n1865), .Y(n900) );
  INVX1 U1161 ( .A(n903), .Y(n901) );
  INVX1 U1162 ( .A(n901), .Y(n902) );
  OR2X1 U1163 ( .A(n1233), .B(n1236), .Y(net89555) );
  INVX1 U1164 ( .A(net89555), .Y(n903) );
  INVX1 U1165 ( .A(n906), .Y(n904) );
  INVX1 U1166 ( .A(n904), .Y(n905) );
  OR2X1 U1167 ( .A(i[27]), .B(i[26]), .Y(n3555) );
  INVX1 U1168 ( .A(n3555), .Y(n906) );
  INVX1 U1169 ( .A(n910), .Y(n908) );
  INVX1 U1170 ( .A(n908), .Y(n909) );
  AND2X1 U1171 ( .A(n1665), .B(n1031), .Y(n2546) );
  INVX1 U1172 ( .A(n2546), .Y(n910) );
  INVX1 U1173 ( .A(n913), .Y(n911) );
  INVX1 U1174 ( .A(n911), .Y(n912) );
  OR2X1 U1175 ( .A(j[11]), .B(j[10]), .Y(n1862) );
  INVX1 U1176 ( .A(n1862), .Y(n913) );
  INVX1 U1177 ( .A(n916), .Y(n914) );
  INVX1 U1178 ( .A(n914), .Y(n915) );
  AND2X1 U1179 ( .A(n1885), .B(n3914), .Y(n4458) );
  INVX1 U1180 ( .A(n4458), .Y(n916) );
  INVX1 U1181 ( .A(n919), .Y(n917) );
  INVX1 U1182 ( .A(n917), .Y(n918) );
  AND2X1 U1183 ( .A(n1886), .B(n3914), .Y(n4464) );
  INVX1 U1184 ( .A(n4464), .Y(n919) );
  INVX1 U1185 ( .A(n922), .Y(n920) );
  INVX1 U1186 ( .A(n920), .Y(n921) );
  AND2X1 U1187 ( .A(n1887), .B(n3914), .Y(n4470) );
  INVX1 U1188 ( .A(n4470), .Y(n922) );
  INVX1 U1189 ( .A(n925), .Y(n923) );
  INVX1 U1190 ( .A(n923), .Y(n924) );
  AND2X1 U1191 ( .A(n1888), .B(n3914), .Y(n4475) );
  INVX1 U1192 ( .A(n4475), .Y(n925) );
  INVX1 U1193 ( .A(n928), .Y(n926) );
  INVX1 U1194 ( .A(n926), .Y(n927) );
  AND2X1 U1195 ( .A(n1889), .B(n3914), .Y(n4480) );
  INVX1 U1196 ( .A(n4480), .Y(n928) );
  INVX1 U1197 ( .A(n931), .Y(n929) );
  INVX1 U1198 ( .A(n929), .Y(n930) );
  AND2X1 U1199 ( .A(n1890), .B(n3914), .Y(n4485) );
  INVX1 U1200 ( .A(n4485), .Y(n931) );
  INVX1 U1201 ( .A(n934), .Y(n932) );
  INVX1 U1202 ( .A(n932), .Y(n933) );
  AND2X1 U1203 ( .A(n1891), .B(n3914), .Y(n4490) );
  INVX1 U1204 ( .A(n4490), .Y(n934) );
  INVX1 U1205 ( .A(n937), .Y(n935) );
  INVX1 U1206 ( .A(n935), .Y(n936) );
  AND2X1 U1207 ( .A(n1892), .B(n3914), .Y(n4495) );
  INVX1 U1208 ( .A(n4495), .Y(n937) );
  INVX1 U1209 ( .A(n940), .Y(n938) );
  INVX1 U1210 ( .A(n938), .Y(n939) );
  AND2X1 U1211 ( .A(n1893), .B(n3914), .Y(n4500) );
  INVX1 U1212 ( .A(n4500), .Y(n940) );
  AND2X2 U1213 ( .A(n635), .B(n3641), .Y(n3748) );
  INVX1 U1214 ( .A(n3748), .Y(n941) );
  INVX4 U1215 ( .A(n3749), .Y(n3641) );
  AND2X2 U1216 ( .A(n2081), .B(n3925), .Y(n3924) );
  INVX1 U1217 ( .A(n3924), .Y(n943) );
  AND2X2 U1218 ( .A(n2082), .B(n3925), .Y(n3926) );
  INVX1 U1219 ( .A(n3926), .Y(n944) );
  AND2X2 U1220 ( .A(n2083), .B(n3925), .Y(n3927) );
  INVX1 U1221 ( .A(n3927), .Y(n945) );
  AND2X2 U1222 ( .A(n2084), .B(n3925), .Y(net66328) );
  INVX1 U1223 ( .A(net66328), .Y(n946) );
  AND2X2 U1224 ( .A(n2085), .B(n3925), .Y(net66330) );
  INVX1 U1225 ( .A(net66330), .Y(n947) );
  AND2X2 U1226 ( .A(n2086), .B(n3925), .Y(n3929) );
  INVX1 U1227 ( .A(n3929), .Y(n948) );
  AND2X2 U1228 ( .A(n2087), .B(n3925), .Y(n3931) );
  INVX1 U1229 ( .A(n3931), .Y(n949) );
  AND2X2 U1230 ( .A(n2088), .B(n3925), .Y(net66336) );
  INVX1 U1231 ( .A(net66336), .Y(n950) );
  AND2X2 U1232 ( .A(n2089), .B(n3925), .Y(net66338) );
  INVX1 U1233 ( .A(net66338), .Y(n951) );
  AND2X2 U1234 ( .A(n2090), .B(n3925), .Y(n3932) );
  INVX1 U1235 ( .A(n3932), .Y(n952) );
  AND2X2 U1236 ( .A(n2091), .B(n3925), .Y(net66342) );
  INVX1 U1237 ( .A(net66342), .Y(n953) );
  AND2X2 U1238 ( .A(n2092), .B(n3925), .Y(net66344) );
  INVX1 U1239 ( .A(net66344), .Y(n954) );
  AND2X2 U1240 ( .A(n2093), .B(n3925), .Y(net66346) );
  INVX1 U1241 ( .A(net66346), .Y(n955) );
  AND2X2 U1242 ( .A(n2094), .B(n3925), .Y(net66348) );
  INVX1 U1243 ( .A(net66348), .Y(n956) );
  AND2X2 U1244 ( .A(n2095), .B(n3925), .Y(net66350) );
  INVX1 U1245 ( .A(net66350), .Y(n957) );
  AND2X2 U1246 ( .A(n2096), .B(n3925), .Y(net66352) );
  INVX1 U1247 ( .A(net66352), .Y(n958) );
  AND2X2 U1248 ( .A(n2097), .B(n3925), .Y(n3934) );
  INVX1 U1249 ( .A(n3934), .Y(n959) );
  AND2X2 U1250 ( .A(n2098), .B(n3925), .Y(n3936) );
  INVX1 U1251 ( .A(n3936), .Y(n960) );
  AND2X2 U1252 ( .A(n2099), .B(n3925), .Y(n3938) );
  INVX1 U1253 ( .A(n3938), .Y(n961) );
  AND2X2 U1254 ( .A(n2100), .B(n3925), .Y(n3940) );
  INVX1 U1255 ( .A(n3940), .Y(n962) );
  AND2X2 U1256 ( .A(n2101), .B(n3925), .Y(n3942) );
  INVX1 U1257 ( .A(n3942), .Y(n963) );
  AND2X2 U1258 ( .A(n2102), .B(n3925), .Y(n3944) );
  INVX1 U1259 ( .A(n3944), .Y(n964) );
  AND2X2 U1260 ( .A(n2103), .B(n3925), .Y(n3946) );
  INVX1 U1261 ( .A(n3946), .Y(n965) );
  AND2X2 U1262 ( .A(n2104), .B(n3925), .Y(net66368) );
  INVX1 U1263 ( .A(net66368), .Y(n966) );
  AND2X2 U1264 ( .A(n2105), .B(n3925), .Y(net66370) );
  INVX1 U1265 ( .A(net66370), .Y(n967) );
  AND2X2 U1266 ( .A(n2106), .B(n3925), .Y(net66372) );
  INVX1 U1267 ( .A(net66372), .Y(n968) );
  AND2X2 U1268 ( .A(n2107), .B(n3925), .Y(net66374) );
  INVX1 U1269 ( .A(net66374), .Y(n969) );
  AND2X2 U1270 ( .A(n2108), .B(n3925), .Y(net66376) );
  INVX1 U1271 ( .A(net66376), .Y(n970) );
  AND2X2 U1272 ( .A(n2109), .B(n3925), .Y(net66378) );
  INVX1 U1273 ( .A(net66378), .Y(n971) );
  AND2X1 U1274 ( .A(net79482), .B(net66140), .Y(n4041) );
  INVX1 U1275 ( .A(n4041), .Y(n972) );
  INVX1 U1276 ( .A(n975), .Y(n973) );
  INVX1 U1277 ( .A(n973), .Y(n974) );
  AND2X1 U1278 ( .A(DQ_out[15]), .B(n4391), .Y(n4390) );
  INVX1 U1279 ( .A(n4390), .Y(n975) );
  INVX1 U1280 ( .A(n987), .Y(n985) );
  INVX1 U1281 ( .A(n985), .Y(n986) );
  AND2X1 U1282 ( .A(DQ_out[14]), .B(n4391), .Y(n4395) );
  INVX1 U1283 ( .A(n4395), .Y(n987) );
  INVX1 U1284 ( .A(n990), .Y(n988) );
  INVX1 U1285 ( .A(n988), .Y(n989) );
  AND2X1 U1286 ( .A(DQ_out[13]), .B(n4391), .Y(n4397) );
  INVX1 U1287 ( .A(n4397), .Y(n990) );
  INVX1 U1288 ( .A(n993), .Y(n991) );
  INVX1 U1289 ( .A(n991), .Y(n992) );
  AND2X1 U1290 ( .A(DQ_out[12]), .B(n4391), .Y(n4399) );
  INVX1 U1291 ( .A(n4399), .Y(n993) );
  INVX1 U1292 ( .A(n996), .Y(n994) );
  INVX1 U1293 ( .A(n994), .Y(n995) );
  AND2X1 U1294 ( .A(DQ_out[11]), .B(n4391), .Y(n4401) );
  INVX1 U1295 ( .A(n4401), .Y(n996) );
  INVX1 U1296 ( .A(n999), .Y(n997) );
  INVX1 U1297 ( .A(n997), .Y(n998) );
  AND2X1 U1298 ( .A(DQ_out[10]), .B(n4391), .Y(n4403) );
  INVX1 U1299 ( .A(n4403), .Y(n999) );
  INVX1 U1300 ( .A(n1002), .Y(n1000) );
  INVX1 U1301 ( .A(n1000), .Y(n1001) );
  AND2X1 U1302 ( .A(DQ_out[9]), .B(n4391), .Y(n4405) );
  INVX1 U1303 ( .A(n4405), .Y(n1002) );
  INVX1 U1304 ( .A(n1005), .Y(n1003) );
  INVX1 U1305 ( .A(n1003), .Y(n1004) );
  AND2X1 U1306 ( .A(DQ_out[8]), .B(n4391), .Y(n4407) );
  INVX1 U1307 ( .A(n4407), .Y(n1005) );
  INVX1 U1308 ( .A(n1008), .Y(n1006) );
  INVX1 U1309 ( .A(n1006), .Y(n1007) );
  AND2X1 U1310 ( .A(DQ_out[7]), .B(n4391), .Y(n4409) );
  INVX1 U1311 ( .A(n4409), .Y(n1008) );
  INVX1 U1312 ( .A(n1011), .Y(n1009) );
  INVX1 U1313 ( .A(n1009), .Y(n1010) );
  AND2X1 U1314 ( .A(DQ_out[6]), .B(n4391), .Y(n4411) );
  INVX1 U1315 ( .A(n4411), .Y(n1011) );
  INVX1 U1316 ( .A(n1014), .Y(n1012) );
  INVX1 U1317 ( .A(n1012), .Y(n1013) );
  AND2X1 U1318 ( .A(DQ_out[5]), .B(n4391), .Y(n4413) );
  INVX1 U1319 ( .A(n4413), .Y(n1014) );
  INVX1 U1320 ( .A(n1017), .Y(n1015) );
  INVX1 U1321 ( .A(n1015), .Y(n1016) );
  AND2X1 U1322 ( .A(DQ_out[4]), .B(n4391), .Y(n4415) );
  INVX1 U1323 ( .A(n4415), .Y(n1017) );
  INVX1 U1324 ( .A(n1020), .Y(n1018) );
  INVX1 U1325 ( .A(n1018), .Y(n1019) );
  AND2X1 U1326 ( .A(DQ_out[3]), .B(n4391), .Y(n4417) );
  INVX1 U1327 ( .A(n4417), .Y(n1020) );
  INVX1 U1328 ( .A(n1023), .Y(n1021) );
  INVX1 U1329 ( .A(n1021), .Y(n1022) );
  AND2X1 U1330 ( .A(DQ_out[2]), .B(n4391), .Y(n4419) );
  INVX1 U1331 ( .A(n4419), .Y(n1023) );
  INVX1 U1332 ( .A(n1026), .Y(n1024) );
  INVX1 U1333 ( .A(n1024), .Y(n1025) );
  AND2X1 U1334 ( .A(DQ_out[1]), .B(n4391), .Y(n4421) );
  INVX1 U1335 ( .A(n4421), .Y(n1026) );
  INVX1 U1336 ( .A(n1029), .Y(n1027) );
  INVX1 U1337 ( .A(n1027), .Y(n1028) );
  AND2X1 U1338 ( .A(DQ_out[0]), .B(n4391), .Y(n4423) );
  INVX1 U1339 ( .A(n4423), .Y(n1029) );
  INVX1 U1340 ( .A(n1032), .Y(n1030) );
  INVX1 U1341 ( .A(n1030), .Y(n1031) );
  AND2X1 U1342 ( .A(ts_con), .B(n4581), .Y(n4580) );
  INVX1 U1343 ( .A(n4580), .Y(n1032) );
  OR2X1 U1344 ( .A(n1041), .B(n1042), .Y(n1039) );
  INVX1 U1345 ( .A(n1039), .Y(n1033) );
  INVX1 U1346 ( .A(n1036), .Y(n1034) );
  INVX1 U1347 ( .A(n1034), .Y(n1035) );
  OR2X1 U1348 ( .A(n1043), .B(n1044), .Y(n1040) );
  INVX1 U1349 ( .A(n1040), .Y(n1036) );
  INVX1 U1350 ( .A(n448), .Y(n1037) );
  INVX1 U1351 ( .A(n1037), .Y(n1038) );
  INVX1 U1352 ( .A(n575), .Y(n1041) );
  INVX8 U1353 ( .A(n1782), .Y(n1042) );
  INVX1 U1354 ( .A(n1785), .Y(n1043) );
  INVX1 U1355 ( .A(n233), .Y(n1044) );
  INVX1 U1356 ( .A(n3511), .Y(n233) );
  INVX1 U1357 ( .A(n1047), .Y(n1045) );
  INVX1 U1358 ( .A(n1045), .Y(n1046) );
  OR2X1 U1359 ( .A(n1055), .B(n1056), .Y(n1053) );
  INVX1 U1360 ( .A(n1053), .Y(n1047) );
  INVX1 U1361 ( .A(n1050), .Y(n1048) );
  INVX1 U1362 ( .A(n1048), .Y(n1049) );
  OR2X1 U1363 ( .A(n1057), .B(n1058), .Y(n1054) );
  INVX1 U1364 ( .A(n1054), .Y(n1050) );
  INVX1 U1365 ( .A(n449), .Y(n1051) );
  INVX1 U1366 ( .A(n1051), .Y(n1052) );
  INVX1 U1367 ( .A(n567), .Y(n1055) );
  INVX1 U1368 ( .A(n1782), .Y(n1056) );
  INVX1 U1369 ( .A(n1785), .Y(n1057) );
  INVX1 U1370 ( .A(n234), .Y(n1058) );
  INVX1 U1371 ( .A(n3510), .Y(n234) );
  OR2X1 U1372 ( .A(n1065), .B(n1066), .Y(n1063) );
  INVX1 U1373 ( .A(n1063), .Y(n1059) );
  INVX1 U1374 ( .A(n1062), .Y(n1060) );
  INVX1 U1375 ( .A(n1060), .Y(n1061) );
  OR2X1 U1376 ( .A(n1067), .B(n1068), .Y(n1064) );
  INVX1 U1377 ( .A(n1064), .Y(n1062) );
  INVX1 U1378 ( .A(n579), .Y(n1065) );
  INVX2 U1379 ( .A(n1782), .Y(n1066) );
  INVX1 U1380 ( .A(n1785), .Y(n1067) );
  INVX1 U1381 ( .A(n235), .Y(n1068) );
  INVX1 U1382 ( .A(n3509), .Y(n235) );
  INVX1 U1383 ( .A(n1071), .Y(n1069) );
  INVX1 U1384 ( .A(n1069), .Y(n1070) );
  OR2X1 U1385 ( .A(n1079), .B(n1080), .Y(n1077) );
  INVX1 U1386 ( .A(n1077), .Y(n1071) );
  INVX1 U1387 ( .A(n1074), .Y(n1072) );
  INVX1 U1388 ( .A(n1072), .Y(n1073) );
  OR2X1 U1389 ( .A(n1081), .B(n1082), .Y(n1078) );
  INVX1 U1390 ( .A(n1078), .Y(n1074) );
  INVX1 U1391 ( .A(n451), .Y(n1075) );
  INVX1 U1392 ( .A(n1075), .Y(n1076) );
  INVX1 U1393 ( .A(n572), .Y(n1079) );
  INVX1 U1394 ( .A(n1782), .Y(n1080) );
  INVX1 U1395 ( .A(n1785), .Y(n1081) );
  INVX1 U1396 ( .A(n236), .Y(n1082) );
  INVX1 U1397 ( .A(n3508), .Y(n236) );
  INVX1 U1398 ( .A(n1085), .Y(n1083) );
  INVX1 U1399 ( .A(n1083), .Y(n1084) );
  OR2X1 U1400 ( .A(n1093), .B(n1094), .Y(n1091) );
  INVX1 U1401 ( .A(n1091), .Y(n1085) );
  INVX1 U1402 ( .A(n1088), .Y(n1086) );
  INVX1 U1403 ( .A(n1086), .Y(n1087) );
  OR2X1 U1404 ( .A(n1095), .B(n1096), .Y(n1092) );
  INVX1 U1405 ( .A(n1092), .Y(n1088) );
  INVX1 U1406 ( .A(n452), .Y(n1089) );
  INVX1 U1407 ( .A(n1089), .Y(n1090) );
  INVX1 U1408 ( .A(n571), .Y(n1093) );
  INVX1 U1409 ( .A(n1782), .Y(n1094) );
  INVX1 U1410 ( .A(n1785), .Y(n1095) );
  INVX1 U1411 ( .A(n237), .Y(n1096) );
  INVX1 U1412 ( .A(n3507), .Y(n237) );
  INVX1 U1413 ( .A(n1099), .Y(n1097) );
  INVX1 U1414 ( .A(n1097), .Y(n1098) );
  OR2X1 U1415 ( .A(n1107), .B(n1108), .Y(n1105) );
  INVX1 U1416 ( .A(n1105), .Y(n1099) );
  INVX1 U1417 ( .A(n1102), .Y(n1100) );
  INVX1 U1418 ( .A(n1100), .Y(n1101) );
  OR2X1 U1419 ( .A(n1109), .B(n1110), .Y(n1106) );
  INVX1 U1420 ( .A(n1106), .Y(n1102) );
  INVX1 U1421 ( .A(n453), .Y(n1103) );
  INVX1 U1422 ( .A(n1103), .Y(n1104) );
  INVX1 U1423 ( .A(n564), .Y(n1107) );
  INVX1 U1424 ( .A(n1782), .Y(n1108) );
  INVX1 U1425 ( .A(n1785), .Y(n1109) );
  INVX1 U1426 ( .A(n238), .Y(n1110) );
  INVX1 U1427 ( .A(n3506), .Y(n238) );
  INVX1 U1428 ( .A(n1113), .Y(n1111) );
  INVX1 U1429 ( .A(n1111), .Y(n1112) );
  OR2X1 U1430 ( .A(n1121), .B(n1122), .Y(n1119) );
  INVX1 U1431 ( .A(n1119), .Y(n1113) );
  INVX1 U1432 ( .A(n1116), .Y(n1114) );
  INVX1 U1433 ( .A(n1114), .Y(n1115) );
  OR2X1 U1434 ( .A(n1123), .B(n1124), .Y(n1120) );
  INVX1 U1435 ( .A(n1120), .Y(n1116) );
  INVX1 U1436 ( .A(n454), .Y(n1117) );
  INVX1 U1437 ( .A(n1117), .Y(n1118) );
  INVX1 U1438 ( .A(n565), .Y(n1121) );
  INVX1 U1439 ( .A(n1782), .Y(n1122) );
  INVX1 U1440 ( .A(n1785), .Y(n1123) );
  INVX1 U1441 ( .A(n239), .Y(n1124) );
  INVX1 U1442 ( .A(n3505), .Y(n239) );
  INVX1 U1443 ( .A(n1127), .Y(n1125) );
  INVX1 U1444 ( .A(n1125), .Y(n1126) );
  OR2X1 U1445 ( .A(n1135), .B(n1136), .Y(n1133) );
  INVX1 U1446 ( .A(n1133), .Y(n1127) );
  INVX1 U1447 ( .A(n1130), .Y(n1128) );
  INVX1 U1448 ( .A(n1128), .Y(n1129) );
  OR2X1 U1449 ( .A(n1137), .B(n1138), .Y(n1134) );
  INVX1 U1450 ( .A(n1134), .Y(n1130) );
  INVX1 U1451 ( .A(n455), .Y(n1131) );
  INVX1 U1452 ( .A(n1131), .Y(n1132) );
  INVX1 U1453 ( .A(n566), .Y(n1135) );
  INVX1 U1454 ( .A(n1782), .Y(n1136) );
  INVX1 U1455 ( .A(n1785), .Y(n1137) );
  INVX1 U1456 ( .A(n240), .Y(n1138) );
  INVX1 U1457 ( .A(n3504), .Y(n240) );
  OR2X1 U1458 ( .A(n1145), .B(n1146), .Y(n1143) );
  INVX1 U1459 ( .A(n1143), .Y(n1139) );
  INVX1 U1460 ( .A(n1142), .Y(n1140) );
  INVX1 U1461 ( .A(n1140), .Y(n1141) );
  OR2X1 U1462 ( .A(n1147), .B(n1148), .Y(n1144) );
  INVX1 U1463 ( .A(n1144), .Y(n1142) );
  INVX1 U1464 ( .A(n578), .Y(n1145) );
  INVX8 U1465 ( .A(n1782), .Y(n1146) );
  INVX1 U1466 ( .A(n1785), .Y(n1147) );
  INVX1 U1467 ( .A(n241), .Y(n1148) );
  INVX1 U1468 ( .A(n3503), .Y(n241) );
  INVX1 U1469 ( .A(n1151), .Y(n1149) );
  INVX1 U1470 ( .A(n1149), .Y(n1150) );
  OR2X1 U1471 ( .A(n1159), .B(n1160), .Y(n1157) );
  INVX1 U1472 ( .A(n1157), .Y(n1151) );
  INVX1 U1473 ( .A(n1154), .Y(n1152) );
  INVX1 U1474 ( .A(n1152), .Y(n1153) );
  OR2X1 U1475 ( .A(n1161), .B(n1162), .Y(n1158) );
  INVX1 U1476 ( .A(n1158), .Y(n1154) );
  INVX1 U1477 ( .A(n457), .Y(n1155) );
  INVX1 U1478 ( .A(n1155), .Y(n1156) );
  INVX1 U1479 ( .A(n570), .Y(n1159) );
  INVX1 U1480 ( .A(n1782), .Y(n1160) );
  INVX1 U1481 ( .A(n1785), .Y(n1161) );
  INVX1 U1482 ( .A(n242), .Y(n1162) );
  INVX1 U1483 ( .A(n3502), .Y(n242) );
  INVX1 U1484 ( .A(n1165), .Y(n1163) );
  INVX1 U1485 ( .A(n1163), .Y(n1164) );
  OR2X1 U1486 ( .A(n1173), .B(n1174), .Y(n1171) );
  INVX1 U1487 ( .A(n1171), .Y(n1165) );
  INVX1 U1488 ( .A(n1168), .Y(n1166) );
  INVX1 U1489 ( .A(n1166), .Y(n1167) );
  OR2X1 U1490 ( .A(n1175), .B(n1176), .Y(n1172) );
  INVX1 U1491 ( .A(n1172), .Y(n1168) );
  INVX1 U1492 ( .A(n458), .Y(n1169) );
  INVX1 U1493 ( .A(n1169), .Y(n1170) );
  INVX1 U1494 ( .A(n569), .Y(n1173) );
  INVX1 U1495 ( .A(n1782), .Y(n1174) );
  INVX1 U1496 ( .A(n1785), .Y(n1175) );
  INVX1 U1497 ( .A(n243), .Y(n1176) );
  INVX1 U1498 ( .A(n3501), .Y(n243) );
  OR2X1 U1499 ( .A(n1183), .B(n1184), .Y(n1181) );
  INVX1 U1500 ( .A(n1181), .Y(n1177) );
  INVX1 U1501 ( .A(n1180), .Y(n1178) );
  INVX1 U1502 ( .A(n1178), .Y(n1179) );
  OR2X1 U1503 ( .A(n1185), .B(n1186), .Y(n1182) );
  INVX1 U1504 ( .A(n1182), .Y(n1180) );
  INVX1 U1505 ( .A(n576), .Y(n1183) );
  INVX2 U1506 ( .A(n1782), .Y(n1184) );
  INVX1 U1507 ( .A(n1785), .Y(n1185) );
  INVX1 U1508 ( .A(n244), .Y(n1186) );
  INVX1 U1509 ( .A(n3500), .Y(n244) );
  INVX1 U1510 ( .A(n1189), .Y(n1187) );
  INVX1 U1511 ( .A(n1187), .Y(n1188) );
  OR2X1 U1512 ( .A(n1197), .B(n1198), .Y(n1195) );
  INVX1 U1513 ( .A(n1195), .Y(n1189) );
  INVX1 U1514 ( .A(n1192), .Y(n1190) );
  INVX1 U1515 ( .A(n1190), .Y(n1191) );
  OR2X1 U1516 ( .A(n1199), .B(n1200), .Y(n1196) );
  INVX1 U1517 ( .A(n1196), .Y(n1192) );
  INVX1 U1518 ( .A(n460), .Y(n1193) );
  INVX1 U1519 ( .A(n1193), .Y(n1194) );
  INVX1 U1520 ( .A(n568), .Y(n1197) );
  INVX1 U1521 ( .A(n1782), .Y(n1198) );
  INVX1 U1522 ( .A(n1785), .Y(n1199) );
  INVX1 U1523 ( .A(n245), .Y(n1200) );
  INVX1 U1524 ( .A(n3499), .Y(n245) );
  OR2X1 U1525 ( .A(n1207), .B(n1208), .Y(n1205) );
  INVX1 U1526 ( .A(n1205), .Y(n1201) );
  INVX1 U1527 ( .A(n1204), .Y(n1202) );
  INVX1 U1528 ( .A(n1202), .Y(n1203) );
  OR2X1 U1529 ( .A(n1209), .B(n1210), .Y(n1206) );
  INVX1 U1530 ( .A(n1206), .Y(n1204) );
  INVX1 U1531 ( .A(n577), .Y(n1207) );
  INVX2 U1532 ( .A(n1782), .Y(n1208) );
  INVX1 U1533 ( .A(n1785), .Y(n1209) );
  INVX1 U1534 ( .A(n247), .Y(n1210) );
  INVX1 U1535 ( .A(n3497), .Y(n247) );
  INVX1 U1536 ( .A(n1213), .Y(n1211) );
  INVX1 U1537 ( .A(n1211), .Y(n1212) );
  AND2X2 U1538 ( .A(BA[0]), .B(n1732), .Y(n4439) );
  INVX1 U1539 ( .A(n4439), .Y(n1213) );
  INVX1 U1540 ( .A(n1216), .Y(n1214) );
  INVX1 U1541 ( .A(n1214), .Y(n1215) );
  AND2X2 U1542 ( .A(BA[1]), .B(n1732), .Y(n4444) );
  INVX1 U1543 ( .A(n4444), .Y(n1216) );
  INVX1 U1544 ( .A(n1219), .Y(n1217) );
  INVX1 U1545 ( .A(n1217), .Y(n1218) );
  AND2X1 U1546 ( .A(BA[2]), .B(n1732), .Y(n4446) );
  INVX1 U1547 ( .A(n4446), .Y(n1219) );
  AND2X2 U1548 ( .A(n1695), .B(n4440), .Y(n4442) );
  AND2X2 U1549 ( .A(n1599), .B(n4440), .Y(n4441) );
  INVX1 U1550 ( .A(n1222), .Y(n1220) );
  INVX1 U1551 ( .A(n1220), .Y(n1221) );
  OR2X1 U1552 ( .A(net79436), .B(net66325), .Y(n1806) );
  INVX1 U1553 ( .A(n1806), .Y(n1222) );
  INVX1 U1554 ( .A(n1225), .Y(n1223) );
  INVX1 U1555 ( .A(n1223), .Y(n1224) );
  OR2X1 U1556 ( .A(n1811), .B(n1572), .Y(n1812) );
  INVX1 U1557 ( .A(n1812), .Y(n1225) );
  INVX1 U1558 ( .A(n1228), .Y(n1226) );
  INVX1 U1559 ( .A(n1226), .Y(n1227) );
  OR2X1 U1560 ( .A(net92738), .B(n1569), .Y(n1844) );
  INVX1 U1561 ( .A(n1844), .Y(n1228) );
  INVX1 U1562 ( .A(n1231), .Y(n1229) );
  INVX1 U1563 ( .A(n1229), .Y(n1230) );
  AND2X1 U1564 ( .A(net89562), .B(n1809), .Y(net89561) );
  INVX1 U1565 ( .A(net89561), .Y(n1231) );
  INVX1 U1566 ( .A(n1234), .Y(n1232) );
  INVX1 U1567 ( .A(n1232), .Y(n1233) );
  AND2X2 U1568 ( .A(n896), .B(n912), .Y(n1864) );
  INVX1 U1569 ( .A(n1864), .Y(n1234) );
  INVX1 U1570 ( .A(n1237), .Y(n1235) );
  INVX1 U1571 ( .A(n1235), .Y(n1236) );
  AND2X2 U1572 ( .A(n899), .B(net66953), .Y(n1866) );
  INVX1 U1573 ( .A(n1866), .Y(n1237) );
  INVX1 U1574 ( .A(n1240), .Y(n1238) );
  INVX1 U1575 ( .A(n1238), .Y(n1239) );
  AND2X2 U1576 ( .A(n653), .B(n3708), .Y(n3706) );
  INVX1 U1577 ( .A(n3706), .Y(n1240) );
  INVX1 U1578 ( .A(n1243), .Y(n1241) );
  INVX1 U1579 ( .A(n1241), .Y(n1242) );
  OR2X1 U1580 ( .A(i[16]), .B(i[15]), .Y(n3548) );
  INVX1 U1581 ( .A(n3548), .Y(n1243) );
  INVX1 U1582 ( .A(n1246), .Y(n1244) );
  INVX1 U1583 ( .A(n1244), .Y(n1245) );
  OR2X2 U1584 ( .A(n792), .B(n811), .Y(n4549) );
  INVX1 U1585 ( .A(n4549), .Y(n1246) );
  INVX1 U1586 ( .A(n1249), .Y(n1247) );
  INVX1 U1587 ( .A(n1247), .Y(n1248) );
  AND2X1 U1588 ( .A(clkcount[3]), .B(clkcount[2]), .Y(n4564) );
  INVX1 U1589 ( .A(n4564), .Y(n1249) );
  INVX1 U1590 ( .A(n465), .Y(n1808) );
  AND2X1 U1591 ( .A(add_576_carry_9_), .B(CMD_data_out[6]), .Y(n3515) );
  INVX1 U1592 ( .A(n3515), .Y(n1250) );
  INVX1 U1593 ( .A(n1250), .Y(add_576_carry_10_) );
  AND2X1 U1594 ( .A(add_576_carry_11_), .B(CMD_data_out[8]), .Y(n3517) );
  INVX1 U1595 ( .A(n3517), .Y(n1251) );
  INVX1 U1596 ( .A(n883), .Y(add_576_carry_11_) );
  INVX1 U1597 ( .A(n1254), .Y(n1252) );
  INVX1 U1598 ( .A(n1252), .Y(n1253) );
  AND2X1 U1599 ( .A(n1875), .B(n1876), .Y(r576_net62619) );
  INVX1 U1600 ( .A(r576_net62619), .Y(n1254) );
  INVX1 U1601 ( .A(n1257), .Y(n1255) );
  INVX1 U1602 ( .A(n1255), .Y(n1256) );
  AND2X1 U1603 ( .A(r576_net62635), .B(r576_net62636), .Y(r576_net62630) );
  INVX1 U1604 ( .A(r576_net62630), .Y(n1257) );
  INVX1 U1605 ( .A(n1260), .Y(n1258) );
  INVX1 U1606 ( .A(n1258), .Y(n1259) );
  AND2X1 U1607 ( .A(n3523), .B(n3522), .Y(n3528) );
  INVX1 U1608 ( .A(n3528), .Y(n1260) );
  INVX1 U1609 ( .A(n1263), .Y(n1261) );
  INVX1 U1610 ( .A(n1261), .Y(n1262) );
  AND2X1 U1611 ( .A(n3532), .B(n3531), .Y(n3538) );
  INVX1 U1612 ( .A(n3538), .Y(n1263) );
  INVX1 U1613 ( .A(n1266), .Y(n1264) );
  INVX1 U1614 ( .A(n1264), .Y(n1265) );
  OR2X1 U1615 ( .A(n3579), .B(net66063), .Y(n3885) );
  INVX1 U1616 ( .A(n3885), .Y(n1266) );
  INVX1 U1617 ( .A(n1269), .Y(n1267) );
  INVX1 U1618 ( .A(n1267), .Y(n1268) );
  AND2X2 U1619 ( .A(n613), .B(n915), .Y(n4456) );
  INVX1 U1620 ( .A(n4456), .Y(n1269) );
  INVX1 U1621 ( .A(n1272), .Y(n1270) );
  INVX1 U1622 ( .A(n1270), .Y(n1271) );
  AND2X2 U1623 ( .A(n615), .B(n918), .Y(n4462) );
  INVX1 U1624 ( .A(n4462), .Y(n1272) );
  INVX1 U1625 ( .A(n1275), .Y(n1273) );
  INVX1 U1626 ( .A(n1273), .Y(n1274) );
  AND2X2 U1627 ( .A(n617), .B(n921), .Y(n4468) );
  INVX1 U1628 ( .A(n4468), .Y(n1275) );
  INVX1 U1629 ( .A(n1278), .Y(n1276) );
  INVX1 U1630 ( .A(n1276), .Y(n1277) );
  AND2X2 U1631 ( .A(n619), .B(n924), .Y(n4473) );
  INVX1 U1632 ( .A(n4473), .Y(n1278) );
  INVX1 U1633 ( .A(n1281), .Y(n1279) );
  INVX1 U1634 ( .A(n1279), .Y(n1280) );
  AND2X2 U1635 ( .A(n621), .B(n927), .Y(n4478) );
  INVX1 U1636 ( .A(n4478), .Y(n1281) );
  INVX1 U1637 ( .A(n1284), .Y(n1282) );
  INVX1 U1638 ( .A(n1282), .Y(n1283) );
  AND2X2 U1639 ( .A(n623), .B(n930), .Y(n4483) );
  INVX1 U1640 ( .A(n4483), .Y(n1284) );
  INVX1 U1641 ( .A(n1287), .Y(n1285) );
  INVX1 U1642 ( .A(n1285), .Y(n1286) );
  AND2X2 U1643 ( .A(n629), .B(n933), .Y(n4488) );
  INVX1 U1644 ( .A(n4488), .Y(n1287) );
  INVX1 U1645 ( .A(n1290), .Y(n1288) );
  INVX1 U1646 ( .A(n1288), .Y(n1289) );
  AND2X2 U1647 ( .A(n631), .B(n936), .Y(n4493) );
  INVX1 U1648 ( .A(n4493), .Y(n1290) );
  INVX1 U1649 ( .A(n1293), .Y(n1291) );
  INVX1 U1650 ( .A(n1291), .Y(n1292) );
  AND2X2 U1651 ( .A(n633), .B(n939), .Y(n4498) );
  INVX1 U1652 ( .A(n4498), .Y(n1293) );
  INVX1 U1653 ( .A(n1296), .Y(n1294) );
  INVX1 U1654 ( .A(n1294), .Y(n1295) );
  AND2X1 U1655 ( .A(clkcount[7]), .B(clkcount[6]), .Y(n4563) );
  INVX1 U1656 ( .A(n4563), .Y(n1296) );
  INVX1 U1657 ( .A(n1299), .Y(n1297) );
  INVX1 U1658 ( .A(n1297), .Y(n1298) );
  BUFX2 U1659 ( .A(n3896), .Y(n1299) );
  INVX1 U1660 ( .A(n1302), .Y(n1300) );
  INVX1 U1661 ( .A(n1300), .Y(n1301) );
  BUFX2 U1662 ( .A(n4517), .Y(n1302) );
  INVX1 U1663 ( .A(n1305), .Y(n1303) );
  INVX1 U1664 ( .A(n1303), .Y(n1304) );
  BUFX2 U1665 ( .A(n3761), .Y(n1305) );
  INVX1 U1666 ( .A(n1307), .Y(n1306) );
  BUFX2 U1667 ( .A(n4525), .Y(n1307) );
  INVX1 U1668 ( .A(n1310), .Y(n1308) );
  INVX1 U1669 ( .A(n1308), .Y(n1309) );
  OR2X1 U1670 ( .A(i[18]), .B(i[17]), .Y(n3547) );
  INVX1 U1671 ( .A(n3547), .Y(n1310) );
  INVX1 U1672 ( .A(n1313), .Y(n1311) );
  INVX1 U1673 ( .A(n1311), .Y(n1312) );
  OR2X2 U1674 ( .A(n789), .B(n808), .Y(n4550) );
  INVX1 U1675 ( .A(n4550), .Y(n1313) );
  INVX1 U1676 ( .A(n1316), .Y(n1314) );
  INVX1 U1677 ( .A(n1314), .Y(n1315) );
  BUFX2 U1678 ( .A(r576_net62631), .Y(n1316) );
  INVX1 U1679 ( .A(n868), .Y(r576_net62631) );
  INVX1 U1680 ( .A(n1879), .Y(n1318) );
  INVX1 U1681 ( .A(n885), .Y(n1319) );
  INVX1 U1682 ( .A(n884), .Y(n1320) );
  INVX1 U1683 ( .A(n869), .Y(n1321) );
  INVX1 U1684 ( .A(n1325), .Y(n1323) );
  INVX1 U1685 ( .A(n1323), .Y(n1324) );
  BUFX2 U1686 ( .A(n3527), .Y(n1325) );
  INVX1 U1687 ( .A(n870), .Y(n3527) );
  INVX1 U1688 ( .A(n3524), .Y(n1327) );
  INVX1 U1689 ( .A(n885), .Y(n1328) );
  INVX1 U1690 ( .A(n884), .Y(n1329) );
  INVX1 U1691 ( .A(n871), .Y(n1330) );
  INVX1 U1692 ( .A(n1334), .Y(n1332) );
  INVX1 U1693 ( .A(n1332), .Y(n1333) );
  BUFX2 U1694 ( .A(n3751), .Y(n1334) );
  INVX1 U1695 ( .A(n872), .Y(n3751) );
  INVX1 U1696 ( .A(n1351), .Y(n1336) );
  INVX1 U1697 ( .A(n889), .Y(n1337) );
  INVX1 U1698 ( .A(n3752), .Y(n1338) );
  INVX1 U1699 ( .A(n874), .Y(n1339) );
  INVX1 U1700 ( .A(n1343), .Y(n1341) );
  INVX1 U1701 ( .A(n1341), .Y(n1342) );
  AND2X1 U1702 ( .A(n1871), .B(n1872), .Y(n1869) );
  INVX1 U1703 ( .A(n1869), .Y(n1343) );
  INVX1 U1704 ( .A(n1346), .Y(n1344) );
  INVX1 U1705 ( .A(n1344), .Y(n1345) );
  AND2X1 U1706 ( .A(n3536), .B(n3535), .Y(n3537) );
  INVX1 U1707 ( .A(n3537), .Y(n1346) );
  INVX1 U1708 ( .A(n1349), .Y(n1347) );
  INVX1 U1709 ( .A(n1347), .Y(n1348) );
  BUFX2 U1710 ( .A(n3657), .Y(n1349) );
  INVX1 U1711 ( .A(n1352), .Y(n1350) );
  INVX1 U1712 ( .A(n1350), .Y(n1351) );
  BUFX2 U1713 ( .A(n3754), .Y(n1352) );
  INVX1 U1714 ( .A(n1355), .Y(n1353) );
  INVX1 U1715 ( .A(n1353), .Y(n1354) );
  BUFX2 U1716 ( .A(n3762), .Y(n1355) );
  INVX1 U1717 ( .A(n1358), .Y(n1356) );
  INVX1 U1718 ( .A(n1356), .Y(n1357) );
  BUFX2 U1719 ( .A(n3867), .Y(n1358) );
  INVX1 U1720 ( .A(n1361), .Y(n1359) );
  INVX1 U1721 ( .A(n1359), .Y(n1360) );
  BUFX2 U1722 ( .A(n3890), .Y(n1361) );
  INVX1 U1723 ( .A(n1364), .Y(n1362) );
  INVX1 U1724 ( .A(n1362), .Y(n1363) );
  BUFX2 U1725 ( .A(n3913), .Y(n1364) );
  INVX1 U1726 ( .A(n1367), .Y(n1365) );
  INVX1 U1727 ( .A(n1365), .Y(n1366) );
  BUFX2 U1728 ( .A(n3998), .Y(n1367) );
  INVX1 U1729 ( .A(n1370), .Y(n1368) );
  INVX1 U1730 ( .A(n1368), .Y(n1369) );
  BUFX2 U1731 ( .A(n4589), .Y(n1370) );
  INVX1 U1732 ( .A(n1373), .Y(n1371) );
  INVX1 U1733 ( .A(n1371), .Y(n1372) );
  OR2X1 U1734 ( .A(n1590), .B(n1605), .Y(n3560) );
  INVX1 U1735 ( .A(n3560), .Y(n1373) );
  INVX1 U1736 ( .A(n1376), .Y(n1374) );
  INVX1 U1737 ( .A(n1374), .Y(n1375) );
  OR2X1 U1738 ( .A(n3564), .B(i[31]), .Y(n2077) );
  INVX1 U1739 ( .A(n2077), .Y(n1376) );
  INVX1 U1740 ( .A(n1379), .Y(n1377) );
  INVX1 U1741 ( .A(n1377), .Y(n1378) );
  OR2X1 U1742 ( .A(n1695), .B(n3846), .Y(n3845) );
  INVX1 U1743 ( .A(n3845), .Y(n1379) );
  INVX1 U1744 ( .A(n1382), .Y(n1380) );
  INVX1 U1745 ( .A(n1380), .Y(n1381) );
  OR2X1 U1746 ( .A(n3914), .B(n3579), .Y(n4449) );
  INVX1 U1747 ( .A(n4449), .Y(n1382) );
  INVX1 U1748 ( .A(n1385), .Y(n1383) );
  INVX1 U1749 ( .A(n1383), .Y(n1384) );
  AND2X1 U1750 ( .A(n3631), .B(n4435), .Y(n4510) );
  INVX1 U1751 ( .A(n4510), .Y(n1385) );
  INVX1 U1752 ( .A(n1388), .Y(n1386) );
  INVX1 U1753 ( .A(n1386), .Y(n1387) );
  OR2X1 U1754 ( .A(n3923), .B(n3631), .Y(n4514) );
  INVX1 U1755 ( .A(n4514), .Y(n1388) );
  INVX1 U1756 ( .A(n1391), .Y(n1389) );
  INVX1 U1757 ( .A(n1389), .Y(n1390) );
  OR2X1 U1758 ( .A(i[2]), .B(n1557), .Y(n4567) );
  INVX1 U1759 ( .A(n4567), .Y(n1391) );
  INVX1 U1760 ( .A(n1394), .Y(n1392) );
  INVX1 U1761 ( .A(n1392), .Y(n1393) );
  AND2X1 U1762 ( .A(n3631), .B(n1657), .Y(n4574) );
  INVX1 U1763 ( .A(n4574), .Y(n1394) );
  INVX1 U1764 ( .A(n891), .Y(n1395) );
  INVX1 U1765 ( .A(n1395), .Y(n1396) );
  INVX1 U1766 ( .A(n1399), .Y(n1397) );
  INVX1 U1767 ( .A(n1397), .Y(n1398) );
  OR2X1 U1768 ( .A(i[5]), .B(n1557), .Y(n4614) );
  INVX1 U1769 ( .A(n4614), .Y(n1399) );
  INVX1 U1770 ( .A(n1402), .Y(n1400) );
  INVX1 U1771 ( .A(n1400), .Y(n1401) );
  BUFX2 U1772 ( .A(n3556), .Y(n1402) );
  INVX1 U1773 ( .A(n1405), .Y(n1403) );
  INVX1 U1774 ( .A(n1403), .Y(n1404) );
  BUFX2 U1775 ( .A(n3648), .Y(n1405) );
  INVX1 U1776 ( .A(n1408), .Y(n1406) );
  INVX1 U1777 ( .A(n1406), .Y(n1407) );
  BUFX2 U1778 ( .A(n3665), .Y(n1408) );
  INVX1 U1779 ( .A(n875), .Y(n3665) );
  INVX1 U1780 ( .A(n888), .Y(n1410) );
  INVX1 U1781 ( .A(n1651), .Y(n1411) );
  INVX1 U1782 ( .A(n3671), .Y(n1412) );
  INVX1 U1783 ( .A(n876), .Y(n1413) );
  INVX1 U1784 ( .A(n1417), .Y(n1415) );
  INVX1 U1785 ( .A(n1415), .Y(n1416) );
  BUFX2 U1786 ( .A(n3683), .Y(n1417) );
  INVX1 U1787 ( .A(n1420), .Y(n1418) );
  INVX1 U1788 ( .A(n1418), .Y(n1419) );
  BUFX2 U1789 ( .A(n4386), .Y(n1420) );
  INVX1 U1790 ( .A(n1423), .Y(n1421) );
  INVX1 U1791 ( .A(n1421), .Y(n1422) );
  BUFX2 U1792 ( .A(n4603), .Y(n1423) );
  INVX1 U1793 ( .A(n1426), .Y(n1424) );
  INVX1 U1794 ( .A(n1424), .Y(n1425) );
  BUFX2 U1795 ( .A(n4606), .Y(n1426) );
  INVX1 U1796 ( .A(n1429), .Y(n1427) );
  INVX1 U1797 ( .A(n1427), .Y(n1428) );
  BUFX2 U1798 ( .A(n4620), .Y(n1429) );
  INVX1 U1799 ( .A(n1432), .Y(n1430) );
  INVX1 U1800 ( .A(n1430), .Y(n1431) );
  AND2X1 U1801 ( .A(n1897), .B(n1898), .Y(net66955) );
  INVX1 U1802 ( .A(net66955), .Y(n1432) );
  INVX1 U1803 ( .A(n1435), .Y(n1433) );
  INVX1 U1804 ( .A(n1433), .Y(n1434) );
  AND2X1 U1805 ( .A(n1880), .B(n1881), .Y(n1899) );
  INVX1 U1806 ( .A(n1899), .Y(n1435) );
  INVX1 U1807 ( .A(n1438), .Y(n1436) );
  INVX1 U1808 ( .A(n1436), .Y(n1437) );
  AND2X1 U1809 ( .A(net66031), .B(n3681), .Y(n3852) );
  INVX1 U1810 ( .A(n3852), .Y(n1438) );
  INVX1 U1811 ( .A(n1441), .Y(n1439) );
  INVX1 U1812 ( .A(n1439), .Y(n1440) );
  AND2X1 U1813 ( .A(n3928), .B(n3930), .Y(net66962) );
  INVX1 U1814 ( .A(net66962), .Y(n1441) );
  INVX1 U1815 ( .A(n1444), .Y(n1442) );
  INVX1 U1816 ( .A(n1442), .Y(n1443) );
  AND2X1 U1817 ( .A(net65992), .B(net66084), .Y(n4428) );
  INVX1 U1818 ( .A(n4428), .Y(n1444) );
  INVX1 U1819 ( .A(n1447), .Y(n1445) );
  INVX1 U1820 ( .A(n1445), .Y(n1446) );
  AND2X1 U1821 ( .A(n1633), .B(n4434), .Y(n4430) );
  INVX1 U1822 ( .A(n4430), .Y(n1447) );
  INVX1 U1823 ( .A(n1450), .Y(n1448) );
  INVX1 U1824 ( .A(n1448), .Y(n1449) );
  AND2X1 U1825 ( .A(n1747), .B(n1735), .Y(n4519) );
  INVX1 U1826 ( .A(n4519), .Y(n1450) );
  INVX1 U1827 ( .A(n1453), .Y(n1451) );
  INVX1 U1828 ( .A(n1451), .Y(n1452) );
  AND2X1 U1829 ( .A(n4599), .B(n4600), .Y(n4595) );
  INVX1 U1830 ( .A(n4595), .Y(n1453) );
  INVX1 U1831 ( .A(n1456), .Y(n1454) );
  INVX1 U1832 ( .A(n1454), .Y(n1455) );
  AND2X1 U1833 ( .A(n3584), .B(n3586), .Y(n4601) );
  INVX1 U1834 ( .A(n4601), .Y(n1456) );
  INVX1 U1835 ( .A(n1459), .Y(n1457) );
  INVX1 U1836 ( .A(n1457), .Y(n1458) );
  AND2X1 U1837 ( .A(n3573), .B(n3576), .Y(n4602) );
  INVX1 U1838 ( .A(n4602), .Y(n1459) );
  INVX1 U1839 ( .A(n1462), .Y(n1460) );
  INVX1 U1840 ( .A(n1460), .Y(n1461) );
  BUFX2 U1841 ( .A(net66956), .Y(n1462) );
  INVX1 U1842 ( .A(n1465), .Y(n1463) );
  INVX1 U1843 ( .A(n1463), .Y(n1464) );
  BUFX2 U1844 ( .A(n4553), .Y(n1465) );
  INVX1 U1845 ( .A(n1468), .Y(n1466) );
  INVX1 U1846 ( .A(n1466), .Y(n1467) );
  BUFX2 U1847 ( .A(n4596), .Y(n1468) );
  INVX1 U1848 ( .A(n1471), .Y(n1469) );
  INVX1 U1849 ( .A(n1469), .Y(n1470) );
  AND2X1 U1850 ( .A(n1707), .B(n1704), .Y(n3649) );
  INVX1 U1851 ( .A(n3649), .Y(n1471) );
  INVX1 U1852 ( .A(n1474), .Y(n1472) );
  INVX1 U1853 ( .A(n1472), .Y(n1473) );
  AND2X1 U1854 ( .A(n1704), .B(n1618), .Y(n3684) );
  INVX1 U1855 ( .A(n3684), .Y(n1474) );
  INVX1 U1856 ( .A(n1477), .Y(n1475) );
  INVX1 U1857 ( .A(n1475), .Y(n1476) );
  AND2X1 U1858 ( .A(n3943), .B(n3945), .Y(n4387) );
  INVX1 U1859 ( .A(n4387), .Y(n1477) );
  INVX1 U1860 ( .A(n1480), .Y(n1478) );
  INVX1 U1861 ( .A(n1478), .Y(n1479) );
  AND2X1 U1862 ( .A(n3612), .B(n3614), .Y(n4604) );
  INVX1 U1863 ( .A(n4604), .Y(n1480) );
  INVX1 U1864 ( .A(n1483), .Y(n1481) );
  INVX1 U1865 ( .A(n1481), .Y(n1482) );
  AND2X1 U1866 ( .A(n3598), .B(n3600), .Y(n4607) );
  INVX1 U1867 ( .A(n4607), .Y(n1483) );
  INVX1 U1868 ( .A(n1486), .Y(n1484) );
  INVX1 U1869 ( .A(n1484), .Y(n1485) );
  BUFX2 U1870 ( .A(n1854), .Y(n1486) );
  INVX1 U1871 ( .A(n1489), .Y(n1487) );
  INVX1 U1872 ( .A(n1487), .Y(n1488) );
  BUFX2 U1873 ( .A(n4554), .Y(n1489) );
  INVX1 U1874 ( .A(n1492), .Y(n1490) );
  INVX1 U1875 ( .A(n1490), .Y(n1491) );
  BUFX2 U1876 ( .A(n4597), .Y(n1492) );
  INVX1 U1877 ( .A(n1495), .Y(n1493) );
  INVX1 U1878 ( .A(n1493), .Y(n1494) );
  AND2X2 U1879 ( .A(n650), .B(n1528), .Y(n1999) );
  INVX1 U1880 ( .A(n1999), .Y(n1495) );
  INVX1 U1881 ( .A(n1498), .Y(n1496) );
  INVX1 U1882 ( .A(n1496), .Y(n1497) );
  AND2X1 U1883 ( .A(n1692), .B(n1624), .Y(n3685) );
  INVX1 U1884 ( .A(n3685), .Y(n1498) );
  INVX1 U1885 ( .A(n1501), .Y(n1499) );
  INVX1 U1886 ( .A(n1499), .Y(n1500) );
  AND2X1 U1887 ( .A(n3939), .B(n3941), .Y(n4388) );
  INVX1 U1888 ( .A(n4388), .Y(n1501) );
  INVX1 U1889 ( .A(n1504), .Y(n1502) );
  INVX1 U1890 ( .A(n1502), .Y(n1503) );
  AND2X1 U1891 ( .A(n3608), .B(n3610), .Y(n4605) );
  INVX1 U1892 ( .A(n4605), .Y(n1504) );
  INVX1 U1893 ( .A(n1507), .Y(n1505) );
  INVX1 U1894 ( .A(n1505), .Y(n1506) );
  AND2X1 U1895 ( .A(n3594), .B(n3596), .Y(n4608) );
  INVX1 U1896 ( .A(n4608), .Y(n1507) );
  INVX1 U1897 ( .A(n1510), .Y(n1508) );
  INVX1 U1898 ( .A(n1508), .Y(n1509) );
  BUFX2 U1899 ( .A(n4000), .Y(n1510) );
  INVX1 U1900 ( .A(n1513), .Y(n1511) );
  INVX1 U1901 ( .A(n1511), .Y(n1512) );
  BUFX2 U1902 ( .A(n3901), .Y(n1513) );
  INVX1 U1903 ( .A(n1516), .Y(n1514) );
  INVX1 U1904 ( .A(n1514), .Y(n1515) );
  BUFX2 U1905 ( .A(n3690), .Y(n1516) );
  INVX1 U1906 ( .A(n1519), .Y(n1517) );
  INVX1 U1907 ( .A(n1517), .Y(n1518) );
  BUFX2 U1908 ( .A(n3655), .Y(n1519) );
  INVX1 U1909 ( .A(n1522), .Y(n1520) );
  INVX1 U1910 ( .A(n1520), .Y(n1521) );
  BUFX2 U1911 ( .A(n3900), .Y(n1522) );
  INVX1 U1912 ( .A(n3776), .Y(n1523) );
  INVX1 U1913 ( .A(n1526), .Y(n1524) );
  INVX1 U1914 ( .A(n1524), .Y(n1525) );
  AND2X1 U1915 ( .A(net66078), .B(net66073), .Y(n4529) );
  INVX1 U1916 ( .A(n4529), .Y(n1526) );
  INVX1 U1917 ( .A(n1529), .Y(n1527) );
  INVX1 U1918 ( .A(n1527), .Y(n1528) );
  BUFX2 U1919 ( .A(n3635), .Y(n1529) );
  INVX1 U1920 ( .A(n1532), .Y(n1530) );
  INVX1 U1921 ( .A(n1530), .Y(n1531) );
  BUFX2 U1922 ( .A(n3766), .Y(n1532) );
  INVX1 U1923 ( .A(n1535), .Y(n1533) );
  INVX1 U1924 ( .A(n1533), .Y(n1534) );
  BUFX2 U1925 ( .A(n3842), .Y(n1535) );
  INVX1 U1926 ( .A(n1538), .Y(n1536) );
  INVX1 U1927 ( .A(n1536), .Y(n1537) );
  AND2X1 U1928 ( .A(n3769), .B(net65987), .Y(n4530) );
  INVX1 U1929 ( .A(n4530), .Y(n1538) );
  INVX1 U1930 ( .A(n3774), .Y(n1539) );
  INVX1 U1931 ( .A(n1542), .Y(n1540) );
  INVX1 U1932 ( .A(n1540), .Y(n1541) );
  AND2X1 U1933 ( .A(n3769), .B(n3855), .Y(n3908) );
  INVX1 U1934 ( .A(n3908), .Y(n1542) );
  BUFX2 U1935 ( .A(n4611), .Y(n1543) );
  INVX4 U1936 ( .A(CMD_data_out[32]), .Y(net66975) );
  INVX1 U1937 ( .A(n1546), .Y(n1544) );
  INVX1 U1938 ( .A(n1544), .Y(n1545) );
  BUFX2 U1939 ( .A(n3757), .Y(n1546) );
  INVX1 U1940 ( .A(n1549), .Y(n1547) );
  INVX1 U1941 ( .A(n1547), .Y(n1548) );
  BUFX2 U1942 ( .A(n4527), .Y(n1549) );
  INVX1 U1943 ( .A(n1552), .Y(n1550) );
  INVX1 U1944 ( .A(n1550), .Y(n1551) );
  BUFX2 U1945 ( .A(n3678), .Y(n1552) );
  INVX1 U1946 ( .A(n1555), .Y(n1553) );
  INVX1 U1947 ( .A(n1553), .Y(n1554) );
  BUFX2 U1948 ( .A(n4431), .Y(n1555) );
  INVX1 U1949 ( .A(n1558), .Y(n1556) );
  INVX1 U1950 ( .A(n1556), .Y(n1557) );
  BUFX2 U1951 ( .A(n4568), .Y(n1558) );
  INVX1 U1952 ( .A(n1561), .Y(n1559) );
  INVX1 U1953 ( .A(n1559), .Y(n1560) );
  OR2X2 U1954 ( .A(n795), .B(n814), .Y(n4583) );
  INVX1 U1955 ( .A(n4583), .Y(n1561) );
  INVX1 U1956 ( .A(n1564), .Y(n1562) );
  INVX1 U1957 ( .A(n1562), .Y(n1563) );
  AND2X1 U1958 ( .A(net66082), .B(net66086), .Y(n4432) );
  INVX1 U1959 ( .A(n4432), .Y(n1564) );
  INVX1 U1960 ( .A(n1567), .Y(n1565) );
  INVX1 U1961 ( .A(n1565), .Y(n1566) );
  BUFX2 U1962 ( .A(n3848), .Y(n1567) );
  INVX1 U1963 ( .A(n1570), .Y(n1568) );
  INVX1 U1964 ( .A(n1568), .Y(n1569) );
  AND2X2 U1965 ( .A(n893), .B(n229), .Y(net92731) );
  INVX1 U1966 ( .A(net92731), .Y(n1570) );
  INVX1 U1967 ( .A(n1573), .Y(n1571) );
  INVX1 U1968 ( .A(n1571), .Y(n1572) );
  AND2X2 U1969 ( .A(n902), .B(net66954), .Y(net89554) );
  INVX1 U1970 ( .A(net89554), .Y(n1573) );
  OR2X1 U1971 ( .A(n231), .B(net66329), .Y(net82454) );
  INVX1 U1972 ( .A(net82454), .Y(n1574) );
  INVX1 U1973 ( .A(n1574), .Y(net82455) );
  OR2X1 U1974 ( .A(net66327), .B(net66329), .Y(net80708) );
  INVX1 U1975 ( .A(net80708), .Y(n1575) );
  INVX1 U1976 ( .A(n1575), .Y(net80709) );
  OR2X1 U1977 ( .A(net66327), .B(n232), .Y(net80717) );
  INVX1 U1978 ( .A(net80717), .Y(n1576) );
  INVX1 U1979 ( .A(n1576), .Y(net80718) );
  INVX1 U1980 ( .A(n1579), .Y(n1577) );
  INVX1 U1981 ( .A(n1577), .Y(n1578) );
  AND2X1 U1982 ( .A(net66063), .B(n4511), .Y(n3686) );
  INVX1 U1983 ( .A(n3686), .Y(n1579) );
  INVX1 U1984 ( .A(n1582), .Y(n1580) );
  INVX1 U1985 ( .A(n1580), .Y(n1581) );
  BUFX2 U1986 ( .A(n4523), .Y(n1582) );
  INVX1 U1987 ( .A(n1585), .Y(n1583) );
  INVX1 U1988 ( .A(n1583), .Y(n1584) );
  BUFX2 U1989 ( .A(n3889), .Y(n1585) );
  INVX1 U1990 ( .A(n1588), .Y(n1586) );
  INVX1 U1991 ( .A(n1586), .Y(n1587) );
  OR2X1 U1992 ( .A(i[31]), .B(n3557), .Y(n3126) );
  INVX1 U1993 ( .A(n3126), .Y(n1588) );
  INVX1 U1994 ( .A(n1591), .Y(n1589) );
  INVX1 U1995 ( .A(n1589), .Y(n1590) );
  BUFX2 U1996 ( .A(n3559), .Y(n1591) );
  INVX1 U1997 ( .A(n877), .Y(n3559) );
  INVX1 U1998 ( .A(n3551), .Y(n1593) );
  INVX1 U1999 ( .A(n887), .Y(n1594) );
  INVX1 U2000 ( .A(n886), .Y(n1595) );
  INVX1 U2001 ( .A(n878), .Y(n1596) );
  INVX1 U2002 ( .A(n1600), .Y(n1598) );
  INVX1 U2003 ( .A(n1598), .Y(n1599) );
  BUFX2 U2004 ( .A(n3849), .Y(n1600) );
  INVX1 U2005 ( .A(n1603), .Y(n1601) );
  INVX1 U2006 ( .A(n1601), .Y(n1602) );
  AND2X1 U2007 ( .A(n3861), .B(ring_ptr[0]), .Y(n3858) );
  INVX1 U2008 ( .A(n3858), .Y(n1603) );
  INVX1 U2009 ( .A(n1606), .Y(n1604) );
  INVX1 U2010 ( .A(n1604), .Y(n1605) );
  AND2X2 U2011 ( .A(n905), .B(n3554), .Y(n3558) );
  INVX1 U2012 ( .A(n3558), .Y(n1606) );
  INVX1 U2013 ( .A(n1610), .Y(n1608) );
  INVX1 U2014 ( .A(n1608), .Y(n1609) );
  AND2X1 U2015 ( .A(n3920), .B(n3639), .Y(n3704) );
  INVX1 U2016 ( .A(n3704), .Y(n1610) );
  INVX1 U2017 ( .A(n1613), .Y(n1611) );
  INVX1 U2018 ( .A(n1611), .Y(n1612) );
  BUFX2 U2019 ( .A(n3949), .Y(n1613) );
  INVX1 U2020 ( .A(n1616), .Y(n1614) );
  INVX1 U2021 ( .A(n1614), .Y(n1615) );
  AND2X2 U2022 ( .A(n3639), .B(n656), .Y(n3921) );
  INVX1 U2023 ( .A(n3921), .Y(n1616) );
  INVX1 U2024 ( .A(n1619), .Y(n1617) );
  INVX1 U2025 ( .A(n1617), .Y(n1618) );
  BUFX2 U2026 ( .A(n3662), .Y(n1619) );
  INVX1 U2027 ( .A(n1622), .Y(n1620) );
  INVX1 U2028 ( .A(n1620), .Y(n1621) );
  BUFX2 U2029 ( .A(n3862), .Y(n1622) );
  INVX1 U2030 ( .A(n1625), .Y(n1623) );
  INVX1 U2031 ( .A(n1623), .Y(n1624) );
  AND2X1 U2032 ( .A(n4531), .B(state[2]), .Y(net66042) );
  INVX1 U2033 ( .A(net66042), .Y(n1625) );
  INVX1 U2034 ( .A(n1628), .Y(n1626) );
  INVX1 U2035 ( .A(n1626), .Y(n1627) );
  AND2X2 U2036 ( .A(n3661), .B(n1541), .Y(n3773) );
  INVX1 U2037 ( .A(n3773), .Y(n1628) );
  INVX1 U2038 ( .A(n1631), .Y(n1629) );
  INVX1 U2039 ( .A(n1629), .Y(n1630) );
  BUFX2 U2040 ( .A(n3909), .Y(n1631) );
  INVX1 U2041 ( .A(n1634), .Y(n1632) );
  INVX1 U2042 ( .A(n1632), .Y(n1633) );
  OR2X2 U2043 ( .A(n798), .B(n820), .Y(n4433) );
  INVX1 U2044 ( .A(n4433), .Y(n1634) );
  INVX1 U2045 ( .A(n1637), .Y(n1635) );
  INVX1 U2046 ( .A(n1635), .Y(n1636) );
  OR2X1 U2047 ( .A(n1698), .B(n1657), .Y(n3702) );
  INVX1 U2048 ( .A(n3702), .Y(n1637) );
  INVX1 U2049 ( .A(n1640), .Y(n1638) );
  INVX1 U2050 ( .A(n1638), .Y(n1639) );
  AND2X2 U2051 ( .A(n3914), .B(n1509), .Y(n3863) );
  INVX1 U2052 ( .A(n3863), .Y(n1640) );
  INVX1 U2053 ( .A(n1643), .Y(n1641) );
  INVX1 U2054 ( .A(n1641), .Y(n1642) );
  AND2X2 U2055 ( .A(net67172), .B(n659), .Y(n4578) );
  INVX1 U2056 ( .A(n4578), .Y(n1643) );
  INVX1 U2057 ( .A(n1646), .Y(n1644) );
  INVX1 U2058 ( .A(n1644), .Y(n1645) );
  OR2X2 U2059 ( .A(n786), .B(n804), .Y(net66061) );
  INVX1 U2061 ( .A(net66061), .Y(n1646) );
  INVX1 U2062 ( .A(n1649), .Y(n1647) );
  INVX1 U2233 ( .A(n1647), .Y(n1648) );
  AND2X1 U2234 ( .A(n1867), .B(n1868), .Y(r576_GE_LT_GT_LE) );
  INVX1 U2236 ( .A(r576_GE_LT_GT_LE), .Y(n1649) );
  INVX1 U2237 ( .A(n1652), .Y(n1650) );
  INVX1 U2238 ( .A(n1650), .Y(n1651) );
  AND2X1 U2239 ( .A(n3914), .B(n4538), .Y(n3672) );
  INVX1 U2240 ( .A(n3672), .Y(n1652) );
  INVX1 U2241 ( .A(n1655), .Y(n1653) );
  INVX1 U2242 ( .A(n1653), .Y(n1654) );
  BUFX2 U2243 ( .A(net66151), .Y(n1655) );
  INVX1 U2244 ( .A(n1658), .Y(n1656) );
  INVX1 U2245 ( .A(n1656), .Y(n1657) );
  BUFX2 U2246 ( .A(n3759), .Y(n1658) );
  INVX1 U2247 ( .A(n1661), .Y(n1659) );
  INVX1 U2248 ( .A(n1659), .Y(n1660) );
  BUFX2 U2249 ( .A(n3922), .Y(n1661) );
  AND2X2 U2250 ( .A(n1716), .B(n1543), .Y(n3705) );
  INVX1 U2251 ( .A(n3705), .Y(n1662) );
  INVX1 U2252 ( .A(n3705), .Y(n1663) );
  INVX1 U2253 ( .A(n1666), .Y(n1664) );
  INVX1 U2254 ( .A(n1664), .Y(n1665) );
  BUFX2 U2255 ( .A(n4579), .Y(n1666) );
  INVX1 U2256 ( .A(n1669), .Y(n1667) );
  INVX1 U2257 ( .A(n1667), .Y(n1668) );
  OR2X2 U2258 ( .A(n801), .B(n817), .Y(n3856) );
  INVX1 U2259 ( .A(n3856), .Y(n1669) );
  BUFX2 U2260 ( .A(n545), .Y(n1818) );
  BUFX2 U2261 ( .A(n545), .Y(n1819) );
  BUFX2 U2262 ( .A(n545), .Y(n1820) );
  INVX1 U2263 ( .A(n3894), .Y(n1670) );
  INVX1 U2264 ( .A(n1670), .Y(n1671) );
  INVX1 U2265 ( .A(n1670), .Y(n1672) );
  INVX1 U2266 ( .A(n1675), .Y(n1673) );
  INVX1 U2267 ( .A(n1673), .Y(n1674) );
  BUFX2 U2268 ( .A(n3674), .Y(n1675) );
  INVX1 U2269 ( .A(n1678), .Y(n1676) );
  INVX1 U2270 ( .A(n1676), .Y(n1677) );
  BUFX2 U2271 ( .A(n3915), .Y(n1678) );
  INVX1 U2272 ( .A(n1681), .Y(n1679) );
  INVX1 U2273 ( .A(n1679), .Y(n1680) );
  AND2X1 U2274 ( .A(n1735), .B(n1707), .Y(n3666) );
  INVX1 U2275 ( .A(n3666), .Y(n1681) );
  INVX1 U2276 ( .A(n1684), .Y(n1682) );
  INVX1 U2277 ( .A(n1682), .Y(n1683) );
  AND2X1 U2278 ( .A(n1692), .B(n1710), .Y(n3758) );
  INVX1 U2279 ( .A(n3758), .Y(n1684) );
  INVX1 U2280 ( .A(n1687), .Y(n1685) );
  INVX1 U2281 ( .A(n1685), .Y(n1686) );
  AND2X1 U2282 ( .A(n3540), .B(n3539), .Y(r577_GE_LT_GT_LE) );
  INVX1 U2283 ( .A(r577_GE_LT_GT_LE), .Y(n1687) );
  INVX1 U2284 ( .A(n3633), .Y(n1688) );
  INVX1 U2285 ( .A(n1688), .Y(n1689) );
  INVX1 U2286 ( .A(n1688), .Y(n1690) );
  INVX1 U2287 ( .A(n1693), .Y(n1691) );
  INVX1 U2288 ( .A(n1691), .Y(n1692) );
  BUFX2 U2289 ( .A(n3652), .Y(n1693) );
  INVX1 U2290 ( .A(n1696), .Y(n1694) );
  INVX1 U2291 ( .A(n1694), .Y(n1695) );
  AND2X1 U2292 ( .A(n1735), .B(n1738), .Y(n3632) );
  INVX1 U2293 ( .A(n3632), .Y(n1696) );
  INVX1 U2294 ( .A(n1699), .Y(n1697) );
  INVX1 U2295 ( .A(n1697), .Y(n1698) );
  BUFX2 U2296 ( .A(n3912), .Y(n1699) );
  INVX1 U2297 ( .A(n1702), .Y(n1700) );
  INVX1 U2298 ( .A(n1700), .Y(n1701) );
  AND2X1 U2299 ( .A(n4533), .B(net65987), .Y(n3699) );
  INVX1 U2300 ( .A(n3699), .Y(n1702) );
  INVX1 U2301 ( .A(n1705), .Y(n1703) );
  INVX1 U2302 ( .A(n1703), .Y(n1704) );
  BUFX2 U2303 ( .A(n3654), .Y(n1705) );
  INVX1 U2304 ( .A(n1708), .Y(n1706) );
  INVX1 U2305 ( .A(n1706), .Y(n1707) );
  BUFX2 U2306 ( .A(n3653), .Y(n1708) );
  INVX1 U2307 ( .A(n1711), .Y(n1709) );
  INVX1 U2308 ( .A(n1709), .Y(n1710) );
  AND2X1 U2309 ( .A(n4531), .B(net66031), .Y(n3700) );
  INVX1 U2310 ( .A(n3700), .Y(n1711) );
  INVX1 U2311 ( .A(n1714), .Y(n1712) );
  INVX1 U2312 ( .A(n1712), .Y(n1713) );
  BUFX2 U2313 ( .A(net66283), .Y(n1714) );
  INVX1 U2314 ( .A(n879), .Y(n1715) );
  INVX1 U2315 ( .A(n1715), .Y(n1716) );
  INVX1 U2316 ( .A(n1715), .Y(n1717) );
  INVX1 U2317 ( .A(n880), .Y(n1718) );
  INVX1 U2318 ( .A(n3647), .Y(n1720) );
  INVX1 U2319 ( .A(n1720), .Y(n1721) );
  INVX1 U2320 ( .A(n1720), .Y(n1722) );
  INVX1 U2321 ( .A(n1720), .Y(n1723) );
  INVX1 U2322 ( .A(n1727), .Y(n1724) );
  INVX1 U2323 ( .A(n1724), .Y(n1725) );
  INVX1 U2324 ( .A(n1724), .Y(n1726) );
  AND2X2 U2325 ( .A(CMD_data_out[33]), .B(n1662), .Y(n3669) );
  INVX1 U2326 ( .A(n3669), .Y(n1727) );
  INVX1 U2327 ( .A(n1730), .Y(n1728) );
  INVX1 U2328 ( .A(n1728), .Y(n1729) );
  BUFX2 U2329 ( .A(net66166), .Y(n1730) );
  INVX1 U2330 ( .A(n1733), .Y(n1731) );
  INVX1 U2331 ( .A(n1731), .Y(n1732) );
  BUFX2 U2332 ( .A(n447), .Y(n1733) );
  INVX1 U2333 ( .A(n1736), .Y(n1734) );
  INVX1 U2334 ( .A(n1734), .Y(n1735) );
  AND2X1 U2335 ( .A(n3847), .B(net67122), .Y(n3680) );
  INVX1 U2336 ( .A(n3680), .Y(n1736) );
  INVX1 U2337 ( .A(n1739), .Y(n1737) );
  INVX1 U2338 ( .A(n1737), .Y(n1738) );
  BUFX2 U2339 ( .A(net66046), .Y(n1739) );
  INVX1 U2340 ( .A(n1742), .Y(n1740) );
  BUFX2 U2341 ( .A(n3675), .Y(n1742) );
  INVX1 U2342 ( .A(n1745), .Y(n1743) );
  INVX1 U2343 ( .A(n1743), .Y(n1744) );
  AND2X2 U2344 ( .A(n1738), .B(n1615), .Y(n4465) );
  INVX1 U2345 ( .A(n4465), .Y(n1745) );
  INVX1 U2346 ( .A(n1748), .Y(n1746) );
  INVX1 U2347 ( .A(n1746), .Y(n1747) );
  BUFX2 U2348 ( .A(n3668), .Y(n1748) );
  INVX1 U2349 ( .A(n1751), .Y(n1749) );
  INVX4 U2350 ( .A(n1749), .Y(n1750) );
  OR2X2 U2351 ( .A(n1689), .B(reset), .Y(n3872) );
  INVX1 U2352 ( .A(n3872), .Y(n1751) );
  INVX1 U2353 ( .A(n1783), .Y(n1781) );
  INVX1 U2354 ( .A(n1781), .Y(n1782) );
  OR2X2 U2355 ( .A(n1707), .B(n4391), .Y(n4392) );
  INVX1 U2356 ( .A(n4392), .Y(n1783) );
  INVX1 U2357 ( .A(n1786), .Y(n1784) );
  INVX1 U2358 ( .A(n1784), .Y(n1785) );
  OR2X2 U2359 ( .A(n1735), .B(n4391), .Y(n4393) );
  INVX1 U2360 ( .A(n4393), .Y(n1786) );
  INVX1 U2361 ( .A(n1789), .Y(n1787) );
  INVX8 U2362 ( .A(n1787), .Y(n1788) );
  BUFX2 U2363 ( .A(n3645), .Y(n1789) );
  INVX1 U2364 ( .A(n1792), .Y(n1790) );
  INVX1 U2365 ( .A(n1790), .Y(n1791) );
  BUFX2 U2366 ( .A(net66319), .Y(n1792) );
  INVX1 U2367 ( .A(n881), .Y(net66319) );
  INVX1 U2368 ( .A(n1738), .Y(n1794) );
  INVX1 U2369 ( .A(n1609), .Y(n1795) );
  INVX1 U2370 ( .A(n1612), .Y(n1796) );
  INVX1 U2371 ( .A(n882), .Y(n1797) );
  INVX1 U2372 ( .A(n546), .Y(n1799) );
  INVX1 U2373 ( .A(net92933), .Y(n1800) );
  INVX1 U2374 ( .A(n535), .Y(net80595) );
  MUX2X1 U2375 ( .B(buff_data[430]), .A(n567), .S(net93057), .Y(n1805) );
  INVX8 U2376 ( .A(n1805), .Y(n2698) );
  INVX1 U2377 ( .A(n462), .Y(net92836) );
  AND2X2 U2378 ( .A(n547), .B(net66441), .Y(net66714) );
  INVX1 U2379 ( .A(n230), .Y(net66325) );
  INVX8 U2380 ( .A(net79438), .Y(net79436) );
  INVX8 U2381 ( .A(n229), .Y(net79438) );
  NOR3X1 U2382 ( .A(net79438), .B(net79414), .C(net66325), .Y(net66423) );
  INVX8 U2383 ( .A(net79438), .Y(net79432) );
  INVX8 U2384 ( .A(net79438), .Y(net79434) );
  MUX2X1 U2385 ( .B(buff_data[446]), .A(buff_data[430]), .S(net79414), .Y(
        C25909_net2920) );
  AND2X2 U2386 ( .A(net92619), .B(net66423), .Y(net66834) );
  INVX2 U2387 ( .A(net92738), .Y(net92651) );
  AND2X2 U2388 ( .A(net92747), .B(net92651), .Y(net92619) );
  OAI21X1 U2389 ( .A(n555), .B(n1807), .C(net92773), .Y(net92747) );
  OAI21X1 U2390 ( .A(net92789), .B(n555), .C(n442), .Y(net92761) );
  INVX1 U2391 ( .A(n464), .Y(n1813) );
  INVX1 U2392 ( .A(n1654), .Y(net66007) );
  NAND3X1 U2393 ( .A(net66974), .B(net66975), .C(CMD_data_out[33]), .Y(
        net66970) );
  INVX2 U2394 ( .A(n1648), .Y(n1811) );
  INVX2 U2395 ( .A(n1738), .Y(n1809) );
  NOR3X1 U2396 ( .A(net66290), .B(n1809), .C(net66160), .Y(net66289) );
  MUX2X1 U2397 ( .B(buff_data[424]), .A(n566), .S(net79538), .Y(n1814) );
  INVX8 U2398 ( .A(n1814), .Y(n2704) );
  MUX2X1 U2399 ( .B(buff_data[440]), .A(buff_data[424]), .S(net79402), .Y(
        C25909_net2740) );
  INVX1 U2400 ( .A(net79794), .Y(net93077) );
  INVX1 U2401 ( .A(n610), .Y(net93072) );
  INVX1 U2402 ( .A(n2129), .Y(n1829) );
  INVX1 U2403 ( .A(n2129), .Y(n1833) );
  INVX1 U2404 ( .A(n4), .Y(n1816) );
  INVX1 U2405 ( .A(net92789), .Y(net93022) );
  INVX1 U2406 ( .A(n2194), .Y(n1817) );
  MUX2X1 U2407 ( .B(n1823), .A(n1822), .S(n543), .Y(n1821) );
  INVX8 U2408 ( .A(buff_data[109]), .Y(n1822) );
  INVX8 U2409 ( .A(n579), .Y(n1823) );
  INVX1 U2410 ( .A(n4356), .Y(n1912) );
  INVX1 U2411 ( .A(n556), .Y(n2027) );
  MUX2X1 U2412 ( .B(n565), .A(buff_data[201]), .S(n404), .Y(n4127) );
  INVX1 U2413 ( .A(n373), .Y(net92933) );
  INVX1 U2414 ( .A(n373), .Y(net79794) );
  MUX2X1 U2415 ( .B(n1828), .A(n1827), .S(n1829), .Y(n1826) );
  INVX8 U2416 ( .A(buff_data[103]), .Y(n1827) );
  INVX8 U2417 ( .A(n578), .Y(n1828) );
  MUX2X1 U2418 ( .B(n1832), .A(n1831), .S(n1833), .Y(n1830) );
  INVX8 U2419 ( .A(buff_data[97]), .Y(n1831) );
  INVX8 U2420 ( .A(n577), .Y(n1832) );
  INVX1 U2421 ( .A(net80718), .Y(n1847) );
  INVX1 U2422 ( .A(n100), .Y(n2037) );
  INVX1 U2423 ( .A(n187), .Y(n1835) );
  INVX1 U2424 ( .A(n4218), .Y(n1836) );
  INVX1 U2425 ( .A(n4218), .Y(n1837) );
  INVX1 U2426 ( .A(n317), .Y(net92856) );
  MUX2X1 U2427 ( .B(n1840), .A(n1839), .S(n86), .Y(n1838) );
  INVX8 U2428 ( .A(buff_data[276]), .Y(n1839) );
  INVX8 U2429 ( .A(n576), .Y(n1840) );
  INVX1 U2430 ( .A(n466), .Y(n4356) );
  AOI21X1 U2431 ( .A(n442), .B(n385), .C(net82455), .Y(net66558) );
  MUX2X1 U2432 ( .B(buff_data[468]), .A(buff_data[452]), .S(net79412), .Y(
        C25909_net2624) );
  INVX2 U2433 ( .A(net80709), .Y(net92748) );
  INVX1 U2434 ( .A(n563), .Y(n1850) );
  INVX1 U2435 ( .A(n424), .Y(net92789) );
  INVX8 U2436 ( .A(n1847), .Y(n1849) );
  OR2X2 U2437 ( .A(net92773), .B(n1849), .Y(n1845) );
  INVX2 U2438 ( .A(n1572), .Y(net89562) );
  BUFX2 U2439 ( .A(net93022), .Y(net82506) );
  NOR3X1 U2440 ( .A(n1431), .B(n1461), .C(n1485), .Y(net66954) );
  NAND3X1 U2441 ( .A(n1852), .B(n1853), .C(n1851), .Y(n1854) );
  INVX1 U2442 ( .A(j[23]), .Y(n1851) );
  OAI21X1 U2443 ( .A(n1791), .B(n1851), .C(n966), .Y(n3154) );
  INVX1 U2444 ( .A(j[25]), .Y(n1853) );
  OAI21X1 U2445 ( .A(n1791), .B(n1853), .C(n968), .Y(n3150) );
  INVX1 U2446 ( .A(j[24]), .Y(n1852) );
  OAI21X1 U2447 ( .A(n1791), .B(n1852), .C(n967), .Y(n3152) );
  INVX1 U2448 ( .A(net92867), .Y(net89705) );
  OR2X2 U2449 ( .A(n1738), .B(n1855), .Y(net65981) );
  OAI21X1 U2450 ( .A(n1791), .B(n1856), .C(n954), .Y(n3178) );
  OAI21X1 U2451 ( .A(n1791), .B(n1857), .C(n953), .Y(n3180) );
  OAI21X1 U2452 ( .A(n1791), .B(n1858), .C(n957), .Y(n3172) );
  OAI21X1 U2453 ( .A(n1791), .B(n1859), .C(n958), .Y(n3170) );
  OAI21X1 U2454 ( .A(n1791), .B(n1860), .C(n955), .Y(n3176) );
  OAI21X1 U2455 ( .A(n1791), .B(n1861), .C(n956), .Y(n3174) );
  INVX2 U2456 ( .A(j[10]), .Y(n1857) );
  INVX2 U2457 ( .A(j[11]), .Y(n1856) );
  INVX2 U2458 ( .A(j[12]), .Y(n1860) );
  INVX2 U2459 ( .A(j[13]), .Y(n1861) );
  INVX2 U2460 ( .A(j[14]), .Y(n1858) );
  INVX2 U2461 ( .A(j[15]), .Y(n1859) );
  INVX8 U2462 ( .A(net79414), .Y(net79422) );
  INVX8 U2463 ( .A(net79414), .Y(net79416) );
  INVX8 U2464 ( .A(net79414), .Y(net79420) );
  INVX1 U2465 ( .A(n1648), .Y(net66140) );
  AOI22X1 U2466 ( .A(n1645), .B(net66062), .C(n1648), .D(net66063), .Y(
        net66060) );
  OAI21X1 U2467 ( .A(n1253), .B(n1342), .C(n1870), .Y(n1868) );
  INVX1 U2468 ( .A(i[31]), .Y(n1870) );
  OAI21X1 U2469 ( .A(n1256), .B(n1315), .C(n1870), .Y(n1867) );
  NOR3X1 U2470 ( .A(n1873), .B(i[14]), .C(i[13]), .Y(n1872) );
  OR2X1 U2471 ( .A(i[1]), .B(i[15]), .Y(n1873) );
  NOR3X1 U2472 ( .A(n1874), .B(i[10]), .C(i[0]), .Y(n1871) );
  OR2X1 U2473 ( .A(i[12]), .B(i[11]), .Y(n1874) );
  NOR3X1 U2474 ( .A(n1877), .B(i[7]), .C(i[6]), .Y(n1876) );
  OR2X1 U2475 ( .A(i[9]), .B(i[8]), .Y(n1877) );
  NOR3X1 U2476 ( .A(n1878), .B(i[3]), .C(i[2]), .Y(n1875) );
  OR2X1 U2477 ( .A(i[5]), .B(i[4]), .Y(n1878) );
  NOR3X1 U2478 ( .A(i[16]), .B(i[18]), .C(i[17]), .Y(n1879) );
  INVX1 U2479 ( .A(n166), .Y(net66499) );
  NAND3X1 U2480 ( .A(net67122), .B(state[0]), .C(state[2]), .Y(net66046) );
  NAND3X1 U2481 ( .A(n1882), .B(n1883), .C(n1896), .Y(net66956) );
  AND2X1 U2482 ( .A(n1895), .B(n1884), .Y(n1896) );
  INVX1 U2483 ( .A(j[28]), .Y(n1884) );
  OAI21X1 U2484 ( .A(n1791), .B(n1884), .C(n971), .Y(n3144) );
  INVX1 U2485 ( .A(j[29]), .Y(n1895) );
  OAI21X1 U2486 ( .A(n1791), .B(n1895), .C(n513), .Y(n3142) );
  INVX1 U2487 ( .A(j[27]), .Y(n1883) );
  OAI21X1 U2488 ( .A(n1791), .B(n1883), .C(n970), .Y(n3146) );
  INVX1 U2489 ( .A(j[26]), .Y(n1882) );
  OAI21X1 U2490 ( .A(n1791), .B(n1882), .C(n969), .Y(n3148) );
  NOR3X1 U2491 ( .A(n1434), .B(reset), .C(j[9]), .Y(n1898) );
  INVX1 U2492 ( .A(j[8]), .Y(n1881) );
  OAI21X1 U2493 ( .A(n1791), .B(n1881), .C(n951), .Y(n3184) );
  INVX1 U2494 ( .A(j[7]), .Y(n1880) );
  OAI21X1 U2495 ( .A(n1791), .B(n1880), .C(n950), .Y(n3186) );
  NOR3X1 U2496 ( .A(n1440), .B(j[31]), .C(j[30]), .Y(n1897) );
  INVX1 U2497 ( .A(n2000), .Y(n1992) );
  INVX8 U2498 ( .A(buff_data[476]), .Y(n1901) );
  MUX2X1 U2499 ( .B(net84792), .A(n1903), .S(n2041), .Y(n1902) );
  INVX8 U2500 ( .A(buff_data[366]), .Y(n1903) );
  INVX8 U2501 ( .A(n567), .Y(net84792) );
  INVX1 U2502 ( .A(n2192), .Y(n1904) );
  INVX8 U2503 ( .A(buff_data[405]), .Y(n1906) );
  MUX2X1 U2504 ( .B(n1910), .A(n579), .S(n206), .Y(n1909) );
  INVX8 U2505 ( .A(n1909), .Y(net80914) );
  OAI21X1 U2506 ( .A(n1791), .B(net66329), .C(n947), .Y(n3192) );
  INVX8 U2507 ( .A(n1908), .Y(n1910) );
  INVX8 U2508 ( .A(buff_data[253]), .Y(n1908) );
  NOR3X1 U2509 ( .A(net79436), .B(n230), .C(net79414), .Y(net66539) );
  MUX2X1 U2510 ( .B(net82576), .A(n1914), .S(n1815), .Y(n1913) );
  INVX8 U2511 ( .A(buff_data[244]), .Y(n1914) );
  INVX8 U2512 ( .A(n576), .Y(net82576) );
  MUX2X1 U2513 ( .B(net82567), .A(n1916), .S(net80464), .Y(n1915) );
  INVX8 U2514 ( .A(buff_data[173]), .Y(n1916) );
  INVX8 U2515 ( .A(n579), .Y(net82567) );
  INVX8 U2516 ( .A(buff_data[168]), .Y(n1918) );
  INVX8 U2517 ( .A(buff_data[255]), .Y(n1920) );
  INVX1 U2518 ( .A(n1912), .Y(n1921) );
  INVX1 U2519 ( .A(n19), .Y(n2028) );
  MUX2X1 U2520 ( .B(n566), .A(buff_data[200]), .S(n404), .Y(n4126) );
  MUX2X1 U2521 ( .B(n1925), .A(n1924), .S(n384), .Y(n1923) );
  INVX8 U2522 ( .A(buff_data[199]), .Y(n1924) );
  INVX8 U2523 ( .A(n578), .Y(n1925) );
  INVX1 U2524 ( .A(n445), .Y(n2116) );
  INVX1 U2525 ( .A(n341), .Y(net82472) );
  INVX8 U2526 ( .A(buff_data[18]), .Y(n1930) );
  INVX1 U2527 ( .A(n210), .Y(n2022) );
  INVX8 U2528 ( .A(buff_data[234]), .Y(n1933) );
  INVX1 U2529 ( .A(n52), .Y(n2126) );
  INVX8 U2530 ( .A(buff_data[233]), .Y(n1935) );
  MUX2X1 U2531 ( .B(net82435), .A(n1937), .S(n552), .Y(n1936) );
  INVX8 U2532 ( .A(buff_data[29]), .Y(n1937) );
  INVX8 U2533 ( .A(n579), .Y(net82435) );
  INVX1 U2534 ( .A(n404), .Y(net82427) );
  INVX1 U2535 ( .A(n404), .Y(net82428) );
  INVX8 U2536 ( .A(buff_data[14]), .Y(n1939) );
  MUX2X1 U2537 ( .B(n1942), .A(n1941), .S(n552), .Y(n1940) );
  INVX8 U2538 ( .A(buff_data[25]), .Y(n1941) );
  INVX8 U2539 ( .A(n565), .Y(n1942) );
  MUX2X1 U2540 ( .B(n1945), .A(n1944), .S(n2), .Y(n1943) );
  INVX8 U2541 ( .A(buff_data[225]), .Y(n1944) );
  INVX8 U2542 ( .A(n577), .Y(n1945) );
  INVX8 U2543 ( .A(buff_data[172]), .Y(n1947) );
  INVX8 U2544 ( .A(buff_data[238]), .Y(n1950) );
  INVX8 U2545 ( .A(buff_data[176]), .Y(n1952) );
  INVX8 U2546 ( .A(n4051), .Y(n3023) );
  INVX8 U2547 ( .A(n4046), .Y(n3029) );
  INVX1 U2548 ( .A(net82506), .Y(net82348) );
  INVX1 U2549 ( .A(net82348), .Y(net82349) );
  MUX2X1 U2550 ( .B(n1957), .A(n1956), .S(n563), .Y(n1955) );
  INVX8 U2551 ( .A(buff_data[473]), .Y(n1956) );
  INVX8 U2552 ( .A(n565), .Y(n1957) );
  INVX1 U2553 ( .A(n610), .Y(net82336) );
  INVX8 U2554 ( .A(buff_data[250]), .Y(n1959) );
  INVX8 U2555 ( .A(buff_data[278]), .Y(n1962) );
  INVX8 U2556 ( .A(buff_data[69]), .Y(n1965) );
  INVX8 U2557 ( .A(buff_data[178]), .Y(n1968) );
  MUX2X1 U2558 ( .B(n1971), .A(n1970), .S(n7), .Y(n1969) );
  INVX8 U2559 ( .A(buff_data[177]), .Y(n1970) );
  INVX8 U2560 ( .A(n577), .Y(n1971) );
  INVX8 U2561 ( .A(buff_data[280]), .Y(n1975) );
  MUX2X1 U2562 ( .B(n1978), .A(n1977), .S(net80839), .Y(n1976) );
  INVX8 U2563 ( .A(buff_data[379]), .Y(n1977) );
  INVX8 U2564 ( .A(n571), .Y(n1978) );
  INVX8 U2565 ( .A(buff_data[416]), .Y(n1980) );
  MUX2X1 U2566 ( .B(n1983), .A(n1982), .S(n414), .Y(n1981) );
  INVX8 U2567 ( .A(buff_data[279]), .Y(n1982) );
  INVX8 U2568 ( .A(n578), .Y(n1983) );
  MUX2X1 U2569 ( .B(net82215), .A(n1985), .S(n2036), .Y(n1984) );
  INVX8 U2570 ( .A(buff_data[333]), .Y(n1985) );
  INVX8 U2571 ( .A(n579), .Y(net82215) );
  MUX2X1 U2572 ( .B(net82209), .A(n1987), .S(net80682), .Y(n1986) );
  INVX8 U2573 ( .A(buff_data[301]), .Y(n1987) );
  INVX8 U2574 ( .A(n579), .Y(net82209) );
  INVX1 U2575 ( .A(n1992), .Y(n1988) );
  INVX8 U2576 ( .A(buff_data[457]), .Y(n1990) );
  INVX1 U2577 ( .A(n216), .Y(n1991) );
  INVX1 U2578 ( .A(n417), .Y(net82191) );
  INVX4 U2579 ( .A(n434), .Y(n4447) );
  AND2X2 U2580 ( .A(n4503), .B(n4440), .Y(n4451) );
  INVX1 U2581 ( .A(n341), .Y(net82138) );
  MUX2X1 U2582 ( .B(net82125), .A(n1994), .S(net80839), .Y(n1993) );
  INVX8 U2583 ( .A(buff_data[372]), .Y(n1994) );
  INVX8 U2584 ( .A(n576), .Y(net82125) );
  AND2X2 U2585 ( .A(net82472), .B(net66503), .Y(n1995) );
  INVX1 U2586 ( .A(n371), .Y(n1996) );
  NOR3X1 U2587 ( .A(net82094), .B(n1998), .C(n1494), .Y(n1997) );
  INVX8 U2588 ( .A(n1690), .Y(n1998) );
  MUX2X1 U2589 ( .B(buff_data[377]), .A(n565), .S(net79518), .Y(n2001) );
  INVX8 U2590 ( .A(n2001), .Y(n2750) );
  AND2X2 U2591 ( .A(n548), .B(net66539), .Y(n2000) );
  MUX2X1 U2592 ( .B(buff_data[377]), .A(buff_data[361]), .S(net79402), .Y(
        C25909_net2767) );
  INVX1 U2593 ( .A(n231), .Y(net66327) );
  OAI21X1 U2594 ( .A(n1791), .B(net66327), .C(n946), .Y(n3194) );
  MUX2X1 U2595 ( .B(n2005), .A(n2004), .S(n2160), .Y(n2003) );
  INVX8 U2596 ( .A(buff_data[316]), .Y(n2004) );
  INVX8 U2597 ( .A(n572), .Y(n2005) );
  INVX8 U2598 ( .A(buff_data[376]), .Y(n2007) );
  INVX8 U2599 ( .A(n558), .Y(net79605) );
  INVX8 U2600 ( .A(buff_data[328]), .Y(n2009) );
  MUX2X1 U2601 ( .B(n2012), .A(n2011), .S(n178), .Y(n2010) );
  INVX8 U2602 ( .A(buff_data[295]), .Y(n2011) );
  INVX8 U2603 ( .A(n578), .Y(n2012) );
  INVX1 U2604 ( .A(n387), .Y(net80872) );
  INVX1 U2605 ( .A(n341), .Y(net80862) );
  INVX1 U2606 ( .A(n1836), .Y(n2013) );
  INVX1 U2607 ( .A(n1912), .Y(n2014) );
  AND2X2 U2608 ( .A(n320), .B(n3963), .Y(n2015) );
  INVX1 U2609 ( .A(n371), .Y(n2016) );
  INVX1 U2610 ( .A(net79533), .Y(net80723) );
  INVX8 U2611 ( .A(buff_data[315]), .Y(n2018) );
  MUX2X1 U2612 ( .B(n2021), .A(n2020), .S(n419), .Y(n2019) );
  INVX8 U2613 ( .A(buff_data[311]), .Y(n2020) );
  INVX8 U2614 ( .A(n578), .Y(n2021) );
  INVX8 U2615 ( .A(buff_data[358]), .Y(n2024) );
  INVX8 U2616 ( .A(buff_data[163]), .Y(n2026) );
  INVX1 U2617 ( .A(n561), .Y(net80781) );
  INVX1 U2618 ( .A(n3), .Y(net80747) );
  INVX1 U2619 ( .A(n103), .Y(net80382) );
  MUX2X1 U2620 ( .B(net80736), .A(n2032), .S(n334), .Y(n2031) );
  INVX8 U2621 ( .A(buff_data[237]), .Y(n2032) );
  INVX8 U2622 ( .A(n579), .Y(net80736) );
  INVX8 U2623 ( .A(buff_data[232]), .Y(n2034) );
  INVX1 U2624 ( .A(net79533), .Y(net79534) );
  INVX1 U2625 ( .A(n1837), .Y(n2038) );
  INVX1 U2626 ( .A(n216), .Y(n2039) );
  INVX1 U2627 ( .A(net79541), .Y(net80661) );
  MUX2X1 U2628 ( .B(n2044), .A(n2043), .S(n328), .Y(n2042) );
  INVX8 U2629 ( .A(buff_data[236]), .Y(n2043) );
  INVX8 U2630 ( .A(n572), .Y(n2044) );
  MUX2X1 U2631 ( .B(n2047), .A(n2046), .S(n335), .Y(n2045) );
  INVX8 U2632 ( .A(buff_data[231]), .Y(n2046) );
  INVX8 U2633 ( .A(n578), .Y(n2047) );
  INVX8 U2634 ( .A(n3990), .Y(n3087) );
  INVX1 U2635 ( .A(net92867), .Y(net80596) );
  INVX1 U2636 ( .A(net80595), .Y(net80598) );
  INVX8 U2637 ( .A(buff_data[198]), .Y(n2051) );
  INVX8 U2638 ( .A(buff_data[230]), .Y(n2055) );
  MUX2X1 U2639 ( .B(net80561), .A(n2057), .S(n384), .Y(n2056) );
  INVX8 U2640 ( .A(buff_data[196]), .Y(n2057) );
  INVX8 U2641 ( .A(n576), .Y(net80561) );
  MUX2X1 U2642 ( .B(n2060), .A(n2059), .S(n462), .Y(n2058) );
  INVX8 U2643 ( .A(buff_data[422]), .Y(n2059) );
  INVX8 U2644 ( .A(n570), .Y(n2060) );
  INVX8 U2645 ( .A(buff_data[229]), .Y(n2062) );
  INVX8 U2646 ( .A(buff_data[197]), .Y(n2064) );
  INVX1 U2647 ( .A(n538), .Y(net80518) );
  INVX1 U2648 ( .A(net92933), .Y(net80519) );
  INVX8 U2649 ( .A(buff_data[235]), .Y(n2066) );
  INVX8 U2650 ( .A(buff_data[203]), .Y(n2068) );
  INVX8 U2651 ( .A(buff_data[170]), .Y(n2070) );
  INVX8 U2652 ( .A(buff_data[154]), .Y(n2072) );
  INVX1 U2653 ( .A(n1802), .Y(n2074) );
  INVX1 U2654 ( .A(n103), .Y(net80463) );
  INVX1 U2655 ( .A(n207), .Y(n2076) );
  MUX2X1 U2656 ( .B(net80435), .A(n2080), .S(n552), .Y(n2079) );
  INVX8 U2657 ( .A(buff_data[20]), .Y(n2080) );
  INVX8 U2658 ( .A(n576), .Y(net80435) );
  MUX2X1 U2659 ( .B(n2115), .A(n2114), .S(n344), .Y(n2113) );
  INVX8 U2660 ( .A(n2113), .Y(n2168) );
  INVX8 U2661 ( .A(n2170), .Y(n2114) );
  INVX8 U2662 ( .A(n2169), .Y(n2115) );
  INVX8 U2663 ( .A(buff_data[499]), .Y(n2119) );
  INVX8 U2664 ( .A(n562), .Y(net79514) );
  INVX8 U2665 ( .A(buff_data[484]), .Y(n2121) );
  INVX8 U2666 ( .A(buff_data[467]), .Y(n2123) );
  INVX8 U2667 ( .A(buff_data[402]), .Y(n2125) );
  AND2X2 U2668 ( .A(net80519), .B(n4056), .Y(n2129) );
  MUX2X1 U2669 ( .B(n2132), .A(n2131), .S(net80839), .Y(n2130) );
  INVX8 U2670 ( .A(buff_data[368]), .Y(n2131) );
  INVX8 U2671 ( .A(n573), .Y(n2132) );
  INVX8 U2672 ( .A(buff_data[323]), .Y(n2134) );
  INVX8 U2673 ( .A(buff_data[288]), .Y(n2136) );
  MUX2X1 U2674 ( .B(n2139), .A(n2138), .S(n2041), .Y(n2137) );
  INVX8 U2675 ( .A(buff_data[352]), .Y(n2138) );
  INVX8 U2676 ( .A(n573), .Y(n2139) );
  INVX8 U2677 ( .A(buff_data[284]), .Y(n2141) );
  MUX2X1 U2678 ( .B(n2144), .A(n2143), .S(n552), .Y(n2142) );
  INVX8 U2679 ( .A(buff_data[31]), .Y(n2143) );
  INVX8 U2680 ( .A(n575), .Y(n2144) );
  INVX8 U2681 ( .A(buff_data[186]), .Y(n2146) );
  INVX8 U2682 ( .A(buff_data[242]), .Y(n2148) );
  MUX2X1 U2683 ( .B(n2151), .A(n2150), .S(n94), .Y(n2149) );
  INVX8 U2684 ( .A(buff_data[145]), .Y(n2150) );
  INVX8 U2685 ( .A(n577), .Y(n2151) );
  INVX8 U2686 ( .A(buff_data[226]), .Y(n2153) );
  MUX2X1 U2687 ( .B(n2156), .A(n2155), .S(n9), .Y(n2154) );
  INVX8 U2688 ( .A(buff_data[193]), .Y(n2155) );
  INVX8 U2689 ( .A(n577), .Y(n2156) );
  MUX2X1 U2690 ( .B(n2159), .A(n2158), .S(n327), .Y(n2157) );
  INVX8 U2691 ( .A(buff_data[161]), .Y(n2158) );
  INVX8 U2692 ( .A(n577), .Y(n2159) );
  INVX8 U2693 ( .A(n4279), .Y(n2736) );
  INVX8 U2694 ( .A(n4277), .Y(n2738) );
  INVX8 U2695 ( .A(n4275), .Y(n2740) );
  INVX8 U2696 ( .A(n4273), .Y(n2742) );
  INVX8 U2697 ( .A(n4271), .Y(n2744) );
  INVX8 U2698 ( .A(n4280), .Y(n2735) );
  INVX8 U2699 ( .A(n4278), .Y(n2737) );
  INVX8 U2700 ( .A(n4276), .Y(n2739) );
  INVX8 U2701 ( .A(n4274), .Y(n2741) );
  INVX8 U2702 ( .A(n4272), .Y(n2743) );
  INVX8 U2703 ( .A(n4285), .Y(n2730) );
  INVX8 U2704 ( .A(n4284), .Y(n2731) );
  INVX8 U2705 ( .A(n4283), .Y(n2732) );
  INVX8 U2706 ( .A(n4282), .Y(n2733) );
  INVX8 U2707 ( .A(n4281), .Y(n2734) );
  INVX8 U2708 ( .A(n4286), .Y(n2729) );
  INVX8 U2709 ( .A(n4054), .Y(n3019) );
  INVX8 U2710 ( .A(n4052), .Y(n3022) );
  INVX8 U2711 ( .A(n4049), .Y(n3025) );
  INVX8 U2712 ( .A(n4047), .Y(n3028) );
  INVX8 U2713 ( .A(n4044), .Y(n3032) );
  MUX2X1 U2714 ( .B(n2164), .A(n575), .S(n287), .Y(n2163) );
  INVX8 U2715 ( .A(n2163), .Y(n2166) );
  INVX8 U2716 ( .A(n2167), .Y(n2164) );
  INVX8 U2717 ( .A(n4053), .Y(n3021) );
  INVX8 U2718 ( .A(n4050), .Y(n3024) );
  INVX8 U2719 ( .A(n4048), .Y(n3027) );
  INVX8 U2720 ( .A(n4045), .Y(n3031) );
  INVX8 U2721 ( .A(n4042), .Y(n3034) );
  INVX8 U2722 ( .A(n4055), .Y(n3018) );
  INVX8 U2723 ( .A(n4174), .Y(n2863) );
  INVX8 U2724 ( .A(n4173), .Y(n2864) );
  INVX8 U2725 ( .A(n4172), .Y(n2865) );
  INVX8 U2726 ( .A(n4171), .Y(n2866) );
  INVX8 U2727 ( .A(n4170), .Y(n2867) );
  INVX8 U2728 ( .A(n4169), .Y(n2868) );
  INVX8 U2729 ( .A(n4168), .Y(n2869) );
  INVX8 U2730 ( .A(n4167), .Y(n2870) );
  INVX8 U2731 ( .A(n4166), .Y(n2871) );
  INVX8 U2732 ( .A(n4164), .Y(n2872) );
  INVX8 U2733 ( .A(n4245), .Y(n2778) );
  INVX8 U2734 ( .A(n4244), .Y(n2779) );
  INVX8 U2735 ( .A(n4242), .Y(n2781) );
  INVX8 U2736 ( .A(n4241), .Y(n2782) );
  INVX8 U2737 ( .A(n4239), .Y(n2784) );
  INVX8 U2738 ( .A(n4238), .Y(n2785) );
  INVX8 U2739 ( .A(n4236), .Y(n2787) );
  INVX8 U2740 ( .A(n4235), .Y(n2788) );
  INVX8 U2741 ( .A(n4233), .Y(n2790) );
  INVX8 U2742 ( .A(n4232), .Y(n2791) );
  INVX8 U2743 ( .A(n4081), .Y(n2991) );
  INVX8 U2744 ( .A(n4080), .Y(n2992) );
  INVX8 U2745 ( .A(n4079), .Y(n2993) );
  INVX8 U2746 ( .A(n4078), .Y(n2994) );
  INVX8 U2747 ( .A(n4077), .Y(n2995) );
  INVX8 U2748 ( .A(n4076), .Y(n2996) );
  INVX8 U2749 ( .A(n4075), .Y(n2998) );
  INVX8 U2750 ( .A(n4074), .Y(n2999) );
  INVX8 U2751 ( .A(n4073), .Y(n3000) );
  INVX8 U2752 ( .A(n4072), .Y(n3001) );
  INVX8 U2753 ( .A(n4147), .Y(n2906) );
  INVX8 U2754 ( .A(n4146), .Y(n2907) );
  INVX8 U2755 ( .A(n4144), .Y(n2909) );
  INVX8 U2756 ( .A(n4143), .Y(n2910) );
  INVX8 U2757 ( .A(n4141), .Y(n2912) );
  INVX8 U2758 ( .A(n4140), .Y(n2913) );
  INVX8 U2759 ( .A(n4138), .Y(n2915) );
  INVX8 U2760 ( .A(n4137), .Y(n2916) );
  INVX8 U2761 ( .A(n4135), .Y(n2918) );
  INVX8 U2762 ( .A(n4134), .Y(n2919) );
  INVX8 U2763 ( .A(n4179), .Y(n2858) );
  INVX8 U2764 ( .A(n4178), .Y(n2859) );
  INVX8 U2765 ( .A(n4177), .Y(n2860) );
  INVX8 U2766 ( .A(n4176), .Y(n2861) );
  INVX8 U2767 ( .A(n4175), .Y(n2862) );
  INVX8 U2768 ( .A(n4243), .Y(n2780) );
  INVX8 U2769 ( .A(n4240), .Y(n2783) );
  INVX8 U2770 ( .A(n4237), .Y(n2786) );
  INVX8 U2771 ( .A(n4234), .Y(n2789) );
  INVX8 U2772 ( .A(n4230), .Y(n2792) );
  INVX8 U2773 ( .A(n4246), .Y(n2777) );
  INVX8 U2774 ( .A(n4180), .Y(n2857) );
  INVX8 U2775 ( .A(n4310), .Y(n2699) );
  INVX8 U2776 ( .A(n4309), .Y(n2700) );
  INVX8 U2777 ( .A(n4308), .Y(n2701) );
  INVX8 U2778 ( .A(n4307), .Y(n2702) );
  INVX8 U2779 ( .A(n4306), .Y(n2703) );
  INVX8 U2780 ( .A(n4305), .Y(n2705) );
  INVX8 U2781 ( .A(n4304), .Y(n2707) );
  INVX8 U2782 ( .A(n4303), .Y(n2708) );
  INVX8 U2783 ( .A(n4302), .Y(n2709) );
  INVX8 U2784 ( .A(n4301), .Y(n2710) );
  INVX8 U2785 ( .A(n4300), .Y(n2711) );
  INVX8 U2786 ( .A(n4311), .Y(n2697) );
  INVX8 U2787 ( .A(n4086), .Y(n2986) );
  INVX8 U2788 ( .A(n4085), .Y(n2987) );
  INVX8 U2789 ( .A(n4084), .Y(n2988) );
  INVX8 U2790 ( .A(n4083), .Y(n2989) );
  INVX8 U2791 ( .A(n4082), .Y(n2990) );
  INVX8 U2792 ( .A(n4145), .Y(n2908) );
  INVX8 U2793 ( .A(n4142), .Y(n2911) );
  INVX8 U2794 ( .A(n4139), .Y(n2914) );
  INVX8 U2795 ( .A(n4136), .Y(n2917) );
  INVX8 U2796 ( .A(n4148), .Y(n2905) );
  INVX8 U2797 ( .A(n4087), .Y(n2985) );
  INVX8 U2798 ( .A(n4341), .Y(n2666) );
  INVX8 U2799 ( .A(n4340), .Y(n2667) );
  INVX8 U2800 ( .A(n4339), .Y(n2668) );
  INVX8 U2801 ( .A(n4338), .Y(n2669) );
  INVX8 U2802 ( .A(n4337), .Y(n2670) );
  INVX8 U2803 ( .A(n4336), .Y(n2672) );
  INVX8 U2804 ( .A(n4335), .Y(n2673) );
  INVX8 U2805 ( .A(n4334), .Y(n2674) );
  INVX8 U2806 ( .A(n4333), .Y(n2675) );
  INVX8 U2807 ( .A(n4332), .Y(n2676) );
  INVX8 U2808 ( .A(n4331), .Y(n2677) );
  INVX8 U2809 ( .A(n4330), .Y(n2678) );
  INVX8 U2810 ( .A(n4329), .Y(n2679) );
  INVX8 U2811 ( .A(n4328), .Y(n2680) );
  INVX8 U2812 ( .A(n4342), .Y(n2665) );
  INVX8 U2813 ( .A(n4326), .Y(n2682) );
  INVX8 U2814 ( .A(n4325), .Y(n2683) );
  INVX8 U2815 ( .A(n4324), .Y(n2684) );
  INVX8 U2816 ( .A(n4323), .Y(n2685) );
  INVX8 U2817 ( .A(n4322), .Y(n2686) );
  INVX8 U2818 ( .A(n4321), .Y(n2687) );
  INVX8 U2819 ( .A(n4320), .Y(n2688) );
  INVX8 U2820 ( .A(n4319), .Y(n2689) );
  INVX8 U2821 ( .A(n4318), .Y(n2690) );
  INVX8 U2822 ( .A(n4317), .Y(n2691) );
  INVX8 U2823 ( .A(n4316), .Y(n2692) );
  INVX8 U2824 ( .A(n4315), .Y(n2693) );
  INVX8 U2825 ( .A(n4314), .Y(n2694) );
  INVX8 U2826 ( .A(n4313), .Y(n2695) );
  INVX8 U2827 ( .A(n4312), .Y(n2696) );
  INVX8 U2828 ( .A(n4327), .Y(n2681) );
  INVX8 U2829 ( .A(n4298), .Y(n2715) );
  INVX8 U2830 ( .A(n4297), .Y(n2716) );
  INVX8 U2831 ( .A(n4296), .Y(n2717) );
  INVX8 U2832 ( .A(n4295), .Y(n2718) );
  INVX8 U2833 ( .A(n4294), .Y(n2719) );
  INVX8 U2834 ( .A(n4293), .Y(n2720) );
  INVX8 U2835 ( .A(n4292), .Y(n2721) );
  INVX8 U2836 ( .A(n4291), .Y(n2722) );
  INVX8 U2837 ( .A(n4290), .Y(n2724) );
  INVX8 U2838 ( .A(n4289), .Y(n2725) );
  INVX8 U2839 ( .A(n4288), .Y(n2727) );
  INVX8 U2840 ( .A(n4287), .Y(n2728) );
  INVX8 U2841 ( .A(n4299), .Y(n2713) );
  INVX8 U2842 ( .A(n4384), .Y(n2618) );
  INVX8 U2843 ( .A(n4383), .Y(n2619) );
  INVX8 U2844 ( .A(n4382), .Y(n2620) );
  INVX8 U2845 ( .A(n4381), .Y(n2621) );
  INVX8 U2846 ( .A(n4380), .Y(n2622) );
  INVX8 U2847 ( .A(n4379), .Y(n2623) );
  INVX8 U2848 ( .A(n4378), .Y(n2624) );
  INVX8 U2849 ( .A(n4377), .Y(n2625) );
  INVX8 U2850 ( .A(n4376), .Y(n2626) );
  INVX8 U2851 ( .A(n4375), .Y(n2627) );
  INVX8 U2852 ( .A(n4374), .Y(n2628) );
  INVX8 U2853 ( .A(n4373), .Y(n2630) );
  INVX8 U2854 ( .A(n4372), .Y(n2631) );
  INVX8 U2855 ( .A(n4371), .Y(n2632) );
  INVX8 U2856 ( .A(n4385), .Y(n2617) );
  INVX8 U2857 ( .A(n4025), .Y(n3053) );
  INVX8 U2858 ( .A(n4024), .Y(n3054) );
  INVX8 U2859 ( .A(n4023), .Y(n3055) );
  INVX8 U2860 ( .A(n4022), .Y(n3056) );
  INVX8 U2861 ( .A(n4021), .Y(n3057) );
  INVX8 U2862 ( .A(n4020), .Y(n3058) );
  INVX8 U2863 ( .A(n4019), .Y(n3059) );
  INVX8 U2864 ( .A(n4018), .Y(n3060) );
  INVX8 U2865 ( .A(n4017), .Y(n3061) );
  INVX8 U2866 ( .A(n4016), .Y(n3063) );
  INVX8 U2867 ( .A(n4015), .Y(n3064) );
  INVX8 U2868 ( .A(n4014), .Y(n3065) );
  INVX8 U2869 ( .A(n4013), .Y(n3066) );
  INVX8 U2870 ( .A(n4012), .Y(n3067) );
  INVX8 U2871 ( .A(n3989), .Y(n3088) );
  INVX8 U2872 ( .A(n3988), .Y(n3089) );
  INVX8 U2873 ( .A(n3987), .Y(n3090) );
  INVX8 U2874 ( .A(n3986), .Y(n3091) );
  INVX8 U2875 ( .A(n3985), .Y(n3092) );
  INVX8 U2876 ( .A(n3984), .Y(n3093) );
  INVX8 U2877 ( .A(n3983), .Y(n3094) );
  INVX8 U2878 ( .A(n3982), .Y(n3095) );
  INVX8 U2879 ( .A(n3981), .Y(n3096) );
  INVX8 U2880 ( .A(n3980), .Y(n3097) );
  INVX8 U2881 ( .A(n3979), .Y(n3098) );
  INVX8 U2882 ( .A(n3978), .Y(n3099) );
  INVX8 U2883 ( .A(n3977), .Y(n3100) );
  INVX8 U2884 ( .A(n3976), .Y(n3101) );
  INVX8 U2885 ( .A(n3975), .Y(n3102) );
  INVX8 U2886 ( .A(n3974), .Y(n3104) );
  INVX8 U2887 ( .A(n3973), .Y(n3106) );
  INVX8 U2888 ( .A(n3972), .Y(n3107) );
  INVX8 U2889 ( .A(n3971), .Y(n3108) );
  INVX8 U2890 ( .A(n3970), .Y(n3110) );
  INVX8 U2891 ( .A(n3969), .Y(n3111) );
  INVX8 U2892 ( .A(n3968), .Y(n3112) );
  INVX8 U2893 ( .A(n3967), .Y(n3113) );
  INVX8 U2894 ( .A(n3966), .Y(n3115) );
  INVX8 U2895 ( .A(n3965), .Y(n3117) );
  INVX8 U2896 ( .A(n3964), .Y(n3118) );
  INVX8 U2897 ( .A(n4370), .Y(n2633) );
  INVX8 U2898 ( .A(n4369), .Y(n2634) );
  INVX8 U2899 ( .A(n4368), .Y(n2635) );
  INVX8 U2900 ( .A(n4367), .Y(n2636) );
  INVX8 U2901 ( .A(n4366), .Y(n2637) );
  INVX8 U2902 ( .A(n4365), .Y(n2638) );
  INVX8 U2903 ( .A(n4364), .Y(n2639) );
  INVX8 U2904 ( .A(n4363), .Y(n2640) );
  INVX8 U2905 ( .A(n4362), .Y(n2641) );
  INVX8 U2906 ( .A(n4361), .Y(n2642) );
  INVX8 U2907 ( .A(n4360), .Y(n2643) );
  INVX8 U2908 ( .A(n4359), .Y(n2644) );
  INVX8 U2909 ( .A(n4358), .Y(n2645) );
  INVX8 U2910 ( .A(n4357), .Y(n2647) );
  INVX8 U2911 ( .A(n4355), .Y(n2648) );
  INVX8 U2912 ( .A(n4354), .Y(n2649) );
  INVX8 U2913 ( .A(n4353), .Y(n2650) );
  INVX8 U2914 ( .A(n4352), .Y(n2651) );
  INVX8 U2915 ( .A(n4351), .Y(n2653) );
  INVX8 U2916 ( .A(n4350), .Y(n2654) );
  INVX8 U2917 ( .A(n4349), .Y(n2656) );
  INVX8 U2918 ( .A(n4348), .Y(n2657) );
  INVX8 U2919 ( .A(n4347), .Y(n2658) );
  INVX8 U2920 ( .A(n4346), .Y(n2659) );
  INVX8 U2921 ( .A(n4345), .Y(n2662) );
  INVX8 U2922 ( .A(n4344), .Y(n2663) );
  INVX8 U2923 ( .A(n4343), .Y(n2664) );
  INVX8 U2924 ( .A(n4071), .Y(n3003) );
  INVX8 U2925 ( .A(n4070), .Y(n3004) );
  INVX8 U2926 ( .A(n4069), .Y(n3005) );
  INVX8 U2927 ( .A(n4068), .Y(n3006) );
  INVX8 U2928 ( .A(n4067), .Y(n3007) );
  INVX8 U2929 ( .A(n4066), .Y(n3008) );
  INVX8 U2930 ( .A(n4065), .Y(n3009) );
  INVX8 U2931 ( .A(n4064), .Y(n3010) );
  INVX8 U2932 ( .A(n4063), .Y(n3011) );
  INVX8 U2933 ( .A(n4062), .Y(n3012) );
  INVX8 U2934 ( .A(n4061), .Y(n3013) );
  INVX8 U2935 ( .A(n4060), .Y(n3014) );
  INVX8 U2936 ( .A(n4059), .Y(n3015) );
  INVX8 U2937 ( .A(n4058), .Y(n3016) );
  INVX8 U2938 ( .A(n4057), .Y(n3017) );
  INVX8 U2939 ( .A(buff_data[127]), .Y(n2167) );
  INVX1 U2940 ( .A(n575), .Y(n2170) );
  INVX8 U2941 ( .A(buff_data[63]), .Y(n2169) );
  INVX8 U2942 ( .A(n4010), .Y(n3069) );
  INVX8 U2943 ( .A(n4009), .Y(n3070) );
  INVX8 U2944 ( .A(n4008), .Y(n3071) );
  INVX8 U2945 ( .A(n4007), .Y(n3072) );
  INVX8 U2946 ( .A(n4005), .Y(n3075) );
  INVX8 U2947 ( .A(n4004), .Y(n3076) );
  INVX8 U2948 ( .A(n4003), .Y(n3077) );
  INVX8 U2949 ( .A(n4002), .Y(n3078) );
  INVX8 U2950 ( .A(n3997), .Y(n3080) );
  INVX8 U2951 ( .A(n3996), .Y(n3081) );
  INVX8 U2952 ( .A(n3995), .Y(n3082) );
  INVX8 U2953 ( .A(n3994), .Y(n3083) );
  INVX8 U2954 ( .A(n3993), .Y(n3084) );
  INVX8 U2955 ( .A(n3992), .Y(n3085) );
  INVX8 U2956 ( .A(n3991), .Y(n3086) );
  INVX8 U2957 ( .A(buff_data[85]), .Y(n2172) );
  INVX8 U2958 ( .A(n4040), .Y(n3037) );
  INVX8 U2959 ( .A(n4039), .Y(n3038) );
  INVX8 U2960 ( .A(n4038), .Y(n3039) );
  INVX8 U2961 ( .A(n4037), .Y(n3040) );
  INVX8 U2962 ( .A(n4036), .Y(n3041) );
  INVX8 U2963 ( .A(n4035), .Y(n3042) );
  INVX8 U2964 ( .A(n4034), .Y(n3043) );
  INVX8 U2965 ( .A(n4033), .Y(n3044) );
  INVX8 U2966 ( .A(n4032), .Y(n3045) );
  INVX8 U2967 ( .A(n4031), .Y(n3046) );
  INVX8 U2968 ( .A(n4030), .Y(n3047) );
  INVX8 U2969 ( .A(n4029), .Y(n3048) );
  INVX8 U2970 ( .A(n4028), .Y(n3049) );
  INVX8 U2971 ( .A(n4027), .Y(n3050) );
  INVX8 U2972 ( .A(n4026), .Y(n3051) );
  INVX8 U2973 ( .A(buff_data[15]), .Y(n2174) );
  INVX8 U2974 ( .A(n3962), .Y(n3121) );
  INVX8 U2975 ( .A(n3961), .Y(n3122) );
  INVX8 U2976 ( .A(n3960), .Y(n3123) );
  INVX8 U2977 ( .A(n3959), .Y(n3124) );
  INVX8 U2978 ( .A(n3958), .Y(n3128) );
  INVX8 U2979 ( .A(n3957), .Y(n3129) );
  INVX8 U2980 ( .A(n3956), .Y(n3130) );
  INVX8 U2981 ( .A(n3955), .Y(n3131) );
  INVX8 U2982 ( .A(n3954), .Y(n3132) );
  INVX8 U2983 ( .A(n3953), .Y(n3134) );
  INVX8 U2984 ( .A(n3952), .Y(n3135) );
  INVX8 U2985 ( .A(n3951), .Y(n3136) );
  INVX8 U2986 ( .A(n3950), .Y(n3137) );
  INVX8 U2987 ( .A(n4123), .Y(n2937) );
  INVX8 U2988 ( .A(n4122), .Y(n2938) );
  INVX8 U2989 ( .A(n4121), .Y(n2939) );
  INVX8 U2990 ( .A(n4120), .Y(n2940) );
  INVX8 U2991 ( .A(n4119), .Y(n2941) );
  INVX8 U2992 ( .A(n4118), .Y(n2942) );
  INVX8 U2993 ( .A(n4117), .Y(n2946) );
  INVX8 U2994 ( .A(n4116), .Y(n2947) );
  INVX8 U2995 ( .A(n4115), .Y(n2948) );
  INVX8 U2996 ( .A(n4114), .Y(n2949) );
  INVX8 U2997 ( .A(n4113), .Y(n2950) );
  INVX8 U2998 ( .A(n4112), .Y(n2952) );
  INVX8 U2999 ( .A(n4259), .Y(n2761) );
  INVX8 U3000 ( .A(n4258), .Y(n2763) );
  INVX8 U3001 ( .A(n4257), .Y(n2764) );
  INVX8 U3002 ( .A(n4256), .Y(n2765) );
  INVX8 U3003 ( .A(n4255), .Y(n2766) );
  INVX8 U3004 ( .A(n4254), .Y(n2767) );
  INVX8 U3005 ( .A(n4253), .Y(n2768) );
  INVX8 U3006 ( .A(n4252), .Y(n2769) );
  INVX8 U3007 ( .A(n4251), .Y(n2771) );
  INVX8 U3008 ( .A(n4250), .Y(n2772) );
  INVX8 U3009 ( .A(n4249), .Y(n2773) );
  INVX8 U3010 ( .A(n4248), .Y(n2774) );
  INVX8 U3011 ( .A(n4247), .Y(n2775) );
  INVX8 U3012 ( .A(n4229), .Y(n2793) );
  INVX8 U3013 ( .A(n4228), .Y(n2794) );
  INVX8 U3014 ( .A(n4227), .Y(n2796) );
  INVX8 U3015 ( .A(n4226), .Y(n2798) );
  INVX8 U3016 ( .A(n4225), .Y(n2799) );
  INVX8 U3017 ( .A(n4224), .Y(n2801) );
  INVX8 U3018 ( .A(n4223), .Y(n2802) );
  INVX8 U3019 ( .A(n4222), .Y(n2803) );
  INVX8 U3020 ( .A(n4221), .Y(n2804) );
  INVX8 U3021 ( .A(n4220), .Y(n2806) );
  INVX8 U3022 ( .A(n4219), .Y(n2807) );
  INVX8 U3023 ( .A(n4217), .Y(n2808) );
  INVX8 U3024 ( .A(n4203), .Y(n2825) );
  INVX8 U3025 ( .A(n4202), .Y(n2826) );
  INVX8 U3026 ( .A(n4201), .Y(n2828) );
  INVX8 U3027 ( .A(n4200), .Y(n2829) );
  INVX8 U3028 ( .A(n4199), .Y(n2830) );
  INVX8 U3029 ( .A(n4198), .Y(n2831) );
  INVX8 U3030 ( .A(n4197), .Y(n2832) );
  INVX8 U3031 ( .A(n4196), .Y(n2834) );
  INVX8 U3032 ( .A(n4195), .Y(n2835) );
  INVX8 U3033 ( .A(n4194), .Y(n2836) );
  INVX8 U3034 ( .A(n4193), .Y(n2837) );
  INVX8 U3035 ( .A(n4192), .Y(n2838) );
  INVX8 U3036 ( .A(n4191), .Y(n2839) );
  INVX8 U3037 ( .A(n4270), .Y(n2745) );
  INVX8 U3038 ( .A(n4269), .Y(n2746) );
  INVX8 U3039 ( .A(n4268), .Y(n2747) );
  INVX8 U3040 ( .A(n4267), .Y(n2749) );
  INVX8 U3041 ( .A(n4266), .Y(n2752) );
  INVX8 U3042 ( .A(n4265), .Y(n2753) );
  INVX8 U3043 ( .A(n4264), .Y(n2754) );
  INVX8 U3044 ( .A(n4263), .Y(n2756) );
  INVX8 U3045 ( .A(n4262), .Y(n2757) );
  INVX8 U3046 ( .A(n4261), .Y(n2758) );
  INVX8 U3047 ( .A(n4260), .Y(n2760) );
  INVX8 U3048 ( .A(n4190), .Y(n2841) );
  INVX8 U3049 ( .A(n4189), .Y(n2842) );
  INVX8 U3050 ( .A(n4188), .Y(n2843) );
  INVX8 U3051 ( .A(n4187), .Y(n2847) );
  INVX8 U3052 ( .A(n4186), .Y(n2849) );
  INVX8 U3053 ( .A(n4185), .Y(n2850) );
  INVX8 U3054 ( .A(n4184), .Y(n2851) );
  INVX8 U3055 ( .A(n4183), .Y(n2852) );
  INVX8 U3056 ( .A(n4182), .Y(n2854) );
  INVX8 U3057 ( .A(n4181), .Y(n2855) );
  MUX2X1 U3058 ( .B(n2177), .A(n2176), .S(n418), .Y(n2175) );
  INVX8 U3059 ( .A(buff_data[319]), .Y(n2176) );
  INVX8 U3060 ( .A(n575), .Y(n2177) );
  INVX8 U3061 ( .A(n4216), .Y(n2810) );
  INVX8 U3062 ( .A(n4215), .Y(n2811) );
  INVX8 U3063 ( .A(n4214), .Y(n2814) );
  INVX8 U3064 ( .A(n4213), .Y(n2815) );
  INVX8 U3065 ( .A(n4212), .Y(n2816) );
  INVX8 U3066 ( .A(n4211), .Y(n2818) );
  INVX8 U3067 ( .A(n4210), .Y(n2819) );
  INVX8 U3068 ( .A(n4209), .Y(n2820) );
  INVX8 U3069 ( .A(n4208), .Y(n2821) );
  INVX8 U3070 ( .A(n4207), .Y(n2822) );
  INVX8 U3071 ( .A(n4206), .Y(n2823) );
  INVX8 U3072 ( .A(n4204), .Y(n2824) );
  INVX8 U3073 ( .A(n4152), .Y(n2889) );
  INVX8 U3074 ( .A(n4151), .Y(n2900) );
  INVX8 U3075 ( .A(n4150), .Y(n2901) );
  INVX8 U3076 ( .A(n4149), .Y(n2904) );
  INVX8 U3077 ( .A(n4131), .Y(n2921) );
  INVX8 U3078 ( .A(n4130), .Y(n2923) );
  INVX8 U3079 ( .A(n4129), .Y(n2924) );
  INVX8 U3080 ( .A(n4128), .Y(n2926) );
  INVX8 U3081 ( .A(n4127), .Y(n2927) );
  INVX8 U3082 ( .A(n4126), .Y(n2928) );
  INVX8 U3083 ( .A(n4125), .Y(n2934) );
  INVX8 U3084 ( .A(n4124), .Y(n2936) );
  INVX8 U3085 ( .A(n4111), .Y(n2953) );
  INVX8 U3086 ( .A(n4110), .Y(n2954) );
  INVX8 U3087 ( .A(n4109), .Y(n2957) );
  INVX8 U3088 ( .A(n4108), .Y(n2959) );
  INVX8 U3089 ( .A(n4107), .Y(n2961) );
  INVX8 U3090 ( .A(n4106), .Y(n2962) );
  INVX8 U3091 ( .A(n4105), .Y(n2963) );
  INVX8 U3092 ( .A(n4104), .Y(n2964) );
  INVX8 U3093 ( .A(n4103), .Y(n2966) );
  INVX8 U3094 ( .A(n4102), .Y(n2968) );
  INVX8 U3095 ( .A(n4163), .Y(n2874) );
  INVX8 U3096 ( .A(n4162), .Y(n2876) );
  INVX8 U3097 ( .A(n4161), .Y(n2877) );
  INVX8 U3098 ( .A(n4160), .Y(n2879) );
  INVX8 U3099 ( .A(n4159), .Y(n2880) );
  INVX8 U3100 ( .A(n4158), .Y(n2881) );
  INVX8 U3101 ( .A(n4157), .Y(n2882) );
  INVX8 U3102 ( .A(n4156), .Y(n2883) );
  INVX8 U3103 ( .A(n4155), .Y(n2885) );
  INVX8 U3104 ( .A(n4154), .Y(n2887) );
  INVX8 U3105 ( .A(n4153), .Y(n2888) );
  INVX8 U3106 ( .A(n4101), .Y(n2969) );
  INVX8 U3107 ( .A(n4100), .Y(n2970) );
  INVX8 U3108 ( .A(n4099), .Y(n2971) );
  INVX8 U3109 ( .A(n4098), .Y(n2972) );
  INVX8 U3110 ( .A(n4097), .Y(n2973) );
  INVX8 U3111 ( .A(n4096), .Y(n2975) );
  INVX8 U3112 ( .A(n4095), .Y(n2976) );
  INVX8 U3113 ( .A(n4094), .Y(n2977) );
  INVX8 U3114 ( .A(n4093), .Y(n2978) );
  INVX8 U3115 ( .A(n4092), .Y(n2979) );
  INVX8 U3116 ( .A(n4091), .Y(n2980) );
  INVX8 U3117 ( .A(n4090), .Y(n2981) );
  INVX8 U3118 ( .A(n4089), .Y(n2982) );
  INVX8 U3119 ( .A(n4088), .Y(n2984) );
  INVX8 U3120 ( .A(n559), .Y(n2180) );
  AND2X2 U3121 ( .A(n82), .B(net66503), .Y(n2182) );
  AND2X2 U3122 ( .A(net66503), .B(net82138), .Y(n2183) );
  AND2X2 U3123 ( .A(net80872), .B(net66503), .Y(n2186) );
  AND2X2 U3124 ( .A(net80872), .B(net66503), .Y(n2187) );
  NAND3X1 U3125 ( .A(n1729), .B(n1735), .C(n3777), .Y(n2188) );
  AND2X2 U3126 ( .A(n541), .B(n3778), .Y(n3777) );
  AND2X2 U3127 ( .A(net80862), .B(n3963), .Y(n2189) );
  AND2X2 U3128 ( .A(net80862), .B(n3963), .Y(n2190) );
  AND2X2 U3129 ( .A(net82472), .B(n3963), .Y(n4165) );
  AND2X2 U3130 ( .A(n547), .B(net66482), .Y(n4218) );
  AND2X2 U3131 ( .A(net66503), .B(net80598), .Y(n4133) );
  INVX8 U3132 ( .A(n4132), .Y(n2920) );
  INVX1 U3133 ( .A(n542), .Y(net79482) );
  AND2X2 U3134 ( .A(n547), .B(n4011), .Y(n4205) );
  AND2X2 U3135 ( .A(n82), .B(net66503), .Y(n4231) );
  INVX8 U3136 ( .A(net79440), .Y(net79428) );
  INVX8 U3137 ( .A(net79440), .Y(net79430) );
  INVX8 U3138 ( .A(net79420), .Y(net79408) );
  INVX8 U3139 ( .A(net79420), .Y(net79410) );
  INVX8 U3140 ( .A(net79420), .Y(net79412) );
  MUX2X1 U3141 ( .B(n2202), .A(n2203), .S(net79430), .Y(n2201) );
  MUX2X1 U3142 ( .B(n2205), .A(n2206), .S(net79430), .Y(n2204) );
  MUX2X1 U3143 ( .B(n2208), .A(n2209), .S(net79430), .Y(n2207) );
  MUX2X1 U3144 ( .B(n2211), .A(n2212), .S(net79430), .Y(n2210) );
  MUX2X1 U3145 ( .B(n2214), .A(n2215), .S(n231), .Y(n2213) );
  MUX2X1 U3146 ( .B(n2217), .A(n2218), .S(net79430), .Y(n2216) );
  MUX2X1 U3147 ( .B(n2220), .A(n2221), .S(net79430), .Y(n2219) );
  MUX2X1 U3148 ( .B(n2223), .A(n2224), .S(net79430), .Y(n2222) );
  MUX2X1 U3149 ( .B(n2226), .A(n2227), .S(net79430), .Y(n2225) );
  MUX2X1 U3150 ( .B(n2229), .A(n2230), .S(n231), .Y(n2228) );
  MUX2X1 U3151 ( .B(n2232), .A(n2233), .S(net79430), .Y(n2231) );
  MUX2X1 U3152 ( .B(n2235), .A(n2236), .S(net79430), .Y(n2234) );
  MUX2X1 U3153 ( .B(n2238), .A(n2239), .S(net79430), .Y(n2237) );
  MUX2X1 U3154 ( .B(n2241), .A(n2242), .S(net79430), .Y(n2240) );
  MUX2X1 U3155 ( .B(n2244), .A(n2245), .S(n231), .Y(n2243) );
  MUX2X1 U3156 ( .B(n2247), .A(n2248), .S(net79430), .Y(n2246) );
  MUX2X1 U3157 ( .B(n2250), .A(n2251), .S(net79430), .Y(n2249) );
  MUX2X1 U3158 ( .B(n2253), .A(n2254), .S(net79430), .Y(n2252) );
  MUX2X1 U3159 ( .B(n2256), .A(n2257), .S(net79430), .Y(n2255) );
  MUX2X1 U3160 ( .B(n2259), .A(n2260), .S(n231), .Y(n2258) );
  MUX2X1 U3161 ( .B(n2262), .A(n2263), .S(net79430), .Y(n2261) );
  MUX2X1 U3162 ( .B(n2265), .A(n2266), .S(net79430), .Y(n2264) );
  MUX2X1 U3163 ( .B(n2268), .A(n2269), .S(net79430), .Y(n2267) );
  MUX2X1 U3164 ( .B(n2271), .A(n2272), .S(net79430), .Y(n2270) );
  MUX2X1 U3165 ( .B(n2274), .A(n2275), .S(n231), .Y(n2273) );
  MUX2X1 U3166 ( .B(n2277), .A(n2278), .S(net79430), .Y(n2276) );
  MUX2X1 U3167 ( .B(n2280), .A(n2281), .S(net79430), .Y(n2279) );
  MUX2X1 U3168 ( .B(n2283), .A(n2284), .S(net79430), .Y(n2282) );
  MUX2X1 U3169 ( .B(n2286), .A(n2287), .S(net79430), .Y(n2285) );
  MUX2X1 U3170 ( .B(n2289), .A(n2290), .S(n231), .Y(n2288) );
  MUX2X1 U3171 ( .B(n2292), .A(n2293), .S(net79430), .Y(n2291) );
  MUX2X1 U3172 ( .B(n2295), .A(n2296), .S(net79430), .Y(n2294) );
  MUX2X1 U3173 ( .B(n2298), .A(n2299), .S(net79430), .Y(n2297) );
  MUX2X1 U3174 ( .B(n2301), .A(n2302), .S(net79430), .Y(n2300) );
  MUX2X1 U3175 ( .B(n2304), .A(n2305), .S(n231), .Y(n2303) );
  MUX2X1 U3176 ( .B(n2307), .A(n2308), .S(net79430), .Y(n2306) );
  MUX2X1 U3177 ( .B(n2310), .A(n2311), .S(net79430), .Y(n2309) );
  MUX2X1 U3178 ( .B(n2313), .A(n2314), .S(net79430), .Y(n2312) );
  MUX2X1 U3179 ( .B(n2316), .A(n2317), .S(net79430), .Y(n2315) );
  MUX2X1 U3180 ( .B(n2319), .A(n2320), .S(n231), .Y(n2318) );
  MUX2X1 U3181 ( .B(n2322), .A(n2323), .S(net79430), .Y(n2321) );
  MUX2X1 U3182 ( .B(n2325), .A(n2326), .S(net79430), .Y(n2324) );
  MUX2X1 U3183 ( .B(n2328), .A(n2329), .S(net79430), .Y(n2327) );
  MUX2X1 U3184 ( .B(n2331), .A(n2332), .S(net79430), .Y(n2330) );
  MUX2X1 U3185 ( .B(n2334), .A(n2335), .S(n231), .Y(n2333) );
  MUX2X1 U3186 ( .B(n2337), .A(n2338), .S(net79430), .Y(n2336) );
  MUX2X1 U3187 ( .B(n2340), .A(n2341), .S(net79430), .Y(n2339) );
  MUX2X1 U3188 ( .B(n2343), .A(n2344), .S(net79430), .Y(n2342) );
  MUX2X1 U3189 ( .B(n2346), .A(C25909_net2624), .S(net79430), .Y(n2345) );
  MUX2X1 U3190 ( .B(n2348), .A(n2349), .S(n231), .Y(n2347) );
  MUX2X1 U3191 ( .B(n2351), .A(n2352), .S(net79430), .Y(n2350) );
  MUX2X1 U3192 ( .B(n2354), .A(n2355), .S(net79430), .Y(n2353) );
  MUX2X1 U3193 ( .B(n2357), .A(n2358), .S(net79430), .Y(n2356) );
  MUX2X1 U3194 ( .B(n2360), .A(n2361), .S(net79430), .Y(n2359) );
  MUX2X1 U3195 ( .B(n2363), .A(n2364), .S(n231), .Y(n2362) );
  MUX2X1 U3196 ( .B(n2366), .A(n2367), .S(net79430), .Y(n2365) );
  MUX2X1 U3197 ( .B(n2369), .A(n2370), .S(net79430), .Y(n2368) );
  MUX2X1 U3198 ( .B(n2372), .A(n2373), .S(net79430), .Y(n2371) );
  MUX2X1 U3199 ( .B(n2376), .A(n2377), .S(net79430), .Y(n2374) );
  MUX2X1 U3200 ( .B(n2409), .A(n2410), .S(n231), .Y(n2408) );
  MUX2X1 U3201 ( .B(n2412), .A(n2413), .S(net79430), .Y(n2411) );
  MUX2X1 U3202 ( .B(n2415), .A(n2416), .S(net79430), .Y(n2414) );
  MUX2X1 U3203 ( .B(n2418), .A(n2419), .S(net79430), .Y(n2417) );
  MUX2X1 U3204 ( .B(n2421), .A(n2422), .S(net79430), .Y(n2420) );
  MUX2X1 U3205 ( .B(n2424), .A(n2425), .S(n231), .Y(n2423) );
  MUX2X1 U3206 ( .B(n2427), .A(n2428), .S(net79430), .Y(n2426) );
  MUX2X1 U3207 ( .B(n2430), .A(n2431), .S(net79430), .Y(n2429) );
  MUX2X1 U3208 ( .B(n2433), .A(n2434), .S(net79432), .Y(n2432) );
  MUX2X1 U3209 ( .B(n2436), .A(n2437), .S(net79432), .Y(n2435) );
  MUX2X1 U3210 ( .B(n2440), .A(n2441), .S(n231), .Y(n2438) );
  MUX2X1 U3211 ( .B(n2444), .A(n2445), .S(net79432), .Y(n2443) );
  MUX2X1 U3212 ( .B(n2447), .A(n2448), .S(net79432), .Y(n2446) );
  MUX2X1 U3213 ( .B(n2450), .A(n2451), .S(net79432), .Y(n2449) );
  MUX2X1 U3214 ( .B(n2453), .A(n2454), .S(net79432), .Y(n2452) );
  MUX2X1 U3215 ( .B(n2456), .A(n2457), .S(n231), .Y(n2455) );
  MUX2X1 U3216 ( .B(n2459), .A(n2460), .S(net79432), .Y(n2458) );
  MUX2X1 U3217 ( .B(n2462), .A(n2463), .S(net79432), .Y(n2461) );
  MUX2X1 U3218 ( .B(n2465), .A(n2466), .S(net79432), .Y(n2464) );
  MUX2X1 U3219 ( .B(n2468), .A(n2469), .S(net79432), .Y(n2467) );
  MUX2X1 U3220 ( .B(n2471), .A(n2472), .S(n231), .Y(n2470) );
  MUX2X1 U3221 ( .B(n2474), .A(n2475), .S(net79432), .Y(n2473) );
  MUX2X1 U3222 ( .B(n2477), .A(n2478), .S(net79432), .Y(n2476) );
  MUX2X1 U3223 ( .B(n2480), .A(n2481), .S(net79432), .Y(n2479) );
  MUX2X1 U3224 ( .B(n2483), .A(n2484), .S(net79432), .Y(n2482) );
  MUX2X1 U3225 ( .B(n2486), .A(n2487), .S(n231), .Y(n2485) );
  MUX2X1 U3226 ( .B(n2489), .A(n2490), .S(net79432), .Y(n2488) );
  MUX2X1 U3227 ( .B(n2492), .A(n2493), .S(net79432), .Y(n2491) );
  MUX2X1 U3228 ( .B(C25909_net2740), .A(n2495), .S(net79432), .Y(n2494) );
  MUX2X1 U3229 ( .B(n2497), .A(n2498), .S(net79432), .Y(n2496) );
  MUX2X1 U3230 ( .B(n2500), .A(n2501), .S(n231), .Y(n2499) );
  MUX2X1 U3231 ( .B(n2503), .A(n2504), .S(net79432), .Y(n2502) );
  MUX2X1 U3232 ( .B(n2506), .A(n2507), .S(net79432), .Y(n2505) );
  MUX2X1 U3233 ( .B(n2510), .A(n2511), .S(net79432), .Y(n2508) );
  MUX2X1 U3234 ( .B(n2513), .A(n2514), .S(net79432), .Y(n2512) );
  MUX2X1 U3235 ( .B(n2516), .A(n2517), .S(n231), .Y(n2515) );
  MUX2X1 U3236 ( .B(n2519), .A(n2520), .S(net79432), .Y(n2518) );
  MUX2X1 U3237 ( .B(C25909_net2767), .A(n2522), .S(net79432), .Y(n2521) );
  MUX2X1 U3238 ( .B(n2524), .A(n2525), .S(net79432), .Y(n2523) );
  MUX2X1 U3239 ( .B(n2527), .A(n2528), .S(net79432), .Y(n2526) );
  MUX2X1 U3240 ( .B(n2530), .A(n2531), .S(n231), .Y(n2529) );
  MUX2X1 U3241 ( .B(n2533), .A(n2534), .S(net79432), .Y(n2532) );
  MUX2X1 U3242 ( .B(n2536), .A(n2537), .S(net79432), .Y(n2535) );
  MUX2X1 U3243 ( .B(n2539), .A(n2540), .S(net79432), .Y(n2538) );
  MUX2X1 U3244 ( .B(n2542), .A(n2543), .S(net79432), .Y(n2541) );
  MUX2X1 U3245 ( .B(n2545), .A(n2549), .S(n231), .Y(n2544) );
  MUX2X1 U3246 ( .B(n2646), .A(n2652), .S(net79434), .Y(n2629) );
  MUX2X1 U3247 ( .B(n2661), .A(n2671), .S(net79434), .Y(n2655) );
  MUX2X1 U3248 ( .B(n2712), .A(n2714), .S(net79434), .Y(n2706) );
  MUX2X1 U3249 ( .B(n2726), .A(n2748), .S(net79434), .Y(n2723) );
  MUX2X1 U3250 ( .B(n2755), .A(n2759), .S(n231), .Y(n2751) );
  MUX2X1 U3251 ( .B(n2770), .A(n2776), .S(net79434), .Y(n2762) );
  MUX2X1 U3252 ( .B(n2797), .A(n2800), .S(net79434), .Y(n2795) );
  MUX2X1 U3253 ( .B(n2809), .A(n2812), .S(net79434), .Y(n2805) );
  MUX2X1 U3254 ( .B(n2817), .A(n2827), .S(net79434), .Y(n2813) );
  MUX2X1 U3255 ( .B(n2840), .A(n2844), .S(n231), .Y(n2833) );
  MUX2X1 U3256 ( .B(n2846), .A(n2848), .S(net79434), .Y(n2845) );
  MUX2X1 U3257 ( .B(n2856), .A(n2873), .S(net79434), .Y(n2853) );
  MUX2X1 U3258 ( .B(n2878), .A(n2884), .S(net79434), .Y(n2875) );
  MUX2X1 U3259 ( .B(n2890), .A(n2891), .S(net79434), .Y(n2886) );
  MUX2X1 U3260 ( .B(n2893), .A(n2894), .S(n231), .Y(n2892) );
  MUX2X1 U3261 ( .B(n2896), .A(n2897), .S(net79434), .Y(n2895) );
  MUX2X1 U3262 ( .B(n2899), .A(n2902), .S(net79434), .Y(n2898) );
  MUX2X1 U3263 ( .B(n2922), .A(n2925), .S(net79434), .Y(n2903) );
  MUX2X1 U3264 ( .B(n2930), .A(n2931), .S(net79434), .Y(n2929) );
  MUX2X1 U3265 ( .B(n2933), .A(n2935), .S(n231), .Y(n2932) );
  MUX2X1 U3266 ( .B(n2944), .A(n2945), .S(net79434), .Y(n2943) );
  MUX2X1 U3267 ( .B(n2955), .A(n2956), .S(net79434), .Y(n2951) );
  MUX2X1 U3268 ( .B(n2960), .A(n2965), .S(net79434), .Y(n2958) );
  MUX2X1 U3269 ( .B(n2974), .A(n2983), .S(net79434), .Y(n2967) );
  MUX2X1 U3270 ( .B(n3002), .A(n3020), .S(n231), .Y(n2997) );
  MUX2X1 U3271 ( .B(n3030), .A(n3033), .S(net79434), .Y(n3026) );
  MUX2X1 U3272 ( .B(n3052), .A(n3062), .S(net79434), .Y(n3035) );
  MUX2X1 U3273 ( .B(n3074), .A(n3103), .S(net79434), .Y(n3068) );
  MUX2X1 U3274 ( .B(n3109), .A(n3114), .S(net79434), .Y(n3105) );
  MUX2X1 U3275 ( .B(n3119), .A(n3120), .S(n231), .Y(n3116) );
  MUX2X1 U3276 ( .B(n3127), .A(n3133), .S(net79434), .Y(n3125) );
  MUX2X1 U3277 ( .B(n3424), .A(n3425), .S(net79434), .Y(n3423) );
  MUX2X1 U3278 ( .B(n3429), .A(n3430), .S(net79434), .Y(n3426) );
  MUX2X1 U3279 ( .B(n3432), .A(n3433), .S(net79434), .Y(n3431) );
  MUX2X1 U3280 ( .B(n3435), .A(n3436), .S(n231), .Y(n3434) );
  MUX2X1 U3281 ( .B(n3438), .A(n3439), .S(net79434), .Y(n3437) );
  MUX2X1 U3282 ( .B(n3441), .A(n3442), .S(net79434), .Y(n3440) );
  MUX2X1 U3283 ( .B(n3444), .A(n3445), .S(net79436), .Y(n3443) );
  MUX2X1 U3284 ( .B(n3447), .A(n3448), .S(net79436), .Y(n3446) );
  MUX2X1 U3285 ( .B(n3450), .A(n3451), .S(n231), .Y(n3449) );
  MUX2X1 U3286 ( .B(n3453), .A(n3454), .S(net79436), .Y(n3452) );
  MUX2X1 U3287 ( .B(n3456), .A(n3457), .S(net79436), .Y(n3455) );
  MUX2X1 U3288 ( .B(C25909_net2920), .A(n3459), .S(net79436), .Y(n3458) );
  MUX2X1 U3289 ( .B(n3461), .A(n3462), .S(net79436), .Y(n3460) );
  MUX2X1 U3290 ( .B(n3464), .A(n3465), .S(n231), .Y(n3463) );
  MUX2X1 U3291 ( .B(n3467), .A(n3468), .S(net79436), .Y(n3466) );
  MUX2X1 U3292 ( .B(n3470), .A(n3471), .S(net79436), .Y(n3469) );
  MUX2X1 U3293 ( .B(n3473), .A(n3474), .S(net79436), .Y(n3472) );
  MUX2X1 U3294 ( .B(n3476), .A(n3477), .S(net79436), .Y(n3475) );
  MUX2X1 U3295 ( .B(n3479), .A(n3480), .S(n231), .Y(n3478) );
  MUX2X1 U3296 ( .B(n3482), .A(n3483), .S(net79436), .Y(n3481) );
  MUX2X1 U3297 ( .B(n3485), .A(n3486), .S(net79436), .Y(n3484) );
  MUX2X1 U3298 ( .B(n3488), .A(n3489), .S(net79436), .Y(n3487) );
  MUX2X1 U3299 ( .B(n3491), .A(n3492), .S(net79436), .Y(n3490) );
  MUX2X1 U3300 ( .B(n3494), .A(n3495), .S(n231), .Y(n3493) );
  MUX2X1 U3301 ( .B(buff_data[16]), .A(buff_data[0]), .S(net79402), .Y(n2203)
         );
  MUX2X1 U3302 ( .B(buff_data[48]), .A(buff_data[32]), .S(net79410), .Y(n2202)
         );
  MUX2X1 U3303 ( .B(buff_data[80]), .A(buff_data[64]), .S(net79414), .Y(n2206)
         );
  MUX2X1 U3304 ( .B(buff_data[112]), .A(buff_data[96]), .S(net79414), .Y(n2205) );
  MUX2X1 U3305 ( .B(n2204), .A(n2201), .S(n230), .Y(n2215) );
  MUX2X1 U3306 ( .B(buff_data[144]), .A(buff_data[128]), .S(net79414), .Y(
        n2209) );
  MUX2X1 U3307 ( .B(buff_data[176]), .A(buff_data[160]), .S(net79414), .Y(
        n2208) );
  MUX2X1 U3308 ( .B(buff_data[208]), .A(buff_data[192]), .S(net79414), .Y(
        n2212) );
  MUX2X1 U3309 ( .B(buff_data[240]), .A(buff_data[224]), .S(net79414), .Y(
        n2211) );
  MUX2X1 U3310 ( .B(n2210), .A(n2207), .S(n230), .Y(n2214) );
  MUX2X1 U3311 ( .B(buff_data[272]), .A(buff_data[256]), .S(net79414), .Y(
        n2218) );
  MUX2X1 U3312 ( .B(buff_data[304]), .A(buff_data[288]), .S(net79414), .Y(
        n2217) );
  MUX2X1 U3313 ( .B(buff_data[336]), .A(buff_data[320]), .S(net79414), .Y(
        n2221) );
  MUX2X1 U3314 ( .B(buff_data[368]), .A(buff_data[352]), .S(net79414), .Y(
        n2220) );
  MUX2X1 U3315 ( .B(n2219), .A(n2216), .S(n230), .Y(n2230) );
  MUX2X1 U3316 ( .B(buff_data[400]), .A(buff_data[384]), .S(net79414), .Y(
        n2224) );
  MUX2X1 U3317 ( .B(buff_data[432]), .A(buff_data[416]), .S(net79414), .Y(
        n2223) );
  MUX2X1 U3318 ( .B(buff_data[464]), .A(buff_data[448]), .S(net79414), .Y(
        n2227) );
  MUX2X1 U3319 ( .B(buff_data[496]), .A(buff_data[480]), .S(net79414), .Y(
        n2226) );
  MUX2X1 U3320 ( .B(n2225), .A(n2222), .S(n230), .Y(n2229) );
  MUX2X1 U3321 ( .B(n2228), .A(n2213), .S(n232), .Y(n3496) );
  INVX2 U3322 ( .A(n3496), .Y(n248) );
  MUX2X1 U3323 ( .B(buff_data[17]), .A(buff_data[1]), .S(net79408), .Y(n2233)
         );
  MUX2X1 U3324 ( .B(buff_data[49]), .A(buff_data[33]), .S(net79408), .Y(n2232)
         );
  MUX2X1 U3325 ( .B(buff_data[81]), .A(buff_data[65]), .S(net79408), .Y(n2236)
         );
  MUX2X1 U3326 ( .B(buff_data[113]), .A(buff_data[97]), .S(net79408), .Y(n2235) );
  MUX2X1 U3327 ( .B(n2234), .A(n2231), .S(n230), .Y(n2245) );
  MUX2X1 U3328 ( .B(buff_data[145]), .A(buff_data[129]), .S(net79408), .Y(
        n2239) );
  MUX2X1 U3329 ( .B(buff_data[177]), .A(buff_data[161]), .S(net79408), .Y(
        n2238) );
  MUX2X1 U3330 ( .B(buff_data[209]), .A(buff_data[193]), .S(net79408), .Y(
        n2242) );
  MUX2X1 U3331 ( .B(buff_data[241]), .A(buff_data[225]), .S(net79408), .Y(
        n2241) );
  MUX2X1 U3332 ( .B(n2240), .A(n2237), .S(n230), .Y(n2244) );
  MUX2X1 U3333 ( .B(buff_data[273]), .A(buff_data[257]), .S(net79408), .Y(
        n2248) );
  MUX2X1 U3334 ( .B(buff_data[305]), .A(buff_data[289]), .S(net79408), .Y(
        n2247) );
  MUX2X1 U3335 ( .B(buff_data[337]), .A(buff_data[321]), .S(net79408), .Y(
        n2251) );
  MUX2X1 U3336 ( .B(buff_data[369]), .A(buff_data[353]), .S(net79408), .Y(
        n2250) );
  MUX2X1 U3337 ( .B(n2249), .A(n2246), .S(n230), .Y(n2260) );
  MUX2X1 U3338 ( .B(buff_data[401]), .A(buff_data[385]), .S(net79408), .Y(
        n2254) );
  MUX2X1 U3339 ( .B(buff_data[433]), .A(buff_data[417]), .S(net79408), .Y(
        n2253) );
  MUX2X1 U3340 ( .B(buff_data[465]), .A(buff_data[449]), .S(net79408), .Y(
        n2257) );
  MUX2X1 U3341 ( .B(buff_data[497]), .A(buff_data[481]), .S(net79408), .Y(
        n2256) );
  MUX2X1 U3342 ( .B(n2255), .A(n2252), .S(n230), .Y(n2259) );
  MUX2X1 U3343 ( .B(n2258), .A(n2243), .S(n232), .Y(n3497) );
  MUX2X1 U3344 ( .B(buff_data[18]), .A(buff_data[2]), .S(net79408), .Y(n2263)
         );
  MUX2X1 U3345 ( .B(buff_data[50]), .A(buff_data[34]), .S(net79408), .Y(n2262)
         );
  MUX2X1 U3346 ( .B(buff_data[82]), .A(buff_data[66]), .S(net79408), .Y(n2266)
         );
  MUX2X1 U3347 ( .B(buff_data[114]), .A(buff_data[98]), .S(net79408), .Y(n2265) );
  MUX2X1 U3348 ( .B(n2264), .A(n2261), .S(n230), .Y(n2275) );
  MUX2X1 U3349 ( .B(buff_data[146]), .A(buff_data[130]), .S(net79408), .Y(
        n2269) );
  MUX2X1 U3350 ( .B(buff_data[178]), .A(buff_data[162]), .S(net79408), .Y(
        n2268) );
  MUX2X1 U3351 ( .B(buff_data[210]), .A(buff_data[194]), .S(net79408), .Y(
        n2272) );
  MUX2X1 U3352 ( .B(buff_data[242]), .A(buff_data[226]), .S(net79408), .Y(
        n2271) );
  MUX2X1 U3353 ( .B(n2270), .A(n2267), .S(n230), .Y(n2274) );
  MUX2X1 U3354 ( .B(buff_data[274]), .A(buff_data[258]), .S(net79408), .Y(
        n2278) );
  MUX2X1 U3355 ( .B(buff_data[306]), .A(buff_data[290]), .S(net79408), .Y(
        n2277) );
  MUX2X1 U3356 ( .B(buff_data[338]), .A(buff_data[322]), .S(net79408), .Y(
        n2281) );
  MUX2X1 U3357 ( .B(buff_data[370]), .A(buff_data[354]), .S(net79408), .Y(
        n2280) );
  MUX2X1 U3358 ( .B(n2279), .A(n2276), .S(n230), .Y(n2290) );
  MUX2X1 U3359 ( .B(buff_data[402]), .A(buff_data[386]), .S(net79408), .Y(
        n2284) );
  MUX2X1 U3360 ( .B(buff_data[434]), .A(buff_data[418]), .S(net79408), .Y(
        n2283) );
  MUX2X1 U3361 ( .B(buff_data[466]), .A(buff_data[450]), .S(net79410), .Y(
        n2287) );
  MUX2X1 U3362 ( .B(buff_data[498]), .A(buff_data[482]), .S(net79410), .Y(
        n2286) );
  MUX2X1 U3363 ( .B(n2285), .A(n2282), .S(n230), .Y(n2289) );
  MUX2X1 U3364 ( .B(n2288), .A(n2273), .S(n232), .Y(n3498) );
  INVX2 U3365 ( .A(n3498), .Y(n246) );
  MUX2X1 U3366 ( .B(buff_data[19]), .A(buff_data[3]), .S(net79410), .Y(n2293)
         );
  MUX2X1 U3367 ( .B(buff_data[51]), .A(buff_data[35]), .S(net79410), .Y(n2292)
         );
  MUX2X1 U3368 ( .B(buff_data[83]), .A(buff_data[67]), .S(net79410), .Y(n2296)
         );
  MUX2X1 U3369 ( .B(buff_data[115]), .A(buff_data[99]), .S(net79410), .Y(n2295) );
  MUX2X1 U3370 ( .B(n2294), .A(n2291), .S(n230), .Y(n2305) );
  MUX2X1 U3371 ( .B(buff_data[147]), .A(buff_data[131]), .S(net79410), .Y(
        n2299) );
  MUX2X1 U3372 ( .B(buff_data[179]), .A(buff_data[163]), .S(net79410), .Y(
        n2298) );
  MUX2X1 U3373 ( .B(buff_data[211]), .A(buff_data[195]), .S(net79410), .Y(
        n2302) );
  MUX2X1 U3374 ( .B(buff_data[243]), .A(buff_data[227]), .S(net79410), .Y(
        n2301) );
  MUX2X1 U3375 ( .B(n2300), .A(n2297), .S(n230), .Y(n2304) );
  MUX2X1 U3376 ( .B(buff_data[275]), .A(buff_data[259]), .S(net79410), .Y(
        n2308) );
  MUX2X1 U3377 ( .B(buff_data[307]), .A(buff_data[291]), .S(net79410), .Y(
        n2307) );
  MUX2X1 U3378 ( .B(buff_data[339]), .A(buff_data[323]), .S(net79410), .Y(
        n2311) );
  MUX2X1 U3379 ( .B(buff_data[371]), .A(buff_data[355]), .S(net79410), .Y(
        n2310) );
  MUX2X1 U3380 ( .B(n2309), .A(n2306), .S(n230), .Y(n2320) );
  MUX2X1 U3381 ( .B(buff_data[403]), .A(buff_data[387]), .S(net79410), .Y(
        n2314) );
  MUX2X1 U3382 ( .B(buff_data[435]), .A(buff_data[419]), .S(net79410), .Y(
        n2313) );
  MUX2X1 U3383 ( .B(buff_data[467]), .A(buff_data[451]), .S(net79410), .Y(
        n2317) );
  MUX2X1 U3384 ( .B(buff_data[499]), .A(buff_data[483]), .S(net79410), .Y(
        n2316) );
  MUX2X1 U3385 ( .B(n2315), .A(n2312), .S(n230), .Y(n2319) );
  MUX2X1 U3386 ( .B(n2318), .A(n2303), .S(n232), .Y(n3499) );
  MUX2X1 U3387 ( .B(buff_data[20]), .A(buff_data[4]), .S(net79410), .Y(n2323)
         );
  MUX2X1 U3388 ( .B(buff_data[52]), .A(buff_data[36]), .S(net79410), .Y(n2322)
         );
  MUX2X1 U3389 ( .B(buff_data[84]), .A(buff_data[68]), .S(net79410), .Y(n2326)
         );
  MUX2X1 U3390 ( .B(buff_data[116]), .A(buff_data[100]), .S(net79410), .Y(
        n2325) );
  MUX2X1 U3391 ( .B(n2324), .A(n2321), .S(n230), .Y(n2335) );
  MUX2X1 U3392 ( .B(buff_data[148]), .A(buff_data[132]), .S(net79410), .Y(
        n2329) );
  MUX2X1 U3393 ( .B(buff_data[180]), .A(buff_data[164]), .S(net79410), .Y(
        n2328) );
  MUX2X1 U3394 ( .B(buff_data[212]), .A(buff_data[196]), .S(net79410), .Y(
        n2332) );
  MUX2X1 U3395 ( .B(buff_data[244]), .A(buff_data[228]), .S(net79410), .Y(
        n2331) );
  MUX2X1 U3396 ( .B(n2330), .A(n2327), .S(n230), .Y(n2334) );
  MUX2X1 U3397 ( .B(buff_data[276]), .A(buff_data[260]), .S(net79410), .Y(
        n2338) );
  MUX2X1 U3398 ( .B(buff_data[308]), .A(buff_data[292]), .S(net79410), .Y(
        n2337) );
  MUX2X1 U3399 ( .B(buff_data[340]), .A(buff_data[324]), .S(net79410), .Y(
        n2341) );
  MUX2X1 U3400 ( .B(buff_data[372]), .A(buff_data[356]), .S(net79412), .Y(
        n2340) );
  MUX2X1 U3401 ( .B(n2339), .A(n2336), .S(n230), .Y(n2349) );
  MUX2X1 U3402 ( .B(buff_data[404]), .A(buff_data[388]), .S(net79412), .Y(
        n2344) );
  MUX2X1 U3403 ( .B(buff_data[436]), .A(buff_data[420]), .S(net79412), .Y(
        n2343) );
  MUX2X1 U3404 ( .B(buff_data[500]), .A(buff_data[484]), .S(net79412), .Y(
        n2346) );
  MUX2X1 U3405 ( .B(n2345), .A(n2342), .S(n230), .Y(n2348) );
  MUX2X1 U3406 ( .B(n2347), .A(n2333), .S(n232), .Y(n3500) );
  MUX2X1 U3407 ( .B(buff_data[21]), .A(buff_data[5]), .S(net79412), .Y(n2352)
         );
  MUX2X1 U3408 ( .B(buff_data[53]), .A(buff_data[37]), .S(net79412), .Y(n2351)
         );
  MUX2X1 U3409 ( .B(buff_data[85]), .A(buff_data[69]), .S(net79412), .Y(n2355)
         );
  MUX2X1 U3410 ( .B(buff_data[117]), .A(buff_data[101]), .S(net79412), .Y(
        n2354) );
  MUX2X1 U3411 ( .B(n2353), .A(n2350), .S(n230), .Y(n2364) );
  MUX2X1 U3412 ( .B(buff_data[149]), .A(buff_data[133]), .S(net79412), .Y(
        n2358) );
  MUX2X1 U3413 ( .B(buff_data[181]), .A(buff_data[165]), .S(net79412), .Y(
        n2357) );
  MUX2X1 U3414 ( .B(buff_data[213]), .A(buff_data[197]), .S(net79412), .Y(
        n2361) );
  MUX2X1 U3415 ( .B(buff_data[245]), .A(buff_data[229]), .S(net79412), .Y(
        n2360) );
  MUX2X1 U3416 ( .B(n2359), .A(n2356), .S(n230), .Y(n2363) );
  MUX2X1 U3417 ( .B(buff_data[277]), .A(buff_data[261]), .S(net79412), .Y(
        n2367) );
  MUX2X1 U3418 ( .B(buff_data[309]), .A(buff_data[293]), .S(net79412), .Y(
        n2366) );
  MUX2X1 U3419 ( .B(buff_data[341]), .A(buff_data[325]), .S(net79412), .Y(
        n2370) );
  MUX2X1 U3420 ( .B(buff_data[373]), .A(buff_data[357]), .S(net79412), .Y(
        n2369) );
  MUX2X1 U3421 ( .B(n2368), .A(n2365), .S(n230), .Y(n2410) );
  MUX2X1 U3422 ( .B(buff_data[405]), .A(buff_data[389]), .S(net79412), .Y(
        n2373) );
  MUX2X1 U3423 ( .B(buff_data[437]), .A(buff_data[421]), .S(net79412), .Y(
        n2372) );
  MUX2X1 U3424 ( .B(buff_data[469]), .A(buff_data[453]), .S(net79412), .Y(
        n2377) );
  MUX2X1 U3425 ( .B(buff_data[501]), .A(buff_data[485]), .S(net79412), .Y(
        n2376) );
  MUX2X1 U3426 ( .B(n2374), .A(n2371), .S(n230), .Y(n2409) );
  MUX2X1 U3427 ( .B(n2408), .A(n2362), .S(n232), .Y(n3501) );
  MUX2X1 U3428 ( .B(buff_data[22]), .A(buff_data[6]), .S(net79412), .Y(n2413)
         );
  MUX2X1 U3429 ( .B(buff_data[54]), .A(buff_data[38]), .S(net79412), .Y(n2412)
         );
  MUX2X1 U3430 ( .B(buff_data[86]), .A(buff_data[70]), .S(net79412), .Y(n2416)
         );
  MUX2X1 U3431 ( .B(buff_data[118]), .A(buff_data[102]), .S(net79412), .Y(
        n2415) );
  MUX2X1 U3432 ( .B(n2414), .A(n2411), .S(n230), .Y(n2425) );
  MUX2X1 U3433 ( .B(buff_data[150]), .A(buff_data[134]), .S(net79412), .Y(
        n2419) );
  MUX2X1 U3434 ( .B(buff_data[182]), .A(buff_data[166]), .S(net79412), .Y(
        n2418) );
  MUX2X1 U3435 ( .B(buff_data[214]), .A(buff_data[198]), .S(net79412), .Y(
        n2422) );
  MUX2X1 U3436 ( .B(buff_data[246]), .A(buff_data[230]), .S(net79412), .Y(
        n2421) );
  MUX2X1 U3437 ( .B(n2420), .A(n2417), .S(n230), .Y(n2424) );
  MUX2X1 U3438 ( .B(buff_data[278]), .A(buff_data[262]), .S(net79412), .Y(
        n2428) );
  MUX2X1 U3439 ( .B(buff_data[310]), .A(buff_data[294]), .S(net79414), .Y(
        n2427) );
  MUX2X1 U3440 ( .B(buff_data[342]), .A(buff_data[326]), .S(net79414), .Y(
        n2431) );
  MUX2X1 U3441 ( .B(buff_data[374]), .A(buff_data[358]), .S(net79414), .Y(
        n2430) );
  MUX2X1 U3442 ( .B(n2429), .A(n2426), .S(n230), .Y(n2441) );
  MUX2X1 U3443 ( .B(buff_data[406]), .A(buff_data[390]), .S(net79414), .Y(
        n2434) );
  MUX2X1 U3444 ( .B(buff_data[438]), .A(buff_data[422]), .S(net79414), .Y(
        n2433) );
  MUX2X1 U3445 ( .B(buff_data[470]), .A(buff_data[454]), .S(net79414), .Y(
        n2437) );
  MUX2X1 U3446 ( .B(buff_data[502]), .A(buff_data[486]), .S(net79414), .Y(
        n2436) );
  MUX2X1 U3447 ( .B(n2435), .A(n2432), .S(n230), .Y(n2440) );
  MUX2X1 U3448 ( .B(n2438), .A(n2423), .S(n232), .Y(n3502) );
  MUX2X1 U3449 ( .B(buff_data[23]), .A(buff_data[7]), .S(net79414), .Y(n2445)
         );
  MUX2X1 U3450 ( .B(buff_data[55]), .A(buff_data[39]), .S(net79414), .Y(n2444)
         );
  MUX2X1 U3451 ( .B(buff_data[87]), .A(buff_data[71]), .S(net79414), .Y(n2448)
         );
  MUX2X1 U3452 ( .B(buff_data[119]), .A(buff_data[103]), .S(net79414), .Y(
        n2447) );
  MUX2X1 U3453 ( .B(n2446), .A(n2443), .S(n230), .Y(n2457) );
  MUX2X1 U3454 ( .B(buff_data[151]), .A(buff_data[135]), .S(net79414), .Y(
        n2451) );
  MUX2X1 U3455 ( .B(buff_data[183]), .A(buff_data[167]), .S(net79414), .Y(
        n2450) );
  MUX2X1 U3456 ( .B(buff_data[215]), .A(buff_data[199]), .S(net79414), .Y(
        n2454) );
  MUX2X1 U3457 ( .B(buff_data[247]), .A(buff_data[231]), .S(net79414), .Y(
        n2453) );
  MUX2X1 U3458 ( .B(n2452), .A(n2449), .S(n230), .Y(n2456) );
  MUX2X1 U3459 ( .B(buff_data[279]), .A(buff_data[263]), .S(net79414), .Y(
        n2460) );
  MUX2X1 U3460 ( .B(buff_data[311]), .A(buff_data[295]), .S(net79414), .Y(
        n2459) );
  MUX2X1 U3461 ( .B(buff_data[343]), .A(buff_data[327]), .S(net79414), .Y(
        n2463) );
  MUX2X1 U3462 ( .B(buff_data[375]), .A(buff_data[359]), .S(net79414), .Y(
        n2462) );
  MUX2X1 U3463 ( .B(n2461), .A(n2458), .S(n230), .Y(n2472) );
  MUX2X1 U3464 ( .B(buff_data[407]), .A(buff_data[391]), .S(net79414), .Y(
        n2466) );
  MUX2X1 U3465 ( .B(buff_data[439]), .A(buff_data[423]), .S(net79414), .Y(
        n2465) );
  MUX2X1 U3466 ( .B(buff_data[471]), .A(buff_data[455]), .S(net79414), .Y(
        n2469) );
  MUX2X1 U3467 ( .B(buff_data[503]), .A(buff_data[487]), .S(net79414), .Y(
        n2468) );
  MUX2X1 U3468 ( .B(n2467), .A(n2464), .S(n230), .Y(n2471) );
  MUX2X1 U3469 ( .B(n2470), .A(n2455), .S(n232), .Y(n3503) );
  MUX2X1 U3470 ( .B(buff_data[24]), .A(buff_data[8]), .S(net79402), .Y(n2475)
         );
  MUX2X1 U3471 ( .B(buff_data[56]), .A(buff_data[40]), .S(net79402), .Y(n2474)
         );
  MUX2X1 U3472 ( .B(buff_data[88]), .A(buff_data[72]), .S(net79402), .Y(n2478)
         );
  MUX2X1 U3473 ( .B(buff_data[120]), .A(buff_data[104]), .S(net79402), .Y(
        n2477) );
  MUX2X1 U3474 ( .B(n2476), .A(n2473), .S(n230), .Y(n2487) );
  MUX2X1 U3475 ( .B(buff_data[152]), .A(buff_data[136]), .S(net79402), .Y(
        n2481) );
  MUX2X1 U3476 ( .B(buff_data[184]), .A(buff_data[168]), .S(net79402), .Y(
        n2480) );
  MUX2X1 U3477 ( .B(buff_data[216]), .A(buff_data[200]), .S(net79402), .Y(
        n2484) );
  MUX2X1 U3478 ( .B(buff_data[248]), .A(buff_data[232]), .S(net79402), .Y(
        n2483) );
  MUX2X1 U3479 ( .B(n2482), .A(n2479), .S(n230), .Y(n2486) );
  MUX2X1 U3480 ( .B(buff_data[280]), .A(buff_data[264]), .S(net79402), .Y(
        n2490) );
  MUX2X1 U3481 ( .B(buff_data[312]), .A(buff_data[296]), .S(net79402), .Y(
        n2489) );
  MUX2X1 U3482 ( .B(buff_data[344]), .A(buff_data[328]), .S(net79402), .Y(
        n2493) );
  MUX2X1 U3483 ( .B(buff_data[376]), .A(buff_data[360]), .S(net79402), .Y(
        n2492) );
  MUX2X1 U3484 ( .B(n2491), .A(n2488), .S(n230), .Y(n2501) );
  MUX2X1 U3485 ( .B(buff_data[408]), .A(buff_data[392]), .S(net79402), .Y(
        n2495) );
  MUX2X1 U3486 ( .B(buff_data[472]), .A(buff_data[456]), .S(net79402), .Y(
        n2498) );
  MUX2X1 U3487 ( .B(buff_data[504]), .A(buff_data[488]), .S(net79402), .Y(
        n2497) );
  MUX2X1 U3488 ( .B(n2496), .A(n2494), .S(n230), .Y(n2500) );
  MUX2X1 U3489 ( .B(n2499), .A(n2485), .S(n232), .Y(n3504) );
  MUX2X1 U3490 ( .B(buff_data[25]), .A(buff_data[9]), .S(net79402), .Y(n2504)
         );
  MUX2X1 U3491 ( .B(buff_data[57]), .A(buff_data[41]), .S(net79402), .Y(n2503)
         );
  MUX2X1 U3492 ( .B(buff_data[89]), .A(buff_data[73]), .S(net79402), .Y(n2507)
         );
  MUX2X1 U3493 ( .B(buff_data[121]), .A(buff_data[105]), .S(net79402), .Y(
        n2506) );
  MUX2X1 U3494 ( .B(n2505), .A(n2502), .S(n230), .Y(n2517) );
  MUX2X1 U3495 ( .B(buff_data[153]), .A(buff_data[137]), .S(net79402), .Y(
        n2511) );
  MUX2X1 U3496 ( .B(buff_data[185]), .A(buff_data[169]), .S(net79402), .Y(
        n2510) );
  MUX2X1 U3497 ( .B(buff_data[217]), .A(buff_data[201]), .S(net79402), .Y(
        n2514) );
  MUX2X1 U3498 ( .B(buff_data[249]), .A(buff_data[233]), .S(net79402), .Y(
        n2513) );
  MUX2X1 U3499 ( .B(n2512), .A(n2508), .S(n230), .Y(n2516) );
  MUX2X1 U3500 ( .B(buff_data[281]), .A(buff_data[265]), .S(net79402), .Y(
        n2520) );
  MUX2X1 U3501 ( .B(buff_data[313]), .A(buff_data[297]), .S(net79402), .Y(
        n2519) );
  MUX2X1 U3502 ( .B(buff_data[345]), .A(buff_data[329]), .S(net79402), .Y(
        n2522) );
  MUX2X1 U3503 ( .B(n2521), .A(n2518), .S(n230), .Y(n2531) );
  MUX2X1 U3504 ( .B(buff_data[409]), .A(buff_data[393]), .S(net79402), .Y(
        n2525) );
  MUX2X1 U3505 ( .B(buff_data[441]), .A(buff_data[425]), .S(net79402), .Y(
        n2524) );
  MUX2X1 U3506 ( .B(buff_data[473]), .A(buff_data[457]), .S(net79402), .Y(
        n2528) );
  MUX2X1 U3507 ( .B(buff_data[505]), .A(buff_data[489]), .S(net79402), .Y(
        n2527) );
  MUX2X1 U3508 ( .B(n2526), .A(n2523), .S(n230), .Y(n2530) );
  MUX2X1 U3509 ( .B(n2529), .A(n2515), .S(n232), .Y(n3505) );
  MUX2X1 U3510 ( .B(buff_data[26]), .A(buff_data[10]), .S(net79402), .Y(n2534)
         );
  MUX2X1 U3511 ( .B(buff_data[58]), .A(buff_data[42]), .S(net79402), .Y(n2533)
         );
  MUX2X1 U3512 ( .B(buff_data[90]), .A(buff_data[74]), .S(net79402), .Y(n2537)
         );
  MUX2X1 U3513 ( .B(buff_data[122]), .A(buff_data[106]), .S(net79402), .Y(
        n2536) );
  MUX2X1 U3514 ( .B(n2535), .A(n2532), .S(n230), .Y(n2549) );
  MUX2X1 U3515 ( .B(buff_data[154]), .A(buff_data[138]), .S(net79402), .Y(
        n2540) );
  MUX2X1 U3516 ( .B(buff_data[186]), .A(buff_data[170]), .S(net79402), .Y(
        n2539) );
  MUX2X1 U3517 ( .B(buff_data[218]), .A(buff_data[202]), .S(net79402), .Y(
        n2543) );
  MUX2X1 U3518 ( .B(buff_data[250]), .A(buff_data[234]), .S(net79402), .Y(
        n2542) );
  MUX2X1 U3519 ( .B(n2541), .A(n2538), .S(n230), .Y(n2545) );
  MUX2X1 U3520 ( .B(buff_data[282]), .A(buff_data[266]), .S(net79402), .Y(
        n2652) );
  MUX2X1 U3521 ( .B(buff_data[314]), .A(buff_data[298]), .S(net79402), .Y(
        n2646) );
  MUX2X1 U3522 ( .B(buff_data[346]), .A(buff_data[330]), .S(net79402), .Y(
        n2671) );
  MUX2X1 U3523 ( .B(buff_data[378]), .A(buff_data[362]), .S(net79402), .Y(
        n2661) );
  MUX2X1 U3524 ( .B(n2655), .A(n2629), .S(n230), .Y(n2759) );
  MUX2X1 U3525 ( .B(buff_data[410]), .A(buff_data[394]), .S(net79402), .Y(
        n2714) );
  MUX2X1 U3526 ( .B(buff_data[442]), .A(buff_data[426]), .S(net79402), .Y(
        n2712) );
  MUX2X1 U3527 ( .B(buff_data[474]), .A(buff_data[458]), .S(net79402), .Y(
        n2748) );
  MUX2X1 U3528 ( .B(buff_data[506]), .A(buff_data[490]), .S(net79402), .Y(
        n2726) );
  MUX2X1 U3529 ( .B(n2723), .A(n2706), .S(n230), .Y(n2755) );
  MUX2X1 U3530 ( .B(n2751), .A(n2544), .S(n232), .Y(n3506) );
  MUX2X1 U3531 ( .B(buff_data[27]), .A(buff_data[11]), .S(net79402), .Y(n2776)
         );
  MUX2X1 U3532 ( .B(buff_data[59]), .A(buff_data[43]), .S(net79402), .Y(n2770)
         );
  MUX2X1 U3533 ( .B(buff_data[91]), .A(buff_data[75]), .S(net79402), .Y(n2800)
         );
  MUX2X1 U3534 ( .B(buff_data[123]), .A(buff_data[107]), .S(net79402), .Y(
        n2797) );
  MUX2X1 U3535 ( .B(n2795), .A(n2762), .S(n230), .Y(n2844) );
  MUX2X1 U3536 ( .B(buff_data[155]), .A(buff_data[139]), .S(net79402), .Y(
        n2812) );
  MUX2X1 U3537 ( .B(buff_data[187]), .A(buff_data[171]), .S(net79402), .Y(
        n2809) );
  MUX2X1 U3538 ( .B(buff_data[219]), .A(buff_data[203]), .S(net79402), .Y(
        n2827) );
  MUX2X1 U3539 ( .B(buff_data[251]), .A(buff_data[235]), .S(net79402), .Y(
        n2817) );
  MUX2X1 U3540 ( .B(n2813), .A(n2805), .S(n230), .Y(n2840) );
  MUX2X1 U3541 ( .B(buff_data[283]), .A(buff_data[267]), .S(net79402), .Y(
        n2848) );
  MUX2X1 U3542 ( .B(buff_data[315]), .A(buff_data[299]), .S(net79402), .Y(
        n2846) );
  MUX2X1 U3543 ( .B(buff_data[347]), .A(buff_data[331]), .S(net79402), .Y(
        n2873) );
  MUX2X1 U3544 ( .B(buff_data[379]), .A(buff_data[363]), .S(net79402), .Y(
        n2856) );
  MUX2X1 U3545 ( .B(n2853), .A(n2845), .S(n230), .Y(n2894) );
  MUX2X1 U3546 ( .B(buff_data[411]), .A(buff_data[395]), .S(net79402), .Y(
        n2884) );
  MUX2X1 U3547 ( .B(buff_data[443]), .A(buff_data[427]), .S(net79402), .Y(
        n2878) );
  MUX2X1 U3548 ( .B(buff_data[475]), .A(buff_data[459]), .S(net79402), .Y(
        n2891) );
  MUX2X1 U3549 ( .B(buff_data[507]), .A(buff_data[491]), .S(net79402), .Y(
        n2890) );
  MUX2X1 U3550 ( .B(n2886), .A(n2875), .S(n230), .Y(n2893) );
  MUX2X1 U3551 ( .B(n2892), .A(n2833), .S(n232), .Y(n3507) );
  MUX2X1 U3552 ( .B(buff_data[28]), .A(buff_data[12]), .S(net79402), .Y(n2897)
         );
  MUX2X1 U3553 ( .B(buff_data[60]), .A(buff_data[44]), .S(net79402), .Y(n2896)
         );
  MUX2X1 U3554 ( .B(buff_data[92]), .A(buff_data[76]), .S(net79402), .Y(n2902)
         );
  MUX2X1 U3555 ( .B(buff_data[124]), .A(buff_data[108]), .S(net79414), .Y(
        n2899) );
  MUX2X1 U3556 ( .B(n2898), .A(n2895), .S(n230), .Y(n2935) );
  MUX2X1 U3557 ( .B(buff_data[156]), .A(buff_data[140]), .S(net79402), .Y(
        n2925) );
  MUX2X1 U3558 ( .B(buff_data[188]), .A(buff_data[172]), .S(net79402), .Y(
        n2922) );
  MUX2X1 U3559 ( .B(buff_data[220]), .A(buff_data[204]), .S(net79402), .Y(
        n2931) );
  MUX2X1 U3560 ( .B(buff_data[252]), .A(buff_data[236]), .S(net79402), .Y(
        n2930) );
  MUX2X1 U3561 ( .B(n2929), .A(n2903), .S(n230), .Y(n2933) );
  MUX2X1 U3562 ( .B(buff_data[284]), .A(buff_data[268]), .S(net79402), .Y(
        n2945) );
  MUX2X1 U3563 ( .B(buff_data[316]), .A(buff_data[300]), .S(net79402), .Y(
        n2944) );
  MUX2X1 U3564 ( .B(buff_data[348]), .A(buff_data[332]), .S(net79402), .Y(
        n2956) );
  MUX2X1 U3565 ( .B(buff_data[380]), .A(buff_data[364]), .S(net79402), .Y(
        n2955) );
  MUX2X1 U3566 ( .B(n2951), .A(n2943), .S(n230), .Y(n3020) );
  MUX2X1 U3567 ( .B(buff_data[412]), .A(buff_data[396]), .S(net79402), .Y(
        n2965) );
  MUX2X1 U3568 ( .B(buff_data[444]), .A(buff_data[428]), .S(net79402), .Y(
        n2960) );
  MUX2X1 U3569 ( .B(buff_data[476]), .A(buff_data[460]), .S(net79402), .Y(
        n2983) );
  MUX2X1 U3570 ( .B(buff_data[508]), .A(buff_data[492]), .S(net79402), .Y(
        n2974) );
  MUX2X1 U3571 ( .B(n2967), .A(n2958), .S(n230), .Y(n3002) );
  MUX2X1 U3572 ( .B(n2997), .A(n2932), .S(n232), .Y(n3508) );
  MUX2X1 U3573 ( .B(buff_data[29]), .A(buff_data[13]), .S(net79402), .Y(n3033)
         );
  MUX2X1 U3574 ( .B(buff_data[61]), .A(buff_data[45]), .S(net79402), .Y(n3030)
         );
  MUX2X1 U3575 ( .B(buff_data[93]), .A(buff_data[77]), .S(net79402), .Y(n3062)
         );
  MUX2X1 U3576 ( .B(buff_data[125]), .A(buff_data[109]), .S(net79414), .Y(
        n3052) );
  MUX2X1 U3577 ( .B(n3035), .A(n3026), .S(n230), .Y(n3120) );
  MUX2X1 U3578 ( .B(buff_data[157]), .A(buff_data[141]), .S(net79414), .Y(
        n3103) );
  MUX2X1 U3579 ( .B(buff_data[189]), .A(buff_data[173]), .S(net79414), .Y(
        n3074) );
  MUX2X1 U3580 ( .B(buff_data[221]), .A(buff_data[205]), .S(net79414), .Y(
        n3114) );
  MUX2X1 U3581 ( .B(buff_data[253]), .A(buff_data[237]), .S(net79414), .Y(
        n3109) );
  MUX2X1 U3582 ( .B(n3105), .A(n3068), .S(n230), .Y(n3119) );
  MUX2X1 U3583 ( .B(buff_data[285]), .A(buff_data[269]), .S(net79414), .Y(
        n3133) );
  MUX2X1 U3584 ( .B(buff_data[317]), .A(buff_data[301]), .S(net79414), .Y(
        n3127) );
  MUX2X1 U3585 ( .B(buff_data[349]), .A(buff_data[333]), .S(net79414), .Y(
        n3425) );
  MUX2X1 U3586 ( .B(buff_data[381]), .A(buff_data[365]), .S(net79414), .Y(
        n3424) );
  MUX2X1 U3587 ( .B(n3423), .A(n3125), .S(n230), .Y(n3436) );
  MUX2X1 U3588 ( .B(buff_data[413]), .A(buff_data[397]), .S(net79414), .Y(
        n3430) );
  MUX2X1 U3589 ( .B(buff_data[445]), .A(buff_data[429]), .S(net79414), .Y(
        n3429) );
  MUX2X1 U3590 ( .B(buff_data[477]), .A(buff_data[461]), .S(net79414), .Y(
        n3433) );
  MUX2X1 U3591 ( .B(buff_data[509]), .A(buff_data[493]), .S(net79414), .Y(
        n3432) );
  MUX2X1 U3592 ( .B(n3431), .A(n3426), .S(n230), .Y(n3435) );
  MUX2X1 U3593 ( .B(n3434), .A(n3116), .S(n232), .Y(n3509) );
  MUX2X1 U3594 ( .B(buff_data[30]), .A(buff_data[14]), .S(net79414), .Y(n3439)
         );
  MUX2X1 U3595 ( .B(buff_data[62]), .A(buff_data[46]), .S(net79414), .Y(n3438)
         );
  MUX2X1 U3596 ( .B(buff_data[94]), .A(buff_data[78]), .S(net79414), .Y(n3442)
         );
  MUX2X1 U3597 ( .B(buff_data[126]), .A(buff_data[110]), .S(net79414), .Y(
        n3441) );
  MUX2X1 U3598 ( .B(n3440), .A(n3437), .S(n230), .Y(n3451) );
  MUX2X1 U3599 ( .B(buff_data[158]), .A(buff_data[142]), .S(net79414), .Y(
        n3445) );
  MUX2X1 U3600 ( .B(buff_data[190]), .A(buff_data[174]), .S(net79414), .Y(
        n3444) );
  MUX2X1 U3601 ( .B(buff_data[222]), .A(buff_data[206]), .S(net79414), .Y(
        n3448) );
  MUX2X1 U3602 ( .B(buff_data[254]), .A(buff_data[238]), .S(net79414), .Y(
        n3447) );
  MUX2X1 U3603 ( .B(n3446), .A(n3443), .S(n230), .Y(n3450) );
  MUX2X1 U3604 ( .B(buff_data[286]), .A(buff_data[270]), .S(net79414), .Y(
        n3454) );
  MUX2X1 U3605 ( .B(buff_data[318]), .A(buff_data[302]), .S(net79414), .Y(
        n3453) );
  MUX2X1 U3606 ( .B(buff_data[350]), .A(buff_data[334]), .S(net79414), .Y(
        n3457) );
  MUX2X1 U3607 ( .B(buff_data[382]), .A(buff_data[366]), .S(net79414), .Y(
        n3456) );
  MUX2X1 U3608 ( .B(n3455), .A(n3452), .S(n230), .Y(n3465) );
  MUX2X1 U3609 ( .B(buff_data[414]), .A(buff_data[398]), .S(net79414), .Y(
        n3459) );
  MUX2X1 U3610 ( .B(buff_data[478]), .A(buff_data[462]), .S(net79414), .Y(
        n3462) );
  MUX2X1 U3611 ( .B(buff_data[510]), .A(buff_data[494]), .S(net79414), .Y(
        n3461) );
  MUX2X1 U3612 ( .B(n3460), .A(n3458), .S(n230), .Y(n3464) );
  MUX2X1 U3613 ( .B(n3463), .A(n3449), .S(n232), .Y(n3510) );
  MUX2X1 U3614 ( .B(buff_data[31]), .A(buff_data[15]), .S(net79414), .Y(n3468)
         );
  MUX2X1 U3615 ( .B(buff_data[63]), .A(buff_data[47]), .S(net79414), .Y(n3467)
         );
  MUX2X1 U3616 ( .B(buff_data[95]), .A(buff_data[79]), .S(net79414), .Y(n3471)
         );
  MUX2X1 U3617 ( .B(buff_data[127]), .A(buff_data[111]), .S(net79414), .Y(
        n3470) );
  MUX2X1 U3618 ( .B(n3469), .A(n3466), .S(n230), .Y(n3480) );
  MUX2X1 U3619 ( .B(buff_data[159]), .A(buff_data[143]), .S(net79414), .Y(
        n3474) );
  MUX2X1 U3620 ( .B(buff_data[191]), .A(buff_data[175]), .S(net79414), .Y(
        n3473) );
  MUX2X1 U3621 ( .B(buff_data[223]), .A(buff_data[207]), .S(net79414), .Y(
        n3477) );
  MUX2X1 U3622 ( .B(buff_data[255]), .A(buff_data[239]), .S(net79414), .Y(
        n3476) );
  MUX2X1 U3623 ( .B(n3475), .A(n3472), .S(n230), .Y(n3479) );
  MUX2X1 U3624 ( .B(buff_data[287]), .A(buff_data[271]), .S(net79414), .Y(
        n3483) );
  MUX2X1 U3625 ( .B(buff_data[319]), .A(buff_data[303]), .S(net79414), .Y(
        n3482) );
  MUX2X1 U3626 ( .B(buff_data[351]), .A(buff_data[335]), .S(net79414), .Y(
        n3486) );
  MUX2X1 U3627 ( .B(buff_data[383]), .A(buff_data[367]), .S(net79414), .Y(
        n3485) );
  MUX2X1 U3628 ( .B(n3484), .A(n3481), .S(n230), .Y(n3495) );
  MUX2X1 U3629 ( .B(buff_data[415]), .A(buff_data[399]), .S(net79414), .Y(
        n3489) );
  MUX2X1 U3630 ( .B(buff_data[447]), .A(buff_data[431]), .S(net79414), .Y(
        n3488) );
  MUX2X1 U3631 ( .B(buff_data[479]), .A(buff_data[463]), .S(net79414), .Y(
        n3492) );
  MUX2X1 U3632 ( .B(buff_data[511]), .A(buff_data[495]), .S(net79414), .Y(
        n3491) );
  MUX2X1 U3633 ( .B(n3490), .A(n3487), .S(n230), .Y(n3494) );
  MUX2X1 U3634 ( .B(n3493), .A(n3478), .S(n232), .Y(n3511) );
  INVX2 U3635 ( .A(CMD_data_out[0]), .Y(n1885) );
  XOR2X1 U3636 ( .A(CMD_data_out[0]), .B(CMD_data_out[1]), .Y(n1886) );
  XOR2X1 U3637 ( .A(n581), .B(CMD_data_out[2]), .Y(n1887) );
  XOR2X1 U3638 ( .A(n607), .B(CMD_data_out[3]), .Y(n1888) );
  XOR2X1 U3639 ( .A(n608), .B(CMD_data_out[4]), .Y(n1889) );
  XOR2X1 U3640 ( .A(add_576_carry_8_), .B(CMD_data_out[5]), .Y(n1890) );
  XOR2X1 U3641 ( .A(add_576_carry_9_), .B(CMD_data_out[6]), .Y(n1891) );
  XOR2X1 U3642 ( .A(add_576_carry_10_), .B(CMD_data_out[7]), .Y(n1892) );
  INVX2 U3643 ( .A(n1251), .Y(add_576_carry_12_) );
  XOR2X1 U3644 ( .A(add_576_carry_11_), .B(CMD_data_out[8]), .Y(n1893) );
  XOR2X1 U3645 ( .A(CMD_data_out[9]), .B(add_576_carry_12_), .Y(n1894) );
  OR2X1 U3646 ( .A(i[26]), .B(i[25]), .Y(n3518) );
  NOR3X1 U3647 ( .A(n3518), .B(i[24]), .C(i[23]), .Y(r576_net62635) );
  OR2X1 U3648 ( .A(i[30]), .B(i[29]), .Y(n3519) );
  NOR3X1 U3649 ( .A(n3519), .B(i[28]), .C(i[27]), .Y(r576_net62636) );
  OR2X1 U3650 ( .A(i[26]), .B(i[25]), .Y(n3520) );
  NOR3X1 U3651 ( .A(n3520), .B(i[24]), .C(i[23]), .Y(n3523) );
  OR2X1 U3652 ( .A(i[30]), .B(i[29]), .Y(n3521) );
  NOR3X1 U3653 ( .A(n3521), .B(i[28]), .C(i[27]), .Y(n3522) );
  NOR3X1 U3654 ( .A(i[16]), .B(i[18]), .C(i[17]), .Y(n3524) );
  INVX1 U3655 ( .A(i[31]), .Y(r577_net62534) );
  OAI21X1 U3656 ( .A(n1259), .B(n1324), .C(r577_net62534), .Y(n3540) );
  OR2X1 U3657 ( .A(i[5]), .B(i[4]), .Y(n3529) );
  NOR3X1 U3658 ( .A(n3529), .B(i[3]), .C(i[2]), .Y(n3532) );
  OR2X1 U3659 ( .A(i[9]), .B(i[8]), .Y(n3530) );
  NOR3X1 U3660 ( .A(n3530), .B(i[7]), .C(i[6]), .Y(n3531) );
  OR2X1 U3661 ( .A(i[12]), .B(i[11]), .Y(n3533) );
  NOR3X1 U3662 ( .A(n3533), .B(i[10]), .C(i[0]), .Y(n3536) );
  OR2X1 U3663 ( .A(i[1]), .B(i[15]), .Y(n3534) );
  NOR3X1 U3664 ( .A(n3534), .B(i[14]), .C(i[13]), .Y(n3535) );
  OAI21X1 U3665 ( .A(n1262), .B(n1345), .C(r577_net62534), .Y(n3539) );
  AND2X1 U3666 ( .A(i[1]), .B(i[0]), .Y(n3541) );
  NAND3X1 U3667 ( .A(i[3]), .B(i[2]), .C(n3541), .Y(n3550) );
  OR2X1 U3668 ( .A(i[5]), .B(i[4]), .Y(n3542) );
  NOR3X1 U3669 ( .A(n3542), .B(i[11]), .C(i[10]), .Y(n3545) );
  OR2X1 U3670 ( .A(i[9]), .B(i[8]), .Y(n3543) );
  NOR3X1 U3671 ( .A(n3543), .B(i[7]), .C(i[6]), .Y(n3544) );
  AND2X1 U3672 ( .A(n3545), .B(n3544), .Y(n3561) );
  NOR3X1 U3673 ( .A(i[12]), .B(i[14]), .C(i[13]), .Y(n3546) );
  NAND3X1 U3674 ( .A(n1242), .B(n1309), .C(n3546), .Y(n3549) );
  INVX1 U3675 ( .A(n3549), .Y(n3562) );
  NAND3X1 U3676 ( .A(n838), .B(n3561), .C(n3562), .Y(n3556) );
  NOR3X1 U3677 ( .A(i[19]), .B(i[21]), .C(i[20]), .Y(n3551) );
  NOR3X1 U3678 ( .A(i[28]), .B(i[30]), .C(i[29]), .Y(n3554) );
  NOR3X1 U3679 ( .A(n1401), .B(n1590), .C(n1605), .Y(n3557) );
  NAND3X1 U3680 ( .A(n3562), .B(n3561), .C(n1372), .Y(n3563) );
  INVX1 U3681 ( .A(n3563), .Y(n3564) );
  OAI21X1 U3682 ( .A(n426), .B(n3566), .C(n479), .Y(n3427) );
  INVX1 U3683 ( .A(blk_cnt[31]), .Y(n3566) );
  OAI21X1 U3684 ( .A(n422), .B(n3569), .C(n475), .Y(n3421) );
  AOI22X1 U3685 ( .A(n3571), .B(n3572), .C(n1752), .D(n3568), .Y(n3570) );
  INVX1 U3686 ( .A(blk_cnt[3]), .Y(n3569) );
  OAI21X1 U3687 ( .A(n426), .B(n3573), .C(n476), .Y(n3419) );
  AOI22X1 U3688 ( .A(n3571), .B(n3575), .C(n1753), .D(n3568), .Y(n3574) );
  XNOR2X1 U3689 ( .A(CMD_data_out[30]), .B(n3572), .Y(n3575) );
  INVX1 U3690 ( .A(CMD_data_out[29]), .Y(n3572) );
  OAI21X1 U3691 ( .A(n423), .B(n3576), .C(n477), .Y(n3417) );
  AOI22X1 U3692 ( .A(n3578), .B(CMD_data_out[29]), .C(n1754), .D(n3568), .Y(
        n3577) );
  OAI21X1 U3693 ( .A(n426), .B(n3580), .C(n582), .Y(n3415) );
  INVX1 U3694 ( .A(blk_cnt[6]), .Y(n3580) );
  OAI21X1 U3695 ( .A(n422), .B(n3582), .C(n583), .Y(n3413) );
  INVX1 U3696 ( .A(blk_cnt[7]), .Y(n3582) );
  OAI21X1 U3697 ( .A(n426), .B(n3584), .C(n584), .Y(n3411) );
  OAI21X1 U3698 ( .A(n423), .B(n3586), .C(n585), .Y(n3409) );
  OAI21X1 U3699 ( .A(n426), .B(n3588), .C(n586), .Y(n3407) );
  OAI21X1 U3700 ( .A(n422), .B(n3590), .C(n587), .Y(n3405) );
  OAI21X1 U3701 ( .A(n426), .B(n3592), .C(n588), .Y(n3403) );
  OAI21X1 U3702 ( .A(n423), .B(n3594), .C(n589), .Y(n3401) );
  OAI21X1 U3703 ( .A(n426), .B(n3596), .C(n590), .Y(n3399) );
  OAI21X1 U3704 ( .A(n422), .B(n3598), .C(n591), .Y(n3397) );
  OAI21X1 U3705 ( .A(n426), .B(n3600), .C(n592), .Y(n3395) );
  OAI21X1 U3706 ( .A(n423), .B(n3602), .C(n593), .Y(n3393) );
  OAI21X1 U3707 ( .A(n426), .B(n3604), .C(n594), .Y(n3391) );
  OAI21X1 U3708 ( .A(n422), .B(n3606), .C(n595), .Y(n3389) );
  OAI21X1 U3709 ( .A(n423), .B(n3608), .C(n596), .Y(n3387) );
  OAI21X1 U3710 ( .A(n422), .B(n3610), .C(n597), .Y(n3385) );
  OAI21X1 U3711 ( .A(n423), .B(n3612), .C(n598), .Y(n3383) );
  OAI21X1 U3712 ( .A(n422), .B(n3614), .C(n599), .Y(n3381) );
  OAI21X1 U3713 ( .A(n423), .B(n3616), .C(n600), .Y(n3379) );
  OAI21X1 U3714 ( .A(n422), .B(n3618), .C(n601), .Y(n3377) );
  OAI21X1 U3715 ( .A(n423), .B(n3620), .C(n602), .Y(n3375) );
  OAI21X1 U3716 ( .A(n422), .B(n3622), .C(n603), .Y(n3373) );
  OAI21X1 U3717 ( .A(n423), .B(n3624), .C(n604), .Y(n3371) );
  OAI21X1 U3718 ( .A(n422), .B(n3626), .C(n605), .Y(n3369) );
  OAI21X1 U3719 ( .A(n423), .B(n3628), .C(n606), .Y(n3367) );
  OAI21X1 U3720 ( .A(n3631), .B(n1695), .C(n421), .Y(n3630) );
  NAND3X1 U3721 ( .A(n3636), .B(net65987), .C(n3637), .Y(n3634) );
  AND2X1 U3722 ( .A(n3638), .B(n3639), .Y(n3636) );
  OAI21X1 U3723 ( .A(n1819), .B(net65992), .C(n480), .Y(n3365) );
  OAI21X1 U3724 ( .A(n3642), .B(n3643), .C(n481), .Y(n3363) );
  MUX2X1 U3725 ( .B(net65999), .A(n3646), .S(n1722), .Y(n3361) );
  NOR3X1 U3726 ( .A(n1404), .B(n1470), .C(n540), .Y(n3646) );
  NAND3X1 U3727 ( .A(n609), .B(net66007), .C(net82349), .Y(n3651) );
  NAND3X1 U3728 ( .A(n1518), .B(n3656), .C(n1348), .Y(n3648) );
  AOI22X1 U3729 ( .A(n3658), .B(n1717), .C(n3660), .D(n3661), .Y(n3657) );
  INVX1 U3730 ( .A(n1618), .Y(n3658) );
  INVX1 U3731 ( .A(n1695), .Y(n3656) );
  MUX2X1 U3732 ( .B(n3663), .A(n3664), .S(n1723), .Y(n3359) );
  NOR3X1 U3733 ( .A(n1407), .B(n1680), .C(n3667), .Y(n3664) );
  OAI21X1 U3734 ( .A(n1747), .B(n1726), .C(n3670), .Y(n3667) );
  NAND3X1 U3735 ( .A(n1717), .B(n1674), .C(n1741), .Y(n3671) );
  MUX2X1 U3736 ( .B(net66031), .A(n3676), .S(n1722), .Y(n3357) );
  NOR3X1 U3737 ( .A(n3677), .B(n1551), .C(n3679), .Y(n3676) );
  OAI21X1 U3738 ( .A(n1618), .B(n1717), .C(n1735), .Y(n3677) );
  MUX2X1 U3739 ( .B(n3681), .A(n3682), .S(n1723), .Y(n3355) );
  NOR3X1 U3740 ( .A(n1416), .B(n1473), .C(n1497), .Y(n3682) );
  NAND3X1 U3741 ( .A(n1674), .B(n1726), .C(n1741), .Y(n3662) );
  NAND3X1 U3742 ( .A(n1578), .B(n1651), .C(n3687), .Y(n3683) );
  NAND3X1 U3743 ( .A(n3688), .B(n1738), .C(n3689), .Y(n3353) );
  INVX1 U3744 ( .A(n1515), .Y(n3689) );
  OR2X1 U3745 ( .A(n1721), .B(n3691), .Y(n3688) );
  NAND3X1 U3746 ( .A(n842), .B(n3693), .C(n3694), .Y(n3647) );
  NOR3X1 U3747 ( .A(n3695), .B(n866), .C(n3696), .Y(n3694) );
  OR2X1 U3748 ( .A(n3697), .B(n3698), .Y(n3696) );
  OAI21X1 U3749 ( .A(n1701), .B(n1710), .C(n662), .Y(n3695) );
  NOR3X1 U3750 ( .A(n3701), .B(n1636), .C(n3703), .Y(n3693) );
  INVX1 U3751 ( .A(n1609), .Y(n3703) );
  AOI21X1 U3752 ( .A(n1741), .B(n1663), .C(n1239), .Y(n3692) );
  NAND3X1 U3753 ( .A(ready), .B(net66007), .C(n3709), .Y(n3707) );
  OAI21X1 U3754 ( .A(net66073), .B(n1819), .C(n482), .Y(n3351) );
  OAI21X1 U3755 ( .A(net65987), .B(n1819), .C(n483), .Y(n3349) );
  OAI21X1 U3756 ( .A(net66076), .B(n1820), .C(n484), .Y(n3347) );
  OAI21X1 U3757 ( .A(net66078), .B(n1820), .C(n485), .Y(n3345) );
  OAI21X1 U3758 ( .A(net66080), .B(n1819), .C(n486), .Y(n3343) );
  OAI21X1 U3759 ( .A(net66082), .B(n1819), .C(n487), .Y(n3341) );
  OAI21X1 U3760 ( .A(n1818), .B(net66084), .C(n488), .Y(n3339) );
  OAI21X1 U3761 ( .A(net66086), .B(n1820), .C(n489), .Y(n3337) );
  OAI21X1 U3762 ( .A(n1820), .B(net66088), .C(n490), .Y(n3335) );
  OAI21X1 U3763 ( .A(n1818), .B(net66090), .C(n491), .Y(n3333) );
  OAI21X1 U3764 ( .A(n1819), .B(net66092), .C(n492), .Y(n3331) );
  OAI21X1 U3765 ( .A(n1818), .B(net66094), .C(n493), .Y(n3329) );
  OAI21X1 U3766 ( .A(n1820), .B(net66096), .C(n494), .Y(n3327) );
  INVX1 U3767 ( .A(i[12]), .Y(net66096) );
  OAI21X1 U3768 ( .A(n1818), .B(net66098), .C(n495), .Y(n3325) );
  INVX1 U3769 ( .A(i[13]), .Y(net66098) );
  OAI21X1 U3770 ( .A(n1819), .B(net66100), .C(n496), .Y(n3323) );
  INVX1 U3771 ( .A(i[14]), .Y(net66100) );
  OAI21X1 U3772 ( .A(n1818), .B(net66102), .C(n497), .Y(n3321) );
  OAI21X1 U3773 ( .A(n1820), .B(net66104), .C(n498), .Y(n3319) );
  OAI21X1 U3774 ( .A(n1818), .B(net66106), .C(n499), .Y(n3317) );
  OAI21X1 U3775 ( .A(n1819), .B(net66108), .C(n500), .Y(n3315) );
  OAI21X1 U3776 ( .A(n1818), .B(net66110), .C(n501), .Y(n3313) );
  OAI21X1 U3777 ( .A(n1820), .B(net66112), .C(n502), .Y(n3311) );
  INVX1 U3778 ( .A(i[20]), .Y(net66112) );
  OAI21X1 U3779 ( .A(n1818), .B(net66114), .C(n503), .Y(n3309) );
  INVX1 U3780 ( .A(i[21]), .Y(net66114) );
  OAI21X1 U3781 ( .A(n1819), .B(net66116), .C(n504), .Y(n3307) );
  OAI21X1 U3782 ( .A(n1818), .B(n3733), .C(n505), .Y(n3305) );
  OAI21X1 U3783 ( .A(n1820), .B(n3735), .C(n506), .Y(n3303) );
  OAI21X1 U3784 ( .A(n1818), .B(n3737), .C(n507), .Y(n3301) );
  INVX1 U3785 ( .A(i[25]), .Y(n3737) );
  OAI21X1 U3786 ( .A(n1819), .B(n3739), .C(n508), .Y(n3299) );
  INVX1 U3787 ( .A(i[26]), .Y(n3739) );
  OAI21X1 U3788 ( .A(n1818), .B(n3741), .C(n509), .Y(n3297) );
  INVX1 U3789 ( .A(i[27]), .Y(n3741) );
  OAI21X1 U3790 ( .A(n1820), .B(n3743), .C(n510), .Y(n3295) );
  INVX1 U3791 ( .A(i[28]), .Y(n3743) );
  OAI21X1 U3792 ( .A(n1820), .B(n3745), .C(n511), .Y(n3293) );
  INVX1 U3793 ( .A(i[29]), .Y(n3745) );
  OAI21X1 U3794 ( .A(n1820), .B(n3747), .C(n941), .Y(n3291) );
  OAI21X1 U3795 ( .A(n852), .B(n1333), .C(n545), .Y(n3749) );
  AOI21X1 U3796 ( .A(net66063), .B(net66140), .C(n3755), .Y(n3754) );
  AOI22X1 U3797 ( .A(n1701), .B(n1683), .C(n3631), .D(n1657), .Y(n3752) );
  NAND3X1 U3798 ( .A(n3760), .B(n1304), .C(n1354), .Y(n3750) );
  AOI21X1 U3799 ( .A(net66062), .B(net66149), .C(n3763), .Y(n3762) );
  OAI21X1 U3800 ( .A(n3709), .B(n1654), .C(n668), .Y(n3763) );
  NAND3X1 U3801 ( .A(n3765), .B(n1531), .C(n3767), .Y(n3764) );
  INVX1 U3802 ( .A(n3768), .Y(n3709) );
  NAND3X1 U3803 ( .A(n3769), .B(i[1]), .C(n3770), .Y(n3768) );
  NAND3X1 U3804 ( .A(n3771), .B(n3770), .C(net66160), .Y(n3761) );
  NAND3X1 U3805 ( .A(n3774), .B(n3579), .C(n3775), .Y(n3772) );
  XNOR2X1 U3806 ( .A(n3776), .B(flag_bl_write), .Y(n3775) );
  INVX1 U3807 ( .A(i[30]), .Y(n3747) );
  OAI21X1 U3808 ( .A(n3779), .B(n3642), .C(n675), .Y(n3289) );
  INVX1 U3809 ( .A(clkcount[0]), .Y(n3779) );
  INVX1 U3810 ( .A(n3781), .Y(n3287) );
  AOI22X1 U3811 ( .A(n254), .B(n1788), .C(clkcount[1]), .D(n3782), .Y(n3781)
         );
  OAI21X1 U3812 ( .A(n3642), .B(n3783), .C(n678), .Y(n3285) );
  INVX1 U3813 ( .A(clkcount[2]), .Y(n3783) );
  OAI21X1 U3814 ( .A(n3642), .B(n3785), .C(n681), .Y(n3283) );
  INVX1 U3815 ( .A(clkcount[3]), .Y(n3785) );
  OAI21X1 U3816 ( .A(n3642), .B(n3787), .C(n684), .Y(n3281) );
  OAI21X1 U3817 ( .A(n3642), .B(n3789), .C(n687), .Y(n3279) );
  INVX1 U3818 ( .A(clkcount[5]), .Y(n3789) );
  OAI21X1 U3819 ( .A(n3642), .B(n3791), .C(n690), .Y(n3277) );
  INVX1 U3820 ( .A(clkcount[6]), .Y(n3791) );
  OAI21X1 U3821 ( .A(n3642), .B(n3793), .C(n693), .Y(n3275) );
  INVX1 U3822 ( .A(clkcount[7]), .Y(n3793) );
  OAI21X1 U3823 ( .A(n3642), .B(n3795), .C(n696), .Y(n3273) );
  OAI21X1 U3824 ( .A(n3642), .B(n3797), .C(n699), .Y(n3271) );
  INVX1 U3825 ( .A(clkcount[9]), .Y(n3797) );
  OAI21X1 U3826 ( .A(n3642), .B(n3799), .C(n702), .Y(n3269) );
  OAI21X1 U3827 ( .A(n3642), .B(n3801), .C(n706), .Y(n3267) );
  OAI21X1 U3828 ( .A(n3803), .B(n3642), .C(n709), .Y(n3265) );
  INVX1 U3829 ( .A(clkcount[12]), .Y(n3803) );
  OAI21X1 U3830 ( .A(n3642), .B(n3805), .C(n712), .Y(n3263) );
  OAI21X1 U3831 ( .A(n3642), .B(n3807), .C(n715), .Y(n3261) );
  OAI21X1 U3832 ( .A(n3642), .B(n3809), .C(n718), .Y(n3259) );
  OAI21X1 U3833 ( .A(n3642), .B(n3811), .C(n721), .Y(n3257) );
  OAI21X1 U3834 ( .A(n3642), .B(n3813), .C(n724), .Y(n3255) );
  OAI21X1 U3835 ( .A(n3642), .B(n3815), .C(n727), .Y(n3253) );
  OAI21X1 U3836 ( .A(n3642), .B(n3817), .C(n730), .Y(n3251) );
  OAI21X1 U3837 ( .A(n3642), .B(n3819), .C(n733), .Y(n3249) );
  OAI21X1 U3838 ( .A(n3642), .B(n3821), .C(n736), .Y(n3247) );
  OAI21X1 U3839 ( .A(n3642), .B(n3823), .C(n740), .Y(n3245) );
  OAI21X1 U3840 ( .A(n3642), .B(n3825), .C(n743), .Y(n3243) );
  OAI21X1 U3841 ( .A(n3642), .B(n3827), .C(n746), .Y(n3241) );
  OAI21X1 U3842 ( .A(n3642), .B(n3829), .C(n749), .Y(n3239) );
  OAI21X1 U3843 ( .A(n3642), .B(n3831), .C(n752), .Y(n3237) );
  OAI21X1 U3844 ( .A(n3642), .B(n3833), .C(n755), .Y(n3235) );
  OAI21X1 U3845 ( .A(n3642), .B(n3835), .C(n758), .Y(n3233) );
  OAI21X1 U3846 ( .A(n3642), .B(n3837), .C(n761), .Y(n3231) );
  OAI21X1 U3847 ( .A(n3642), .B(n3839), .C(n512), .Y(n3229) );
  AOI21X1 U3848 ( .A(n3841), .B(n1645), .C(n3782), .Y(n3645) );
  INVX1 U3849 ( .A(n1534), .Y(n3841) );
  OAI21X1 U3850 ( .A(n1729), .B(net66149), .C(n3843), .Y(n3642) );
  OAI21X1 U3851 ( .A(net66062), .B(n1534), .C(ready), .Y(n3843) );
  NAND3X1 U3852 ( .A(n3844), .B(n3778), .C(n1378), .Y(n3842) );
  OAI21X1 U3853 ( .A(state[4]), .B(n3847), .C(n1566), .Y(n3846) );
  NOR3X1 U3854 ( .A(n3756), .B(n3661), .C(n1599), .Y(n3778) );
  INVX1 U3855 ( .A(n1704), .Y(n3756) );
  INVX1 U3856 ( .A(n3698), .Y(n3844) );
  OAI21X1 U3857 ( .A(net66031), .B(n1566), .C(n3850), .Y(n3698) );
  MUX2X1 U3858 ( .B(state[3]), .A(n3851), .S(n3691), .Y(n3850) );
  NOR3X1 U3859 ( .A(n1437), .B(state[0]), .C(n3663), .Y(n3851) );
  NAND3X1 U3860 ( .A(state[4]), .B(state[0]), .C(state[1]), .Y(n3848) );
  INVX1 U3861 ( .A(n1729), .Y(net66062) );
  INVX1 U3862 ( .A(n1645), .Y(net66149) );
  NAND3X1 U3863 ( .A(i[5]), .B(n3855), .C(i[7]), .Y(n3854) );
  NAND3X1 U3864 ( .A(i[4]), .B(net66076), .C(n1668), .Y(n3853) );
  OAI21X1 U3865 ( .A(n3857), .B(n1602), .C(n3859), .Y(n3227) );
  OAI21X1 U3866 ( .A(n3860), .B(n3861), .C(ring_ptr[2]), .Y(n3859) );
  INVX1 U3867 ( .A(n1621), .Y(n3860) );
  MUX2X1 U3868 ( .B(n1639), .A(n1621), .S(ring_ptr[0]), .Y(n3225) );
  MUX2X1 U3869 ( .B(n3864), .A(n1602), .S(n3857), .Y(n3223) );
  INVX1 U3870 ( .A(ring_ptr[1]), .Y(n3857) );
  INVX1 U3871 ( .A(n3865), .Y(n3864) );
  OAI21X1 U3872 ( .A(n1639), .B(ring_ptr[0]), .C(n1621), .Y(n3865) );
  NAND3X1 U3873 ( .A(n1710), .B(n3866), .C(n1357), .Y(n3862) );
  AOI21X1 U3874 ( .A(n3868), .B(n3765), .C(n3861), .Y(n3867) );
  MUX2X1 U3875 ( .B(n1747), .A(n3869), .S(n3870), .Y(n3221) );
  AND2X1 U3876 ( .A(n1609), .B(n1690), .Y(n3870) );
  INVX1 U3877 ( .A(n3871), .Y(n3220) );
  MUX2X1 U3878 ( .B(buff_col_addr[0]), .A(CMD_data_out[0]), .S(n1750), .Y(
        n3871) );
  INVX1 U3879 ( .A(n3873), .Y(n3219) );
  MUX2X1 U3880 ( .B(buff_col_addr[1]), .A(CMD_data_out[1]), .S(n1750), .Y(
        n3873) );
  INVX1 U3881 ( .A(n3874), .Y(n3218) );
  MUX2X1 U3882 ( .B(buff_col_addr[2]), .A(CMD_data_out[2]), .S(n1750), .Y(
        n3874) );
  INVX1 U3883 ( .A(n3875), .Y(n3217) );
  MUX2X1 U3884 ( .B(buff_col_addr[3]), .A(CMD_data_out[3]), .S(n1750), .Y(
        n3875) );
  INVX1 U3885 ( .A(n3876), .Y(n3216) );
  MUX2X1 U3886 ( .B(buff_col_addr[4]), .A(CMD_data_out[4]), .S(n1750), .Y(
        n3876) );
  INVX1 U3887 ( .A(n3877), .Y(n3215) );
  MUX2X1 U3888 ( .B(buff_col_addr[5]), .A(CMD_data_out[5]), .S(n1750), .Y(
        n3877) );
  INVX1 U3889 ( .A(n3878), .Y(n3214) );
  MUX2X1 U3890 ( .B(buff_col_addr[6]), .A(CMD_data_out[6]), .S(n1750), .Y(
        n3878) );
  INVX1 U3891 ( .A(n3879), .Y(n3213) );
  MUX2X1 U3892 ( .B(buff_col_addr[7]), .A(CMD_data_out[7]), .S(n1750), .Y(
        n3879) );
  INVX1 U3893 ( .A(n3880), .Y(n3212) );
  MUX2X1 U3894 ( .B(buff_col_addr[8]), .A(CMD_data_out[8]), .S(n1750), .Y(
        n3880) );
  INVX1 U3895 ( .A(n3881), .Y(n3211) );
  MUX2X1 U3896 ( .B(buff_col_addr[9]), .A(CMD_data_out[9]), .S(n1750), .Y(
        n3881) );
  INVX1 U3897 ( .A(n3882), .Y(n3210) );
  MUX2X1 U3898 ( .B(buff_bank_addr[0]), .A(CMD_data_out[23]), .S(n1750), .Y(
        n3882) );
  INVX1 U3899 ( .A(n3883), .Y(n3209) );
  MUX2X1 U3900 ( .B(buff_bank_addr[1]), .A(CMD_data_out[24]), .S(n1750), .Y(
        n3883) );
  INVX1 U3901 ( .A(n3884), .Y(n3208) );
  MUX2X1 U3902 ( .B(buff_bank_addr[2]), .A(CMD_data_out[25]), .S(n1750), .Y(
        n3884) );
  NAND3X1 U3903 ( .A(n3776), .B(n3869), .C(n3579), .Y(n3633) );
  MUX2X1 U3904 ( .B(n1265), .A(n3886), .S(n3887), .Y(n3206) );
  AND2X1 U3905 ( .A(n783), .B(n1584), .Y(n3887) );
  NAND3X1 U3906 ( .A(CMD_data_out[31]), .B(CMD_data_out[33]), .C(n1360), .Y(
        n3888) );
  AOI21X1 U3907 ( .A(n3891), .B(n1713), .C(CMD_data_out[32]), .Y(n3890) );
  OR2X1 U3908 ( .A(n1726), .B(n1747), .Y(n3891) );
  INVX1 U3909 ( .A(flag_at_read), .Y(n3886) );
  INVX1 U3910 ( .A(n3892), .Y(n3204) );
  MUX2X1 U3911 ( .B(ras_bar), .A(n532), .S(n1671), .Y(n3892) );
  NAND3X1 U3912 ( .A(n530), .B(n1298), .C(net66289), .Y(n3893) );
  OAI21X1 U3913 ( .A(n3660), .B(n3708), .C(n3897), .Y(net66290) );
  AOI22X1 U3914 ( .A(n1686), .B(n858), .C(n1663), .D(n1741), .Y(n3896) );
  NAND3X1 U3915 ( .A(n1627), .B(n3899), .C(n1729), .Y(n3898) );
  INVX1 U3916 ( .A(n1741), .Y(n3899) );
  AOI21X1 U3917 ( .A(n3639), .B(n1521), .C(n1512), .Y(n3895) );
  INVX1 U3918 ( .A(n3902), .Y(n3202) );
  MUX2X1 U3919 ( .B(we_bar), .A(n533), .S(n1672), .Y(n3902) );
  NAND3X1 U3920 ( .A(n835), .B(n3905), .C(n3906), .Y(n3903) );
  INVX1 U3921 ( .A(n3907), .Y(n3906) );
  NAND3X1 U3922 ( .A(n1704), .B(n3708), .C(n1729), .Y(n3907) );
  OR2X1 U3923 ( .A(n1541), .B(n1630), .Y(n3708) );
  INVX1 U3924 ( .A(n1512), .Y(n3905) );
  NAND3X1 U3925 ( .A(n1713), .B(n1654), .C(n863), .Y(n3901) );
  AOI21X1 U3926 ( .A(n3911), .B(n1701), .C(n1515), .Y(n3910) );
  NAND3X1 U3927 ( .A(n1710), .B(n1698), .C(n1363), .Y(n3690) );
  AOI21X1 U3928 ( .A(n3914), .B(n1677), .C(n3697), .Y(n3913) );
  OAI21X1 U3929 ( .A(n1747), .B(n1726), .C(n478), .Y(n3697) );
  AOI21X1 U3930 ( .A(n1741), .B(n3917), .C(n3918), .Y(n3916) );
  AOI22X1 U3931 ( .A(n1686), .B(n3919), .C(n1741), .D(n1717), .Y(n3904) );
  OR2X1 U3932 ( .A(n3755), .B(n3661), .Y(n3919) );
  OAI21X1 U3933 ( .A(n3920), .B(n1615), .C(n3897), .Y(n3755) );
  OAI21X1 U3934 ( .A(net65987), .B(n1660), .C(n3923), .Y(n3897) );
  OAI21X1 U3935 ( .A(n1791), .B(net79420), .C(n943), .Y(n3200) );
  OAI21X1 U3936 ( .A(n1791), .B(net79440), .C(n944), .Y(n3198) );
  OAI21X1 U3937 ( .A(n1791), .B(net66325), .C(n945), .Y(n3196) );
  OAI21X1 U3938 ( .A(n1791), .B(n3928), .C(n948), .Y(n3190) );
  OAI21X1 U3939 ( .A(n1791), .B(n3930), .C(n949), .Y(n3188) );
  OAI21X1 U3940 ( .A(n1791), .B(net66339), .C(n952), .Y(n3182) );
  INVX1 U3941 ( .A(j[9]), .Y(net66339) );
  OAI21X1 U3942 ( .A(n1791), .B(n3933), .C(n959), .Y(n3168) );
  OAI21X1 U3943 ( .A(n1791), .B(n3935), .C(n960), .Y(n3166) );
  OAI21X1 U3944 ( .A(n1791), .B(n3937), .C(n961), .Y(n3164) );
  OAI21X1 U3945 ( .A(n1791), .B(n3939), .C(n962), .Y(n3162) );
  OAI21X1 U3946 ( .A(n1791), .B(n3941), .C(n963), .Y(n3160) );
  OAI21X1 U3947 ( .A(n1791), .B(n3943), .C(n964), .Y(n3158) );
  OAI21X1 U3948 ( .A(n1791), .B(n3945), .C(n965), .Y(n3156) );
  OAI21X1 U3949 ( .A(n1791), .B(net66381), .C(n514), .Y(n3140) );
  INVX1 U3950 ( .A(j[30]), .Y(net66381) );
  OAI21X1 U3951 ( .A(n1791), .B(net66383), .C(n515), .Y(n3138) );
  OAI21X1 U3952 ( .A(net66385), .B(n1738), .C(n1612), .Y(n3925) );
  INVX1 U3953 ( .A(j[31]), .Y(net66383) );
  MUX2X1 U3954 ( .B(buff_data[1]), .A(n577), .S(n2162), .Y(n3951) );
  MUX2X1 U3955 ( .B(buff_data[4]), .A(n576), .S(n2162), .Y(n3954) );
  MUX2X1 U3956 ( .B(buff_data[5]), .A(n569), .S(n2162), .Y(n3955) );
  MUX2X1 U3957 ( .B(buff_data[6]), .A(n570), .S(n2162), .Y(n3956) );
  MUX2X1 U3958 ( .B(buff_data[7]), .A(n578), .S(n2179), .Y(n3957) );
  MUX2X1 U3959 ( .B(buff_data[8]), .A(n566), .S(n2179), .Y(n3958) );
  MUX2X1 U3960 ( .B(buff_data[10]), .A(n564), .S(n2162), .Y(n3959) );
  MUX2X1 U3961 ( .B(buff_data[11]), .A(n571), .S(n2162), .Y(n3960) );
  MUX2X1 U3962 ( .B(buff_data[12]), .A(n572), .S(n2179), .Y(n3961) );
  MUX2X1 U3963 ( .B(buff_data[13]), .A(n579), .S(n2179), .Y(n3962) );
  MUX2X1 U3964 ( .B(buff_data[16]), .A(n573), .S(n190), .Y(n3964) );
  MUX2X1 U3965 ( .B(buff_data[17]), .A(n577), .S(n2181), .Y(n3965) );
  MUX2X1 U3966 ( .B(buff_data[19]), .A(n568), .S(n2049), .Y(n3966) );
  MUX2X1 U3967 ( .B(buff_data[21]), .A(n569), .S(n168), .Y(n3967) );
  MUX2X1 U3968 ( .B(buff_data[22]), .A(n570), .S(n191), .Y(n3968) );
  MUX2X1 U3969 ( .B(buff_data[23]), .A(n578), .S(n192), .Y(n3969) );
  MUX2X1 U3970 ( .B(buff_data[24]), .A(n566), .S(n169), .Y(n3970) );
  MUX2X1 U3971 ( .B(buff_data[26]), .A(n564), .S(n369), .Y(n3971) );
  MUX2X1 U3972 ( .B(buff_data[27]), .A(n571), .S(n2181), .Y(n3972) );
  MUX2X1 U3973 ( .B(buff_data[28]), .A(n572), .S(n189), .Y(n3973) );
  MUX2X1 U3974 ( .B(buff_data[30]), .A(n567), .S(n167), .Y(n3974) );
  MUX2X1 U3975 ( .B(buff_data[32]), .A(n573), .S(net79605), .Y(n3975) );
  MUX2X1 U3976 ( .B(buff_data[33]), .A(n577), .S(net79605), .Y(n3976) );
  MUX2X1 U3977 ( .B(buff_data[34]), .A(n574), .S(n336), .Y(n3977) );
  MUX2X1 U3978 ( .B(buff_data[35]), .A(n568), .S(n194), .Y(n3978) );
  MUX2X1 U3979 ( .B(buff_data[36]), .A(n576), .S(net79605), .Y(n3979) );
  MUX2X1 U3980 ( .B(buff_data[37]), .A(n569), .S(n193), .Y(n3980) );
  MUX2X1 U3981 ( .B(buff_data[38]), .A(n570), .S(n155), .Y(n3981) );
  MUX2X1 U3982 ( .B(buff_data[39]), .A(n578), .S(net79605), .Y(n3982) );
  MUX2X1 U3983 ( .B(buff_data[40]), .A(n566), .S(n53), .Y(n3983) );
  MUX2X1 U3984 ( .B(buff_data[41]), .A(n565), .S(n46), .Y(n3984) );
  MUX2X1 U3985 ( .B(buff_data[42]), .A(n564), .S(n157), .Y(n3985) );
  MUX2X1 U3986 ( .B(buff_data[43]), .A(n571), .S(n68), .Y(n3986) );
  MUX2X1 U3987 ( .B(buff_data[44]), .A(n572), .S(n158), .Y(n3987) );
  MUX2X1 U3988 ( .B(buff_data[45]), .A(n579), .S(n38), .Y(n3988) );
  MUX2X1 U3989 ( .B(buff_data[46]), .A(n567), .S(n156), .Y(n3989) );
  MUX2X1 U3990 ( .B(buff_data[47]), .A(n575), .S(n67), .Y(n3990) );
  MUX2X1 U3991 ( .B(buff_data[48]), .A(n573), .S(n199), .Y(n3991) );
  MUX2X1 U3992 ( .B(buff_data[49]), .A(n577), .S(n2180), .Y(n3992) );
  MUX2X1 U3993 ( .B(buff_data[50]), .A(n574), .S(n182), .Y(n3993) );
  MUX2X1 U3994 ( .B(buff_data[51]), .A(n568), .S(n165), .Y(n3994) );
  MUX2X1 U3995 ( .B(buff_data[52]), .A(n576), .S(n183), .Y(n3995) );
  MUX2X1 U3996 ( .B(buff_data[53]), .A(n569), .S(n196), .Y(n3996) );
  MUX2X1 U3997 ( .B(buff_data[54]), .A(n570), .S(n197), .Y(n3997) );
  NAND3X1 U3998 ( .A(n3866), .B(n1584), .C(n1366), .Y(n3079) );
  AOI21X1 U3999 ( .A(n3911), .B(n3999), .C(n3861), .Y(n3998) );
  INVX1 U4000 ( .A(n1639), .Y(n3861) );
  NAND3X1 U4001 ( .A(n4001), .B(n3999), .C(flag_at_read), .Y(n3889) );
  INVX1 U4002 ( .A(n1710), .Y(n4001) );
  INVX1 U4003 ( .A(n1636), .Y(n3866) );
  MUX2X1 U4004 ( .B(buff_data[55]), .A(n578), .S(n164), .Y(n4002) );
  MUX2X1 U4005 ( .B(buff_data[56]), .A(n566), .S(n198), .Y(n4003) );
  MUX2X1 U4006 ( .B(buff_data[57]), .A(n565), .S(n2180), .Y(n4004) );
  MUX2X1 U4007 ( .B(buff_data[58]), .A(n564), .S(n42), .Y(n4005) );
  OAI21X1 U4008 ( .A(flag_bl_read), .B(n1698), .C(n672), .Y(n3073) );
  AOI21X1 U4009 ( .A(n1701), .B(n1683), .C(n2439), .Y(n4006) );
  MUX2X1 U4010 ( .B(buff_data[59]), .A(n571), .S(n43), .Y(n4007) );
  MUX2X1 U4011 ( .B(buff_data[60]), .A(n572), .S(n2180), .Y(n4008) );
  MUX2X1 U4012 ( .B(buff_data[61]), .A(n579), .S(n2180), .Y(n4009) );
  MUX2X1 U4013 ( .B(buff_data[62]), .A(n567), .S(n2180), .Y(n4010) );
  MUX2X1 U4014 ( .B(buff_data[65]), .A(n577), .S(n124), .Y(n4013) );
  MUX2X1 U4015 ( .B(buff_data[66]), .A(n574), .S(n1953), .Y(n4014) );
  MUX2X1 U4016 ( .B(buff_data[68]), .A(n576), .S(n291), .Y(n4016) );
  MUX2X1 U4017 ( .B(buff_data[70]), .A(n570), .S(n1927), .Y(n4017) );
  MUX2X1 U4018 ( .B(buff_data[72]), .A(n566), .S(n215), .Y(n4019) );
  MUX2X1 U4019 ( .B(buff_data[73]), .A(n565), .S(n360), .Y(n4020) );
  MUX2X1 U4020 ( .B(buff_data[74]), .A(n564), .S(n360), .Y(n4021) );
  MUX2X1 U4021 ( .B(buff_data[75]), .A(n571), .S(n2178), .Y(n4022) );
  MUX2X1 U4022 ( .B(buff_data[76]), .A(n572), .S(n1927), .Y(n4023) );
  MUX2X1 U4023 ( .B(buff_data[77]), .A(n579), .S(n215), .Y(n4024) );
  MUX2X1 U4024 ( .B(buff_data[78]), .A(n567), .S(n1953), .Y(n4025) );
  MUX2X1 U4025 ( .B(buff_data[86]), .A(n570), .S(n223), .Y(n4026) );
  MUX2X1 U4026 ( .B(buff_data[87]), .A(n578), .S(n2078), .Y(n4027) );
  MUX2X1 U4027 ( .B(buff_data[88]), .A(n566), .S(n300), .Y(n4028) );
  MUX2X1 U4028 ( .B(buff_data[89]), .A(n565), .S(n306), .Y(n4029) );
  MUX2X1 U4029 ( .B(buff_data[90]), .A(n564), .S(n71), .Y(n4030) );
  MUX2X1 U4030 ( .B(buff_data[91]), .A(n571), .S(n379), .Y(n4031) );
  MUX2X1 U4031 ( .B(buff_data[92]), .A(n572), .S(n351), .Y(n4032) );
  MUX2X1 U4032 ( .B(buff_data[93]), .A(n579), .S(n222), .Y(n4033) );
  MUX2X1 U4033 ( .B(buff_data[94]), .A(n567), .S(n436), .Y(n4034) );
  MUX2X1 U4034 ( .B(buff_data[95]), .A(n575), .S(n306), .Y(n4035) );
  MUX2X1 U4035 ( .B(buff_data[80]), .A(n573), .S(n352), .Y(n4036) );
  MUX2X1 U4036 ( .B(buff_data[81]), .A(n577), .S(n306), .Y(n4037) );
  MUX2X1 U4037 ( .B(buff_data[82]), .A(n574), .S(n306), .Y(n4038) );
  MUX2X1 U4038 ( .B(buff_data[83]), .A(n568), .S(n435), .Y(n4039) );
  MUX2X1 U4039 ( .B(buff_data[84]), .A(n576), .S(n209), .Y(n4040) );
  OAI21X1 U4040 ( .A(n1738), .B(net66499), .C(n972), .Y(n3036) );
  MUX2X1 U4041 ( .B(buff_data[96]), .A(n573), .S(n368), .Y(n4042) );
  MUX2X1 U4042 ( .B(buff_data[98]), .A(n574), .S(n212), .Y(n4044) );
  MUX2X1 U4043 ( .B(buff_data[99]), .A(n568), .S(n368), .Y(n4045) );
  MUX2X1 U4044 ( .B(buff_data[100]), .A(n576), .S(n186), .Y(n4046) );
  MUX2X1 U4045 ( .B(buff_data[101]), .A(n569), .S(n225), .Y(n4047) );
  MUX2X1 U4046 ( .B(buff_data[102]), .A(n570), .S(n368), .Y(n4048) );
  MUX2X1 U4047 ( .B(buff_data[104]), .A(n566), .S(n4043), .Y(n4049) );
  MUX2X1 U4048 ( .B(buff_data[105]), .A(n565), .S(n368), .Y(n4050) );
  MUX2X1 U4049 ( .B(buff_data[106]), .A(n564), .S(n186), .Y(n4051) );
  MUX2X1 U4050 ( .B(buff_data[107]), .A(n571), .S(n299), .Y(n4052) );
  MUX2X1 U4051 ( .B(buff_data[108]), .A(n572), .S(n368), .Y(n4053) );
  MUX2X1 U4052 ( .B(buff_data[110]), .A(n567), .S(n211), .Y(n4054) );
  MUX2X1 U4053 ( .B(buff_data[111]), .A(n575), .S(n224), .Y(n4055) );
  MUX2X1 U4054 ( .B(buff_data[112]), .A(n573), .S(n290), .Y(n4057) );
  MUX2X1 U4055 ( .B(buff_data[113]), .A(n577), .S(n286), .Y(n4058) );
  MUX2X1 U4056 ( .B(buff_data[114]), .A(n574), .S(net80376), .Y(n4059) );
  MUX2X1 U4057 ( .B(buff_data[115]), .A(n568), .S(n303), .Y(n4060) );
  MUX2X1 U4058 ( .B(buff_data[116]), .A(n576), .S(net80376), .Y(n4061) );
  MUX2X1 U4059 ( .B(buff_data[117]), .A(n569), .S(n289), .Y(n4062) );
  MUX2X1 U4060 ( .B(buff_data[118]), .A(n570), .S(net80376), .Y(n4063) );
  MUX2X1 U4061 ( .B(buff_data[119]), .A(n578), .S(n288), .Y(n4064) );
  MUX2X1 U4062 ( .B(buff_data[120]), .A(n566), .S(n298), .Y(n4065) );
  MUX2X1 U4063 ( .B(buff_data[121]), .A(n565), .S(n304), .Y(n4066) );
  MUX2X1 U4064 ( .B(buff_data[122]), .A(n564), .S(n333), .Y(n4067) );
  MUX2X1 U4065 ( .B(buff_data[123]), .A(n571), .S(net80376), .Y(n4068) );
  MUX2X1 U4066 ( .B(buff_data[124]), .A(n572), .S(n332), .Y(n4069) );
  MUX2X1 U4067 ( .B(buff_data[125]), .A(n579), .S(net80376), .Y(n4070) );
  MUX2X1 U4068 ( .B(buff_data[126]), .A(n567), .S(net79593), .Y(n4071) );
  MUX2X1 U4069 ( .B(buff_data[128]), .A(n573), .S(n1), .Y(n4072) );
  MUX2X1 U4070 ( .B(buff_data[129]), .A(n577), .S(n81), .Y(n4073) );
  MUX2X1 U4071 ( .B(buff_data[130]), .A(n574), .S(n2191), .Y(n4074) );
  MUX2X1 U4072 ( .B(buff_data[131]), .A(n568), .S(n2191), .Y(n4075) );
  MUX2X1 U4073 ( .B(buff_data[132]), .A(n576), .S(n2191), .Y(n4076) );
  MUX2X1 U4074 ( .B(buff_data[133]), .A(n569), .S(n2191), .Y(n4077) );
  MUX2X1 U4075 ( .B(buff_data[134]), .A(n570), .S(n81), .Y(n4078) );
  MUX2X1 U4076 ( .B(buff_data[135]), .A(n578), .S(n2191), .Y(n4079) );
  MUX2X1 U4077 ( .B(buff_data[136]), .A(n566), .S(n2191), .Y(n4080) );
  MUX2X1 U4078 ( .B(buff_data[137]), .A(n565), .S(n2191), .Y(n4081) );
  MUX2X1 U4079 ( .B(buff_data[138]), .A(n564), .S(n1), .Y(n4082) );
  MUX2X1 U4080 ( .B(buff_data[139]), .A(n571), .S(n1607), .Y(n4083) );
  MUX2X1 U4081 ( .B(buff_data[140]), .A(n572), .S(n2191), .Y(n4084) );
  MUX2X1 U4082 ( .B(buff_data[141]), .A(n579), .S(n2191), .Y(n4085) );
  MUX2X1 U4083 ( .B(buff_data[142]), .A(n567), .S(n2191), .Y(n4086) );
  MUX2X1 U4084 ( .B(buff_data[143]), .A(n575), .S(n1607), .Y(n4087) );
  MUX2X1 U4085 ( .B(buff_data[144]), .A(n573), .S(n2128), .Y(n4088) );
  MUX2X1 U4086 ( .B(buff_data[146]), .A(n574), .S(n162), .Y(n4089) );
  MUX2X1 U4087 ( .B(buff_data[147]), .A(n568), .S(n432), .Y(n4090) );
  MUX2X1 U4088 ( .B(buff_data[148]), .A(n576), .S(n133), .Y(n4091) );
  MUX2X1 U4089 ( .B(buff_data[149]), .A(n569), .S(n146), .Y(n4092) );
  MUX2X1 U4090 ( .B(buff_data[150]), .A(n570), .S(n24), .Y(n4093) );
  MUX2X1 U4091 ( .B(buff_data[151]), .A(n578), .S(n176), .Y(n4094) );
  MUX2X1 U4092 ( .B(buff_data[152]), .A(n566), .S(n135), .Y(n4095) );
  MUX2X1 U4093 ( .B(buff_data[153]), .A(n565), .S(n154), .Y(n4096) );
  MUX2X1 U4094 ( .B(buff_data[155]), .A(n571), .S(n134), .Y(n4097) );
  MUX2X1 U4095 ( .B(buff_data[156]), .A(n572), .S(n21), .Y(n4098) );
  MUX2X1 U4096 ( .B(buff_data[157]), .A(n579), .S(n177), .Y(n4099) );
  MUX2X1 U4097 ( .B(buff_data[158]), .A(n567), .S(n161), .Y(n4100) );
  MUX2X1 U4098 ( .B(buff_data[159]), .A(n575), .S(n2197), .Y(n4101) );
  MUX2X1 U4099 ( .B(buff_data[160]), .A(n573), .S(n12), .Y(n4102) );
  MUX2X1 U4100 ( .B(buff_data[162]), .A(n574), .S(net80723), .Y(n4103) );
  MUX2X1 U4101 ( .B(buff_data[164]), .A(n576), .S(net80723), .Y(n4104) );
  MUX2X1 U4102 ( .B(buff_data[165]), .A(n569), .S(net79534), .Y(n4105) );
  MUX2X1 U4103 ( .B(buff_data[166]), .A(n570), .S(net79534), .Y(n4106) );
  MUX2X1 U4104 ( .B(buff_data[167]), .A(n578), .S(n75), .Y(n4107) );
  MUX2X1 U4105 ( .B(buff_data[169]), .A(n565), .S(n76), .Y(n4108) );
  MUX2X1 U4106 ( .B(buff_data[171]), .A(n571), .S(net80382), .Y(n4109) );
  MUX2X1 U4107 ( .B(buff_data[174]), .A(n567), .S(net80463), .Y(n4110) );
  MUX2X1 U4108 ( .B(buff_data[175]), .A(n575), .S(net80747), .Y(n4111) );
  MUX2X1 U4109 ( .B(buff_data[187]), .A(n571), .S(n345), .Y(n4113) );
  MUX2X1 U4110 ( .B(buff_data[188]), .A(n572), .S(n106), .Y(n4114) );
  MUX2X1 U4111 ( .B(buff_data[189]), .A(n579), .S(n84), .Y(n4115) );
  MUX2X1 U4112 ( .B(buff_data[191]), .A(n575), .S(n83), .Y(n4117) );
  MUX2X1 U4113 ( .B(buff_data[179]), .A(n568), .S(n386), .Y(n4118) );
  MUX2X1 U4114 ( .B(buff_data[180]), .A(n576), .S(n345), .Y(n4119) );
  MUX2X1 U4115 ( .B(buff_data[181]), .A(n569), .S(n343), .Y(n4120) );
  MUX2X1 U4116 ( .B(buff_data[182]), .A(n570), .S(n1816), .Y(n4121) );
  MUX2X1 U4117 ( .B(buff_data[183]), .A(n578), .S(n106), .Y(n4122) );
  MUX2X1 U4118 ( .B(buff_data[184]), .A(n566), .S(n342), .Y(n4123) );
  MUX2X1 U4119 ( .B(buff_data[192]), .A(n573), .S(net82427), .Y(n4124) );
  MUX2X1 U4120 ( .B(buff_data[194]), .A(n574), .S(net82428), .Y(n4125) );
  MUX2X1 U4121 ( .B(buff_data[202]), .A(n564), .S(n217), .Y(n4128) );
  MUX2X1 U4122 ( .B(buff_data[204]), .A(n572), .S(n2127), .Y(n4129) );
  MUX2X1 U4123 ( .B(buff_data[205]), .A(n579), .S(n85), .Y(n4130) );
  MUX2X1 U4124 ( .B(buff_data[208]), .A(n573), .S(n97), .Y(n4132) );
  MUX2X1 U4125 ( .B(buff_data[209]), .A(n577), .S(n4133), .Y(n4134) );
  MUX2X1 U4126 ( .B(buff_data[210]), .A(n574), .S(n57), .Y(n4135) );
  MUX2X1 U4127 ( .B(buff_data[211]), .A(n568), .S(n4133), .Y(n4136) );
  MUX2X1 U4128 ( .B(buff_data[212]), .A(n576), .S(n57), .Y(n4137) );
  MUX2X1 U4129 ( .B(buff_data[213]), .A(n569), .S(n2186), .Y(n4138) );
  MUX2X1 U4130 ( .B(buff_data[214]), .A(n570), .S(n4133), .Y(n4139) );
  MUX2X1 U4131 ( .B(buff_data[215]), .A(n578), .S(n97), .Y(n4140) );
  MUX2X1 U4132 ( .B(buff_data[216]), .A(n566), .S(n2186), .Y(n4141) );
  MUX2X1 U4133 ( .B(buff_data[217]), .A(n565), .S(n97), .Y(n4142) );
  MUX2X1 U4134 ( .B(buff_data[218]), .A(n564), .S(n4133), .Y(n4143) );
  MUX2X1 U4135 ( .B(buff_data[219]), .A(n571), .S(n4133), .Y(n4144) );
  MUX2X1 U4136 ( .B(buff_data[220]), .A(n572), .S(n2187), .Y(n4145) );
  MUX2X1 U4137 ( .B(buff_data[221]), .A(n579), .S(n97), .Y(n4146) );
  MUX2X1 U4138 ( .B(buff_data[222]), .A(n567), .S(n2187), .Y(n4147) );
  MUX2X1 U4139 ( .B(buff_data[223]), .A(n575), .S(n97), .Y(n4148) );
  MUX2X1 U4140 ( .B(buff_data[228]), .A(n576), .S(n402), .Y(n4151) );
  MUX2X1 U4141 ( .B(buff_data[239]), .A(n575), .S(n338), .Y(n4152) );
  MUX2X1 U4142 ( .B(buff_data[240]), .A(n573), .S(n35), .Y(n4153) );
  MUX2X1 U4143 ( .B(buff_data[241]), .A(n577), .S(n400), .Y(n4154) );
  MUX2X1 U4144 ( .B(buff_data[243]), .A(n568), .S(n205), .Y(n4155) );
  MUX2X1 U4145 ( .B(buff_data[245]), .A(n569), .S(n91), .Y(n4156) );
  MUX2X1 U4146 ( .B(buff_data[246]), .A(n570), .S(n87), .Y(n4157) );
  MUX2X1 U4147 ( .B(buff_data[247]), .A(n578), .S(n348), .Y(n4158) );
  MUX2X1 U4148 ( .B(buff_data[248]), .A(n566), .S(n305), .Y(n4159) );
  MUX2X1 U4149 ( .B(buff_data[249]), .A(n565), .S(n88), .Y(n4160) );
  MUX2X1 U4150 ( .B(buff_data[251]), .A(n571), .S(net79510), .Y(n4161) );
  MUX2X1 U4151 ( .B(buff_data[252]), .A(n572), .S(n88), .Y(n4162) );
  MUX2X1 U4152 ( .B(buff_data[254]), .A(n567), .S(n87), .Y(n4163) );
  MUX2X1 U4153 ( .B(buff_data[256]), .A(n573), .S(n2190), .Y(n4164) );
  MUX2X1 U4154 ( .B(buff_data[257]), .A(n577), .S(n2189), .Y(n4166) );
  MUX2X1 U4155 ( .B(buff_data[258]), .A(n574), .S(n4165), .Y(n4167) );
  MUX2X1 U4156 ( .B(buff_data[259]), .A(n568), .S(n2015), .Y(n4168) );
  MUX2X1 U4157 ( .B(buff_data[260]), .A(n576), .S(n2189), .Y(n4169) );
  MUX2X1 U4158 ( .B(buff_data[261]), .A(n569), .S(n2015), .Y(n4170) );
  MUX2X1 U4159 ( .B(buff_data[262]), .A(n570), .S(n39), .Y(n4171) );
  MUX2X1 U4160 ( .B(buff_data[263]), .A(n578), .S(n2189), .Y(n4172) );
  MUX2X1 U4161 ( .B(buff_data[264]), .A(n566), .S(n4165), .Y(n4173) );
  MUX2X1 U4162 ( .B(buff_data[265]), .A(n565), .S(n2190), .Y(n4174) );
  MUX2X1 U4163 ( .B(buff_data[266]), .A(n564), .S(n4165), .Y(n4175) );
  MUX2X1 U4164 ( .B(buff_data[267]), .A(n571), .S(n2190), .Y(n4176) );
  MUX2X1 U4165 ( .B(buff_data[268]), .A(n572), .S(n2015), .Y(n4177) );
  MUX2X1 U4166 ( .B(buff_data[269]), .A(n579), .S(n4165), .Y(n4178) );
  MUX2X1 U4167 ( .B(buff_data[270]), .A(n567), .S(n39), .Y(n4179) );
  MUX2X1 U4168 ( .B(buff_data[271]), .A(n575), .S(n39), .Y(n4180) );
  MUX2X1 U4169 ( .B(buff_data[285]), .A(n579), .S(n2016), .Y(n4181) );
  MUX2X1 U4170 ( .B(buff_data[286]), .A(n567), .S(n372), .Y(n4182) );
  MUX2X1 U4171 ( .B(buff_data[273]), .A(n577), .S(n2037), .Y(n4184) );
  MUX2X1 U4172 ( .B(buff_data[275]), .A(n568), .S(n1996), .Y(n4186) );
  MUX2X1 U4173 ( .B(buff_data[277]), .A(n569), .S(n2196), .Y(n4187) );
  MUX2X1 U4174 ( .B(buff_data[281]), .A(n565), .S(n1996), .Y(n4188) );
  MUX2X1 U4175 ( .B(buff_data[282]), .A(n564), .S(n372), .Y(n4189) );
  MUX2X1 U4176 ( .B(buff_data[283]), .A(n571), .S(n2196), .Y(n4190) );
  MUX2X1 U4177 ( .B(buff_data[289]), .A(n577), .S(n367), .Y(n4191) );
  MUX2X1 U4178 ( .B(buff_data[290]), .A(n574), .S(n141), .Y(n4192) );
  MUX2X1 U4179 ( .B(buff_data[291]), .A(n568), .S(n141), .Y(n4193) );
  MUX2X1 U4180 ( .B(buff_data[292]), .A(n576), .S(n171), .Y(n4194) );
  MUX2X1 U4181 ( .B(buff_data[293]), .A(n569), .S(n172), .Y(n4195) );
  MUX2X1 U4182 ( .B(buff_data[294]), .A(n570), .S(net82191), .Y(n4196) );
  MUX2X1 U4183 ( .B(buff_data[296]), .A(n566), .S(n172), .Y(n4197) );
  MUX2X1 U4184 ( .B(buff_data[297]), .A(n565), .S(net82191), .Y(n4198) );
  MUX2X1 U4185 ( .B(buff_data[298]), .A(n564), .S(n171), .Y(n4199) );
  MUX2X1 U4186 ( .B(buff_data[299]), .A(n571), .S(n185), .Y(n4200) );
  MUX2X1 U4187 ( .B(buff_data[300]), .A(n572), .S(n185), .Y(n4201) );
  MUX2X1 U4188 ( .B(buff_data[302]), .A(n567), .S(net80661), .Y(n4202) );
  MUX2X1 U4189 ( .B(buff_data[303]), .A(n575), .S(net80661), .Y(n4203) );
  MUX2X1 U4190 ( .B(buff_data[304]), .A(n573), .S(n204), .Y(n4204) );
  MUX2X1 U4191 ( .B(buff_data[305]), .A(n577), .S(n353), .Y(n4206) );
  MUX2X1 U4192 ( .B(buff_data[306]), .A(n574), .S(n366), .Y(n4207) );
  MUX2X1 U4193 ( .B(buff_data[307]), .A(n568), .S(n308), .Y(n4208) );
  MUX2X1 U4194 ( .B(buff_data[308]), .A(n576), .S(n294), .Y(n4209) );
  MUX2X1 U4195 ( .B(buff_data[309]), .A(n569), .S(n308), .Y(n4210) );
  MUX2X1 U4196 ( .B(buff_data[310]), .A(n570), .S(n174), .Y(n4211) );
  MUX2X1 U4197 ( .B(buff_data[312]), .A(n566), .S(n353), .Y(n4212) );
  MUX2X1 U4198 ( .B(buff_data[313]), .A(n565), .S(n204), .Y(n4213) );
  MUX2X1 U4199 ( .B(buff_data[314]), .A(n564), .S(n366), .Y(n4214) );
  MUX2X1 U4200 ( .B(buff_data[317]), .A(n579), .S(n2185), .Y(n4215) );
  MUX2X1 U4201 ( .B(buff_data[318]), .A(n567), .S(n2185), .Y(n4216) );
  MUX2X1 U4202 ( .B(buff_data[320]), .A(n573), .S(n1991), .Y(n4217) );
  MUX2X1 U4203 ( .B(buff_data[321]), .A(n577), .S(n331), .Y(n4219) );
  MUX2X1 U4204 ( .B(buff_data[322]), .A(n574), .S(n440), .Y(n4220) );
  MUX2X1 U4205 ( .B(buff_data[324]), .A(n576), .S(n2013), .Y(n4221) );
  MUX2X1 U4206 ( .B(buff_data[325]), .A(n569), .S(n2038), .Y(n4222) );
  MUX2X1 U4207 ( .B(buff_data[326]), .A(n570), .S(n1991), .Y(n4223) );
  MUX2X1 U4208 ( .B(buff_data[327]), .A(n578), .S(n2039), .Y(n4224) );
  MUX2X1 U4209 ( .B(buff_data[329]), .A(n565), .S(n1904), .Y(n4225) );
  MUX2X1 U4210 ( .B(buff_data[330]), .A(n564), .S(n2013), .Y(n4226) );
  MUX2X1 U4211 ( .B(buff_data[332]), .A(n572), .S(n1904), .Y(n4227) );
  MUX2X1 U4212 ( .B(buff_data[334]), .A(n567), .S(n331), .Y(n4228) );
  MUX2X1 U4213 ( .B(buff_data[335]), .A(n575), .S(n440), .Y(n4229) );
  MUX2X1 U4214 ( .B(buff_data[336]), .A(n573), .S(n4231), .Y(n4230) );
  MUX2X1 U4215 ( .B(buff_data[337]), .A(n577), .S(n4231), .Y(n4232) );
  MUX2X1 U4216 ( .B(buff_data[338]), .A(n574), .S(n2182), .Y(n4233) );
  MUX2X1 U4217 ( .B(buff_data[339]), .A(n568), .S(n2182), .Y(n4234) );
  MUX2X1 U4218 ( .B(buff_data[340]), .A(n576), .S(n4231), .Y(n4235) );
  MUX2X1 U4219 ( .B(buff_data[341]), .A(n569), .S(n1995), .Y(n4236) );
  MUX2X1 U4220 ( .B(buff_data[342]), .A(n570), .S(n4231), .Y(n4237) );
  MUX2X1 U4221 ( .B(buff_data[343]), .A(n578), .S(n2182), .Y(n4238) );
  MUX2X1 U4222 ( .B(buff_data[344]), .A(n566), .S(n2183), .Y(n4239) );
  MUX2X1 U4223 ( .B(buff_data[345]), .A(n565), .S(n2182), .Y(n4240) );
  MUX2X1 U4224 ( .B(buff_data[346]), .A(n564), .S(n2183), .Y(n4241) );
  MUX2X1 U4225 ( .B(buff_data[347]), .A(n571), .S(n2183), .Y(n4242) );
  MUX2X1 U4226 ( .B(buff_data[348]), .A(n572), .S(n1995), .Y(n4243) );
  MUX2X1 U4227 ( .B(buff_data[349]), .A(n579), .S(n1995), .Y(n4244) );
  MUX2X1 U4228 ( .B(buff_data[350]), .A(n567), .S(n1995), .Y(n4245) );
  MUX2X1 U4229 ( .B(buff_data[351]), .A(n575), .S(n1995), .Y(n4246) );
  MUX2X1 U4230 ( .B(buff_data[353]), .A(n577), .S(n45), .Y(n4247) );
  MUX2X1 U4231 ( .B(buff_data[354]), .A(n574), .S(n2040), .Y(n4248) );
  MUX2X1 U4232 ( .B(buff_data[355]), .A(n568), .S(n125), .Y(n4249) );
  MUX2X1 U4233 ( .B(buff_data[356]), .A(n576), .S(n2022), .Y(n4250) );
  MUX2X1 U4234 ( .B(buff_data[357]), .A(n569), .S(n45), .Y(n4251) );
  MUX2X1 U4235 ( .B(buff_data[359]), .A(n578), .S(n60), .Y(n4252) );
  MUX2X1 U4236 ( .B(buff_data[360]), .A(n566), .S(n2040), .Y(n4253) );
  MUX2X1 U4237 ( .B(buff_data[361]), .A(n565), .S(n23), .Y(n4254) );
  MUX2X1 U4238 ( .B(buff_data[362]), .A(n564), .S(n148), .Y(n4255) );
  MUX2X1 U4239 ( .B(buff_data[363]), .A(n571), .S(n2198), .Y(n4256) );
  MUX2X1 U4240 ( .B(buff_data[364]), .A(n572), .S(n44), .Y(n4257) );
  MUX2X1 U4241 ( .B(buff_data[365]), .A(n579), .S(n44), .Y(n4258) );
  MUX2X1 U4242 ( .B(buff_data[367]), .A(n575), .S(n2198), .Y(n4259) );
  MUX2X1 U4243 ( .B(buff_data[383]), .A(n575), .S(n350), .Y(n4260) );
  MUX2X1 U4244 ( .B(buff_data[369]), .A(n577), .S(net79518), .Y(n4261) );
  MUX2X1 U4245 ( .B(buff_data[370]), .A(n574), .S(n1988), .Y(n4262) );
  MUX2X1 U4246 ( .B(buff_data[371]), .A(n568), .S(n349), .Y(n4263) );
  MUX2X1 U4247 ( .B(buff_data[373]), .A(n569), .S(net79518), .Y(n4264) );
  MUX2X1 U4248 ( .B(buff_data[374]), .A(n570), .S(n349), .Y(n4265) );
  MUX2X1 U4249 ( .B(buff_data[375]), .A(n578), .S(n350), .Y(n4266) );
  MUX2X1 U4250 ( .B(buff_data[378]), .A(n564), .S(n1988), .Y(n4267) );
  MUX2X1 U4251 ( .B(buff_data[380]), .A(n572), .S(n349), .Y(n4268) );
  MUX2X1 U4252 ( .B(buff_data[381]), .A(n579), .S(n184), .Y(n4269) );
  MUX2X1 U4253 ( .B(buff_data[382]), .A(n567), .S(net79518), .Y(n4270) );
  MUX2X1 U4254 ( .B(buff_data[384]), .A(n573), .S(n409), .Y(n4271) );
  MUX2X1 U4255 ( .B(buff_data[385]), .A(n577), .S(n443), .Y(n4272) );
  MUX2X1 U4256 ( .B(buff_data[386]), .A(n574), .S(n49), .Y(n4273) );
  MUX2X1 U4257 ( .B(buff_data[387]), .A(n568), .S(n443), .Y(n4274) );
  MUX2X1 U4258 ( .B(buff_data[388]), .A(n576), .S(n444), .Y(n4275) );
  MUX2X1 U4259 ( .B(buff_data[389]), .A(n569), .S(n444), .Y(n4276) );
  MUX2X1 U4260 ( .B(buff_data[390]), .A(n570), .S(n49), .Y(n4277) );
  MUX2X1 U4261 ( .B(buff_data[391]), .A(n578), .S(n444), .Y(n4278) );
  MUX2X1 U4262 ( .B(buff_data[392]), .A(n566), .S(n409), .Y(n4279) );
  MUX2X1 U4263 ( .B(buff_data[393]), .A(n565), .S(n444), .Y(n4280) );
  MUX2X1 U4264 ( .B(buff_data[394]), .A(n564), .S(n50), .Y(n4281) );
  MUX2X1 U4265 ( .B(buff_data[395]), .A(n571), .S(n408), .Y(n4282) );
  MUX2X1 U4266 ( .B(buff_data[396]), .A(n572), .S(n408), .Y(n4283) );
  MUX2X1 U4267 ( .B(buff_data[397]), .A(n579), .S(n443), .Y(n4284) );
  MUX2X1 U4268 ( .B(buff_data[398]), .A(n567), .S(n443), .Y(n4285) );
  MUX2X1 U4269 ( .B(buff_data[399]), .A(n575), .S(n50), .Y(n4286) );
  NOR3X1 U4270 ( .A(net79440), .B(net79422), .C(net66325), .Y(n3963) );
  MUX2X1 U4271 ( .B(buff_data[401]), .A(n577), .S(n113), .Y(n4288) );
  MUX2X1 U4272 ( .B(buff_data[403]), .A(n568), .S(net66834), .Y(n4289) );
  MUX2X1 U4273 ( .B(buff_data[404]), .A(n576), .S(n1799), .Y(n4290) );
  MUX2X1 U4274 ( .B(buff_data[406]), .A(n570), .S(net82336), .Y(n4291) );
  MUX2X1 U4275 ( .B(buff_data[407]), .A(n578), .S(net66834), .Y(n4292) );
  MUX2X1 U4276 ( .B(buff_data[408]), .A(n566), .S(n611), .Y(n4293) );
  MUX2X1 U4277 ( .B(buff_data[409]), .A(n565), .S(net66834), .Y(n4294) );
  MUX2X1 U4278 ( .B(buff_data[410]), .A(n564), .S(net93072), .Y(n4295) );
  MUX2X1 U4279 ( .B(buff_data[411]), .A(n571), .S(n611), .Y(n4296) );
  MUX2X1 U4280 ( .B(buff_data[412]), .A(n572), .S(n611), .Y(n4297) );
  MUX2X1 U4281 ( .B(buff_data[413]), .A(n579), .S(net66834), .Y(n4298) );
  MUX2X1 U4282 ( .B(buff_data[415]), .A(n575), .S(n611), .Y(n4299) );
  MUX2X1 U4283 ( .B(buff_data[417]), .A(n577), .S(net80783), .Y(n4300) );
  MUX2X1 U4284 ( .B(buff_data[418]), .A(n574), .S(net93057), .Y(n4301) );
  MUX2X1 U4285 ( .B(buff_data[419]), .A(n568), .S(net80783), .Y(n4302) );
  MUX2X1 U4286 ( .B(buff_data[420]), .A(n576), .S(net79538), .Y(n4303) );
  MUX2X1 U4287 ( .B(buff_data[421]), .A(n569), .S(net79538), .Y(n4304) );
  MUX2X1 U4288 ( .B(buff_data[423]), .A(n578), .S(net93057), .Y(n4305) );
  MUX2X1 U4289 ( .B(buff_data[425]), .A(n565), .S(net93057), .Y(n4306) );
  MUX2X1 U4290 ( .B(buff_data[426]), .A(n564), .S(net80783), .Y(n4307) );
  MUX2X1 U4291 ( .B(buff_data[427]), .A(n571), .S(net80783), .Y(n4308) );
  MUX2X1 U4292 ( .B(buff_data[428]), .A(n572), .S(net79538), .Y(n4309) );
  MUX2X1 U4293 ( .B(buff_data[429]), .A(n579), .S(net80783), .Y(n4310) );
  MUX2X1 U4294 ( .B(buff_data[431]), .A(n575), .S(net92836), .Y(n4311) );
  MUX2X1 U4295 ( .B(buff_data[432]), .A(n573), .S(n1928), .Y(n4312) );
  MUX2X1 U4296 ( .B(buff_data[433]), .A(n577), .S(n1928), .Y(n4313) );
  MUX2X1 U4297 ( .B(buff_data[434]), .A(n574), .S(n1928), .Y(n4314) );
  MUX2X1 U4298 ( .B(buff_data[435]), .A(n568), .S(n122), .Y(n4315) );
  MUX2X1 U4299 ( .B(buff_data[436]), .A(n576), .S(n140), .Y(n4316) );
  MUX2X1 U4300 ( .B(buff_data[437]), .A(n569), .S(n145), .Y(n4317) );
  MUX2X1 U4301 ( .B(buff_data[438]), .A(n570), .S(n1928), .Y(n4318) );
  MUX2X1 U4302 ( .B(buff_data[439]), .A(n578), .S(n2200), .Y(n4319) );
  MUX2X1 U4303 ( .B(buff_data[440]), .A(n566), .S(n121), .Y(n4320) );
  MUX2X1 U4304 ( .B(buff_data[441]), .A(n565), .S(n1928), .Y(n4321) );
  MUX2X1 U4305 ( .B(buff_data[442]), .A(n564), .S(n2027), .Y(n4322) );
  MUX2X1 U4306 ( .B(buff_data[443]), .A(n571), .S(n127), .Y(n4323) );
  MUX2X1 U4307 ( .B(buff_data[444]), .A(n572), .S(n126), .Y(n4324) );
  MUX2X1 U4308 ( .B(buff_data[445]), .A(n579), .S(n144), .Y(n4325) );
  MUX2X1 U4309 ( .B(buff_data[446]), .A(n567), .S(n139), .Y(n4326) );
  MUX2X1 U4310 ( .B(buff_data[447]), .A(n575), .S(n147), .Y(n4327) );
  NOR3X1 U4311 ( .A(net79414), .B(net79436), .C(net66325), .Y(n4011) );
  MUX2X1 U4312 ( .B(buff_data[448]), .A(n573), .S(n2195), .Y(n4328) );
  MUX2X1 U4313 ( .B(buff_data[449]), .A(n577), .S(n18), .Y(n4329) );
  MUX2X1 U4314 ( .B(buff_data[450]), .A(n574), .S(n2030), .Y(n4330) );
  MUX2X1 U4315 ( .B(buff_data[451]), .A(n568), .S(n2195), .Y(n4331) );
  MUX2X1 U4316 ( .B(buff_data[453]), .A(n569), .S(n2030), .Y(n4333) );
  MUX2X1 U4317 ( .B(buff_data[454]), .A(n570), .S(n2195), .Y(n4334) );
  MUX2X1 U4318 ( .B(buff_data[455]), .A(n578), .S(n2195), .Y(n4335) );
  MUX2X1 U4319 ( .B(buff_data[456]), .A(n566), .S(n2030), .Y(n4336) );
  MUX2X1 U4320 ( .B(buff_data[458]), .A(n564), .S(n2195), .Y(n4337) );
  MUX2X1 U4321 ( .B(buff_data[459]), .A(n571), .S(n2030), .Y(n4338) );
  MUX2X1 U4322 ( .B(buff_data[460]), .A(n572), .S(n2030), .Y(n4339) );
  MUX2X1 U4323 ( .B(buff_data[461]), .A(n579), .S(n17), .Y(n4340) );
  MUX2X1 U4324 ( .B(buff_data[462]), .A(n567), .S(n2030), .Y(n4341) );
  MUX2X1 U4325 ( .B(buff_data[463]), .A(n575), .S(n2030), .Y(n4342) );
  NOR3X1 U4326 ( .A(net79416), .B(n230), .C(net79440), .Y(net66482) );
  MUX2X1 U4327 ( .B(buff_data[464]), .A(n573), .S(n119), .Y(n4343) );
  MUX2X1 U4328 ( .B(buff_data[465]), .A(n577), .S(n108), .Y(n4344) );
  MUX2X1 U4329 ( .B(buff_data[466]), .A(n574), .S(n13), .Y(n4345) );
  MUX2X1 U4330 ( .B(buff_data[469]), .A(n569), .S(net80760), .Y(n4346) );
  MUX2X1 U4331 ( .B(buff_data[470]), .A(n570), .S(n111), .Y(n4347) );
  MUX2X1 U4332 ( .B(buff_data[471]), .A(n578), .S(n131), .Y(n4348) );
  MUX2X1 U4333 ( .B(buff_data[472]), .A(n566), .S(n110), .Y(n4349) );
  MUX2X1 U4334 ( .B(buff_data[474]), .A(n564), .S(n129), .Y(n4350) );
  MUX2X1 U4335 ( .B(buff_data[475]), .A(n571), .S(n109), .Y(n4351) );
  MUX2X1 U4336 ( .B(buff_data[477]), .A(n579), .S(n128), .Y(n4352) );
  MUX2X1 U4337 ( .B(buff_data[478]), .A(n567), .S(n112), .Y(n4353) );
  MUX2X1 U4338 ( .B(buff_data[479]), .A(n575), .S(n130), .Y(n4354) );
  MUX2X1 U4339 ( .B(buff_data[482]), .A(n574), .S(n2028), .Y(n4355) );
  MUX2X1 U4340 ( .B(buff_data[483]), .A(n568), .S(n2199), .Y(n4357) );
  MUX2X1 U4341 ( .B(buff_data[485]), .A(n569), .S(n138), .Y(n4358) );
  MUX2X1 U4342 ( .B(buff_data[486]), .A(n570), .S(n142), .Y(n4359) );
  MUX2X1 U4343 ( .B(buff_data[487]), .A(n578), .S(n2014), .Y(n4360) );
  MUX2X1 U4344 ( .B(buff_data[488]), .A(n566), .S(n137), .Y(n4361) );
  MUX2X1 U4345 ( .B(buff_data[489]), .A(n565), .S(n27), .Y(n4362) );
  MUX2X1 U4346 ( .B(buff_data[490]), .A(n564), .S(n31), .Y(n4363) );
  MUX2X1 U4347 ( .B(buff_data[491]), .A(n571), .S(n26), .Y(n4364) );
  MUX2X1 U4348 ( .B(buff_data[492]), .A(n572), .S(n180), .Y(n4365) );
  MUX2X1 U4349 ( .B(buff_data[493]), .A(n579), .S(n159), .Y(n4366) );
  MUX2X1 U4350 ( .B(buff_data[494]), .A(n567), .S(n136), .Y(n4367) );
  MUX2X1 U4351 ( .B(buff_data[495]), .A(n575), .S(n132), .Y(n4368) );
  MUX2X1 U4352 ( .B(buff_data[480]), .A(n573), .S(n1921), .Y(n4369) );
  MUX2X1 U4353 ( .B(buff_data[481]), .A(n577), .S(n36), .Y(n4370) );
  NOR3X1 U4354 ( .A(net79436), .B(n230), .C(net79422), .Y(n4056) );
  MUX2X1 U4355 ( .B(buff_data[496]), .A(n573), .S(n34), .Y(n4371) );
  MUX2X1 U4356 ( .B(buff_data[497]), .A(n577), .S(net79514), .Y(n4372) );
  MUX2X1 U4357 ( .B(buff_data[498]), .A(n574), .S(net79514), .Y(n4373) );
  MUX2X1 U4358 ( .B(buff_data[500]), .A(n576), .S(n34), .Y(n4374) );
  MUX2X1 U4359 ( .B(buff_data[501]), .A(n569), .S(n34), .Y(n4375) );
  MUX2X1 U4360 ( .B(buff_data[502]), .A(n570), .S(net79514), .Y(n4376) );
  MUX2X1 U4361 ( .B(buff_data[503]), .A(n578), .S(net79514), .Y(n4377) );
  MUX2X1 U4362 ( .B(buff_data[504]), .A(n566), .S(net79514), .Y(n4378) );
  MUX2X1 U4363 ( .B(buff_data[505]), .A(n565), .S(net79514), .Y(n4379) );
  MUX2X1 U4364 ( .B(buff_data[507]), .A(n571), .S(net79514), .Y(n4381) );
  MUX2X1 U4365 ( .B(buff_data[508]), .A(n572), .S(n34), .Y(n4382) );
  MUX2X1 U4366 ( .B(buff_data[509]), .A(n579), .S(n34), .Y(n4383) );
  MUX2X1 U4367 ( .B(buff_data[510]), .A(n567), .S(n34), .Y(n4384) );
  MUX2X1 U4368 ( .B(buff_data[511]), .A(n575), .S(net80781), .Y(n4385) );
  INVX1 U4369 ( .A(j[6]), .Y(n3930) );
  INVX1 U4370 ( .A(j[5]), .Y(n3928) );
  NOR3X1 U4371 ( .A(n1419), .B(n1476), .C(n1500), .Y(net66953) );
  INVX1 U4372 ( .A(j[20]), .Y(n3941) );
  INVX1 U4373 ( .A(j[19]), .Y(n3939) );
  INVX1 U4374 ( .A(j[22]), .Y(n3945) );
  INVX1 U4375 ( .A(j[21]), .Y(n3943) );
  NAND3X1 U4376 ( .A(n3935), .B(n3937), .C(n3933), .Y(n4386) );
  INVX1 U4377 ( .A(j[16]), .Y(n3933) );
  INVX1 U4378 ( .A(j[18]), .Y(n3937) );
  INVX1 U4379 ( .A(j[17]), .Y(n3935) );
  NAND2X1 U4380 ( .A(n1038), .B(n974), .Y(n2615) );
  NAND2X1 U4381 ( .A(n1052), .B(n986), .Y(n2613) );
  NAND2X1 U4382 ( .A(n772), .B(n989), .Y(n2611) );
  NAND2X1 U4383 ( .A(n1076), .B(n992), .Y(n2609) );
  NAND2X1 U4384 ( .A(n1090), .B(n995), .Y(n2607) );
  NAND2X1 U4385 ( .A(n1104), .B(n998), .Y(n2605) );
  NAND2X1 U4386 ( .A(n1118), .B(n1001), .Y(n2603) );
  NAND2X1 U4387 ( .A(n1132), .B(n1004), .Y(n2601) );
  NAND2X1 U4388 ( .A(n774), .B(n1007), .Y(n2599) );
  NAND2X1 U4389 ( .A(n1156), .B(n1010), .Y(n2597) );
  NAND2X1 U4390 ( .A(n1170), .B(n1013), .Y(n2595) );
  NAND2X1 U4391 ( .A(n776), .B(n1016), .Y(n2593) );
  NAND2X1 U4392 ( .A(n1194), .B(n1019), .Y(n2591) );
  NAND2X1 U4393 ( .A(n764), .B(n1022), .Y(n2589) );
  AOI22X1 U4394 ( .A(n1782), .B(n574), .C(n246), .D(n1785), .Y(n4418) );
  NAND2X1 U4395 ( .A(n778), .B(n1025), .Y(n2587) );
  NAND2X1 U4396 ( .A(n767), .B(n1028), .Y(n2585) );
  AOI22X1 U4397 ( .A(n1782), .B(n573), .C(n248), .D(n1785), .Y(n4422) );
  AND2X1 U4398 ( .A(n1612), .B(n823), .Y(n4391) );
  NAND3X1 U4399 ( .A(n3923), .B(i[4]), .C(n4425), .Y(n4424) );
  NAND3X1 U4400 ( .A(n4425), .B(n3639), .C(n1375), .Y(n3949) );
  AND2X1 U4401 ( .A(n4426), .B(n4427), .Y(n4425) );
  NOR3X1 U4402 ( .A(n1443), .B(i[15]), .C(n4429), .Y(n4427) );
  NOR3X1 U4403 ( .A(n1446), .B(n1554), .C(n1563), .Y(n4426) );
  MUX2X1 U4404 ( .B(n1698), .A(n4435), .S(n4436), .Y(n2583) );
  AND2X1 U4405 ( .A(n1528), .B(n826), .Y(n4436) );
  NAND3X1 U4406 ( .A(n3767), .B(n3765), .C(n3868), .Y(n4437) );
  AOI21X1 U4407 ( .A(n3579), .B(n3917), .C(n1636), .Y(n3635) );
  INVX1 U4408 ( .A(n1674), .Y(n3917) );
  NAND2X1 U4409 ( .A(n1212), .B(n516), .Y(n2581) );
  AOI22X1 U4410 ( .A(n4441), .B(CMD_data_out[23]), .C(n4442), .D(
        buff_bank_addr[0]), .Y(n4438) );
  NAND2X1 U4411 ( .A(n1215), .B(n517), .Y(n2579) );
  AOI22X1 U4412 ( .A(CMD_data_out[24]), .B(n4441), .C(n4442), .D(
        buff_bank_addr[1]), .Y(n4443) );
  NAND2X1 U4413 ( .A(n1218), .B(n518), .Y(n2577) );
  AOI22X1 U4414 ( .A(n4441), .B(CMD_data_out[25]), .C(n4442), .D(
        buff_bank_addr[2]), .Y(n4445) );
  NAND3X1 U4415 ( .A(n4448), .B(n1713), .C(n1381), .Y(n3849) );
  INVX1 U4416 ( .A(n1747), .Y(n3579) );
  INVX1 U4417 ( .A(n4450), .Y(n2575) );
  AOI22X1 U4418 ( .A(CMD_data_out[10]), .B(n4451), .C(A[0]), .D(n1732), .Y(
        n4450) );
  INVX1 U4419 ( .A(n4452), .Y(n2573) );
  AOI22X1 U4420 ( .A(CMD_data_out[11]), .B(n4451), .C(A[1]), .D(n1732), .Y(
        n4452) );
  INVX1 U4421 ( .A(n4453), .Y(n2571) );
  AOI22X1 U4422 ( .A(CMD_data_out[12]), .B(n4451), .C(A[2]), .D(n1732), .Y(
        n4453) );
  NAND2X1 U4423 ( .A(n4454), .B(n519), .Y(n2569) );
  MUX2X1 U4424 ( .B(A[3]), .A(n1268), .S(n4447), .Y(n4454) );
  AOI22X1 U4425 ( .A(buff_col_addr[0]), .B(n1695), .C(CMD_data_out[0]), .D(
        n4459), .Y(n4457) );
  NAND2X1 U4426 ( .A(n4460), .B(n520), .Y(n2567) );
  MUX2X1 U4427 ( .B(A[4]), .A(n1271), .S(n4447), .Y(n4460) );
  AOI22X1 U4428 ( .A(buff_col_addr[1]), .B(n1744), .C(CMD_data_out[1]), .D(
        n4459), .Y(n4463) );
  NAND2X1 U4429 ( .A(n4466), .B(n521), .Y(n2565) );
  MUX2X1 U4430 ( .B(A[5]), .A(n1274), .S(n4447), .Y(n4466) );
  AOI22X1 U4431 ( .A(buff_col_addr[2]), .B(n1744), .C(CMD_data_out[2]), .D(
        n4459), .Y(n4469) );
  NAND2X1 U4432 ( .A(n4471), .B(n522), .Y(n2563) );
  MUX2X1 U4433 ( .B(A[6]), .A(n1277), .S(n4447), .Y(n4471) );
  AOI22X1 U4434 ( .A(buff_col_addr[3]), .B(n1744), .C(CMD_data_out[3]), .D(
        n4459), .Y(n4474) );
  NAND2X1 U4435 ( .A(n4476), .B(n523), .Y(n2561) );
  MUX2X1 U4436 ( .B(A[7]), .A(n1280), .S(n4447), .Y(n4476) );
  AOI22X1 U4437 ( .A(buff_col_addr[4]), .B(n1744), .C(CMD_data_out[4]), .D(
        n4459), .Y(n4479) );
  NAND2X1 U4438 ( .A(n4481), .B(n524), .Y(n2559) );
  MUX2X1 U4439 ( .B(A[8]), .A(n1283), .S(n4447), .Y(n4481) );
  AOI22X1 U4440 ( .A(buff_col_addr[5]), .B(n1744), .C(CMD_data_out[5]), .D(
        n4459), .Y(n4484) );
  NAND2X1 U4441 ( .A(n4486), .B(n525), .Y(n2557) );
  MUX2X1 U4442 ( .B(A[9]), .A(n1286), .S(n4447), .Y(n4486) );
  AOI22X1 U4443 ( .A(buff_col_addr[6]), .B(n1744), .C(CMD_data_out[6]), .D(
        n4459), .Y(n4489) );
  NAND2X1 U4444 ( .A(n4491), .B(n526), .Y(n2555) );
  MUX2X1 U4445 ( .B(A[10]), .A(n1289), .S(n4447), .Y(n4491) );
  AOI22X1 U4446 ( .A(buff_col_addr[7]), .B(n1744), .C(CMD_data_out[7]), .D(
        n4459), .Y(n4494) );
  NAND2X1 U4447 ( .A(n4496), .B(n527), .Y(n2553) );
  MUX2X1 U4448 ( .B(A[11]), .A(n1292), .S(n4447), .Y(n4496) );
  AOI22X1 U4449 ( .A(buff_col_addr[8]), .B(n1744), .C(CMD_data_out[8]), .D(
        n4459), .Y(n4499) );
  NAND2X1 U4450 ( .A(n4501), .B(n528), .Y(n2551) );
  OAI21X1 U4451 ( .A(n1539), .B(n1747), .C(n1713), .Y(n4503) );
  MUX2X1 U4452 ( .B(A[12]), .A(n534), .S(n4447), .Y(n4501) );
  NAND3X1 U4453 ( .A(n3687), .B(n3670), .C(n4508), .Y(n4507) );
  INVX1 U4454 ( .A(n1680), .Y(n3687) );
  INVX1 U4455 ( .A(n4509), .Y(n4508) );
  NAND3X1 U4456 ( .A(n1578), .B(n1747), .C(n1384), .Y(n4506) );
  INVX1 U4457 ( .A(flag_bl_read), .Y(n4435) );
  AOI22X1 U4458 ( .A(buff_col_addr[9]), .B(n1744), .C(CMD_data_out[9]), .D(
        n4459), .Y(n4512) );
  OAI21X1 U4459 ( .A(n3774), .B(n1747), .C(n4448), .Y(n4459) );
  INVX1 U4460 ( .A(n1551), .Y(n4448) );
  NAND3X1 U4461 ( .A(n3670), .B(n1624), .C(n1387), .Y(n3678) );
  INVX1 U4462 ( .A(n1707), .Y(n3923) );
  INVX1 U4463 ( .A(n1683), .Y(n3670) );
  NAND3X1 U4464 ( .A(n845), .B(n1301), .C(n4518), .Y(n3894) );
  NOR3X1 U4465 ( .A(n1449), .B(net66007), .C(n3661), .Y(n4518) );
  AOI22X1 U4466 ( .A(n1686), .B(n4520), .C(n4521), .D(net66063), .Y(n4517) );
  INVX1 U4467 ( .A(n1713), .Y(net66063) );
  INVX1 U4468 ( .A(n4511), .Y(n4521) );
  OAI21X1 U4469 ( .A(CMD_data_out[33]), .B(net66974), .C(n4522), .Y(n4511) );
  MUX2X1 U4470 ( .B(net66974), .A(CMD_data_out[33]), .S(net66975), .Y(n4522)
         );
  OAI21X1 U4471 ( .A(n3999), .B(n1710), .C(n1692), .Y(n4520) );
  AOI21X1 U4472 ( .A(n3911), .B(n3999), .C(n865), .Y(n4526) );
  NAND3X1 U4473 ( .A(n1548), .B(net65981), .C(n4528), .Y(n4509) );
  OAI21X1 U4474 ( .A(n1525), .B(n1537), .C(net66160), .Y(n4528) );
  INVX1 U4475 ( .A(n1624), .Y(net66160) );
  INVX1 U4476 ( .A(net67120), .Y(net66385) );
  NAND3X1 U4477 ( .A(n4532), .B(clkcount[0]), .C(n2509), .Y(net67120) );
  INVX1 U4478 ( .A(n1701), .Y(n3999) );
  INVX1 U4479 ( .A(n1692), .Y(n3911) );
  NAND3X1 U4480 ( .A(n3767), .B(n3914), .C(n3868), .Y(n4525) );
  INVX1 U4481 ( .A(n1531), .Y(n3868) );
  NAND3X1 U4482 ( .A(i[3]), .B(net66073), .C(n3771), .Y(n3766) );
  OR2X1 U4483 ( .A(n1545), .B(n1704), .Y(n4524) );
  NAND3X1 U4484 ( .A(i[0]), .B(net66078), .C(n3771), .Y(n3757) );
  INVX1 U4485 ( .A(n1537), .Y(n3771) );
  NAND3X1 U4486 ( .A(n4534), .B(n4535), .C(n4536), .Y(n4515) );
  NOR3X1 U4487 ( .A(n4537), .B(n1683), .C(n3679), .Y(n4536) );
  INVX1 U4488 ( .A(n1518), .Y(n3679) );
  AOI21X1 U4489 ( .A(n1726), .B(n3918), .C(n3765), .Y(n3655) );
  INVX1 U4490 ( .A(n1651), .Y(n3765) );
  NOR3X1 U4491 ( .A(n1747), .B(n3776), .C(n3869), .Y(n3918) );
  INVX1 U4492 ( .A(flag_bl_write), .Y(n3869) );
  INVX1 U4493 ( .A(n4539), .Y(n3776) );
  INVX1 U4494 ( .A(n4540), .Y(n4531) );
  NAND3X1 U4495 ( .A(state[1]), .B(state[4]), .C(n4541), .Y(n4540) );
  AND2X1 U4496 ( .A(n3681), .B(net65999), .Y(n4541) );
  NAND3X1 U4497 ( .A(state[3]), .B(net66031), .C(n4542), .Y(n3652) );
  OAI21X1 U4498 ( .A(n3660), .B(n1630), .C(n665), .Y(n4537) );
  AOI22X1 U4499 ( .A(n1741), .B(n3774), .C(n3920), .D(n4544), .Y(n4543) );
  INVX1 U4500 ( .A(n1521), .Y(n3920) );
  NAND3X1 U4501 ( .A(n4533), .B(i[1]), .C(n4538), .Y(n3900) );
  INVX1 U4502 ( .A(n1677), .Y(n4538) );
  INVX1 U4503 ( .A(n1660), .Y(n4533) );
  INVX1 U4504 ( .A(n890), .Y(n3774) );
  AOI21X1 U4505 ( .A(flag_bl_write), .B(n1523), .C(n1747), .Y(n3675) );
  NAND3X1 U4506 ( .A(CMD_data_out[33]), .B(n4546), .C(n4547), .Y(n4539) );
  INVX1 U4507 ( .A(n4548), .Y(n3660) );
  NAND3X1 U4508 ( .A(n1245), .B(n1312), .C(n4551), .Y(n4548) );
  NOR3X1 U4509 ( .A(n4552), .B(n1464), .C(n1488), .Y(n4551) );
  NAND3X1 U4510 ( .A(n3821), .B(n3823), .C(n3819), .Y(n4554) );
  INVX1 U4511 ( .A(clkcount[20]), .Y(n3819) );
  INVX1 U4512 ( .A(clkcount[22]), .Y(n3823) );
  INVX1 U4513 ( .A(clkcount[21]), .Y(n3821) );
  NAND3X1 U4514 ( .A(n3827), .B(n3829), .C(n3825), .Y(n4553) );
  INVX1 U4515 ( .A(clkcount[23]), .Y(n3825) );
  INVX1 U4516 ( .A(clkcount[25]), .Y(n3829) );
  INVX1 U4517 ( .A(clkcount[24]), .Y(n3827) );
  OR2X1 U4518 ( .A(n832), .B(n829), .Y(n4552) );
  NAND3X1 U4519 ( .A(n3833), .B(n3835), .C(n3831), .Y(n4556) );
  INVX1 U4520 ( .A(clkcount[26]), .Y(n3831) );
  INVX1 U4521 ( .A(clkcount[28]), .Y(n3835) );
  INVX1 U4522 ( .A(clkcount[27]), .Y(n3833) );
  NAND3X1 U4523 ( .A(n3839), .B(n3643), .C(n3837), .Y(n4555) );
  INVX1 U4524 ( .A(clkcount[29]), .Y(n3837) );
  INVX1 U4525 ( .A(clkcount[31]), .Y(n3643) );
  INVX1 U4526 ( .A(clkcount[30]), .Y(n3839) );
  NAND3X1 U4527 ( .A(n3809), .B(n3811), .C(n3807), .Y(n4558) );
  INVX1 U4528 ( .A(clkcount[14]), .Y(n3807) );
  INVX1 U4529 ( .A(clkcount[16]), .Y(n3811) );
  INVX1 U4530 ( .A(clkcount[15]), .Y(n3809) );
  NAND3X1 U4531 ( .A(n3815), .B(n3817), .C(n3813), .Y(n4557) );
  INVX1 U4532 ( .A(clkcount[17]), .Y(n3813) );
  INVX1 U4533 ( .A(clkcount[19]), .Y(n3817) );
  INVX1 U4534 ( .A(clkcount[18]), .Y(n3815) );
  NAND3X1 U4535 ( .A(clkcount[9]), .B(clkcount[12]), .C(n4561), .Y(n4560) );
  MUX2X1 U4536 ( .B(n855), .A(n1295), .S(n3795), .Y(n4561) );
  INVX1 U4537 ( .A(clkcount[8]), .Y(n3795) );
  NAND3X1 U4538 ( .A(n1248), .B(n3787), .C(n4565), .Y(n4562) );
  NOR3X1 U4539 ( .A(clkcount[5]), .B(clkcount[7]), .C(clkcount[6]), .Y(n4565)
         );
  INVX1 U4540 ( .A(clkcount[4]), .Y(n3787) );
  NAND3X1 U4541 ( .A(n3801), .B(n3805), .C(n3799), .Y(n4559) );
  INVX1 U4542 ( .A(clkcount[10]), .Y(n3799) );
  INVX1 U4543 ( .A(clkcount[13]), .Y(n3805) );
  INVX1 U4544 ( .A(clkcount[11]), .Y(n3801) );
  NOR3X1 U4545 ( .A(net66007), .B(n4566), .C(n3701), .Y(n4535) );
  NOR3X1 U4546 ( .A(n1660), .B(net65987), .C(n1707), .Y(n3701) );
  NAND3X1 U4547 ( .A(i[5]), .B(n3770), .C(n1390), .Y(n3922) );
  INVX1 U4548 ( .A(n1525), .Y(n3770) );
  INVX1 U4549 ( .A(n1627), .Y(n4566) );
  AND2X1 U4550 ( .A(n3637), .B(net66080), .Y(n3769) );
  INVX1 U4551 ( .A(n1630), .Y(n3661) );
  NAND3X1 U4552 ( .A(state[2]), .B(state[3]), .C(n4542), .Y(n3909) );
  NAND3X1 U4553 ( .A(net65999), .B(n3681), .C(n4569), .Y(net66151) );
  INVX1 U4554 ( .A(n4570), .Y(n4534) );
  NAND3X1 U4555 ( .A(n4571), .B(n1704), .C(n1713), .Y(n4570) );
  NAND3X1 U4556 ( .A(n4569), .B(n3681), .C(state[0]), .Y(net66283) );
  NAND3X1 U4557 ( .A(n4569), .B(net65999), .C(state[3]), .Y(n3654) );
  OAI21X1 U4558 ( .A(n1581), .B(n4544), .C(n1686), .Y(n4571) );
  INVX1 U4559 ( .A(n1615), .Y(n4544) );
  NAND3X1 U4560 ( .A(n3637), .B(net65987), .C(n3638), .Y(n4572) );
  INVX1 U4561 ( .A(n4573), .Y(n3638) );
  NAND3X1 U4562 ( .A(i[0]), .B(n1677), .C(n4429), .Y(n4573) );
  INVX1 U4563 ( .A(n1735), .Y(n3639) );
  NAND3X1 U4564 ( .A(n1707), .B(n1729), .C(n1393), .Y(n4523) );
  NAND3X1 U4565 ( .A(n3637), .B(n4429), .C(n4575), .Y(n3759) );
  AND2X1 U4566 ( .A(net65987), .B(net66073), .Y(n4575) );
  INVX1 U4567 ( .A(n4576), .Y(n3637) );
  NAND3X1 U4568 ( .A(n1668), .B(net66076), .C(n4577), .Y(n4576) );
  INVX1 U4569 ( .A(n1698), .Y(n3631) );
  NAND3X1 U4570 ( .A(net65999), .B(net66031), .C(net67122), .Y(n3912) );
  NAND3X1 U4571 ( .A(net66031), .B(n3681), .C(n4542), .Y(net66166) );
  NOR3X1 U4572 ( .A(net65999), .B(state[4]), .C(n3663), .Y(n4542) );
  INVX1 U4573 ( .A(state[1]), .Y(n3663) );
  INVX1 U4574 ( .A(state[3]), .Y(n3681) );
  MUX2X1 U4575 ( .B(n1642), .A(n1665), .S(DQS_bar_out[0]), .Y(n2548) );
  MUX2X1 U4576 ( .B(n1642), .A(n1665), .S(DQS_bar_out[1]), .Y(n2547) );
  INVX1 U4577 ( .A(n1642), .Y(n4581) );
  NAND3X1 U4578 ( .A(n1560), .B(n1680), .C(n1587), .Y(n4582) );
  NAND3X1 U4579 ( .A(n1680), .B(net67172), .C(n4584), .Y(n4579) );
  AND2X1 U4580 ( .A(n1560), .B(n1587), .Y(n4584) );
  NAND3X1 U4581 ( .A(n4577), .B(n4587), .C(n4588), .Y(n4586) );
  AND2X1 U4582 ( .A(n4434), .B(n1633), .Y(n4588) );
  INVX1 U4583 ( .A(n1563), .Y(n4577) );
  INVX1 U4584 ( .A(i[5]), .Y(net66082) );
  NAND3X1 U4585 ( .A(net65992), .B(net66084), .C(n1369), .Y(n4585) );
  AOI21X1 U4586 ( .A(n4429), .B(n849), .C(i[15]), .Y(n4589) );
  NAND3X1 U4587 ( .A(net65987), .B(net66076), .C(net66073), .Y(n4590) );
  INVX1 U4588 ( .A(i[2]), .Y(net66076) );
  AND2X1 U4589 ( .A(i[3]), .B(i[4]), .Y(n4429) );
  INVX1 U4590 ( .A(reset), .Y(net67172) );
  NAND3X1 U4591 ( .A(state[2]), .B(state[3]), .C(n4591), .Y(n3653) );
  NOR3X1 U4592 ( .A(state[0]), .B(state[4]), .C(state[1]), .Y(n4591) );
  AND2X1 U4593 ( .A(state[0]), .B(net66031), .Y(n3847) );
  INVX1 U4594 ( .A(state[2]), .Y(net66031) );
  OAI21X1 U4595 ( .A(n4545), .B(n1747), .C(n1548), .Y(n2439) );
  NAND3X1 U4596 ( .A(n3914), .B(n1677), .C(n3767), .Y(n4527) );
  INVX1 U4597 ( .A(n1509), .Y(n3767) );
  NAND3X1 U4598 ( .A(ring_ptr[1]), .B(ring_ptr[0]), .C(ring_ptr[2]), .Y(n4000)
         );
  NAND3X1 U4599 ( .A(n4592), .B(n4593), .C(n4594), .Y(n3915) );
  NOR3X1 U4600 ( .A(n1452), .B(n1467), .C(n1491), .Y(n4594) );
  NAND3X1 U4601 ( .A(n3618), .B(n3620), .C(n3616), .Y(n4597) );
  INVX1 U4602 ( .A(blk_cnt[24]), .Y(n3616) );
  INVX1 U4603 ( .A(blk_cnt[26]), .Y(n3620) );
  INVX1 U4604 ( .A(blk_cnt[25]), .Y(n3618) );
  NAND3X1 U4605 ( .A(n3622), .B(n3624), .C(n4598), .Y(n4596) );
  AND2X1 U4606 ( .A(n3628), .B(n3626), .Y(n4598) );
  INVX1 U4607 ( .A(blk_cnt[29]), .Y(n3626) );
  INVX1 U4608 ( .A(blk_cnt[30]), .Y(n3628) );
  INVX1 U4609 ( .A(blk_cnt[28]), .Y(n3624) );
  INVX1 U4610 ( .A(blk_cnt[27]), .Y(n3622) );
  NOR3X1 U4611 ( .A(n1455), .B(blk_cnt[7]), .C(blk_cnt[6]), .Y(n4600) );
  INVX1 U4612 ( .A(blk_cnt[9]), .Y(n3586) );
  INVX1 U4613 ( .A(blk_cnt[8]), .Y(n3584) );
  NOR3X1 U4614 ( .A(n1458), .B(blk_cnt[3]), .C(blk_cnt[31]), .Y(n4599) );
  INVX1 U4615 ( .A(blk_cnt[5]), .Y(n3576) );
  INVX1 U4616 ( .A(blk_cnt[4]), .Y(n3573) );
  NOR3X1 U4617 ( .A(n1422), .B(n1479), .C(n1503), .Y(n4593) );
  INVX1 U4618 ( .A(blk_cnt[21]), .Y(n3610) );
  INVX1 U4619 ( .A(blk_cnt[20]), .Y(n3608) );
  INVX1 U4620 ( .A(blk_cnt[23]), .Y(n3614) );
  INVX1 U4621 ( .A(blk_cnt[22]), .Y(n3612) );
  NAND3X1 U4622 ( .A(n3604), .B(n3606), .C(n3602), .Y(n4603) );
  INVX1 U4623 ( .A(blk_cnt[17]), .Y(n3602) );
  INVX1 U4624 ( .A(blk_cnt[19]), .Y(n3606) );
  INVX1 U4625 ( .A(blk_cnt[18]), .Y(n3604) );
  NOR3X1 U4626 ( .A(n1425), .B(n1482), .C(n1506), .Y(n4592) );
  INVX1 U4627 ( .A(blk_cnt[14]), .Y(n3596) );
  INVX1 U4628 ( .A(blk_cnt[13]), .Y(n3594) );
  INVX1 U4629 ( .A(blk_cnt[16]), .Y(n3600) );
  INVX1 U4630 ( .A(blk_cnt[15]), .Y(n3598) );
  NAND3X1 U4631 ( .A(n3590), .B(n3592), .C(n3588), .Y(n4606) );
  INVX1 U4632 ( .A(blk_cnt[10]), .Y(n3588) );
  INVX1 U4633 ( .A(blk_cnt[12]), .Y(n3592) );
  INVX1 U4634 ( .A(blk_cnt[11]), .Y(n3590) );
  INVX1 U4635 ( .A(n4609), .Y(n3914) );
  NAND3X1 U4636 ( .A(net67122), .B(net65999), .C(state[2]), .Y(n4609) );
  INVX1 U4637 ( .A(state[0]), .Y(net65999) );
  NOR3X1 U4638 ( .A(state[1]), .B(state[3]), .C(n3691), .Y(net67122) );
  INVX1 U4639 ( .A(state[4]), .Y(n3691) );
  NAND3X1 U4640 ( .A(state[0]), .B(n4569), .C(state[3]), .Y(n3668) );
  NOR3X1 U4641 ( .A(state[2]), .B(state[4]), .C(state[1]), .Y(n4569) );
  INVX1 U4642 ( .A(n4610), .Y(n4545) );
  NAND3X1 U4643 ( .A(n1543), .B(n1725), .C(n1674), .Y(n4610) );
  NAND3X1 U4644 ( .A(n4546), .B(net67203), .C(n1396), .Y(n3674) );
  INVX1 U4645 ( .A(CMD_data_out[33]), .Y(net67203) );
  NAND3X1 U4646 ( .A(CMD_data_out[31]), .B(net66975), .C(n4546), .Y(n4611) );
  INVX1 U4647 ( .A(n4613), .Y(n4546) );
  NAND3X1 U4648 ( .A(i[2]), .B(n3855), .C(n1398), .Y(n4613) );
  NAND3X1 U4649 ( .A(net66080), .B(net66086), .C(n1668), .Y(n4568) );
  NAND3X1 U4650 ( .A(n1633), .B(n4434), .C(n4587), .Y(n4616) );
  INVX1 U4651 ( .A(n1554), .Y(n4587) );
  NAND3X1 U4652 ( .A(n4617), .B(n4618), .C(n4619), .Y(n4431) );
  NOR3X1 U4653 ( .A(n1428), .B(i[21]), .C(i[20]), .Y(n4619) );
  NAND3X1 U4654 ( .A(n3733), .B(n3735), .C(net66116), .Y(n4620) );
  INVX1 U4655 ( .A(i[22]), .Y(net66116) );
  INVX1 U4656 ( .A(i[24]), .Y(n3735) );
  INVX1 U4657 ( .A(i[23]), .Y(n3733) );
  NOR3X1 U4658 ( .A(i[28]), .B(i[30]), .C(i[29]), .Y(n4618) );
  NOR3X1 U4659 ( .A(i[25]), .B(i[27]), .C(i[26]), .Y(n4617) );
  INVX1 U4660 ( .A(n4621), .Y(n4434) );
  NAND3X1 U4661 ( .A(net66092), .B(net66094), .C(n4622), .Y(n4621) );
  NOR3X1 U4662 ( .A(i[12]), .B(i[14]), .C(i[13]), .Y(n4622) );
  INVX1 U4663 ( .A(i[11]), .Y(net66094) );
  INVX1 U4664 ( .A(i[10]), .Y(net66092) );
  NAND3X1 U4665 ( .A(net66106), .B(net66108), .C(net66104), .Y(n4624) );
  INVX1 U4666 ( .A(i[16]), .Y(net66104) );
  INVX1 U4667 ( .A(i[18]), .Y(net66108) );
  INVX1 U4668 ( .A(i[17]), .Y(net66106) );
  NAND3X1 U4669 ( .A(net66088), .B(net66090), .C(net66110), .Y(n4623) );
  INVX1 U4670 ( .A(i[19]), .Y(net66110) );
  INVX1 U4671 ( .A(i[9]), .Y(net66090) );
  INVX1 U4672 ( .A(i[8]), .Y(net66088) );
  NAND3X1 U4673 ( .A(net65992), .B(net66084), .C(net66102), .Y(n4615) );
  INVX1 U4674 ( .A(i[15]), .Y(net66102) );
  INVX1 U4675 ( .A(i[6]), .Y(net66084) );
  INVX1 U4676 ( .A(i[31]), .Y(net65992) );
  INVX1 U4677 ( .A(i[7]), .Y(net66086) );
  INVX1 U4678 ( .A(i[4]), .Y(net66080) );
  NOR3X1 U4679 ( .A(net65987), .B(net66073), .C(net66078), .Y(n3855) );
  INVX1 U4680 ( .A(i[3]), .Y(net66078) );
  INVX1 U4681 ( .A(i[0]), .Y(net66073) );
  INVX1 U4682 ( .A(i[1]), .Y(net65987) );
  INVX1 U4683 ( .A(DQS_out[1]), .Y(DQS_bar_out[1]) );
  INVX1 U4684 ( .A(DQS_out[0]), .Y(DQS_bar_out[0]) );
endmodule


module SSTL18DDR3DIFF ( PAD, PADN, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD,  PADN;
  wire   n1, n2, n3;

  TBUFX2 b2 ( .A(A), .EN(TS), .Y(PADN) );
  TBUFX2 b1 ( .A(n3), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n3) );
  INVX1 U2 ( .A(n1), .Y(Z) );
  NAND3X1 U3 ( .A(PAD), .B(n2), .C(RI), .Y(n1) );
  INVX1 U4 ( .A(PADN), .Y(n2) );
endmodule


module SSTL18DDR3_44 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n1) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_43 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n2;

  TBUFX2 b1 ( .A(n2), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n2) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_42 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n2;

  TBUFX2 b1 ( .A(n2), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n2) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_41 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n2;

  TBUFX2 b1 ( .A(n2), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n2) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_40 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n2;

  TBUFX2 b1 ( .A(n2), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n2) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_39 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n2;

  TBUFX2 b1 ( .A(n2), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n2) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_38 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n2;

  TBUFX2 b1 ( .A(n2), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n2) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_37 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n2;

  TBUFX2 b1 ( .A(n2), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n2) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_36 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n2;

  TBUFX2 b1 ( .A(n2), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n2) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_35 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n2;

  TBUFX2 b1 ( .A(n2), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n2) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_34 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n2;

  TBUFX2 b1 ( .A(n2), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n2) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_33 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n2;

  TBUFX2 b1 ( .A(n2), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n2) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_32 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n2;

  TBUFX2 b1 ( .A(n2), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n2) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_31 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n2;

  TBUFX2 b1 ( .A(n2), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n2) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_30 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n2;

  TBUFX2 b1 ( .A(n2), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n2) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_29 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n2;

  TBUFX2 b1 ( .A(n2), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n2) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_28 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n2;

  TBUFX2 b1 ( .A(n2), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n2) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_27 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n2;

  TBUFX2 b1 ( .A(n2), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n2) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_26 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n2;

  TBUFX2 b1 ( .A(n2), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n2) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_25 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n2;

  TBUFX2 b1 ( .A(n2), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n2) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_24 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n2;

  TBUFX2 b1 ( .A(n2), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n2) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_23 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n2;

  TBUFX2 b1 ( .A(n2), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n2) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_22 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n2;

  TBUFX2 b1 ( .A(n2), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n2) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_21 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n2;

  TBUFX2 b1 ( .A(n2), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n2) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_20 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n2;

  TBUFX2 b1 ( .A(n2), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n2) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_19 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n2;

  TBUFX2 b1 ( .A(n2), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n2) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_18 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n2;

  TBUFX2 b1 ( .A(n2), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n2) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_17 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n2;

  TBUFX2 b1 ( .A(n2), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n2) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_16 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n2;

  TBUFX2 b1 ( .A(n2), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n2) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_15 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n2;

  TBUFX2 b1 ( .A(n2), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n2) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_14 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n2;

  TBUFX2 b1 ( .A(n2), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n2) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_13 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n2;

  TBUFX2 b1 ( .A(n2), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n2) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_12 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n2;

  TBUFX2 b1 ( .A(n2), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n2) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_11 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n2;

  TBUFX2 b1 ( .A(n2), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n2) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_10 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n2;

  TBUFX2 b1 ( .A(n2), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n2) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_9 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n2;

  TBUFX2 b1 ( .A(n2), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n2) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_8 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n2;

  TBUFX2 b1 ( .A(n2), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n2) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_7 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n2;

  TBUFX2 b1 ( .A(n2), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n2) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_6 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n2;

  TBUFX2 b1 ( .A(n2), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n2) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_5 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n2;

  TBUFX2 b1 ( .A(n2), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n2) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_4 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n2;

  TBUFX2 b1 ( .A(n2), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n2) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_3 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n2;

  TBUFX2 b1 ( .A(n2), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n2) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_2 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n2;

  TBUFX2 b1 ( .A(n2), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n2) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_1 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n2;

  TBUFX2 b1 ( .A(n2), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n2) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_0 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n2;

  TBUFX2 b1 ( .A(n2), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n2) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3INTERFACE ( ck_pad, ckbar_pad, cke_pad, csbar_pad, rasbar_pad, 
        casbar_pad, webar_pad, ba_pad, a_pad, dm_pad, odt_pad, resetbar_pad, 
        dq_o, dqs_o, dqsbar_o, dq_pad, dqs_pad, dqsbar_pad, ri_i, ts_i, ck_i, 
        cke_i, csbar_i, rasbar_i, casbar_i, webar_i, ba_i, a_i, dq_i, dqs_i, 
        dqsbar_i, dm_i, odt_i, resetbar_i );
  output [2:0] ba_pad;
  output [12:0] a_pad;
  output [1:0] dm_pad;
  output [15:0] dq_o;
  output [1:0] dqs_o;
  output [1:0] dqsbar_o;
  inout [15:0] dq_pad;
  inout [1:0] dqs_pad;
  inout [1:0] dqsbar_pad;
  input [2:0] ba_i;
  input [12:0] a_i;
  input [15:0] dq_i;
  input [1:0] dqs_i;
  input [1:0] dqsbar_i;
  input [1:0] dm_i;
  input ri_i, ts_i, ck_i, cke_i, csbar_i, rasbar_i, casbar_i, webar_i, odt_i,
         resetbar_i;
  output ck_pad, ckbar_pad, cke_pad, csbar_pad, rasbar_pad, casbar_pad,
         webar_pad, odt_pad, resetbar_pad;


  SSTL18DDR3DIFF ck_sstl ( .PAD(ck_pad), .PADN(ckbar_pad), .Z(), .A(ck_i), 
        .RI(1'b0), .TS(1'b1) );
  SSTL18DDR3_44 cke_sstl ( .PAD(cke_pad), .Z(), .A(cke_i), .RI(1'b0), .TS(1'b1) );
  SSTL18DDR3_43 casbar_sstl ( .PAD(casbar_pad), .Z(), .A(casbar_i), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_42 rasbar_sstl ( .PAD(rasbar_pad), .Z(), .A(rasbar_i), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_41 csbar_sstl ( .PAD(csbar_pad), .Z(), .A(csbar_i), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_40 webar_sstl ( .PAD(webar_pad), .Z(), .A(webar_i), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_39 odt_sstl ( .PAD(odt_pad), .Z(), .A(odt_i), .RI(1'b0), .TS(1'b1) );
  SSTL18DDR3_38 resetbar_sstl ( .PAD(resetbar_pad), .Z(), .A(resetbar_i), .RI(
        1'b0), .TS(1'b1) );
  SSTL18DDR3_37 BA_0__sstl_ba ( .PAD(ba_pad[0]), .Z(), .A(ba_i[0]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_36 BA_1__sstl_ba ( .PAD(ba_pad[1]), .Z(), .A(ba_i[1]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_35 BA_2__sstl_ba ( .PAD(ba_pad[2]), .Z(), .A(ba_i[2]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_34 A_0__sstl_a ( .PAD(a_pad[0]), .Z(), .A(a_i[0]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_33 A_1__sstl_a ( .PAD(a_pad[1]), .Z(), .A(a_i[1]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_32 A_2__sstl_a ( .PAD(a_pad[2]), .Z(), .A(a_i[2]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_31 A_3__sstl_a ( .PAD(a_pad[3]), .Z(), .A(a_i[3]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_30 A_4__sstl_a ( .PAD(a_pad[4]), .Z(), .A(a_i[4]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_29 A_5__sstl_a ( .PAD(a_pad[5]), .Z(), .A(a_i[5]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_28 A_6__sstl_a ( .PAD(a_pad[6]), .Z(), .A(a_i[6]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_27 A_7__sstl_a ( .PAD(a_pad[7]), .Z(), .A(a_i[7]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_26 A_8__sstl_a ( .PAD(a_pad[8]), .Z(), .A(a_i[8]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_25 A_9__sstl_a ( .PAD(a_pad[9]), .Z(), .A(a_i[9]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_24 A_10__sstl_a ( .PAD(a_pad[10]), .Z(), .A(a_i[10]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_23 A_11__sstl_a ( .PAD(a_pad[11]), .Z(), .A(a_i[11]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_22 A_12__sstl_a ( .PAD(a_pad[12]), .Z(), .A(a_i[12]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_21 DQ_0__sstl_dq ( .PAD(dq_pad[0]), .Z(dq_o[0]), .A(dq_i[0]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_20 DQ_1__sstl_dq ( .PAD(dq_pad[1]), .Z(dq_o[1]), .A(dq_i[1]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_19 DQ_2__sstl_dq ( .PAD(dq_pad[2]), .Z(dq_o[2]), .A(dq_i[2]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_18 DQ_3__sstl_dq ( .PAD(dq_pad[3]), .Z(dq_o[3]), .A(dq_i[3]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_17 DQ_4__sstl_dq ( .PAD(dq_pad[4]), .Z(dq_o[4]), .A(dq_i[4]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_16 DQ_5__sstl_dq ( .PAD(dq_pad[5]), .Z(dq_o[5]), .A(dq_i[5]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_15 DQ_6__sstl_dq ( .PAD(dq_pad[6]), .Z(dq_o[6]), .A(dq_i[6]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_14 DQ_7__sstl_dq ( .PAD(dq_pad[7]), .Z(dq_o[7]), .A(dq_i[7]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_13 DQ_8__sstl_dq ( .PAD(dq_pad[8]), .Z(dq_o[8]), .A(dq_i[8]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_12 DQ_9__sstl_dq ( .PAD(dq_pad[9]), .Z(dq_o[9]), .A(dq_i[9]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_11 DQ_10__sstl_dq ( .PAD(dq_pad[10]), .Z(dq_o[10]), .A(dq_i[10]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_10 DQ_11__sstl_dq ( .PAD(dq_pad[11]), .Z(dq_o[11]), .A(dq_i[11]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_9 DQ_12__sstl_dq ( .PAD(dq_pad[12]), .Z(dq_o[12]), .A(dq_i[12]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_8 DQ_13__sstl_dq ( .PAD(dq_pad[13]), .Z(dq_o[13]), .A(dq_i[13]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_7 DQ_14__sstl_dq ( .PAD(dq_pad[14]), .Z(dq_o[14]), .A(dq_i[14]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_6 DQ_15__sstl_dq ( .PAD(dq_pad[15]), .Z(dq_o[15]), .A(dq_i[15]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_5 DQS_0__sstl_dqs ( .PAD(dqs_pad[0]), .Z(dqs_o[0]), .A(dqs_i[0]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_4 DQS_1__sstl_dqs ( .PAD(dqs_pad[1]), .Z(dqs_o[1]), .A(dqs_i[1]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_3 DQSBAR_0__sstl_dqsbar ( .PAD(dqsbar_pad[0]), .Z(dqsbar_o[0]), 
        .A(dqsbar_i[0]), .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_2 DQSBAR_1__sstl_dqsbar ( .PAD(dqsbar_pad[1]), .Z(dqsbar_o[1]), 
        .A(dqsbar_i[1]), .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_1 DM_0__sstl_dm ( .PAD(dm_pad[0]), .Z(), .A(dm_i[0]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_0 DM_1__sstl_dm ( .PAD(dm_pad[1]), .Z(), .A(dm_i[1]), .RI(1'b0), 
        .TS(1'b1) );
endmodule


module ddr3_controller_DW01_inc_0 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;

  wire   [31:2] carry;

  HAX1 U1_1_30 ( .A(A[30]), .B(carry[30]), .YC(carry[31]), .YS(SUM[30]) );
  HAX1 U1_1_29 ( .A(A[29]), .B(carry[29]), .YC(carry[30]), .YS(SUM[29]) );
  HAX1 U1_1_28 ( .A(A[28]), .B(carry[28]), .YC(carry[29]), .YS(SUM[28]) );
  HAX1 U1_1_27 ( .A(A[27]), .B(carry[27]), .YC(carry[28]), .YS(SUM[27]) );
  HAX1 U1_1_26 ( .A(A[26]), .B(carry[26]), .YC(carry[27]), .YS(SUM[26]) );
  HAX1 U1_1_25 ( .A(A[25]), .B(carry[25]), .YC(carry[26]), .YS(SUM[25]) );
  HAX1 U1_1_24 ( .A(A[24]), .B(carry[24]), .YC(carry[25]), .YS(SUM[24]) );
  HAX1 U1_1_23 ( .A(A[23]), .B(carry[23]), .YC(carry[24]), .YS(SUM[23]) );
  HAX1 U1_1_22 ( .A(A[22]), .B(carry[22]), .YC(carry[23]), .YS(SUM[22]) );
  HAX1 U1_1_21 ( .A(A[21]), .B(carry[21]), .YC(carry[22]), .YS(SUM[21]) );
  HAX1 U1_1_20 ( .A(A[20]), .B(carry[20]), .YC(carry[21]), .YS(SUM[20]) );
  HAX1 U1_1_19 ( .A(A[19]), .B(carry[19]), .YC(carry[20]), .YS(SUM[19]) );
  HAX1 U1_1_18 ( .A(A[18]), .B(carry[18]), .YC(carry[19]), .YS(SUM[18]) );
  HAX1 U1_1_17 ( .A(A[17]), .B(carry[17]), .YC(carry[18]), .YS(SUM[17]) );
  HAX1 U1_1_16 ( .A(A[16]), .B(carry[16]), .YC(carry[17]), .YS(SUM[16]) );
  HAX1 U1_1_15 ( .A(A[15]), .B(carry[15]), .YC(carry[16]), .YS(SUM[15]) );
  HAX1 U1_1_14 ( .A(A[14]), .B(carry[14]), .YC(carry[15]), .YS(SUM[14]) );
  HAX1 U1_1_13 ( .A(A[13]), .B(carry[13]), .YC(carry[14]), .YS(SUM[13]) );
  HAX1 U1_1_12 ( .A(A[12]), .B(carry[12]), .YC(carry[13]), .YS(SUM[12]) );
  HAX1 U1_1_11 ( .A(A[11]), .B(carry[11]), .YC(carry[12]), .YS(SUM[11]) );
  HAX1 U1_1_10 ( .A(A[10]), .B(carry[10]), .YC(carry[11]), .YS(SUM[10]) );
  HAX1 U1_1_9 ( .A(A[9]), .B(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  HAX1 U1_1_8 ( .A(A[8]), .B(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  HAX1 U1_1_7 ( .A(A[7]), .B(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  HAX1 U1_1_6 ( .A(A[6]), .B(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  HAX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry[2]), .YS(SUM[1]) );
  XOR2X1 U1 ( .A(carry[31]), .B(A[31]), .Y(SUM[31]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module ddr3_controller ( dout, raddr, fillcount, notfull, ready, ck_pad, 
        ckbar_pad, cke_pad, csbar_pad, rasbar_pad, casbar_pad, webar_pad, 
        ba_pad, a_pad, dm_pad, odt_pad, resetbar_pad, validout, dq_pad, 
        dqs_pad, dqsbar_pad, clk, reset, read, cmd, din, sz, op, addr, initddr, 
        waiting );
  output [15:0] dout;
  output [25:0] raddr;
  output [5:0] fillcount;
  output [2:0] ba_pad;
  output [12:0] a_pad;
  output [1:0] dm_pad;
  inout [15:0] dq_pad;
  inout [1:0] dqs_pad;
  inout [1:0] dqsbar_pad;
  input [2:0] cmd;
  input [15:0] din;
  input [1:0] sz;
  input [2:0] op;
  input [25:0] addr;
  input clk, reset, read, initddr, waiting;
  output notfull, ready, ck_pad, ckbar_pad, cke_pad, csbar_pad, rasbar_pad,
         casbar_pad, webar_pad, odt_pad, resetbar_pad, validout;
  wire   RETURN_put, RETURN_put_reg, ck_i, CMD_put, DATA_put, RETURN_get, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n139, n176, n183, n185, n186,
         n187, n188, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         reset_out, resetbar_i, DATA_get, CMD_get, CMD_empty, RETURN_full,
         init_rasbar, init_casbar, init_webar, init_cke, rasbar, casbar, webar,
         plogic_ts, plogic_ri, rasbar_i, casbar_i, webar_i, ts_i, ri_i, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, SYNOPSYS_UNCONNECTED_1,
         SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3,
         SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5,
         SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7,
         SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9,
         SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11,
         SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13,
         SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15,
         SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17,
         SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19,
         SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21,
         SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23,
         SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25;
  wire   [31:0] i;
  wire   [41:0] RETURN_data_out;
  wire   [33:0] CMD_data_out;
  wire   [15:0] dataOut;
  wire   [41:0] RETURN_data_in;
  wire   [1:0] init_ba;
  wire   [10:4] init_a;
  wire   [2:0] ba;
  wire   [12:0] a;
  wire   [1:0] dm_i;
  wire   [1:0] dqs_i;
  wire   [1:0] dqsbar_i;
  wire   [15:0] dq_i;
  wire   [1:0] dqs_o;
  wire   [1:0] dqsbar_o;
  wire   [15:0] dq_o;
  wire   [12:0] a_i;
  wire   [2:0] ba_i;

  INVX2 I_17 ( .A(reset), .Y(n360) );
  AND2X2 C983 ( .A(n360), .B(reset_out), .Y(resetbar_i) );
  AND2X2 C978 ( .A(n314), .B(n318), .Y(n139) );
  AND2X2 C973 ( .A(n599), .B(n69), .Y(n359) );
  AND2X2 C972 ( .A(n359), .B(n358), .Y(n70) );
  BUFX2 B_31 ( .A(RETURN_put), .Y(n34) );
  INVX2 I_10 ( .A(n357), .Y(n358) );
  OR2X2 C916 ( .A(n355), .B(n356), .Y(n357) );
  OR2X2 C915 ( .A(n354), .B(CMD_data_out[33]), .Y(n356) );
  INVX2 I_9 ( .A(CMD_data_out[31]), .Y(n355) );
  INVX2 I_8 ( .A(CMD_data_out[32]), .Y(n354) );
  OR2X2 C911 ( .A(n321), .B(n351), .Y(n352) );
  OR2X2 C910 ( .A(n320), .B(n350), .Y(n351) );
  OR2X2 C909 ( .A(i[2]), .B(n349), .Y(n350) );
  OR2X2 C908 ( .A(n319), .B(n348), .Y(n349) );
  OR2X2 C907 ( .A(i[4]), .B(n347), .Y(n348) );
  OR2X2 C906 ( .A(i[5]), .B(n346), .Y(n347) );
  OR2X2 C905 ( .A(i[6]), .B(n345), .Y(n346) );
  OR2X2 C904 ( .A(i[7]), .B(n344), .Y(n345) );
  OR2X2 C903 ( .A(i[8]), .B(n343), .Y(n344) );
  OR2X2 C902 ( .A(i[9]), .B(n342), .Y(n343) );
  OR2X2 C901 ( .A(i[10]), .B(n341), .Y(n342) );
  OR2X2 C900 ( .A(i[11]), .B(n340), .Y(n341) );
  OR2X2 C899 ( .A(i[12]), .B(n339), .Y(n340) );
  OR2X2 C898 ( .A(i[13]), .B(n338), .Y(n339) );
  OR2X2 C897 ( .A(i[14]), .B(n337), .Y(n338) );
  OR2X2 C896 ( .A(i[15]), .B(n336), .Y(n337) );
  OR2X2 C895 ( .A(i[16]), .B(n335), .Y(n336) );
  OR2X2 C894 ( .A(i[17]), .B(n334), .Y(n335) );
  OR2X2 C893 ( .A(i[18]), .B(n333), .Y(n334) );
  OR2X2 C892 ( .A(i[19]), .B(n332), .Y(n333) );
  OR2X2 C891 ( .A(i[20]), .B(n331), .Y(n332) );
  OR2X2 C890 ( .A(i[21]), .B(n330), .Y(n331) );
  OR2X2 C889 ( .A(i[22]), .B(n329), .Y(n330) );
  OR2X2 C888 ( .A(i[23]), .B(n328), .Y(n329) );
  OR2X2 C887 ( .A(i[24]), .B(n327), .Y(n328) );
  OR2X2 C886 ( .A(i[25]), .B(n326), .Y(n327) );
  OR2X2 C885 ( .A(i[26]), .B(n325), .Y(n326) );
  OR2X2 C884 ( .A(i[27]), .B(n324), .Y(n325) );
  OR2X2 C883 ( .A(i[28]), .B(n323), .Y(n324) );
  OR2X2 C882 ( .A(i[29]), .B(n322), .Y(n323) );
  OR2X2 C881 ( .A(i[30]), .B(i[31]), .Y(n322) );
  INVX2 I_6 ( .A(i[0]), .Y(n321) );
  INVX2 I_5 ( .A(i[1]), .Y(n320) );
  INVX2 I_4 ( .A(i[3]), .Y(n319) );
  INVX2 I_3 ( .A(n317), .Y(n318) );
  OR2X2 C876 ( .A(n315), .B(n316), .Y(n317) );
  OR2X2 C875 ( .A(CMD_data_out[32]), .B(CMD_data_out[33]), .Y(n316) );
  INVX2 I_2 ( .A(CMD_data_out[31]), .Y(n315) );
  INVX2 I_1 ( .A(n313), .Y(n314) );
  OR2X2 C872 ( .A(i[0]), .B(n312), .Y(n313) );
  OR2X2 C871 ( .A(i[1]), .B(n311), .Y(n312) );
  OR2X2 C870 ( .A(n282), .B(n310), .Y(n311) );
  OR2X2 C864 ( .A(i[8]), .B(n304), .Y(n305) );
  OR2X2 C863 ( .A(i[9]), .B(n303), .Y(n304) );
  OR2X2 C862 ( .A(i[10]), .B(n302), .Y(n303) );
  OR2X2 C861 ( .A(i[11]), .B(n301), .Y(n302) );
  OR2X2 C860 ( .A(i[12]), .B(n300), .Y(n301) );
  OR2X2 C859 ( .A(i[13]), .B(n299), .Y(n300) );
  OR2X2 C858 ( .A(i[14]), .B(n298), .Y(n299) );
  OR2X2 C857 ( .A(i[15]), .B(n297), .Y(n298) );
  OR2X2 C856 ( .A(i[16]), .B(n296), .Y(n297) );
  OR2X2 C855 ( .A(n566), .B(i[17]), .Y(n296) );
  OR2X2 C852 ( .A(i[20]), .B(n292), .Y(n293) );
  OR2X2 C851 ( .A(i[21]), .B(n291), .Y(n292) );
  OR2X2 C850 ( .A(i[22]), .B(n290), .Y(n291) );
  OR2X2 C849 ( .A(i[23]), .B(n289), .Y(n290) );
  OR2X2 C848 ( .A(i[24]), .B(n288), .Y(n289) );
  OR2X2 C847 ( .A(i[25]), .B(n287), .Y(n288) );
  OR2X2 C846 ( .A(i[26]), .B(n286), .Y(n287) );
  OR2X2 C845 ( .A(i[27]), .B(n285), .Y(n286) );
  OR2X2 C844 ( .A(i[28]), .B(n284), .Y(n285) );
  OR2X2 C843 ( .A(i[29]), .B(n283), .Y(n284) );
  OR2X2 C842 ( .A(i[30]), .B(i[31]), .Y(n283) );
  INVX2 I_0 ( .A(i[2]), .Y(n282) );
  DFFPOSX1 DATA_put_reg ( .D(n185), .CLK(clk), .Q(DATA_put) );
  DFFPOSX1 CMD_put_reg ( .D(n185), .CLK(clk), .Q(CMD_put) );
  DFFPOSX1 ck_i_reg ( .D(n602), .CLK(clk), .Q(ck_i) );
  DFFPOSX1 RETURN_put_reg_reg ( .D(n551), .CLK(clk), .Q(RETURN_put_reg) );
  DFFPOSX1 RETURN_get_reg ( .D(n519), .CLK(clk), .Q(RETURN_get) );
  DFFPOSX1 i_reg_31_ ( .D(n552), .CLK(clk), .Q(i[31]) );
  DFFPOSX1 i_reg_0_ ( .D(n550), .CLK(clk), .Q(i[0]) );
  DFFPOSX1 i_reg_1_ ( .D(n549), .CLK(clk), .Q(i[1]) );
  DFFPOSX1 i_reg_2_ ( .D(n548), .CLK(clk), .Q(i[2]) );
  DFFPOSX1 i_reg_3_ ( .D(n547), .CLK(clk), .Q(i[3]) );
  DFFPOSX1 i_reg_4_ ( .D(n546), .CLK(clk), .Q(i[4]) );
  DFFPOSX1 i_reg_5_ ( .D(n545), .CLK(clk), .Q(i[5]) );
  DFFPOSX1 i_reg_6_ ( .D(n544), .CLK(clk), .Q(i[6]) );
  DFFPOSX1 i_reg_7_ ( .D(n543), .CLK(clk), .Q(i[7]) );
  DFFPOSX1 i_reg_8_ ( .D(n542), .CLK(clk), .Q(i[8]) );
  DFFPOSX1 i_reg_9_ ( .D(n541), .CLK(clk), .Q(i[9]) );
  DFFPOSX1 i_reg_10_ ( .D(n540), .CLK(clk), .Q(i[10]) );
  DFFPOSX1 i_reg_11_ ( .D(n539), .CLK(clk), .Q(i[11]) );
  DFFPOSX1 i_reg_12_ ( .D(n538), .CLK(clk), .Q(i[12]) );
  DFFPOSX1 i_reg_13_ ( .D(n537), .CLK(clk), .Q(i[13]) );
  DFFPOSX1 i_reg_14_ ( .D(n536), .CLK(clk), .Q(i[14]) );
  DFFPOSX1 i_reg_15_ ( .D(n535), .CLK(clk), .Q(i[15]) );
  DFFPOSX1 i_reg_16_ ( .D(n534), .CLK(clk), .Q(i[16]) );
  DFFPOSX1 i_reg_17_ ( .D(n533), .CLK(clk), .Q(i[17]) );
  DFFPOSX1 i_reg_18_ ( .D(n532), .CLK(clk), .Q(i[18]) );
  DFFPOSX1 i_reg_19_ ( .D(n531), .CLK(clk), .Q(i[19]) );
  DFFPOSX1 i_reg_20_ ( .D(n530), .CLK(clk), .Q(i[20]) );
  DFFPOSX1 i_reg_21_ ( .D(n529), .CLK(clk), .Q(i[21]) );
  DFFPOSX1 i_reg_22_ ( .D(n528), .CLK(clk), .Q(i[22]) );
  DFFPOSX1 i_reg_23_ ( .D(n527), .CLK(clk), .Q(i[23]) );
  DFFPOSX1 i_reg_24_ ( .D(n526), .CLK(clk), .Q(i[24]) );
  DFFPOSX1 i_reg_25_ ( .D(n525), .CLK(clk), .Q(i[25]) );
  DFFPOSX1 i_reg_26_ ( .D(n524), .CLK(clk), .Q(i[26]) );
  DFFPOSX1 i_reg_27_ ( .D(n523), .CLK(clk), .Q(i[27]) );
  DFFPOSX1 i_reg_28_ ( .D(n522), .CLK(clk), .Q(i[28]) );
  DFFPOSX1 i_reg_29_ ( .D(n521), .CLK(clk), .Q(i[29]) );
  DFFPOSX1 i_reg_30_ ( .D(n520), .CLK(clk), .Q(i[30]) );
  DFFPOSX1 raddr_reg_25_ ( .D(n477), .CLK(clk), .Q(raddr[25]) );
  DFFPOSX1 raddr_reg_24_ ( .D(n478), .CLK(clk), .Q(raddr[24]) );
  DFFPOSX1 raddr_reg_23_ ( .D(n479), .CLK(clk), .Q(raddr[23]) );
  DFFPOSX1 raddr_reg_22_ ( .D(n480), .CLK(clk), .Q(raddr[22]) );
  DFFPOSX1 raddr_reg_21_ ( .D(n481), .CLK(clk), .Q(raddr[21]) );
  DFFPOSX1 raddr_reg_20_ ( .D(n482), .CLK(clk), .Q(raddr[20]) );
  DFFPOSX1 raddr_reg_19_ ( .D(n483), .CLK(clk), .Q(raddr[19]) );
  DFFPOSX1 raddr_reg_18_ ( .D(n484), .CLK(clk), .Q(raddr[18]) );
  DFFPOSX1 raddr_reg_17_ ( .D(n485), .CLK(clk), .Q(raddr[17]) );
  DFFPOSX1 raddr_reg_16_ ( .D(n486), .CLK(clk), .Q(raddr[16]) );
  DFFPOSX1 raddr_reg_15_ ( .D(n487), .CLK(clk), .Q(raddr[15]) );
  DFFPOSX1 raddr_reg_14_ ( .D(n488), .CLK(clk), .Q(raddr[14]) );
  DFFPOSX1 raddr_reg_13_ ( .D(n489), .CLK(clk), .Q(raddr[13]) );
  DFFPOSX1 raddr_reg_12_ ( .D(n490), .CLK(clk), .Q(raddr[12]) );
  DFFPOSX1 raddr_reg_11_ ( .D(n491), .CLK(clk), .Q(raddr[11]) );
  DFFPOSX1 raddr_reg_10_ ( .D(n492), .CLK(clk), .Q(raddr[10]) );
  DFFPOSX1 raddr_reg_9_ ( .D(n493), .CLK(clk), .Q(raddr[9]) );
  DFFPOSX1 raddr_reg_8_ ( .D(n494), .CLK(clk), .Q(raddr[8]) );
  DFFPOSX1 raddr_reg_7_ ( .D(n495), .CLK(clk), .Q(raddr[7]) );
  DFFPOSX1 raddr_reg_6_ ( .D(n496), .CLK(clk), .Q(raddr[6]) );
  DFFPOSX1 raddr_reg_5_ ( .D(n497), .CLK(clk), .Q(raddr[5]) );
  DFFPOSX1 raddr_reg_4_ ( .D(n498), .CLK(clk), .Q(raddr[4]) );
  DFFPOSX1 raddr_reg_3_ ( .D(n499), .CLK(clk), .Q(raddr[3]) );
  DFFPOSX1 raddr_reg_2_ ( .D(n500), .CLK(clk), .Q(raddr[2]) );
  DFFPOSX1 raddr_reg_1_ ( .D(n501), .CLK(clk), .Q(raddr[1]) );
  DFFPOSX1 raddr_reg_0_ ( .D(n502), .CLK(clk), .Q(raddr[0]) );
  DFFPOSX1 dout_reg_15_ ( .D(n503), .CLK(clk), .Q(dout[15]) );
  DFFPOSX1 dout_reg_14_ ( .D(n504), .CLK(clk), .Q(dout[14]) );
  DFFPOSX1 dout_reg_13_ ( .D(n505), .CLK(clk), .Q(dout[13]) );
  DFFPOSX1 dout_reg_12_ ( .D(n506), .CLK(clk), .Q(dout[12]) );
  DFFPOSX1 dout_reg_11_ ( .D(n507), .CLK(clk), .Q(dout[11]) );
  DFFPOSX1 dout_reg_10_ ( .D(n508), .CLK(clk), .Q(dout[10]) );
  DFFPOSX1 dout_reg_9_ ( .D(n509), .CLK(clk), .Q(dout[9]) );
  DFFPOSX1 dout_reg_8_ ( .D(n510), .CLK(clk), .Q(dout[8]) );
  DFFPOSX1 dout_reg_7_ ( .D(n511), .CLK(clk), .Q(dout[7]) );
  DFFPOSX1 dout_reg_6_ ( .D(n512), .CLK(clk), .Q(dout[6]) );
  DFFPOSX1 dout_reg_5_ ( .D(n513), .CLK(clk), .Q(dout[5]) );
  DFFPOSX1 dout_reg_4_ ( .D(n514), .CLK(clk), .Q(dout[4]) );
  DFFPOSX1 dout_reg_3_ ( .D(n515), .CLK(clk), .Q(dout[3]) );
  DFFPOSX1 dout_reg_2_ ( .D(n516), .CLK(clk), .Q(dout[2]) );
  DFFPOSX1 dout_reg_1_ ( .D(n517), .CLK(clk), .Q(dout[1]) );
  DFFPOSX1 dout_reg_0_ ( .D(n656), .CLK(clk), .Q(dout[0]) );
  DFFPOSX1 validout_reg ( .D(n476), .CLK(clk), .Q(validout) );
  INVX1 U3 ( .A(n367), .Y(webar_i) );
  AOI22X1 U4 ( .A(init_webar), .B(n368), .C(webar), .D(ready), .Y(n367) );
  INVX1 U5 ( .A(n597), .Y(ts_i) );
  AND2X1 U10 ( .A(plogic_ri), .B(ready), .Y(ri_i) );
  INVX1 U11 ( .A(n370), .Y(rasbar_i) );
  AOI22X1 U12 ( .A(init_rasbar), .B(n368), .C(rasbar), .D(ready), .Y(n370) );
  INVX1 U13 ( .A(n371), .Y(n265) );
  OAI21X1 U14 ( .A(n372), .B(n34), .C(n185), .Y(n371) );
  OAI21X1 U15 ( .A(n35), .B(n368), .C(n373), .Y(n264) );
  AND2X1 U16 ( .A(n67), .B(n374), .Y(n263) );
  AND2X1 U17 ( .A(n66), .B(n374), .Y(n262) );
  AND2X1 U18 ( .A(n65), .B(n374), .Y(n261) );
  AND2X1 U19 ( .A(n64), .B(n374), .Y(n260) );
  AND2X1 U20 ( .A(n63), .B(n374), .Y(n259) );
  AND2X1 U21 ( .A(n62), .B(n374), .Y(n258) );
  AND2X1 U22 ( .A(n61), .B(n374), .Y(n257) );
  AND2X1 U23 ( .A(n60), .B(n374), .Y(n256) );
  AND2X1 U24 ( .A(n59), .B(n374), .Y(n255) );
  AND2X1 U25 ( .A(n58), .B(n374), .Y(n254) );
  AND2X1 U26 ( .A(n57), .B(n374), .Y(n253) );
  AND2X1 U27 ( .A(n56), .B(n374), .Y(n252) );
  AND2X1 U28 ( .A(n55), .B(n374), .Y(n251) );
  AND2X1 U29 ( .A(n54), .B(n374), .Y(n250) );
  AND2X1 U30 ( .A(n53), .B(n374), .Y(n249) );
  AND2X1 U31 ( .A(n52), .B(n374), .Y(n248) );
  AND2X1 U32 ( .A(n51), .B(n374), .Y(n247) );
  AND2X1 U33 ( .A(n50), .B(n374), .Y(n246) );
  AND2X1 U34 ( .A(n49), .B(n374), .Y(n245) );
  AND2X1 U35 ( .A(n48), .B(n374), .Y(n244) );
  AND2X1 U36 ( .A(n47), .B(n374), .Y(n243) );
  AND2X1 U37 ( .A(n46), .B(n374), .Y(n242) );
  AND2X1 U38 ( .A(n45), .B(n374), .Y(n241) );
  AND2X1 U39 ( .A(n44), .B(n374), .Y(n240) );
  AND2X1 U40 ( .A(n43), .B(n374), .Y(n239) );
  AND2X1 U41 ( .A(n42), .B(n374), .Y(n238) );
  AND2X1 U42 ( .A(n41), .B(n374), .Y(n237) );
  AND2X1 U43 ( .A(n40), .B(n374), .Y(n236) );
  AND2X1 U44 ( .A(n39), .B(n374), .Y(n235) );
  AND2X1 U45 ( .A(n38), .B(n374), .Y(n234) );
  AND2X1 U46 ( .A(n37), .B(n374), .Y(n233) );
  AND2X1 U50 ( .A(RETURN_data_out[41]), .B(n373), .Y(n231) );
  AND2X1 U51 ( .A(RETURN_data_out[40]), .B(n373), .Y(n230) );
  AND2X1 U52 ( .A(RETURN_data_out[39]), .B(n373), .Y(n229) );
  AND2X1 U53 ( .A(RETURN_data_out[38]), .B(n373), .Y(n228) );
  AND2X1 U54 ( .A(RETURN_data_out[37]), .B(n373), .Y(n227) );
  AND2X1 U55 ( .A(RETURN_data_out[36]), .B(n373), .Y(n226) );
  AND2X1 U56 ( .A(RETURN_data_out[35]), .B(n373), .Y(n225) );
  AND2X1 U57 ( .A(RETURN_data_out[34]), .B(n373), .Y(n224) );
  AND2X1 U58 ( .A(RETURN_data_out[33]), .B(n373), .Y(n223) );
  AND2X1 U59 ( .A(RETURN_data_out[32]), .B(n373), .Y(n222) );
  AND2X1 U60 ( .A(RETURN_data_out[31]), .B(n373), .Y(n221) );
  AND2X1 U61 ( .A(RETURN_data_out[30]), .B(n373), .Y(n220) );
  AND2X1 U62 ( .A(RETURN_data_out[29]), .B(n373), .Y(n219) );
  AND2X1 U63 ( .A(RETURN_data_out[28]), .B(n373), .Y(n218) );
  AND2X1 U64 ( .A(RETURN_data_out[27]), .B(n373), .Y(n217) );
  AND2X1 U65 ( .A(RETURN_data_out[26]), .B(n373), .Y(n216) );
  AND2X1 U66 ( .A(RETURN_data_out[25]), .B(n373), .Y(n215) );
  AND2X1 U67 ( .A(RETURN_data_out[24]), .B(n373), .Y(n214) );
  AND2X1 U68 ( .A(RETURN_data_out[23]), .B(n373), .Y(n213) );
  AND2X1 U69 ( .A(RETURN_data_out[22]), .B(n373), .Y(n212) );
  AND2X1 U70 ( .A(RETURN_data_out[21]), .B(n373), .Y(n211) );
  AND2X1 U71 ( .A(RETURN_data_out[20]), .B(n373), .Y(n210) );
  AND2X1 U72 ( .A(RETURN_data_out[19]), .B(n373), .Y(n209) );
  AND2X1 U73 ( .A(RETURN_data_out[18]), .B(n373), .Y(n208) );
  AND2X1 U74 ( .A(RETURN_data_out[17]), .B(n373), .Y(n207) );
  AND2X1 U75 ( .A(RETURN_data_out[16]), .B(n373), .Y(n206) );
  AND2X1 U76 ( .A(RETURN_data_out[15]), .B(n373), .Y(n205) );
  AND2X1 U77 ( .A(RETURN_data_out[14]), .B(n373), .Y(n204) );
  AND2X1 U78 ( .A(RETURN_data_out[13]), .B(n373), .Y(n203) );
  AND2X1 U79 ( .A(RETURN_data_out[12]), .B(n373), .Y(n202) );
  AND2X1 U80 ( .A(RETURN_data_out[11]), .B(n373), .Y(n201) );
  AND2X1 U81 ( .A(RETURN_data_out[10]), .B(n373), .Y(n200) );
  AND2X1 U82 ( .A(RETURN_data_out[9]), .B(n373), .Y(n199) );
  AND2X1 U83 ( .A(RETURN_data_out[8]), .B(n373), .Y(n198) );
  AND2X1 U84 ( .A(RETURN_data_out[7]), .B(n373), .Y(n197) );
  AND2X1 U85 ( .A(RETURN_data_out[6]), .B(n373), .Y(n196) );
  AND2X1 U86 ( .A(RETURN_data_out[5]), .B(n373), .Y(n195) );
  AND2X1 U87 ( .A(RETURN_data_out[4]), .B(n373), .Y(n194) );
  AND2X1 U88 ( .A(RETURN_data_out[3]), .B(n373), .Y(n193) );
  AND2X1 U89 ( .A(RETURN_data_out[2]), .B(n373), .Y(n192) );
  AND2X1 U90 ( .A(RETURN_data_out[1]), .B(n373), .Y(n191) );
  NAND3X1 U93 ( .A(n379), .B(n380), .C(ready), .Y(n378) );
  AND2X1 U94 ( .A(n186), .B(n379), .Y(n188) );
  AND2X1 U97 ( .A(n380), .B(n373), .Y(n186) );
  INVX1 U98 ( .A(n35), .Y(n380) );
  AND2X1 U99 ( .A(ready), .B(n373), .Y(n185) );
  INVX1 U100 ( .A(reset), .Y(n373) );
  INVX1 U102 ( .A(n372), .Y(n176) );
  INVX1 U105 ( .A(n139), .Y(n376) );
  INVX1 U108 ( .A(n382), .Y(casbar_i) );
  AOI22X1 U109 ( .A(casbar), .B(ready), .C(init_casbar), .D(n368), .Y(n382) );
  INVX1 U110 ( .A(n586), .Y(ba_i[2]) );
  INVX1 U112 ( .A(n384), .Y(ba_i[1]) );
  AOI22X1 U113 ( .A(ba[1]), .B(ready), .C(init_ba[1]), .D(n368), .Y(n384) );
  INVX1 U114 ( .A(n385), .Y(ba_i[0]) );
  AOI22X1 U115 ( .A(ba[0]), .B(ready), .C(init_ba[0]), .D(n368), .Y(n385) );
  INVX1 U116 ( .A(n589), .Y(a_i[9]) );
  INVX1 U118 ( .A(n387), .Y(a_i[8]) );
  AOI22X1 U119 ( .A(a[8]), .B(ready), .C(init_a[8]), .D(n368), .Y(n387) );
  INVX1 U120 ( .A(n590), .Y(a_i[7]) );
  INVX1 U122 ( .A(n591), .Y(a_i[6]) );
  INVX1 U124 ( .A(n592), .Y(a_i[5]) );
  INVX1 U126 ( .A(n391), .Y(a_i[4]) );
  AOI22X1 U127 ( .A(a[4]), .B(ready), .C(init_a[4]), .D(n368), .Y(n391) );
  INVX1 U128 ( .A(n593), .Y(a_i[3]) );
  INVX1 U130 ( .A(n594), .Y(a_i[2]) );
  INVX1 U132 ( .A(n595), .Y(a_i[1]) );
  INVX1 U134 ( .A(n587), .Y(a_i[12]) );
  INVX1 U136 ( .A(n588), .Y(a_i[11]) );
  INVX1 U138 ( .A(n397), .Y(a_i[10]) );
  AOI22X1 U139 ( .A(a[10]), .B(ready), .C(init_a[10]), .D(n368), .Y(n397) );
  INVX1 U140 ( .A(n596), .Y(a_i[0]) );
  INVX1 U142 ( .A(ready), .Y(n368) );
  MUX2X1 U143 ( .B(n558), .A(n263), .S(n264), .Y(n399) );
  INVX2 U144 ( .A(n399), .Y(n552) );
  MUX2X1 U145 ( .B(RETURN_put_reg), .A(n176), .S(n265), .Y(n400) );
  INVX2 U146 ( .A(n400), .Y(n551) );
  MUX2X1 U147 ( .B(i[0]), .A(n232), .S(n264), .Y(n401) );
  INVX2 U148 ( .A(n401), .Y(n550) );
  MUX2X1 U149 ( .B(i[1]), .A(n233), .S(n264), .Y(n402) );
  INVX2 U150 ( .A(n402), .Y(n549) );
  MUX2X1 U151 ( .B(i[2]), .A(n234), .S(n264), .Y(n403) );
  INVX2 U152 ( .A(n403), .Y(n548) );
  MUX2X1 U153 ( .B(i[3]), .A(n235), .S(n264), .Y(n404) );
  INVX2 U154 ( .A(n404), .Y(n547) );
  MUX2X1 U155 ( .B(i[4]), .A(n236), .S(n264), .Y(n405) );
  INVX2 U156 ( .A(n405), .Y(n546) );
  MUX2X1 U157 ( .B(i[5]), .A(n237), .S(n264), .Y(n406) );
  INVX2 U158 ( .A(n406), .Y(n545) );
  MUX2X1 U159 ( .B(i[6]), .A(n238), .S(n264), .Y(n407) );
  INVX2 U160 ( .A(n407), .Y(n544) );
  MUX2X1 U161 ( .B(i[7]), .A(n239), .S(n264), .Y(n408) );
  INVX2 U162 ( .A(n408), .Y(n543) );
  MUX2X1 U163 ( .B(i[8]), .A(n240), .S(n264), .Y(n409) );
  INVX2 U164 ( .A(n409), .Y(n542) );
  MUX2X1 U165 ( .B(i[9]), .A(n241), .S(n264), .Y(n410) );
  INVX2 U166 ( .A(n410), .Y(n541) );
  MUX2X1 U167 ( .B(i[10]), .A(n242), .S(n264), .Y(n411) );
  INVX2 U168 ( .A(n411), .Y(n540) );
  MUX2X1 U169 ( .B(i[11]), .A(n243), .S(n264), .Y(n412) );
  INVX2 U170 ( .A(n412), .Y(n539) );
  MUX2X1 U171 ( .B(i[12]), .A(n244), .S(n264), .Y(n413) );
  INVX2 U172 ( .A(n413), .Y(n538) );
  MUX2X1 U173 ( .B(i[13]), .A(n245), .S(n264), .Y(n414) );
  INVX2 U174 ( .A(n414), .Y(n537) );
  MUX2X1 U175 ( .B(i[14]), .A(n246), .S(n264), .Y(n415) );
  INVX2 U176 ( .A(n415), .Y(n536) );
  MUX2X1 U177 ( .B(i[15]), .A(n247), .S(n264), .Y(n416) );
  INVX2 U178 ( .A(n416), .Y(n535) );
  MUX2X1 U179 ( .B(i[16]), .A(n248), .S(n264), .Y(n417) );
  INVX2 U180 ( .A(n417), .Y(n534) );
  MUX2X1 U181 ( .B(i[17]), .A(n249), .S(n264), .Y(n418) );
  INVX2 U182 ( .A(n418), .Y(n533) );
  MUX2X1 U183 ( .B(i[18]), .A(n250), .S(n264), .Y(n419) );
  INVX2 U184 ( .A(n419), .Y(n532) );
  MUX2X1 U185 ( .B(i[19]), .A(n251), .S(n264), .Y(n420) );
  INVX2 U186 ( .A(n420), .Y(n531) );
  MUX2X1 U187 ( .B(i[20]), .A(n252), .S(n264), .Y(n421) );
  INVX2 U188 ( .A(n421), .Y(n530) );
  MUX2X1 U189 ( .B(i[21]), .A(n253), .S(n264), .Y(n422) );
  INVX2 U190 ( .A(n422), .Y(n529) );
  MUX2X1 U191 ( .B(i[22]), .A(n254), .S(n264), .Y(n423) );
  INVX2 U192 ( .A(n423), .Y(n528) );
  MUX2X1 U193 ( .B(i[23]), .A(n255), .S(n264), .Y(n424) );
  INVX2 U194 ( .A(n424), .Y(n527) );
  MUX2X1 U195 ( .B(i[24]), .A(n256), .S(n264), .Y(n425) );
  INVX2 U196 ( .A(n425), .Y(n526) );
  MUX2X1 U197 ( .B(i[25]), .A(n257), .S(n264), .Y(n426) );
  INVX2 U198 ( .A(n426), .Y(n525) );
  MUX2X1 U199 ( .B(i[26]), .A(n258), .S(n264), .Y(n427) );
  INVX2 U200 ( .A(n427), .Y(n524) );
  MUX2X1 U201 ( .B(i[27]), .A(n259), .S(n264), .Y(n428) );
  INVX2 U202 ( .A(n428), .Y(n523) );
  MUX2X1 U203 ( .B(i[28]), .A(n260), .S(n264), .Y(n429) );
  INVX2 U204 ( .A(n429), .Y(n522) );
  MUX2X1 U205 ( .B(i[29]), .A(n261), .S(n264), .Y(n430) );
  INVX2 U206 ( .A(n430), .Y(n521) );
  MUX2X1 U207 ( .B(n557), .A(n262), .S(n264), .Y(n431) );
  INVX2 U208 ( .A(n431), .Y(n520) );
  MUX2X1 U209 ( .B(RETURN_get), .A(n186), .S(n650), .Y(n432) );
  INVX2 U210 ( .A(n432), .Y(n519) );
  MUX2X1 U213 ( .B(dout[1]), .A(n191), .S(n568), .Y(n434) );
  MUX2X1 U215 ( .B(dout[2]), .A(n192), .S(n568), .Y(n435) );
  INVX2 U216 ( .A(n435), .Y(n516) );
  MUX2X1 U217 ( .B(dout[3]), .A(n193), .S(n568), .Y(n436) );
  INVX2 U218 ( .A(n436), .Y(n515) );
  MUX2X1 U219 ( .B(dout[4]), .A(n194), .S(n568), .Y(n437) );
  INVX2 U220 ( .A(n437), .Y(n514) );
  MUX2X1 U221 ( .B(dout[5]), .A(n195), .S(n568), .Y(n438) );
  INVX2 U222 ( .A(n438), .Y(n513) );
  MUX2X1 U223 ( .B(dout[6]), .A(n196), .S(n568), .Y(n439) );
  INVX2 U224 ( .A(n439), .Y(n512) );
  MUX2X1 U225 ( .B(dout[7]), .A(n197), .S(n568), .Y(n440) );
  INVX2 U226 ( .A(n440), .Y(n511) );
  MUX2X1 U227 ( .B(dout[8]), .A(n198), .S(n568), .Y(n441) );
  INVX2 U228 ( .A(n441), .Y(n510) );
  MUX2X1 U229 ( .B(dout[9]), .A(n199), .S(n568), .Y(n442) );
  INVX2 U230 ( .A(n442), .Y(n509) );
  MUX2X1 U231 ( .B(dout[10]), .A(n200), .S(n568), .Y(n443) );
  INVX2 U232 ( .A(n443), .Y(n508) );
  MUX2X1 U233 ( .B(dout[11]), .A(n201), .S(n568), .Y(n444) );
  INVX2 U234 ( .A(n444), .Y(n507) );
  MUX2X1 U235 ( .B(dout[12]), .A(n202), .S(n568), .Y(n445) );
  INVX2 U236 ( .A(n445), .Y(n506) );
  MUX2X1 U237 ( .B(dout[13]), .A(n203), .S(n568), .Y(n446) );
  INVX2 U238 ( .A(n446), .Y(n505) );
  MUX2X1 U239 ( .B(dout[14]), .A(n204), .S(n568), .Y(n447) );
  INVX2 U240 ( .A(n447), .Y(n504) );
  MUX2X1 U241 ( .B(dout[15]), .A(n205), .S(n568), .Y(n448) );
  INVX2 U242 ( .A(n448), .Y(n503) );
  MUX2X1 U243 ( .B(raddr[0]), .A(n206), .S(n568), .Y(n449) );
  INVX2 U244 ( .A(n449), .Y(n502) );
  MUX2X1 U245 ( .B(raddr[1]), .A(n207), .S(n568), .Y(n450) );
  INVX2 U246 ( .A(n450), .Y(n501) );
  MUX2X1 U247 ( .B(raddr[2]), .A(n208), .S(n568), .Y(n451) );
  INVX2 U248 ( .A(n451), .Y(n500) );
  MUX2X1 U249 ( .B(raddr[3]), .A(n209), .S(n568), .Y(n452) );
  INVX2 U250 ( .A(n452), .Y(n499) );
  MUX2X1 U251 ( .B(raddr[4]), .A(n210), .S(n568), .Y(n453) );
  INVX2 U252 ( .A(n453), .Y(n498) );
  MUX2X1 U253 ( .B(raddr[5]), .A(n211), .S(n568), .Y(n454) );
  INVX2 U254 ( .A(n454), .Y(n497) );
  MUX2X1 U255 ( .B(raddr[6]), .A(n212), .S(n568), .Y(n455) );
  INVX2 U256 ( .A(n455), .Y(n496) );
  MUX2X1 U257 ( .B(raddr[7]), .A(n213), .S(n568), .Y(n456) );
  INVX2 U258 ( .A(n456), .Y(n495) );
  MUX2X1 U259 ( .B(raddr[8]), .A(n214), .S(n568), .Y(n457) );
  INVX2 U260 ( .A(n457), .Y(n494) );
  MUX2X1 U261 ( .B(raddr[9]), .A(n215), .S(n568), .Y(n458) );
  INVX2 U262 ( .A(n458), .Y(n493) );
  MUX2X1 U263 ( .B(raddr[10]), .A(n216), .S(n568), .Y(n459) );
  INVX2 U264 ( .A(n459), .Y(n492) );
  MUX2X1 U265 ( .B(raddr[11]), .A(n217), .S(n568), .Y(n460) );
  INVX2 U266 ( .A(n460), .Y(n491) );
  MUX2X1 U267 ( .B(raddr[12]), .A(n218), .S(n568), .Y(n461) );
  INVX2 U268 ( .A(n461), .Y(n490) );
  MUX2X1 U269 ( .B(raddr[13]), .A(n219), .S(n568), .Y(n462) );
  INVX2 U270 ( .A(n462), .Y(n489) );
  MUX2X1 U271 ( .B(raddr[14]), .A(n220), .S(n568), .Y(n463) );
  INVX2 U272 ( .A(n463), .Y(n488) );
  MUX2X1 U273 ( .B(raddr[15]), .A(n221), .S(n568), .Y(n464) );
  INVX2 U274 ( .A(n464), .Y(n487) );
  MUX2X1 U275 ( .B(raddr[16]), .A(n222), .S(n568), .Y(n465) );
  INVX2 U276 ( .A(n465), .Y(n486) );
  MUX2X1 U277 ( .B(raddr[17]), .A(n223), .S(n568), .Y(n466) );
  INVX2 U278 ( .A(n466), .Y(n485) );
  MUX2X1 U279 ( .B(raddr[18]), .A(n224), .S(n568), .Y(n467) );
  INVX2 U280 ( .A(n467), .Y(n484) );
  MUX2X1 U281 ( .B(raddr[19]), .A(n225), .S(n568), .Y(n468) );
  INVX2 U282 ( .A(n468), .Y(n483) );
  MUX2X1 U283 ( .B(raddr[20]), .A(n226), .S(n568), .Y(n469) );
  INVX2 U284 ( .A(n469), .Y(n482) );
  MUX2X1 U285 ( .B(raddr[21]), .A(n227), .S(n568), .Y(n470) );
  INVX2 U286 ( .A(n470), .Y(n481) );
  MUX2X1 U287 ( .B(raddr[22]), .A(n228), .S(n568), .Y(n471) );
  INVX2 U288 ( .A(n471), .Y(n480) );
  MUX2X1 U289 ( .B(raddr[23]), .A(n229), .S(n568), .Y(n472) );
  INVX2 U290 ( .A(n472), .Y(n479) );
  MUX2X1 U291 ( .B(raddr[24]), .A(n230), .S(n568), .Y(n473) );
  INVX2 U292 ( .A(n473), .Y(n478) );
  MUX2X1 U293 ( .B(raddr[25]), .A(n231), .S(n568), .Y(n474) );
  INVX2 U294 ( .A(n474), .Y(n477) );
  MUX2X1 U295 ( .B(validout), .A(n188), .S(n650), .Y(n475) );
  INVX2 U296 ( .A(n475), .Y(n476) );
  FIFO_2clk_DATA_WIDTH16_FIFO_DEPTH32_PTR_WIDTH6 FIFO_DATA ( .rclk(clk), 
        .wclk(clk), .reset(reset), .we(DATA_put), .re(DATA_get), .data_in(din), 
        .empty_bar(), .full_bar(), .data_out(dataOut), .fillcount(fillcount)
         );
  FIFO_2clk_DATA_WIDTH34_FIFO_DEPTH32_PTR_WIDTH6 FIFO_CMD ( .rclk(clk), .wclk(
        clk), .reset(reset), .we(CMD_put), .re(CMD_get), .data_in({cmd, sz, op, 
        addr}), .empty_bar(CMD_empty), .full_bar(notfull), .data_out(
        CMD_data_out), .fillcount({SYNOPSYS_UNCONNECTED_1, 
        SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, 
        SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6}) );
  FIFO_2clk_DATA_WIDTH42_FIFO_DEPTH32_PTR_WIDTH6 FIFO_RETURN ( .rclk(clk), 
        .wclk(clk), .reset(reset), .we(RETURN_put), .re(RETURN_get), .data_in(
        RETURN_data_in), .empty_bar(), .full_bar(RETURN_full), .data_out(
        RETURN_data_out), .fillcount({SYNOPSYS_UNCONNECTED_7, 
        SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12}) );
  ddr3_init_engine XINIT ( .ready(ready), .csbar(), .rasbar(init_rasbar), 
        .casbar(init_casbar), .webar(init_webar), .ba({SYNOPSYS_UNCONNECTED_13, 
        init_ba}), .a({SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        init_a[10], SYNOPSYS_UNCONNECTED_16, init_a[8], 
        SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18, 
        SYNOPSYS_UNCONNECTED_19, init_a[4], SYNOPSYS_UNCONNECTED_20, 
        SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22, 
        SYNOPSYS_UNCONNECTED_23}), .odt(), .ts_con(), .cke(init_cke), .clk(clk), .reset(reset), .init(initddr), .ck(1'b0), .reset_out(reset_out) );
  Processing_logic PLOGIC ( .clk(clk), .ck(ck_i), .reset(reset), .ready(ready), 
        .DATA_data_out(dataOut), .DATA_get(DATA_get), .CMD_empty(CMD_empty), 
        .CMD_data_out(CMD_data_out), .CMD_get(CMD_get), .RETURN_full(
        RETURN_full), .RETURN_put(RETURN_put), .RETURN_address(
        RETURN_data_in[41:16]), .RETURN_data(RETURN_data_in[15:0]), .DQ_in(
        dq_o), .DQS_in(dqs_o), .DQS_bar_in(dqsbar_o), .cs_bar(), .ras_bar(
        rasbar), .cas_bar(casbar), .we_bar(webar), .DQ_out(dq_i), .DQS_out(
        dqs_i), .DQS_bar_out(dqsbar_i), .BA(ba), .A(a), .DM({
        SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25}), .ts_con(plogic_ts), 
        .ri_o(plogic_ri) );
  SSTL18DDR3INTERFACE XSSTL ( .ck_pad(ck_pad), .ckbar_pad(ckbar_pad), 
        .cke_pad(cke_pad), .csbar_pad(csbar_pad), .rasbar_pad(rasbar_pad), 
        .casbar_pad(casbar_pad), .webar_pad(webar_pad), .ba_pad(ba_pad), 
        .a_pad(a_pad), .dm_pad(dm_pad), .odt_pad(odt_pad), .resetbar_pad(
        resetbar_pad), .dq_o(dq_o), .dqs_o(dqs_o), .dqsbar_o(dqsbar_o), 
        .dq_pad(dq_pad), .dqs_pad(dqs_pad), .dqsbar_pad(dqsbar_pad), .ri_i(
        ri_i), .ts_i(ts_i), .ck_i(ck_i), .cke_i(init_cke), .csbar_i(1'b0), 
        .rasbar_i(rasbar_i), .casbar_i(casbar_i), .webar_i(webar_i), .ba_i(
        ba_i), .a_i(a_i), .dq_i(dq_i), .dqs_i(dqs_i), .dqsbar_i(dqsbar_i), 
        .dm_i({1'b0, 1'b0}), .odt_i(1'b0), .resetbar_i(resetbar_i) );
  ddr3_controller_DW01_inc_0 add_144 ( .A({n558, n557, i[29:0]}), .SUM({n67, 
        n66, n65, n64, n63, n62, n61, n60, n59, n58, n57, n56, n55, n54, n53, 
        n52, n51, n50, n49, n48, n47, n46, n45, n44, n43, n42, n41, n40, n39, 
        n38, n37, n36}) );
  OR2X2 U297 ( .A(n305), .B(i[7]), .Y(n553) );
  OR2X2 U298 ( .A(i[5]), .B(i[6]), .Y(n554) );
  OR2X2 U299 ( .A(n553), .B(n554), .Y(n555) );
  OR2X2 U300 ( .A(n555), .B(n556), .Y(n310) );
  OR2X2 U301 ( .A(i[3]), .B(i[4]), .Y(n556) );
  INVX1 U302 ( .A(n434), .Y(n517) );
  INVX2 U303 ( .A(n568), .Y(n655) );
  INVX8 U304 ( .A(n654), .Y(n568) );
  BUFX2 U305 ( .A(i[30]), .Y(n557) );
  INVX1 U306 ( .A(n692), .Y(n558) );
  AND2X1 U307 ( .A(n373), .B(n564), .Y(n654) );
  OR2X2 U308 ( .A(i[28]), .B(i[27]), .Y(n679) );
  INVX1 U309 ( .A(n679), .Y(n559) );
  OR2X2 U310 ( .A(i[30]), .B(i[29]), .Y(n678) );
  INVX1 U311 ( .A(n678), .Y(n560) );
  OR2X2 U312 ( .A(n571), .B(n567), .Y(n640) );
  INVX1 U313 ( .A(n640), .Y(n561) );
  OR2X2 U314 ( .A(n646), .B(n647), .Y(n643) );
  INVX1 U315 ( .A(n643), .Y(n562) );
  OR2X2 U316 ( .A(n644), .B(n645), .Y(n648) );
  INVX1 U317 ( .A(n648), .Y(n563) );
  BUFX2 U318 ( .A(n378), .Y(n564) );
  OR2X2 U319 ( .A(i[19]), .B(n293), .Y(n653) );
  INVX1 U320 ( .A(n653), .Y(n565) );
  AND2X2 U321 ( .A(n652), .B(n565), .Y(n295) );
  INVX1 U322 ( .A(n295), .Y(n566) );
  OR2X2 U323 ( .A(n569), .B(n35), .Y(n641) );
  INVX1 U324 ( .A(n641), .Y(n567) );
  AND2X2 U325 ( .A(n70), .B(n353), .Y(n377) );
  INVX1 U326 ( .A(n377), .Y(n569) );
  INVX1 U327 ( .A(n377), .Y(n570) );
  OR2X2 U328 ( .A(n376), .B(n35), .Y(n642) );
  INVX1 U329 ( .A(n642), .Y(n571) );
  INVX1 U330 ( .A(n574), .Y(n572) );
  INVX1 U331 ( .A(n572), .Y(n573) );
  BUFX2 U332 ( .A(n559), .Y(n574) );
  INVX1 U333 ( .A(n577), .Y(n575) );
  INVX1 U334 ( .A(n575), .Y(n576) );
  BUFX2 U335 ( .A(n683), .Y(n577) );
  OR2X1 U336 ( .A(n628), .B(n629), .Y(n625) );
  INVX1 U337 ( .A(n625), .Y(n578) );
  OR2X1 U338 ( .A(n626), .B(n627), .Y(n630) );
  INVX1 U339 ( .A(n630), .Y(n579) );
  OR2X1 U340 ( .A(n637), .B(n638), .Y(n634) );
  INVX1 U341 ( .A(n634), .Y(n580) );
  OR2X1 U342 ( .A(n635), .B(n636), .Y(n639) );
  INVX1 U343 ( .A(n639), .Y(n581) );
  OR2X1 U344 ( .A(i[20]), .B(i[19]), .Y(n668) );
  INVX1 U345 ( .A(n668), .Y(n582) );
  OR2X1 U346 ( .A(i[22]), .B(i[21]), .Y(n667) );
  INVX1 U347 ( .A(n667), .Y(n583) );
  OR2X1 U348 ( .A(i[11]), .B(i[10]), .Y(n672) );
  INVX1 U349 ( .A(n672), .Y(n584) );
  AND2X2 U350 ( .A(i[3]), .B(i[2]), .Y(n671) );
  INVX1 U351 ( .A(n671), .Y(n585) );
  AND2X2 U352 ( .A(ba[2]), .B(ready), .Y(n383) );
  INVX1 U353 ( .A(n383), .Y(n586) );
  AND2X2 U354 ( .A(a[12]), .B(ready), .Y(n395) );
  INVX1 U355 ( .A(n395), .Y(n587) );
  AND2X2 U356 ( .A(a[11]), .B(ready), .Y(n396) );
  INVX1 U357 ( .A(n396), .Y(n588) );
  AND2X2 U358 ( .A(a[9]), .B(ready), .Y(n386) );
  INVX1 U359 ( .A(n386), .Y(n589) );
  AND2X2 U360 ( .A(a[7]), .B(ready), .Y(n388) );
  INVX1 U361 ( .A(n388), .Y(n590) );
  AND2X2 U362 ( .A(a[6]), .B(ready), .Y(n389) );
  INVX1 U363 ( .A(n389), .Y(n591) );
  AND2X2 U364 ( .A(a[5]), .B(ready), .Y(n390) );
  INVX1 U365 ( .A(n390), .Y(n592) );
  AND2X2 U366 ( .A(a[3]), .B(ready), .Y(n392) );
  INVX1 U367 ( .A(n392), .Y(n593) );
  AND2X2 U368 ( .A(a[2]), .B(ready), .Y(n393) );
  INVX1 U369 ( .A(n393), .Y(n594) );
  AND2X2 U370 ( .A(a[1]), .B(ready), .Y(n394) );
  INVX1 U371 ( .A(n394), .Y(n595) );
  AND2X2 U372 ( .A(a[0]), .B(ready), .Y(n398) );
  INVX1 U373 ( .A(n398), .Y(n596) );
  AND2X2 U374 ( .A(plogic_ts), .B(ready), .Y(n369) );
  INVX1 U375 ( .A(n369), .Y(n597) );
  INVX1 U376 ( .A(n600), .Y(n598) );
  INVX1 U377 ( .A(n598), .Y(n599) );
  AND2X1 U378 ( .A(n696), .B(n695), .Y(n68) );
  INVX1 U379 ( .A(n68), .Y(n600) );
  INVX1 U380 ( .A(n603), .Y(n601) );
  INVX1 U381 ( .A(n601), .Y(n602) );
  OR2X1 U382 ( .A(reset), .B(ck_i), .Y(n183) );
  INVX1 U383 ( .A(n183), .Y(n603) );
  OR2X2 U384 ( .A(n70), .B(n139), .Y(n379) );
  INVX1 U385 ( .A(n606), .Y(n604) );
  INVX1 U386 ( .A(n604), .Y(n605) );
  AND2X1 U387 ( .A(n687), .B(n686), .Y(n694) );
  INVX1 U388 ( .A(n694), .Y(n606) );
  INVX1 U389 ( .A(n609), .Y(n607) );
  INVX1 U390 ( .A(n607), .Y(n608) );
  AND2X1 U391 ( .A(RETURN_data_out[0]), .B(n373), .Y(n658) );
  INVX1 U392 ( .A(n658), .Y(n609) );
  INVX1 U393 ( .A(n612), .Y(n610) );
  INVX1 U394 ( .A(n610), .Y(n611) );
  BUFX2 U395 ( .A(n560), .Y(n612) );
  INVX1 U396 ( .A(n615), .Y(n613) );
  INVX1 U397 ( .A(n613), .Y(n614) );
  AND2X1 U398 ( .A(n681), .B(n680), .Y(n682) );
  INVX1 U399 ( .A(n682), .Y(n615) );
  INVX1 U400 ( .A(n618), .Y(n616) );
  INVX1 U401 ( .A(n616), .Y(n617) );
  AND2X1 U402 ( .A(n691), .B(n690), .Y(n693) );
  INVX1 U403 ( .A(n693), .Y(n618) );
  INVX1 U404 ( .A(n621), .Y(n619) );
  INVX1 U405 ( .A(n619), .Y(n620) );
  BUFX2 U406 ( .A(n675), .Y(n621) );
  INVX1 U407 ( .A(n624), .Y(n622) );
  INVX1 U408 ( .A(n622), .Y(n623) );
  BUFX2 U409 ( .A(n674), .Y(n624) );
  INVX1 U410 ( .A(n578), .Y(n674) );
  INVX1 U411 ( .A(n666), .Y(n626) );
  INVX1 U412 ( .A(n583), .Y(n627) );
  INVX1 U413 ( .A(n582), .Y(n628) );
  INVX1 U414 ( .A(n579), .Y(n629) );
  INVX1 U415 ( .A(n633), .Y(n631) );
  INVX1 U416 ( .A(n631), .Y(n632) );
  BUFX2 U417 ( .A(n673), .Y(n633) );
  INVX1 U418 ( .A(n580), .Y(n673) );
  INVX1 U419 ( .A(n670), .Y(n635) );
  INVX1 U420 ( .A(n585), .Y(n636) );
  INVX1 U421 ( .A(n584), .Y(n637) );
  INVX1 U422 ( .A(n581), .Y(n638) );
  INVX1 U423 ( .A(n561), .Y(n372) );
  INVX1 U424 ( .A(RETURN_put_reg), .Y(n35) );
  INVX1 U425 ( .A(n562), .Y(n375) );
  INVX1 U426 ( .A(n570), .Y(n644) );
  INVX1 U427 ( .A(n373), .Y(n645) );
  INVX1 U428 ( .A(n376), .Y(n646) );
  INVX1 U429 ( .A(n563), .Y(n647) );
  INVX1 U430 ( .A(n352), .Y(n353) );
  INVX1 U431 ( .A(n651), .Y(n649) );
  INVX1 U432 ( .A(n649), .Y(n650) );
  AND2X1 U433 ( .A(n373), .B(n368), .Y(n187) );
  INVX1 U434 ( .A(n187), .Y(n651) );
  INVX8 U435 ( .A(i[18]), .Y(n652) );
  INVX8 U436 ( .A(n375), .Y(n374) );
  AND2X2 U437 ( .A(n36), .B(n374), .Y(n232) );
  MUX2X1 U438 ( .B(n608), .A(n657), .S(n655), .Y(n656) );
  INVX8 U439 ( .A(dout[0]), .Y(n657) );
  OR2X2 U440 ( .A(n558), .B(n676), .Y(n69) );
  NOR3X1 U441 ( .A(i[23]), .B(i[25]), .C(i[24]), .Y(n665) );
  OR2X1 U442 ( .A(i[29]), .B(i[28]), .Y(n659) );
  NOR3X1 U443 ( .A(n659), .B(i[27]), .C(i[26]), .Y(n664) );
  NOR3X1 U444 ( .A(i[30]), .B(i[5]), .C(i[4]), .Y(n662) );
  OR2X1 U445 ( .A(i[9]), .B(i[8]), .Y(n660) );
  NOR3X1 U446 ( .A(n660), .B(i[7]), .C(i[6]), .Y(n661) );
  AND2X1 U447 ( .A(n662), .B(n661), .Y(n663) );
  NAND3X1 U448 ( .A(n665), .B(n664), .C(n663), .Y(n675) );
  NOR3X1 U449 ( .A(i[16]), .B(i[18]), .C(i[17]), .Y(n666) );
  OR2X1 U450 ( .A(i[15]), .B(i[14]), .Y(n669) );
  NOR3X1 U451 ( .A(n669), .B(i[13]), .C(i[12]), .Y(n670) );
  NOR3X1 U452 ( .A(n620), .B(n623), .C(n632), .Y(n676) );
  NOR3X1 U453 ( .A(i[24]), .B(i[26]), .C(i[25]), .Y(n677) );
  NAND3X1 U454 ( .A(n573), .B(n611), .C(n677), .Y(n683) );
  NOR3X1 U455 ( .A(i[18]), .B(i[20]), .C(i[19]), .Y(n681) );
  NOR3X1 U456 ( .A(i[21]), .B(i[23]), .C(i[22]), .Y(n680) );
  INVX1 U457 ( .A(i[31]), .Y(n692) );
  OAI21X1 U458 ( .A(n576), .B(n614), .C(n692), .Y(n696) );
  OR2X1 U459 ( .A(i[5]), .B(i[4]), .Y(n684) );
  NOR3X1 U460 ( .A(n684), .B(i[3]), .C(i[2]), .Y(n687) );
  OR2X1 U461 ( .A(i[9]), .B(i[8]), .Y(n685) );
  NOR3X1 U462 ( .A(n685), .B(i[7]), .C(i[6]), .Y(n686) );
  OR2X1 U463 ( .A(i[13]), .B(i[12]), .Y(n688) );
  NOR3X1 U464 ( .A(n688), .B(i[11]), .C(i[10]), .Y(n691) );
  OR2X1 U465 ( .A(i[17]), .B(i[16]), .Y(n689) );
  NOR3X1 U466 ( .A(n689), .B(i[15]), .C(i[14]), .Y(n690) );
  OAI21X1 U467 ( .A(n605), .B(n617), .C(n692), .Y(n695) );
endmodule

