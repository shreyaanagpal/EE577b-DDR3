
module FIFO_DEPTH_P25_WIDTH16 ( clk, reset, data_in, put, get, data_out, 
        empty_bar, full_bar, fillcount );
  input [15:0] data_in;
  output [15:0] data_out;
  output [5:0] fillcount;
  input clk, reset, put, get;
  output empty_bar, full_bar;
  wire   n12, n13, n14, n15, n16, n2314, n2315, n20, n21, n22, n23, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n73, n74, n75, n76, n281, n283, n285, n287, n289, n291, n293, n295,
         n297, n299, n301, n303, n305, n307, n309, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n17, n18, n19, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n72, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n282, n284, n286, n288, n290, n292, n294, n296, n298, n300, n302,
         n304, n306, n308, n310, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313;
  wire   [4:0] wr_ptr;
  wire   [511:0] mem;
  wire   [4:2] add_57_carry;
  wire   [4:2] add_51_carry;
  wire   [5:1] sub_93_carry;

  DFFPOSX1 wr_ptr_reg_0_ ( .D(n1413), .CLK(clk), .Q(wr_ptr[0]) );
  DFFPOSX1 rd_ptr_reg_4_ ( .D(n1412), .CLK(clk), .Q(n16) );
  DFFPOSX1 rd_ptr_reg_0_ ( .D(n1411), .CLK(clk), .Q(n12) );
  DFFPOSX1 rd_ptr_reg_1_ ( .D(n1410), .CLK(clk), .Q(n13) );
  DFFPOSX1 rd_ptr_reg_2_ ( .D(n1409), .CLK(clk), .Q(n14) );
  DFFPOSX1 rd_ptr_reg_3_ ( .D(n1408), .CLK(clk), .Q(n15) );
  DFFPOSX1 wr_ptr_reg_4_ ( .D(n1407), .CLK(clk), .Q(wr_ptr[4]) );
  DFFPOSX1 wr_ptr_reg_1_ ( .D(n1406), .CLK(clk), .Q(wr_ptr[1]) );
  DFFPOSX1 wr_ptr_reg_2_ ( .D(n1405), .CLK(clk), .Q(wr_ptr[2]) );
  DFFPOSX1 wr_ptr_reg_3_ ( .D(n1404), .CLK(clk), .Q(wr_ptr[3]) );
  DFFPOSX1 data_out_reg_15_ ( .D(n2308), .CLK(clk), .Q(data_out[15]) );
  DFFPOSX1 data_out_reg_14_ ( .D(n2307), .CLK(clk), .Q(data_out[14]) );
  DFFPOSX1 data_out_reg_13_ ( .D(n2306), .CLK(clk), .Q(data_out[13]) );
  DFFPOSX1 data_out_reg_12_ ( .D(n2305), .CLK(clk), .Q(data_out[12]) );
  DFFPOSX1 data_out_reg_11_ ( .D(n2304), .CLK(clk), .Q(data_out[11]) );
  DFFPOSX1 data_out_reg_10_ ( .D(n2303), .CLK(clk), .Q(data_out[10]) );
  DFFPOSX1 data_out_reg_9_ ( .D(n2302), .CLK(clk), .Q(data_out[9]) );
  DFFPOSX1 data_out_reg_8_ ( .D(n2301), .CLK(clk), .Q(data_out[8]) );
  DFFPOSX1 data_out_reg_7_ ( .D(n2300), .CLK(clk), .Q(data_out[7]) );
  DFFPOSX1 data_out_reg_6_ ( .D(n2299), .CLK(clk), .Q(data_out[6]) );
  DFFPOSX1 data_out_reg_5_ ( .D(n2298), .CLK(clk), .Q(data_out[5]) );
  DFFPOSX1 data_out_reg_4_ ( .D(n2297), .CLK(clk), .Q(data_out[4]) );
  DFFPOSX1 data_out_reg_3_ ( .D(n2296), .CLK(clk), .Q(data_out[3]) );
  DFFPOSX1 data_out_reg_2_ ( .D(n2295), .CLK(clk), .Q(data_out[2]) );
  DFFPOSX1 data_out_reg_1_ ( .D(n2294), .CLK(clk), .Q(data_out[1]) );
  DFFPOSX1 data_out_reg_0_ ( .D(n2293), .CLK(clk), .Q(data_out[0]) );
  DFFPOSX1 mem_reg_31__15_ ( .D(n1403), .CLK(clk), .Q(mem[511]) );
  DFFPOSX1 mem_reg_31__14_ ( .D(n1402), .CLK(clk), .Q(mem[510]) );
  DFFPOSX1 mem_reg_31__13_ ( .D(n1401), .CLK(clk), .Q(mem[509]) );
  DFFPOSX1 mem_reg_31__12_ ( .D(n1400), .CLK(clk), .Q(mem[508]) );
  DFFPOSX1 mem_reg_31__11_ ( .D(n1399), .CLK(clk), .Q(mem[507]) );
  DFFPOSX1 mem_reg_31__10_ ( .D(n1398), .CLK(clk), .Q(mem[506]) );
  DFFPOSX1 mem_reg_31__9_ ( .D(n1397), .CLK(clk), .Q(mem[505]) );
  DFFPOSX1 mem_reg_31__8_ ( .D(n1396), .CLK(clk), .Q(mem[504]) );
  DFFPOSX1 mem_reg_31__7_ ( .D(n1395), .CLK(clk), .Q(mem[503]) );
  DFFPOSX1 mem_reg_31__6_ ( .D(n1394), .CLK(clk), .Q(mem[502]) );
  DFFPOSX1 mem_reg_31__5_ ( .D(n1393), .CLK(clk), .Q(mem[501]) );
  DFFPOSX1 mem_reg_31__4_ ( .D(n1392), .CLK(clk), .Q(mem[500]) );
  DFFPOSX1 mem_reg_31__3_ ( .D(n1391), .CLK(clk), .Q(mem[499]) );
  DFFPOSX1 mem_reg_31__2_ ( .D(n1390), .CLK(clk), .Q(mem[498]) );
  DFFPOSX1 mem_reg_31__1_ ( .D(n1389), .CLK(clk), .Q(mem[497]) );
  DFFPOSX1 mem_reg_31__0_ ( .D(n1388), .CLK(clk), .Q(mem[496]) );
  DFFPOSX1 mem_reg_30__15_ ( .D(n1387), .CLK(clk), .Q(mem[495]) );
  DFFPOSX1 mem_reg_30__14_ ( .D(n1386), .CLK(clk), .Q(mem[494]) );
  DFFPOSX1 mem_reg_30__13_ ( .D(n1385), .CLK(clk), .Q(mem[493]) );
  DFFPOSX1 mem_reg_30__12_ ( .D(n1384), .CLK(clk), .Q(mem[492]) );
  DFFPOSX1 mem_reg_30__11_ ( .D(n1383), .CLK(clk), .Q(mem[491]) );
  DFFPOSX1 mem_reg_30__10_ ( .D(n1382), .CLK(clk), .Q(mem[490]) );
  DFFPOSX1 mem_reg_30__9_ ( .D(n1381), .CLK(clk), .Q(mem[489]) );
  DFFPOSX1 mem_reg_30__8_ ( .D(n1380), .CLK(clk), .Q(mem[488]) );
  DFFPOSX1 mem_reg_30__7_ ( .D(n1379), .CLK(clk), .Q(mem[487]) );
  DFFPOSX1 mem_reg_30__6_ ( .D(n1378), .CLK(clk), .Q(mem[486]) );
  DFFPOSX1 mem_reg_30__5_ ( .D(n1377), .CLK(clk), .Q(mem[485]) );
  DFFPOSX1 mem_reg_30__4_ ( .D(n1376), .CLK(clk), .Q(mem[484]) );
  DFFPOSX1 mem_reg_30__3_ ( .D(n1375), .CLK(clk), .Q(mem[483]) );
  DFFPOSX1 mem_reg_30__2_ ( .D(n1374), .CLK(clk), .Q(mem[482]) );
  DFFPOSX1 mem_reg_30__1_ ( .D(n1373), .CLK(clk), .Q(mem[481]) );
  DFFPOSX1 mem_reg_30__0_ ( .D(n1372), .CLK(clk), .Q(mem[480]) );
  DFFPOSX1 mem_reg_29__15_ ( .D(n1371), .CLK(clk), .Q(mem[479]) );
  DFFPOSX1 mem_reg_29__14_ ( .D(n1370), .CLK(clk), .Q(mem[478]) );
  DFFPOSX1 mem_reg_29__13_ ( .D(n1369), .CLK(clk), .Q(mem[477]) );
  DFFPOSX1 mem_reg_29__12_ ( .D(n1368), .CLK(clk), .Q(mem[476]) );
  DFFPOSX1 mem_reg_29__11_ ( .D(n1367), .CLK(clk), .Q(mem[475]) );
  DFFPOSX1 mem_reg_29__10_ ( .D(n1366), .CLK(clk), .Q(mem[474]) );
  DFFPOSX1 mem_reg_29__9_ ( .D(n1365), .CLK(clk), .Q(mem[473]) );
  DFFPOSX1 mem_reg_29__8_ ( .D(n1364), .CLK(clk), .Q(mem[472]) );
  DFFPOSX1 mem_reg_29__7_ ( .D(n1363), .CLK(clk), .Q(mem[471]) );
  DFFPOSX1 mem_reg_29__6_ ( .D(n1362), .CLK(clk), .Q(mem[470]) );
  DFFPOSX1 mem_reg_29__5_ ( .D(n1361), .CLK(clk), .Q(mem[469]) );
  DFFPOSX1 mem_reg_29__4_ ( .D(n1360), .CLK(clk), .Q(mem[468]) );
  DFFPOSX1 mem_reg_29__3_ ( .D(n1359), .CLK(clk), .Q(mem[467]) );
  DFFPOSX1 mem_reg_29__2_ ( .D(n1358), .CLK(clk), .Q(mem[466]) );
  DFFPOSX1 mem_reg_29__1_ ( .D(n1357), .CLK(clk), .Q(mem[465]) );
  DFFPOSX1 mem_reg_29__0_ ( .D(n1356), .CLK(clk), .Q(mem[464]) );
  DFFPOSX1 mem_reg_28__15_ ( .D(n1355), .CLK(clk), .Q(mem[463]) );
  DFFPOSX1 mem_reg_28__14_ ( .D(n1354), .CLK(clk), .Q(mem[462]) );
  DFFPOSX1 mem_reg_28__13_ ( .D(n1353), .CLK(clk), .Q(mem[461]) );
  DFFPOSX1 mem_reg_28__12_ ( .D(n1352), .CLK(clk), .Q(mem[460]) );
  DFFPOSX1 mem_reg_28__11_ ( .D(n1351), .CLK(clk), .Q(mem[459]) );
  DFFPOSX1 mem_reg_28__10_ ( .D(n1350), .CLK(clk), .Q(mem[458]) );
  DFFPOSX1 mem_reg_28__9_ ( .D(n1349), .CLK(clk), .Q(mem[457]) );
  DFFPOSX1 mem_reg_28__8_ ( .D(n1348), .CLK(clk), .Q(mem[456]) );
  DFFPOSX1 mem_reg_28__7_ ( .D(n1347), .CLK(clk), .Q(mem[455]) );
  DFFPOSX1 mem_reg_28__6_ ( .D(n1346), .CLK(clk), .Q(mem[454]) );
  DFFPOSX1 mem_reg_28__5_ ( .D(n1345), .CLK(clk), .Q(mem[453]) );
  DFFPOSX1 mem_reg_28__4_ ( .D(n1344), .CLK(clk), .Q(mem[452]) );
  DFFPOSX1 mem_reg_28__3_ ( .D(n1343), .CLK(clk), .Q(mem[451]) );
  DFFPOSX1 mem_reg_28__2_ ( .D(n1342), .CLK(clk), .Q(mem[450]) );
  DFFPOSX1 mem_reg_28__1_ ( .D(n1341), .CLK(clk), .Q(mem[449]) );
  DFFPOSX1 mem_reg_28__0_ ( .D(n1340), .CLK(clk), .Q(mem[448]) );
  DFFPOSX1 mem_reg_27__15_ ( .D(n1339), .CLK(clk), .Q(mem[447]) );
  DFFPOSX1 mem_reg_27__14_ ( .D(n1338), .CLK(clk), .Q(mem[446]) );
  DFFPOSX1 mem_reg_27__13_ ( .D(n1337), .CLK(clk), .Q(mem[445]) );
  DFFPOSX1 mem_reg_27__12_ ( .D(n1336), .CLK(clk), .Q(mem[444]) );
  DFFPOSX1 mem_reg_27__11_ ( .D(n1335), .CLK(clk), .Q(mem[443]) );
  DFFPOSX1 mem_reg_27__10_ ( .D(n1334), .CLK(clk), .Q(mem[442]) );
  DFFPOSX1 mem_reg_27__9_ ( .D(n1333), .CLK(clk), .Q(mem[441]) );
  DFFPOSX1 mem_reg_27__8_ ( .D(n1332), .CLK(clk), .Q(mem[440]) );
  DFFPOSX1 mem_reg_27__7_ ( .D(n1331), .CLK(clk), .Q(mem[439]) );
  DFFPOSX1 mem_reg_27__6_ ( .D(n1330), .CLK(clk), .Q(mem[438]) );
  DFFPOSX1 mem_reg_27__5_ ( .D(n1329), .CLK(clk), .Q(mem[437]) );
  DFFPOSX1 mem_reg_27__4_ ( .D(n1328), .CLK(clk), .Q(mem[436]) );
  DFFPOSX1 mem_reg_27__3_ ( .D(n1327), .CLK(clk), .Q(mem[435]) );
  DFFPOSX1 mem_reg_27__2_ ( .D(n1326), .CLK(clk), .Q(mem[434]) );
  DFFPOSX1 mem_reg_27__1_ ( .D(n1325), .CLK(clk), .Q(mem[433]) );
  DFFPOSX1 mem_reg_27__0_ ( .D(n1324), .CLK(clk), .Q(mem[432]) );
  DFFPOSX1 mem_reg_26__15_ ( .D(n1323), .CLK(clk), .Q(mem[431]) );
  DFFPOSX1 mem_reg_26__14_ ( .D(n1322), .CLK(clk), .Q(mem[430]) );
  DFFPOSX1 mem_reg_26__13_ ( .D(n1321), .CLK(clk), .Q(mem[429]) );
  DFFPOSX1 mem_reg_26__12_ ( .D(n1320), .CLK(clk), .Q(mem[428]) );
  DFFPOSX1 mem_reg_26__11_ ( .D(n1319), .CLK(clk), .Q(mem[427]) );
  DFFPOSX1 mem_reg_26__10_ ( .D(n1318), .CLK(clk), .Q(mem[426]) );
  DFFPOSX1 mem_reg_26__9_ ( .D(n1317), .CLK(clk), .Q(mem[425]) );
  DFFPOSX1 mem_reg_26__8_ ( .D(n1316), .CLK(clk), .Q(mem[424]) );
  DFFPOSX1 mem_reg_26__7_ ( .D(n1315), .CLK(clk), .Q(mem[423]) );
  DFFPOSX1 mem_reg_26__6_ ( .D(n1314), .CLK(clk), .Q(mem[422]) );
  DFFPOSX1 mem_reg_26__5_ ( .D(n1313), .CLK(clk), .Q(mem[421]) );
  DFFPOSX1 mem_reg_26__4_ ( .D(n1312), .CLK(clk), .Q(mem[420]) );
  DFFPOSX1 mem_reg_26__3_ ( .D(n1311), .CLK(clk), .Q(mem[419]) );
  DFFPOSX1 mem_reg_26__2_ ( .D(n1310), .CLK(clk), .Q(mem[418]) );
  DFFPOSX1 mem_reg_26__1_ ( .D(n1309), .CLK(clk), .Q(mem[417]) );
  DFFPOSX1 mem_reg_26__0_ ( .D(n1308), .CLK(clk), .Q(mem[416]) );
  DFFPOSX1 mem_reg_25__15_ ( .D(n1307), .CLK(clk), .Q(mem[415]) );
  DFFPOSX1 mem_reg_25__14_ ( .D(n1306), .CLK(clk), .Q(mem[414]) );
  DFFPOSX1 mem_reg_25__13_ ( .D(n1305), .CLK(clk), .Q(mem[413]) );
  DFFPOSX1 mem_reg_25__12_ ( .D(n1304), .CLK(clk), .Q(mem[412]) );
  DFFPOSX1 mem_reg_25__11_ ( .D(n1303), .CLK(clk), .Q(mem[411]) );
  DFFPOSX1 mem_reg_25__10_ ( .D(n1302), .CLK(clk), .Q(mem[410]) );
  DFFPOSX1 mem_reg_25__9_ ( .D(n1301), .CLK(clk), .Q(mem[409]) );
  DFFPOSX1 mem_reg_25__8_ ( .D(n1300), .CLK(clk), .Q(mem[408]) );
  DFFPOSX1 mem_reg_25__7_ ( .D(n1299), .CLK(clk), .Q(mem[407]) );
  DFFPOSX1 mem_reg_25__6_ ( .D(n1298), .CLK(clk), .Q(mem[406]) );
  DFFPOSX1 mem_reg_25__5_ ( .D(n1297), .CLK(clk), .Q(mem[405]) );
  DFFPOSX1 mem_reg_25__4_ ( .D(n1296), .CLK(clk), .Q(mem[404]) );
  DFFPOSX1 mem_reg_25__3_ ( .D(n1295), .CLK(clk), .Q(mem[403]) );
  DFFPOSX1 mem_reg_25__2_ ( .D(n1294), .CLK(clk), .Q(mem[402]) );
  DFFPOSX1 mem_reg_25__1_ ( .D(n1293), .CLK(clk), .Q(mem[401]) );
  DFFPOSX1 mem_reg_25__0_ ( .D(n1292), .CLK(clk), .Q(mem[400]) );
  DFFPOSX1 mem_reg_24__15_ ( .D(n1291), .CLK(clk), .Q(mem[399]) );
  DFFPOSX1 mem_reg_24__14_ ( .D(n1290), .CLK(clk), .Q(mem[398]) );
  DFFPOSX1 mem_reg_24__13_ ( .D(n1289), .CLK(clk), .Q(mem[397]) );
  DFFPOSX1 mem_reg_24__12_ ( .D(n1288), .CLK(clk), .Q(mem[396]) );
  DFFPOSX1 mem_reg_24__11_ ( .D(n1287), .CLK(clk), .Q(mem[395]) );
  DFFPOSX1 mem_reg_24__10_ ( .D(n1286), .CLK(clk), .Q(mem[394]) );
  DFFPOSX1 mem_reg_24__9_ ( .D(n1285), .CLK(clk), .Q(mem[393]) );
  DFFPOSX1 mem_reg_24__8_ ( .D(n1284), .CLK(clk), .Q(mem[392]) );
  DFFPOSX1 mem_reg_24__7_ ( .D(n1283), .CLK(clk), .Q(mem[391]) );
  DFFPOSX1 mem_reg_24__6_ ( .D(n1282), .CLK(clk), .Q(mem[390]) );
  DFFPOSX1 mem_reg_24__5_ ( .D(n1281), .CLK(clk), .Q(mem[389]) );
  DFFPOSX1 mem_reg_24__4_ ( .D(n1280), .CLK(clk), .Q(mem[388]) );
  DFFPOSX1 mem_reg_24__3_ ( .D(n1279), .CLK(clk), .Q(mem[387]) );
  DFFPOSX1 mem_reg_24__2_ ( .D(n1278), .CLK(clk), .Q(mem[386]) );
  DFFPOSX1 mem_reg_24__1_ ( .D(n1277), .CLK(clk), .Q(mem[385]) );
  DFFPOSX1 mem_reg_24__0_ ( .D(n1276), .CLK(clk), .Q(mem[384]) );
  DFFPOSX1 mem_reg_23__15_ ( .D(n1275), .CLK(clk), .Q(mem[383]) );
  DFFPOSX1 mem_reg_23__14_ ( .D(n1274), .CLK(clk), .Q(mem[382]) );
  DFFPOSX1 mem_reg_23__13_ ( .D(n1273), .CLK(clk), .Q(mem[381]) );
  DFFPOSX1 mem_reg_23__12_ ( .D(n1272), .CLK(clk), .Q(mem[380]) );
  DFFPOSX1 mem_reg_23__11_ ( .D(n1271), .CLK(clk), .Q(mem[379]) );
  DFFPOSX1 mem_reg_23__10_ ( .D(n1270), .CLK(clk), .Q(mem[378]) );
  DFFPOSX1 mem_reg_23__9_ ( .D(n1269), .CLK(clk), .Q(mem[377]) );
  DFFPOSX1 mem_reg_23__8_ ( .D(n1268), .CLK(clk), .Q(mem[376]) );
  DFFPOSX1 mem_reg_23__7_ ( .D(n1267), .CLK(clk), .Q(mem[375]) );
  DFFPOSX1 mem_reg_23__6_ ( .D(n1266), .CLK(clk), .Q(mem[374]) );
  DFFPOSX1 mem_reg_23__5_ ( .D(n1265), .CLK(clk), .Q(mem[373]) );
  DFFPOSX1 mem_reg_23__4_ ( .D(n1264), .CLK(clk), .Q(mem[372]) );
  DFFPOSX1 mem_reg_23__3_ ( .D(n1263), .CLK(clk), .Q(mem[371]) );
  DFFPOSX1 mem_reg_23__2_ ( .D(n1262), .CLK(clk), .Q(mem[370]) );
  DFFPOSX1 mem_reg_23__1_ ( .D(n1261), .CLK(clk), .Q(mem[369]) );
  DFFPOSX1 mem_reg_23__0_ ( .D(n1260), .CLK(clk), .Q(mem[368]) );
  DFFPOSX1 mem_reg_22__15_ ( .D(n1259), .CLK(clk), .Q(mem[367]) );
  DFFPOSX1 mem_reg_22__14_ ( .D(n1258), .CLK(clk), .Q(mem[366]) );
  DFFPOSX1 mem_reg_22__13_ ( .D(n1257), .CLK(clk), .Q(mem[365]) );
  DFFPOSX1 mem_reg_22__12_ ( .D(n1256), .CLK(clk), .Q(mem[364]) );
  DFFPOSX1 mem_reg_22__11_ ( .D(n1255), .CLK(clk), .Q(mem[363]) );
  DFFPOSX1 mem_reg_22__10_ ( .D(n1254), .CLK(clk), .Q(mem[362]) );
  DFFPOSX1 mem_reg_22__9_ ( .D(n1253), .CLK(clk), .Q(mem[361]) );
  DFFPOSX1 mem_reg_22__8_ ( .D(n1252), .CLK(clk), .Q(mem[360]) );
  DFFPOSX1 mem_reg_22__7_ ( .D(n1251), .CLK(clk), .Q(mem[359]) );
  DFFPOSX1 mem_reg_22__6_ ( .D(n1250), .CLK(clk), .Q(mem[358]) );
  DFFPOSX1 mem_reg_22__5_ ( .D(n1249), .CLK(clk), .Q(mem[357]) );
  DFFPOSX1 mem_reg_22__4_ ( .D(n1248), .CLK(clk), .Q(mem[356]) );
  DFFPOSX1 mem_reg_22__3_ ( .D(n1247), .CLK(clk), .Q(mem[355]) );
  DFFPOSX1 mem_reg_22__2_ ( .D(n1246), .CLK(clk), .Q(mem[354]) );
  DFFPOSX1 mem_reg_22__1_ ( .D(n1245), .CLK(clk), .Q(mem[353]) );
  DFFPOSX1 mem_reg_22__0_ ( .D(n1244), .CLK(clk), .Q(mem[352]) );
  DFFPOSX1 mem_reg_21__15_ ( .D(n1243), .CLK(clk), .Q(mem[351]) );
  DFFPOSX1 mem_reg_21__14_ ( .D(n1242), .CLK(clk), .Q(mem[350]) );
  DFFPOSX1 mem_reg_21__13_ ( .D(n1241), .CLK(clk), .Q(mem[349]) );
  DFFPOSX1 mem_reg_21__12_ ( .D(n1240), .CLK(clk), .Q(mem[348]) );
  DFFPOSX1 mem_reg_21__11_ ( .D(n1239), .CLK(clk), .Q(mem[347]) );
  DFFPOSX1 mem_reg_21__10_ ( .D(n1238), .CLK(clk), .Q(mem[346]) );
  DFFPOSX1 mem_reg_21__9_ ( .D(n1237), .CLK(clk), .Q(mem[345]) );
  DFFPOSX1 mem_reg_21__8_ ( .D(n1236), .CLK(clk), .Q(mem[344]) );
  DFFPOSX1 mem_reg_21__7_ ( .D(n1235), .CLK(clk), .Q(mem[343]) );
  DFFPOSX1 mem_reg_21__6_ ( .D(n1234), .CLK(clk), .Q(mem[342]) );
  DFFPOSX1 mem_reg_21__5_ ( .D(n1233), .CLK(clk), .Q(mem[341]) );
  DFFPOSX1 mem_reg_21__4_ ( .D(n1232), .CLK(clk), .Q(mem[340]) );
  DFFPOSX1 mem_reg_21__3_ ( .D(n1231), .CLK(clk), .Q(mem[339]) );
  DFFPOSX1 mem_reg_21__2_ ( .D(n1230), .CLK(clk), .Q(mem[338]) );
  DFFPOSX1 mem_reg_21__1_ ( .D(n1229), .CLK(clk), .Q(mem[337]) );
  DFFPOSX1 mem_reg_21__0_ ( .D(n1228), .CLK(clk), .Q(mem[336]) );
  DFFPOSX1 mem_reg_20__15_ ( .D(n1227), .CLK(clk), .Q(mem[335]) );
  DFFPOSX1 mem_reg_20__14_ ( .D(n1226), .CLK(clk), .Q(mem[334]) );
  DFFPOSX1 mem_reg_20__13_ ( .D(n1225), .CLK(clk), .Q(mem[333]) );
  DFFPOSX1 mem_reg_20__12_ ( .D(n1224), .CLK(clk), .Q(mem[332]) );
  DFFPOSX1 mem_reg_20__11_ ( .D(n1223), .CLK(clk), .Q(mem[331]) );
  DFFPOSX1 mem_reg_20__10_ ( .D(n1222), .CLK(clk), .Q(mem[330]) );
  DFFPOSX1 mem_reg_20__9_ ( .D(n1221), .CLK(clk), .Q(mem[329]) );
  DFFPOSX1 mem_reg_20__8_ ( .D(n1220), .CLK(clk), .Q(mem[328]) );
  DFFPOSX1 mem_reg_20__7_ ( .D(n1219), .CLK(clk), .Q(mem[327]) );
  DFFPOSX1 mem_reg_20__6_ ( .D(n1218), .CLK(clk), .Q(mem[326]) );
  DFFPOSX1 mem_reg_20__5_ ( .D(n1217), .CLK(clk), .Q(mem[325]) );
  DFFPOSX1 mem_reg_20__4_ ( .D(n1216), .CLK(clk), .Q(mem[324]) );
  DFFPOSX1 mem_reg_20__3_ ( .D(n1215), .CLK(clk), .Q(mem[323]) );
  DFFPOSX1 mem_reg_20__2_ ( .D(n1214), .CLK(clk), .Q(mem[322]) );
  DFFPOSX1 mem_reg_20__1_ ( .D(n1213), .CLK(clk), .Q(mem[321]) );
  DFFPOSX1 mem_reg_20__0_ ( .D(n1212), .CLK(clk), .Q(mem[320]) );
  DFFPOSX1 mem_reg_19__15_ ( .D(n1211), .CLK(clk), .Q(mem[319]) );
  DFFPOSX1 mem_reg_19__14_ ( .D(n1210), .CLK(clk), .Q(mem[318]) );
  DFFPOSX1 mem_reg_19__13_ ( .D(n1209), .CLK(clk), .Q(mem[317]) );
  DFFPOSX1 mem_reg_19__12_ ( .D(n1208), .CLK(clk), .Q(mem[316]) );
  DFFPOSX1 mem_reg_19__11_ ( .D(n1207), .CLK(clk), .Q(mem[315]) );
  DFFPOSX1 mem_reg_19__10_ ( .D(n1206), .CLK(clk), .Q(mem[314]) );
  DFFPOSX1 mem_reg_19__9_ ( .D(n1205), .CLK(clk), .Q(mem[313]) );
  DFFPOSX1 mem_reg_19__8_ ( .D(n1204), .CLK(clk), .Q(mem[312]) );
  DFFPOSX1 mem_reg_19__7_ ( .D(n1203), .CLK(clk), .Q(mem[311]) );
  DFFPOSX1 mem_reg_19__6_ ( .D(n1202), .CLK(clk), .Q(mem[310]) );
  DFFPOSX1 mem_reg_19__5_ ( .D(n1201), .CLK(clk), .Q(mem[309]) );
  DFFPOSX1 mem_reg_19__4_ ( .D(n1200), .CLK(clk), .Q(mem[308]) );
  DFFPOSX1 mem_reg_19__3_ ( .D(n1199), .CLK(clk), .Q(mem[307]) );
  DFFPOSX1 mem_reg_19__2_ ( .D(n1198), .CLK(clk), .Q(mem[306]) );
  DFFPOSX1 mem_reg_19__1_ ( .D(n1197), .CLK(clk), .Q(mem[305]) );
  DFFPOSX1 mem_reg_19__0_ ( .D(n1196), .CLK(clk), .Q(mem[304]) );
  DFFPOSX1 mem_reg_18__15_ ( .D(n1195), .CLK(clk), .Q(mem[303]) );
  DFFPOSX1 mem_reg_18__14_ ( .D(n1194), .CLK(clk), .Q(mem[302]) );
  DFFPOSX1 mem_reg_18__13_ ( .D(n1193), .CLK(clk), .Q(mem[301]) );
  DFFPOSX1 mem_reg_18__12_ ( .D(n1192), .CLK(clk), .Q(mem[300]) );
  DFFPOSX1 mem_reg_18__11_ ( .D(n1191), .CLK(clk), .Q(mem[299]) );
  DFFPOSX1 mem_reg_18__10_ ( .D(n1190), .CLK(clk), .Q(mem[298]) );
  DFFPOSX1 mem_reg_18__9_ ( .D(n1189), .CLK(clk), .Q(mem[297]) );
  DFFPOSX1 mem_reg_18__8_ ( .D(n1188), .CLK(clk), .Q(mem[296]) );
  DFFPOSX1 mem_reg_18__7_ ( .D(n1187), .CLK(clk), .Q(mem[295]) );
  DFFPOSX1 mem_reg_18__6_ ( .D(n1186), .CLK(clk), .Q(mem[294]) );
  DFFPOSX1 mem_reg_18__5_ ( .D(n1185), .CLK(clk), .Q(mem[293]) );
  DFFPOSX1 mem_reg_18__4_ ( .D(n1184), .CLK(clk), .Q(mem[292]) );
  DFFPOSX1 mem_reg_18__3_ ( .D(n1183), .CLK(clk), .Q(mem[291]) );
  DFFPOSX1 mem_reg_18__2_ ( .D(n1182), .CLK(clk), .Q(mem[290]) );
  DFFPOSX1 mem_reg_18__1_ ( .D(n1181), .CLK(clk), .Q(mem[289]) );
  DFFPOSX1 mem_reg_18__0_ ( .D(n1180), .CLK(clk), .Q(mem[288]) );
  DFFPOSX1 mem_reg_17__15_ ( .D(n1179), .CLK(clk), .Q(mem[287]) );
  DFFPOSX1 mem_reg_17__14_ ( .D(n1178), .CLK(clk), .Q(mem[286]) );
  DFFPOSX1 mem_reg_17__13_ ( .D(n1177), .CLK(clk), .Q(mem[285]) );
  DFFPOSX1 mem_reg_17__12_ ( .D(n1176), .CLK(clk), .Q(mem[284]) );
  DFFPOSX1 mem_reg_17__11_ ( .D(n1175), .CLK(clk), .Q(mem[283]) );
  DFFPOSX1 mem_reg_17__10_ ( .D(n1174), .CLK(clk), .Q(mem[282]) );
  DFFPOSX1 mem_reg_17__9_ ( .D(n1173), .CLK(clk), .Q(mem[281]) );
  DFFPOSX1 mem_reg_17__8_ ( .D(n1172), .CLK(clk), .Q(mem[280]) );
  DFFPOSX1 mem_reg_17__7_ ( .D(n1171), .CLK(clk), .Q(mem[279]) );
  DFFPOSX1 mem_reg_17__6_ ( .D(n1170), .CLK(clk), .Q(mem[278]) );
  DFFPOSX1 mem_reg_17__5_ ( .D(n1169), .CLK(clk), .Q(mem[277]) );
  DFFPOSX1 mem_reg_17__4_ ( .D(n1168), .CLK(clk), .Q(mem[276]) );
  DFFPOSX1 mem_reg_17__3_ ( .D(n1167), .CLK(clk), .Q(mem[275]) );
  DFFPOSX1 mem_reg_17__2_ ( .D(n1166), .CLK(clk), .Q(mem[274]) );
  DFFPOSX1 mem_reg_17__1_ ( .D(n1165), .CLK(clk), .Q(mem[273]) );
  DFFPOSX1 mem_reg_17__0_ ( .D(n1164), .CLK(clk), .Q(mem[272]) );
  DFFPOSX1 mem_reg_16__15_ ( .D(n1163), .CLK(clk), .Q(mem[271]) );
  DFFPOSX1 mem_reg_16__14_ ( .D(n1162), .CLK(clk), .Q(mem[270]) );
  DFFPOSX1 mem_reg_16__13_ ( .D(n1161), .CLK(clk), .Q(mem[269]) );
  DFFPOSX1 mem_reg_16__12_ ( .D(n1160), .CLK(clk), .Q(mem[268]) );
  DFFPOSX1 mem_reg_16__11_ ( .D(n1159), .CLK(clk), .Q(mem[267]) );
  DFFPOSX1 mem_reg_16__10_ ( .D(n1158), .CLK(clk), .Q(mem[266]) );
  DFFPOSX1 mem_reg_16__9_ ( .D(n1157), .CLK(clk), .Q(mem[265]) );
  DFFPOSX1 mem_reg_16__8_ ( .D(n1156), .CLK(clk), .Q(mem[264]) );
  DFFPOSX1 mem_reg_16__7_ ( .D(n1155), .CLK(clk), .Q(mem[263]) );
  DFFPOSX1 mem_reg_16__6_ ( .D(n1154), .CLK(clk), .Q(mem[262]) );
  DFFPOSX1 mem_reg_16__5_ ( .D(n1153), .CLK(clk), .Q(mem[261]) );
  DFFPOSX1 mem_reg_16__4_ ( .D(n1152), .CLK(clk), .Q(mem[260]) );
  DFFPOSX1 mem_reg_16__3_ ( .D(n1151), .CLK(clk), .Q(mem[259]) );
  DFFPOSX1 mem_reg_16__2_ ( .D(n1150), .CLK(clk), .Q(mem[258]) );
  DFFPOSX1 mem_reg_16__1_ ( .D(n1149), .CLK(clk), .Q(mem[257]) );
  DFFPOSX1 mem_reg_16__0_ ( .D(n1148), .CLK(clk), .Q(mem[256]) );
  DFFPOSX1 mem_reg_15__15_ ( .D(n1147), .CLK(clk), .Q(mem[255]) );
  DFFPOSX1 mem_reg_15__14_ ( .D(n1146), .CLK(clk), .Q(mem[254]) );
  DFFPOSX1 mem_reg_15__13_ ( .D(n1145), .CLK(clk), .Q(mem[253]) );
  DFFPOSX1 mem_reg_15__12_ ( .D(n1144), .CLK(clk), .Q(mem[252]) );
  DFFPOSX1 mem_reg_15__11_ ( .D(n1143), .CLK(clk), .Q(mem[251]) );
  DFFPOSX1 mem_reg_15__10_ ( .D(n1142), .CLK(clk), .Q(mem[250]) );
  DFFPOSX1 mem_reg_15__9_ ( .D(n1141), .CLK(clk), .Q(mem[249]) );
  DFFPOSX1 mem_reg_15__8_ ( .D(n1140), .CLK(clk), .Q(mem[248]) );
  DFFPOSX1 mem_reg_15__7_ ( .D(n1139), .CLK(clk), .Q(mem[247]) );
  DFFPOSX1 mem_reg_15__6_ ( .D(n1138), .CLK(clk), .Q(mem[246]) );
  DFFPOSX1 mem_reg_15__5_ ( .D(n1137), .CLK(clk), .Q(mem[245]) );
  DFFPOSX1 mem_reg_15__4_ ( .D(n1136), .CLK(clk), .Q(mem[244]) );
  DFFPOSX1 mem_reg_15__3_ ( .D(n1135), .CLK(clk), .Q(mem[243]) );
  DFFPOSX1 mem_reg_15__2_ ( .D(n1134), .CLK(clk), .Q(mem[242]) );
  DFFPOSX1 mem_reg_15__1_ ( .D(n1133), .CLK(clk), .Q(mem[241]) );
  DFFPOSX1 mem_reg_15__0_ ( .D(n1132), .CLK(clk), .Q(mem[240]) );
  DFFPOSX1 mem_reg_14__15_ ( .D(n1131), .CLK(clk), .Q(mem[239]) );
  DFFPOSX1 mem_reg_14__14_ ( .D(n1130), .CLK(clk), .Q(mem[238]) );
  DFFPOSX1 mem_reg_14__13_ ( .D(n1129), .CLK(clk), .Q(mem[237]) );
  DFFPOSX1 mem_reg_14__12_ ( .D(n1128), .CLK(clk), .Q(mem[236]) );
  DFFPOSX1 mem_reg_14__11_ ( .D(n1127), .CLK(clk), .Q(mem[235]) );
  DFFPOSX1 mem_reg_14__10_ ( .D(n1126), .CLK(clk), .Q(mem[234]) );
  DFFPOSX1 mem_reg_14__9_ ( .D(n1125), .CLK(clk), .Q(mem[233]) );
  DFFPOSX1 mem_reg_14__8_ ( .D(n1124), .CLK(clk), .Q(mem[232]) );
  DFFPOSX1 mem_reg_14__7_ ( .D(n1123), .CLK(clk), .Q(mem[231]) );
  DFFPOSX1 mem_reg_14__6_ ( .D(n1122), .CLK(clk), .Q(mem[230]) );
  DFFPOSX1 mem_reg_14__5_ ( .D(n1121), .CLK(clk), .Q(mem[229]) );
  DFFPOSX1 mem_reg_14__4_ ( .D(n1120), .CLK(clk), .Q(mem[228]) );
  DFFPOSX1 mem_reg_14__3_ ( .D(n1119), .CLK(clk), .Q(mem[227]) );
  DFFPOSX1 mem_reg_14__2_ ( .D(n1118), .CLK(clk), .Q(mem[226]) );
  DFFPOSX1 mem_reg_14__1_ ( .D(n1117), .CLK(clk), .Q(mem[225]) );
  DFFPOSX1 mem_reg_14__0_ ( .D(n1116), .CLK(clk), .Q(mem[224]) );
  DFFPOSX1 mem_reg_13__15_ ( .D(n1115), .CLK(clk), .Q(mem[223]) );
  DFFPOSX1 mem_reg_13__14_ ( .D(n1114), .CLK(clk), .Q(mem[222]) );
  DFFPOSX1 mem_reg_13__13_ ( .D(n1113), .CLK(clk), .Q(mem[221]) );
  DFFPOSX1 mem_reg_13__12_ ( .D(n1112), .CLK(clk), .Q(mem[220]) );
  DFFPOSX1 mem_reg_13__11_ ( .D(n1111), .CLK(clk), .Q(mem[219]) );
  DFFPOSX1 mem_reg_13__10_ ( .D(n1110), .CLK(clk), .Q(mem[218]) );
  DFFPOSX1 mem_reg_13__9_ ( .D(n1109), .CLK(clk), .Q(mem[217]) );
  DFFPOSX1 mem_reg_13__8_ ( .D(n1108), .CLK(clk), .Q(mem[216]) );
  DFFPOSX1 mem_reg_13__7_ ( .D(n1107), .CLK(clk), .Q(mem[215]) );
  DFFPOSX1 mem_reg_13__6_ ( .D(n1106), .CLK(clk), .Q(mem[214]) );
  DFFPOSX1 mem_reg_13__5_ ( .D(n1105), .CLK(clk), .Q(mem[213]) );
  DFFPOSX1 mem_reg_13__4_ ( .D(n1104), .CLK(clk), .Q(mem[212]) );
  DFFPOSX1 mem_reg_13__3_ ( .D(n1103), .CLK(clk), .Q(mem[211]) );
  DFFPOSX1 mem_reg_13__2_ ( .D(n1102), .CLK(clk), .Q(mem[210]) );
  DFFPOSX1 mem_reg_13__1_ ( .D(n1101), .CLK(clk), .Q(mem[209]) );
  DFFPOSX1 mem_reg_13__0_ ( .D(n1100), .CLK(clk), .Q(mem[208]) );
  DFFPOSX1 mem_reg_12__15_ ( .D(n1099), .CLK(clk), .Q(mem[207]) );
  DFFPOSX1 mem_reg_12__14_ ( .D(n1098), .CLK(clk), .Q(mem[206]) );
  DFFPOSX1 mem_reg_12__13_ ( .D(n1097), .CLK(clk), .Q(mem[205]) );
  DFFPOSX1 mem_reg_12__12_ ( .D(n1096), .CLK(clk), .Q(mem[204]) );
  DFFPOSX1 mem_reg_12__11_ ( .D(n1095), .CLK(clk), .Q(mem[203]) );
  DFFPOSX1 mem_reg_12__10_ ( .D(n1094), .CLK(clk), .Q(mem[202]) );
  DFFPOSX1 mem_reg_12__9_ ( .D(n1093), .CLK(clk), .Q(mem[201]) );
  DFFPOSX1 mem_reg_12__8_ ( .D(n1092), .CLK(clk), .Q(mem[200]) );
  DFFPOSX1 mem_reg_12__7_ ( .D(n1091), .CLK(clk), .Q(mem[199]) );
  DFFPOSX1 mem_reg_12__6_ ( .D(n1090), .CLK(clk), .Q(mem[198]) );
  DFFPOSX1 mem_reg_12__5_ ( .D(n1089), .CLK(clk), .Q(mem[197]) );
  DFFPOSX1 mem_reg_12__4_ ( .D(n1088), .CLK(clk), .Q(mem[196]) );
  DFFPOSX1 mem_reg_12__3_ ( .D(n1087), .CLK(clk), .Q(mem[195]) );
  DFFPOSX1 mem_reg_12__2_ ( .D(n1086), .CLK(clk), .Q(mem[194]) );
  DFFPOSX1 mem_reg_12__1_ ( .D(n1085), .CLK(clk), .Q(mem[193]) );
  DFFPOSX1 mem_reg_12__0_ ( .D(n1084), .CLK(clk), .Q(mem[192]) );
  DFFPOSX1 mem_reg_11__15_ ( .D(n1083), .CLK(clk), .Q(mem[191]) );
  DFFPOSX1 mem_reg_11__14_ ( .D(n1082), .CLK(clk), .Q(mem[190]) );
  DFFPOSX1 mem_reg_11__13_ ( .D(n1081), .CLK(clk), .Q(mem[189]) );
  DFFPOSX1 mem_reg_11__12_ ( .D(n1080), .CLK(clk), .Q(mem[188]) );
  DFFPOSX1 mem_reg_11__11_ ( .D(n1079), .CLK(clk), .Q(mem[187]) );
  DFFPOSX1 mem_reg_11__10_ ( .D(n1078), .CLK(clk), .Q(mem[186]) );
  DFFPOSX1 mem_reg_11__9_ ( .D(n1077), .CLK(clk), .Q(mem[185]) );
  DFFPOSX1 mem_reg_11__8_ ( .D(n1076), .CLK(clk), .Q(mem[184]) );
  DFFPOSX1 mem_reg_11__7_ ( .D(n1075), .CLK(clk), .Q(mem[183]) );
  DFFPOSX1 mem_reg_11__6_ ( .D(n1074), .CLK(clk), .Q(mem[182]) );
  DFFPOSX1 mem_reg_11__5_ ( .D(n1073), .CLK(clk), .Q(mem[181]) );
  DFFPOSX1 mem_reg_11__4_ ( .D(n1072), .CLK(clk), .Q(mem[180]) );
  DFFPOSX1 mem_reg_11__3_ ( .D(n1071), .CLK(clk), .Q(mem[179]) );
  DFFPOSX1 mem_reg_11__2_ ( .D(n1070), .CLK(clk), .Q(mem[178]) );
  DFFPOSX1 mem_reg_11__1_ ( .D(n1069), .CLK(clk), .Q(mem[177]) );
  DFFPOSX1 mem_reg_11__0_ ( .D(n1068), .CLK(clk), .Q(mem[176]) );
  DFFPOSX1 mem_reg_10__15_ ( .D(n1067), .CLK(clk), .Q(mem[175]) );
  DFFPOSX1 mem_reg_10__14_ ( .D(n1066), .CLK(clk), .Q(mem[174]) );
  DFFPOSX1 mem_reg_10__13_ ( .D(n1065), .CLK(clk), .Q(mem[173]) );
  DFFPOSX1 mem_reg_10__12_ ( .D(n1064), .CLK(clk), .Q(mem[172]) );
  DFFPOSX1 mem_reg_10__11_ ( .D(n1063), .CLK(clk), .Q(mem[171]) );
  DFFPOSX1 mem_reg_10__10_ ( .D(n1062), .CLK(clk), .Q(mem[170]) );
  DFFPOSX1 mem_reg_10__9_ ( .D(n1061), .CLK(clk), .Q(mem[169]) );
  DFFPOSX1 mem_reg_10__8_ ( .D(n1060), .CLK(clk), .Q(mem[168]) );
  DFFPOSX1 mem_reg_10__7_ ( .D(n1059), .CLK(clk), .Q(mem[167]) );
  DFFPOSX1 mem_reg_10__6_ ( .D(n1058), .CLK(clk), .Q(mem[166]) );
  DFFPOSX1 mem_reg_10__5_ ( .D(n1057), .CLK(clk), .Q(mem[165]) );
  DFFPOSX1 mem_reg_10__4_ ( .D(n1056), .CLK(clk), .Q(mem[164]) );
  DFFPOSX1 mem_reg_10__3_ ( .D(n1055), .CLK(clk), .Q(mem[163]) );
  DFFPOSX1 mem_reg_10__2_ ( .D(n1054), .CLK(clk), .Q(mem[162]) );
  DFFPOSX1 mem_reg_10__1_ ( .D(n1053), .CLK(clk), .Q(mem[161]) );
  DFFPOSX1 mem_reg_10__0_ ( .D(n1052), .CLK(clk), .Q(mem[160]) );
  DFFPOSX1 mem_reg_9__15_ ( .D(n1051), .CLK(clk), .Q(mem[159]) );
  DFFPOSX1 mem_reg_9__14_ ( .D(n1050), .CLK(clk), .Q(mem[158]) );
  DFFPOSX1 mem_reg_9__13_ ( .D(n1049), .CLK(clk), .Q(mem[157]) );
  DFFPOSX1 mem_reg_9__12_ ( .D(n1048), .CLK(clk), .Q(mem[156]) );
  DFFPOSX1 mem_reg_9__11_ ( .D(n1047), .CLK(clk), .Q(mem[155]) );
  DFFPOSX1 mem_reg_9__10_ ( .D(n1046), .CLK(clk), .Q(mem[154]) );
  DFFPOSX1 mem_reg_9__9_ ( .D(n1045), .CLK(clk), .Q(mem[153]) );
  DFFPOSX1 mem_reg_9__8_ ( .D(n1044), .CLK(clk), .Q(mem[152]) );
  DFFPOSX1 mem_reg_9__7_ ( .D(n1043), .CLK(clk), .Q(mem[151]) );
  DFFPOSX1 mem_reg_9__6_ ( .D(n1042), .CLK(clk), .Q(mem[150]) );
  DFFPOSX1 mem_reg_9__5_ ( .D(n1041), .CLK(clk), .Q(mem[149]) );
  DFFPOSX1 mem_reg_9__4_ ( .D(n1040), .CLK(clk), .Q(mem[148]) );
  DFFPOSX1 mem_reg_9__3_ ( .D(n1039), .CLK(clk), .Q(mem[147]) );
  DFFPOSX1 mem_reg_9__2_ ( .D(n1038), .CLK(clk), .Q(mem[146]) );
  DFFPOSX1 mem_reg_9__1_ ( .D(n1037), .CLK(clk), .Q(mem[145]) );
  DFFPOSX1 mem_reg_9__0_ ( .D(n1036), .CLK(clk), .Q(mem[144]) );
  DFFPOSX1 mem_reg_8__15_ ( .D(n1035), .CLK(clk), .Q(mem[143]) );
  DFFPOSX1 mem_reg_8__14_ ( .D(n1034), .CLK(clk), .Q(mem[142]) );
  DFFPOSX1 mem_reg_8__13_ ( .D(n1033), .CLK(clk), .Q(mem[141]) );
  DFFPOSX1 mem_reg_8__12_ ( .D(n1032), .CLK(clk), .Q(mem[140]) );
  DFFPOSX1 mem_reg_8__11_ ( .D(n1031), .CLK(clk), .Q(mem[139]) );
  DFFPOSX1 mem_reg_8__10_ ( .D(n1030), .CLK(clk), .Q(mem[138]) );
  DFFPOSX1 mem_reg_8__9_ ( .D(n1029), .CLK(clk), .Q(mem[137]) );
  DFFPOSX1 mem_reg_8__8_ ( .D(n1028), .CLK(clk), .Q(mem[136]) );
  DFFPOSX1 mem_reg_8__7_ ( .D(n1027), .CLK(clk), .Q(mem[135]) );
  DFFPOSX1 mem_reg_8__6_ ( .D(n1026), .CLK(clk), .Q(mem[134]) );
  DFFPOSX1 mem_reg_8__5_ ( .D(n1025), .CLK(clk), .Q(mem[133]) );
  DFFPOSX1 mem_reg_8__4_ ( .D(n1024), .CLK(clk), .Q(mem[132]) );
  DFFPOSX1 mem_reg_8__3_ ( .D(n1023), .CLK(clk), .Q(mem[131]) );
  DFFPOSX1 mem_reg_8__2_ ( .D(n1022), .CLK(clk), .Q(mem[130]) );
  DFFPOSX1 mem_reg_8__1_ ( .D(n1021), .CLK(clk), .Q(mem[129]) );
  DFFPOSX1 mem_reg_8__0_ ( .D(n1020), .CLK(clk), .Q(mem[128]) );
  DFFPOSX1 mem_reg_7__15_ ( .D(n1019), .CLK(clk), .Q(mem[127]) );
  DFFPOSX1 mem_reg_7__14_ ( .D(n1018), .CLK(clk), .Q(mem[126]) );
  DFFPOSX1 mem_reg_7__13_ ( .D(n1017), .CLK(clk), .Q(mem[125]) );
  DFFPOSX1 mem_reg_7__12_ ( .D(n1016), .CLK(clk), .Q(mem[124]) );
  DFFPOSX1 mem_reg_7__11_ ( .D(n1015), .CLK(clk), .Q(mem[123]) );
  DFFPOSX1 mem_reg_7__10_ ( .D(n1014), .CLK(clk), .Q(mem[122]) );
  DFFPOSX1 mem_reg_7__9_ ( .D(n1013), .CLK(clk), .Q(mem[121]) );
  DFFPOSX1 mem_reg_7__8_ ( .D(n1012), .CLK(clk), .Q(mem[120]) );
  DFFPOSX1 mem_reg_7__7_ ( .D(n1011), .CLK(clk), .Q(mem[119]) );
  DFFPOSX1 mem_reg_7__6_ ( .D(n1010), .CLK(clk), .Q(mem[118]) );
  DFFPOSX1 mem_reg_7__5_ ( .D(n1009), .CLK(clk), .Q(mem[117]) );
  DFFPOSX1 mem_reg_7__4_ ( .D(n1008), .CLK(clk), .Q(mem[116]) );
  DFFPOSX1 mem_reg_7__3_ ( .D(n1007), .CLK(clk), .Q(mem[115]) );
  DFFPOSX1 mem_reg_7__2_ ( .D(n1006), .CLK(clk), .Q(mem[114]) );
  DFFPOSX1 mem_reg_7__1_ ( .D(n1005), .CLK(clk), .Q(mem[113]) );
  DFFPOSX1 mem_reg_7__0_ ( .D(n1004), .CLK(clk), .Q(mem[112]) );
  DFFPOSX1 mem_reg_6__15_ ( .D(n1003), .CLK(clk), .Q(mem[111]) );
  DFFPOSX1 mem_reg_6__14_ ( .D(n1002), .CLK(clk), .Q(mem[110]) );
  DFFPOSX1 mem_reg_6__13_ ( .D(n1001), .CLK(clk), .Q(mem[109]) );
  DFFPOSX1 mem_reg_6__12_ ( .D(n1000), .CLK(clk), .Q(mem[108]) );
  DFFPOSX1 mem_reg_6__11_ ( .D(n999), .CLK(clk), .Q(mem[107]) );
  DFFPOSX1 mem_reg_6__10_ ( .D(n998), .CLK(clk), .Q(mem[106]) );
  DFFPOSX1 mem_reg_6__9_ ( .D(n997), .CLK(clk), .Q(mem[105]) );
  DFFPOSX1 mem_reg_6__8_ ( .D(n996), .CLK(clk), .Q(mem[104]) );
  DFFPOSX1 mem_reg_6__7_ ( .D(n995), .CLK(clk), .Q(mem[103]) );
  DFFPOSX1 mem_reg_6__6_ ( .D(n994), .CLK(clk), .Q(mem[102]) );
  DFFPOSX1 mem_reg_6__5_ ( .D(n993), .CLK(clk), .Q(mem[101]) );
  DFFPOSX1 mem_reg_6__4_ ( .D(n992), .CLK(clk), .Q(mem[100]) );
  DFFPOSX1 mem_reg_6__3_ ( .D(n991), .CLK(clk), .Q(mem[99]) );
  DFFPOSX1 mem_reg_6__2_ ( .D(n990), .CLK(clk), .Q(mem[98]) );
  DFFPOSX1 mem_reg_6__1_ ( .D(n989), .CLK(clk), .Q(mem[97]) );
  DFFPOSX1 mem_reg_6__0_ ( .D(n988), .CLK(clk), .Q(mem[96]) );
  DFFPOSX1 mem_reg_5__15_ ( .D(n987), .CLK(clk), .Q(mem[95]) );
  DFFPOSX1 mem_reg_5__14_ ( .D(n986), .CLK(clk), .Q(mem[94]) );
  DFFPOSX1 mem_reg_5__13_ ( .D(n985), .CLK(clk), .Q(mem[93]) );
  DFFPOSX1 mem_reg_5__12_ ( .D(n984), .CLK(clk), .Q(mem[92]) );
  DFFPOSX1 mem_reg_5__11_ ( .D(n983), .CLK(clk), .Q(mem[91]) );
  DFFPOSX1 mem_reg_5__10_ ( .D(n982), .CLK(clk), .Q(mem[90]) );
  DFFPOSX1 mem_reg_5__9_ ( .D(n981), .CLK(clk), .Q(mem[89]) );
  DFFPOSX1 mem_reg_5__8_ ( .D(n980), .CLK(clk), .Q(mem[88]) );
  DFFPOSX1 mem_reg_5__7_ ( .D(n979), .CLK(clk), .Q(mem[87]) );
  DFFPOSX1 mem_reg_5__6_ ( .D(n978), .CLK(clk), .Q(mem[86]) );
  DFFPOSX1 mem_reg_5__5_ ( .D(n977), .CLK(clk), .Q(mem[85]) );
  DFFPOSX1 mem_reg_5__4_ ( .D(n976), .CLK(clk), .Q(mem[84]) );
  DFFPOSX1 mem_reg_5__3_ ( .D(n975), .CLK(clk), .Q(mem[83]) );
  DFFPOSX1 mem_reg_5__2_ ( .D(n974), .CLK(clk), .Q(mem[82]) );
  DFFPOSX1 mem_reg_5__1_ ( .D(n973), .CLK(clk), .Q(mem[81]) );
  DFFPOSX1 mem_reg_5__0_ ( .D(n972), .CLK(clk), .Q(mem[80]) );
  DFFPOSX1 mem_reg_4__15_ ( .D(n971), .CLK(clk), .Q(mem[79]) );
  DFFPOSX1 mem_reg_4__14_ ( .D(n970), .CLK(clk), .Q(mem[78]) );
  DFFPOSX1 mem_reg_4__13_ ( .D(n969), .CLK(clk), .Q(mem[77]) );
  DFFPOSX1 mem_reg_4__12_ ( .D(n968), .CLK(clk), .Q(mem[76]) );
  DFFPOSX1 mem_reg_4__11_ ( .D(n967), .CLK(clk), .Q(mem[75]) );
  DFFPOSX1 mem_reg_4__10_ ( .D(n966), .CLK(clk), .Q(mem[74]) );
  DFFPOSX1 mem_reg_4__9_ ( .D(n965), .CLK(clk), .Q(mem[73]) );
  DFFPOSX1 mem_reg_4__8_ ( .D(n964), .CLK(clk), .Q(mem[72]) );
  DFFPOSX1 mem_reg_4__7_ ( .D(n963), .CLK(clk), .Q(mem[71]) );
  DFFPOSX1 mem_reg_4__6_ ( .D(n962), .CLK(clk), .Q(mem[70]) );
  DFFPOSX1 mem_reg_4__5_ ( .D(n961), .CLK(clk), .Q(mem[69]) );
  DFFPOSX1 mem_reg_4__4_ ( .D(n960), .CLK(clk), .Q(mem[68]) );
  DFFPOSX1 mem_reg_4__3_ ( .D(n959), .CLK(clk), .Q(mem[67]) );
  DFFPOSX1 mem_reg_4__2_ ( .D(n958), .CLK(clk), .Q(mem[66]) );
  DFFPOSX1 mem_reg_4__1_ ( .D(n957), .CLK(clk), .Q(mem[65]) );
  DFFPOSX1 mem_reg_4__0_ ( .D(n956), .CLK(clk), .Q(mem[64]) );
  DFFPOSX1 mem_reg_3__15_ ( .D(n955), .CLK(clk), .Q(mem[63]) );
  DFFPOSX1 mem_reg_3__14_ ( .D(n954), .CLK(clk), .Q(mem[62]) );
  DFFPOSX1 mem_reg_3__13_ ( .D(n953), .CLK(clk), .Q(mem[61]) );
  DFFPOSX1 mem_reg_3__12_ ( .D(n952), .CLK(clk), .Q(mem[60]) );
  DFFPOSX1 mem_reg_3__11_ ( .D(n951), .CLK(clk), .Q(mem[59]) );
  DFFPOSX1 mem_reg_3__10_ ( .D(n950), .CLK(clk), .Q(mem[58]) );
  DFFPOSX1 mem_reg_3__9_ ( .D(n949), .CLK(clk), .Q(mem[57]) );
  DFFPOSX1 mem_reg_3__8_ ( .D(n948), .CLK(clk), .Q(mem[56]) );
  DFFPOSX1 mem_reg_3__7_ ( .D(n947), .CLK(clk), .Q(mem[55]) );
  DFFPOSX1 mem_reg_3__6_ ( .D(n946), .CLK(clk), .Q(mem[54]) );
  DFFPOSX1 mem_reg_3__5_ ( .D(n945), .CLK(clk), .Q(mem[53]) );
  DFFPOSX1 mem_reg_3__4_ ( .D(n944), .CLK(clk), .Q(mem[52]) );
  DFFPOSX1 mem_reg_3__3_ ( .D(n943), .CLK(clk), .Q(mem[51]) );
  DFFPOSX1 mem_reg_3__2_ ( .D(n942), .CLK(clk), .Q(mem[50]) );
  DFFPOSX1 mem_reg_3__1_ ( .D(n941), .CLK(clk), .Q(mem[49]) );
  DFFPOSX1 mem_reg_3__0_ ( .D(n940), .CLK(clk), .Q(mem[48]) );
  DFFPOSX1 mem_reg_2__15_ ( .D(n939), .CLK(clk), .Q(mem[47]) );
  DFFPOSX1 mem_reg_2__14_ ( .D(n938), .CLK(clk), .Q(mem[46]) );
  DFFPOSX1 mem_reg_2__13_ ( .D(n937), .CLK(clk), .Q(mem[45]) );
  DFFPOSX1 mem_reg_2__12_ ( .D(n936), .CLK(clk), .Q(mem[44]) );
  DFFPOSX1 mem_reg_2__11_ ( .D(n935), .CLK(clk), .Q(mem[43]) );
  DFFPOSX1 mem_reg_2__10_ ( .D(n934), .CLK(clk), .Q(mem[42]) );
  DFFPOSX1 mem_reg_2__9_ ( .D(n933), .CLK(clk), .Q(mem[41]) );
  DFFPOSX1 mem_reg_2__8_ ( .D(n932), .CLK(clk), .Q(mem[40]) );
  DFFPOSX1 mem_reg_2__7_ ( .D(n931), .CLK(clk), .Q(mem[39]) );
  DFFPOSX1 mem_reg_2__6_ ( .D(n930), .CLK(clk), .Q(mem[38]) );
  DFFPOSX1 mem_reg_2__5_ ( .D(n929), .CLK(clk), .Q(mem[37]) );
  DFFPOSX1 mem_reg_2__4_ ( .D(n928), .CLK(clk), .Q(mem[36]) );
  DFFPOSX1 mem_reg_2__3_ ( .D(n927), .CLK(clk), .Q(mem[35]) );
  DFFPOSX1 mem_reg_2__2_ ( .D(n926), .CLK(clk), .Q(mem[34]) );
  DFFPOSX1 mem_reg_2__1_ ( .D(n925), .CLK(clk), .Q(mem[33]) );
  DFFPOSX1 mem_reg_2__0_ ( .D(n924), .CLK(clk), .Q(mem[32]) );
  DFFPOSX1 mem_reg_1__15_ ( .D(n923), .CLK(clk), .Q(mem[31]) );
  DFFPOSX1 mem_reg_1__14_ ( .D(n922), .CLK(clk), .Q(mem[30]) );
  DFFPOSX1 mem_reg_1__13_ ( .D(n921), .CLK(clk), .Q(mem[29]) );
  DFFPOSX1 mem_reg_1__12_ ( .D(n920), .CLK(clk), .Q(mem[28]) );
  DFFPOSX1 mem_reg_1__11_ ( .D(n919), .CLK(clk), .Q(mem[27]) );
  DFFPOSX1 mem_reg_1__10_ ( .D(n918), .CLK(clk), .Q(mem[26]) );
  DFFPOSX1 mem_reg_1__9_ ( .D(n917), .CLK(clk), .Q(mem[25]) );
  DFFPOSX1 mem_reg_1__8_ ( .D(n916), .CLK(clk), .Q(mem[24]) );
  DFFPOSX1 mem_reg_1__7_ ( .D(n915), .CLK(clk), .Q(mem[23]) );
  DFFPOSX1 mem_reg_1__6_ ( .D(n914), .CLK(clk), .Q(mem[22]) );
  DFFPOSX1 mem_reg_1__5_ ( .D(n913), .CLK(clk), .Q(mem[21]) );
  DFFPOSX1 mem_reg_1__4_ ( .D(n912), .CLK(clk), .Q(mem[20]) );
  DFFPOSX1 mem_reg_1__3_ ( .D(n911), .CLK(clk), .Q(mem[19]) );
  DFFPOSX1 mem_reg_1__2_ ( .D(n910), .CLK(clk), .Q(mem[18]) );
  DFFPOSX1 mem_reg_1__1_ ( .D(n909), .CLK(clk), .Q(mem[17]) );
  DFFPOSX1 mem_reg_1__0_ ( .D(n908), .CLK(clk), .Q(mem[16]) );
  DFFPOSX1 mem_reg_0__15_ ( .D(n907), .CLK(clk), .Q(mem[15]) );
  DFFPOSX1 mem_reg_0__14_ ( .D(n906), .CLK(clk), .Q(mem[14]) );
  DFFPOSX1 mem_reg_0__13_ ( .D(n905), .CLK(clk), .Q(mem[13]) );
  DFFPOSX1 mem_reg_0__12_ ( .D(n904), .CLK(clk), .Q(mem[12]) );
  DFFPOSX1 mem_reg_0__11_ ( .D(n903), .CLK(clk), .Q(mem[11]) );
  DFFPOSX1 mem_reg_0__10_ ( .D(n902), .CLK(clk), .Q(mem[10]) );
  DFFPOSX1 mem_reg_0__9_ ( .D(n901), .CLK(clk), .Q(mem[9]) );
  DFFPOSX1 mem_reg_0__8_ ( .D(n900), .CLK(clk), .Q(mem[8]) );
  DFFPOSX1 mem_reg_0__7_ ( .D(n899), .CLK(clk), .Q(mem[7]) );
  DFFPOSX1 mem_reg_0__6_ ( .D(n898), .CLK(clk), .Q(mem[6]) );
  DFFPOSX1 mem_reg_0__5_ ( .D(n897), .CLK(clk), .Q(mem[5]) );
  DFFPOSX1 mem_reg_0__4_ ( .D(n896), .CLK(clk), .Q(mem[4]) );
  DFFPOSX1 mem_reg_0__3_ ( .D(n895), .CLK(clk), .Q(mem[3]) );
  DFFPOSX1 mem_reg_0__2_ ( .D(n894), .CLK(clk), .Q(mem[2]) );
  DFFPOSX1 mem_reg_0__1_ ( .D(n893), .CLK(clk), .Q(mem[1]) );
  DFFPOSX1 mem_reg_0__0_ ( .D(n892), .CLK(clk), .Q(mem[0]) );
  OAI21X1 U66 ( .A(n2271), .B(n2287), .C(n1699), .Y(n892) );
  OAI21X1 U68 ( .A(n2271), .B(n2286), .C(n1659), .Y(n893) );
  OAI21X1 U70 ( .A(n2271), .B(n2285), .C(n1619), .Y(n894) );
  OAI21X1 U72 ( .A(n2271), .B(n2284), .C(n1577), .Y(n895) );
  OAI21X1 U74 ( .A(n2271), .B(n2283), .C(n1535), .Y(n896) );
  OAI21X1 U76 ( .A(n2271), .B(n2282), .C(n1498), .Y(n897) );
  OAI21X1 U78 ( .A(n2271), .B(n2281), .C(n1460), .Y(n898) );
  OAI21X1 U80 ( .A(n2271), .B(n2280), .C(n1422), .Y(n899) );
  OAI21X1 U82 ( .A(n2271), .B(n2279), .C(n270), .Y(n900) );
  OAI21X1 U84 ( .A(n2271), .B(n2278), .C(n239), .Y(n901) );
  OAI21X1 U86 ( .A(n2271), .B(n2277), .C(n209), .Y(n902) );
  OAI21X1 U88 ( .A(n2271), .B(n2276), .C(n179), .Y(n903) );
  OAI21X1 U90 ( .A(n2271), .B(n2275), .C(n1698), .Y(n904) );
  OAI21X1 U92 ( .A(n2271), .B(n2274), .C(n1658), .Y(n905) );
  OAI21X1 U94 ( .A(n2271), .B(n2273), .C(n149), .Y(n906) );
  OAI21X1 U96 ( .A(n2271), .B(n2272), .C(n123), .Y(n907) );
  OAI21X1 U98 ( .A(n1579), .B(n1538), .C(reset), .Y(n312) );
  OAI21X1 U99 ( .A(n2270), .B(n2287), .C(n1657), .Y(n908) );
  OAI21X1 U101 ( .A(n2270), .B(n2286), .C(n1697), .Y(n909) );
  OAI21X1 U103 ( .A(n2270), .B(n2285), .C(n1576), .Y(n910) );
  OAI21X1 U105 ( .A(n2270), .B(n2284), .C(n1618), .Y(n911) );
  OAI21X1 U107 ( .A(n2270), .B(n2283), .C(n1497), .Y(n912) );
  OAI21X1 U109 ( .A(n2270), .B(n2282), .C(n1534), .Y(n913) );
  OAI21X1 U111 ( .A(n2270), .B(n2281), .C(n1421), .Y(n914) );
  OAI21X1 U113 ( .A(n2270), .B(n2280), .C(n1459), .Y(n915) );
  OAI21X1 U115 ( .A(n2270), .B(n2279), .C(n238), .Y(n916) );
  OAI21X1 U117 ( .A(n2270), .B(n2278), .C(n269), .Y(n917) );
  OAI21X1 U119 ( .A(n2270), .B(n2277), .C(n178), .Y(n918) );
  OAI21X1 U121 ( .A(n2270), .B(n2276), .C(n208), .Y(n919) );
  OAI21X1 U123 ( .A(n2270), .B(n2275), .C(n1656), .Y(n920) );
  OAI21X1 U125 ( .A(n2270), .B(n2274), .C(n1696), .Y(n921) );
  OAI21X1 U127 ( .A(n2270), .B(n2273), .C(n122), .Y(n922) );
  OAI21X1 U129 ( .A(n2270), .B(n2272), .C(n148), .Y(n923) );
  OAI21X1 U131 ( .A(n1579), .B(n1500), .C(reset), .Y(n331) );
  OAI21X1 U132 ( .A(n2269), .B(n2287), .C(n1617), .Y(n924) );
  OAI21X1 U134 ( .A(n2269), .B(n2286), .C(n1575), .Y(n925) );
  OAI21X1 U136 ( .A(n2269), .B(n2285), .C(n1695), .Y(n926) );
  OAI21X1 U138 ( .A(n2269), .B(n2284), .C(n1655), .Y(n927) );
  OAI21X1 U140 ( .A(n2269), .B(n2283), .C(n1458), .Y(n928) );
  OAI21X1 U142 ( .A(n2269), .B(n2282), .C(n1420), .Y(n929) );
  OAI21X1 U144 ( .A(n2269), .B(n2281), .C(n1533), .Y(n930) );
  OAI21X1 U146 ( .A(n2269), .B(n2280), .C(n1496), .Y(n931) );
  OAI21X1 U148 ( .A(n2269), .B(n2279), .C(n207), .Y(n932) );
  OAI21X1 U150 ( .A(n2269), .B(n2278), .C(n177), .Y(n933) );
  OAI21X1 U152 ( .A(n2269), .B(n2277), .C(n268), .Y(n934) );
  OAI21X1 U154 ( .A(n2269), .B(n2276), .C(n237), .Y(n935) );
  OAI21X1 U156 ( .A(n2269), .B(n2275), .C(n1616), .Y(n936) );
  OAI21X1 U158 ( .A(n2269), .B(n2274), .C(n1574), .Y(n937) );
  OAI21X1 U160 ( .A(n2269), .B(n2273), .C(n97), .Y(n938) );
  OAI21X1 U162 ( .A(n2269), .B(n2272), .C(n51), .Y(n939) );
  OAI21X1 U164 ( .A(n1579), .B(n1462), .C(reset), .Y(n349) );
  OAI21X1 U165 ( .A(n2268), .B(n2287), .C(n1573), .Y(n940) );
  OAI21X1 U167 ( .A(n2268), .B(n2286), .C(n1615), .Y(n941) );
  OAI21X1 U169 ( .A(n2268), .B(n2285), .C(n1654), .Y(n942) );
  OAI21X1 U171 ( .A(n2268), .B(n2284), .C(n1694), .Y(n943) );
  OAI21X1 U173 ( .A(n2268), .B(n2283), .C(n1419), .Y(n944) );
  OAI21X1 U175 ( .A(n2268), .B(n2282), .C(n1457), .Y(n945) );
  OAI21X1 U177 ( .A(n2268), .B(n2281), .C(n1495), .Y(n946) );
  OAI21X1 U179 ( .A(n2268), .B(n2280), .C(n1532), .Y(n947) );
  OAI21X1 U181 ( .A(n2268), .B(n2279), .C(n176), .Y(n948) );
  OAI21X1 U183 ( .A(n2268), .B(n2278), .C(n206), .Y(n949) );
  OAI21X1 U185 ( .A(n2268), .B(n2277), .C(n236), .Y(n950) );
  OAI21X1 U187 ( .A(n2268), .B(n2276), .C(n267), .Y(n951) );
  OAI21X1 U189 ( .A(n2268), .B(n2275), .C(n1572), .Y(n952) );
  OAI21X1 U191 ( .A(n2268), .B(n2274), .C(n1614), .Y(n953) );
  OAI21X1 U193 ( .A(n2268), .B(n2273), .C(n50), .Y(n954) );
  OAI21X1 U195 ( .A(n2268), .B(n2272), .C(n96), .Y(n955) );
  OAI21X1 U197 ( .A(n1579), .B(n1424), .C(reset), .Y(n367) );
  OAI21X1 U198 ( .A(n2267), .B(n2287), .C(n1531), .Y(n956) );
  OAI21X1 U200 ( .A(n2267), .B(n2286), .C(n1494), .Y(n957) );
  OAI21X1 U202 ( .A(n2267), .B(n2285), .C(n1456), .Y(n958) );
  OAI21X1 U204 ( .A(n2267), .B(n2284), .C(n1418), .Y(n959) );
  OAI21X1 U206 ( .A(n2267), .B(n2283), .C(n1693), .Y(n960) );
  OAI21X1 U208 ( .A(n2267), .B(n2282), .C(n1653), .Y(n961) );
  OAI21X1 U210 ( .A(n2267), .B(n2281), .C(n1613), .Y(n962) );
  OAI21X1 U212 ( .A(n2267), .B(n2280), .C(n1571), .Y(n963) );
  OAI21X1 U214 ( .A(n2267), .B(n2279), .C(n147), .Y(n964) );
  OAI21X1 U216 ( .A(n2267), .B(n2278), .C(n121), .Y(n965) );
  OAI21X1 U218 ( .A(n2267), .B(n2277), .C(n95), .Y(n966) );
  OAI21X1 U220 ( .A(n2267), .B(n2276), .C(n49), .Y(n967) );
  OAI21X1 U222 ( .A(n2267), .B(n2275), .C(n1530), .Y(n968) );
  OAI21X1 U224 ( .A(n2267), .B(n2274), .C(n1493), .Y(n969) );
  OAI21X1 U226 ( .A(n2267), .B(n2273), .C(n266), .Y(n970) );
  OAI21X1 U228 ( .A(n2267), .B(n2272), .C(n235), .Y(n971) );
  OAI21X1 U230 ( .A(n1579), .B(n1423), .C(reset), .Y(n385) );
  OAI21X1 U231 ( .A(n2266), .B(n2287), .C(n1492), .Y(n972) );
  OAI21X1 U233 ( .A(n2266), .B(n2286), .C(n1529), .Y(n973) );
  OAI21X1 U235 ( .A(n2266), .B(n2285), .C(n1417), .Y(n974) );
  OAI21X1 U237 ( .A(n2266), .B(n2284), .C(n1455), .Y(n975) );
  OAI21X1 U239 ( .A(n2266), .B(n2283), .C(n1652), .Y(n976) );
  OAI21X1 U241 ( .A(n2266), .B(n2282), .C(n1692), .Y(n977) );
  OAI21X1 U243 ( .A(n2266), .B(n2281), .C(n1570), .Y(n978) );
  OAI21X1 U245 ( .A(n2266), .B(n2280), .C(n1612), .Y(n979) );
  OAI21X1 U247 ( .A(n2266), .B(n2279), .C(n120), .Y(n980) );
  OAI21X1 U249 ( .A(n2266), .B(n2278), .C(n146), .Y(n981) );
  OAI21X1 U251 ( .A(n2266), .B(n2277), .C(n48), .Y(n982) );
  OAI21X1 U253 ( .A(n2266), .B(n2276), .C(n94), .Y(n983) );
  OAI21X1 U255 ( .A(n2266), .B(n2275), .C(n1491), .Y(n984) );
  OAI21X1 U257 ( .A(n2266), .B(n2274), .C(n1528), .Y(n985) );
  OAI21X1 U259 ( .A(n2266), .B(n2273), .C(n234), .Y(n986) );
  OAI21X1 U261 ( .A(n2266), .B(n2272), .C(n265), .Y(n987) );
  OAI21X1 U263 ( .A(n1579), .B(n1461), .C(reset), .Y(n403) );
  OAI21X1 U264 ( .A(n2265), .B(n2287), .C(n1454), .Y(n988) );
  OAI21X1 U266 ( .A(n2265), .B(n2286), .C(n1416), .Y(n989) );
  OAI21X1 U268 ( .A(n2265), .B(n2285), .C(n1527), .Y(n990) );
  OAI21X1 U270 ( .A(n2265), .B(n2284), .C(n1490), .Y(n991) );
  OAI21X1 U272 ( .A(n2265), .B(n2283), .C(n1611), .Y(n992) );
  OAI21X1 U274 ( .A(n2265), .B(n2282), .C(n1569), .Y(n993) );
  OAI21X1 U276 ( .A(n2265), .B(n2281), .C(n1691), .Y(n994) );
  OAI21X1 U278 ( .A(n2265), .B(n2280), .C(n1651), .Y(n995) );
  OAI21X1 U280 ( .A(n2265), .B(n2279), .C(n93), .Y(n996) );
  OAI21X1 U282 ( .A(n2265), .B(n2278), .C(n47), .Y(n997) );
  OAI21X1 U284 ( .A(n2265), .B(n2277), .C(n145), .Y(n998) );
  OAI21X1 U286 ( .A(n2265), .B(n2276), .C(n119), .Y(n999) );
  OAI21X1 U288 ( .A(n2265), .B(n2275), .C(n1453), .Y(n1000) );
  OAI21X1 U290 ( .A(n2265), .B(n2274), .C(n1415), .Y(n1001) );
  OAI21X1 U292 ( .A(n2265), .B(n2273), .C(n205), .Y(n1002) );
  OAI21X1 U294 ( .A(n2265), .B(n2272), .C(n175), .Y(n1003) );
  OAI21X1 U296 ( .A(n1579), .B(n1499), .C(reset), .Y(n421) );
  OAI21X1 U297 ( .A(n2264), .B(n2287), .C(n1414), .Y(n1004) );
  OAI21X1 U299 ( .A(n2264), .B(n2286), .C(n1452), .Y(n1005) );
  OAI21X1 U301 ( .A(n2264), .B(n2285), .C(n1489), .Y(n1006) );
  OAI21X1 U303 ( .A(n2264), .B(n2284), .C(n1526), .Y(n1007) );
  OAI21X1 U305 ( .A(n2264), .B(n2283), .C(n1568), .Y(n1008) );
  OAI21X1 U307 ( .A(n2264), .B(n2282), .C(n1610), .Y(n1009) );
  OAI21X1 U309 ( .A(n2264), .B(n2281), .C(n1650), .Y(n1010) );
  OAI21X1 U311 ( .A(n2264), .B(n2280), .C(n1690), .Y(n1011) );
  OAI21X1 U313 ( .A(n2264), .B(n2279), .C(n46), .Y(n1012) );
  OAI21X1 U315 ( .A(n2264), .B(n2278), .C(n92), .Y(n1013) );
  OAI21X1 U317 ( .A(n2264), .B(n2277), .C(n118), .Y(n1014) );
  OAI21X1 U319 ( .A(n2264), .B(n2276), .C(n144), .Y(n1015) );
  OAI21X1 U321 ( .A(n2264), .B(n2275), .C(n310), .Y(n1016) );
  OAI21X1 U323 ( .A(n2264), .B(n2274), .C(n1451), .Y(n1017) );
  OAI21X1 U325 ( .A(n2264), .B(n2273), .C(n174), .Y(n1018) );
  OAI21X1 U327 ( .A(n2264), .B(n2272), .C(n204), .Y(n1019) );
  OAI21X1 U329 ( .A(n1579), .B(n1537), .C(reset), .Y(n439) );
  NAND3X1 U330 ( .A(n2313), .B(n2310), .C(n852), .Y(n313) );
  OAI21X1 U331 ( .A(n2263), .B(n2287), .C(n1689), .Y(n1020) );
  OAI21X1 U333 ( .A(n2263), .B(n2286), .C(n1649), .Y(n1021) );
  OAI21X1 U335 ( .A(n2263), .B(n2285), .C(n1609), .Y(n1022) );
  OAI21X1 U337 ( .A(n2263), .B(n2284), .C(n1567), .Y(n1023) );
  OAI21X1 U339 ( .A(n2263), .B(n2283), .C(n1525), .Y(n1024) );
  OAI21X1 U341 ( .A(n2263), .B(n2282), .C(n1488), .Y(n1025) );
  OAI21X1 U343 ( .A(n2263), .B(n2281), .C(n1450), .Y(n1026) );
  OAI21X1 U345 ( .A(n2263), .B(n2280), .C(n308), .Y(n1027) );
  OAI21X1 U347 ( .A(n2263), .B(n2279), .C(n264), .Y(n1028) );
  OAI21X1 U349 ( .A(n2263), .B(n2278), .C(n233), .Y(n1029) );
  OAI21X1 U351 ( .A(n2263), .B(n2277), .C(n203), .Y(n1030) );
  OAI21X1 U353 ( .A(n2263), .B(n2276), .C(n173), .Y(n1031) );
  OAI21X1 U355 ( .A(n2263), .B(n2275), .C(n1688), .Y(n1032) );
  OAI21X1 U357 ( .A(n2263), .B(n2274), .C(n1648), .Y(n1033) );
  OAI21X1 U359 ( .A(n2263), .B(n2273), .C(n143), .Y(n1034) );
  OAI21X1 U361 ( .A(n2263), .B(n2272), .C(n117), .Y(n1035) );
  OAI21X1 U363 ( .A(n1538), .B(n1702), .C(reset), .Y(n457) );
  OAI21X1 U364 ( .A(n2262), .B(n2287), .C(n1647), .Y(n1036) );
  OAI21X1 U366 ( .A(n2262), .B(n2286), .C(n1687), .Y(n1037) );
  OAI21X1 U368 ( .A(n2262), .B(n2285), .C(n1566), .Y(n1038) );
  OAI21X1 U370 ( .A(n2262), .B(n2284), .C(n1608), .Y(n1039) );
  OAI21X1 U372 ( .A(n2262), .B(n2283), .C(n1487), .Y(n1040) );
  OAI21X1 U374 ( .A(n2262), .B(n2282), .C(n1524), .Y(n1041) );
  OAI21X1 U376 ( .A(n2262), .B(n2281), .C(n306), .Y(n1042) );
  OAI21X1 U378 ( .A(n2262), .B(n2280), .C(n1449), .Y(n1043) );
  OAI21X1 U380 ( .A(n2262), .B(n2279), .C(n232), .Y(n1044) );
  OAI21X1 U382 ( .A(n2262), .B(n2278), .C(n263), .Y(n1045) );
  OAI21X1 U384 ( .A(n2262), .B(n2277), .C(n172), .Y(n1046) );
  OAI21X1 U386 ( .A(n2262), .B(n2276), .C(n202), .Y(n1047) );
  OAI21X1 U388 ( .A(n2262), .B(n2275), .C(n1646), .Y(n1048) );
  OAI21X1 U390 ( .A(n2262), .B(n2274), .C(n1686), .Y(n1049) );
  OAI21X1 U392 ( .A(n2262), .B(n2273), .C(n116), .Y(n1050) );
  OAI21X1 U394 ( .A(n2262), .B(n2272), .C(n142), .Y(n1051) );
  OAI21X1 U396 ( .A(n1500), .B(n1702), .C(reset), .Y(n475) );
  OAI21X1 U397 ( .A(n2261), .B(n2287), .C(n1607), .Y(n1052) );
  OAI21X1 U399 ( .A(n2261), .B(n2286), .C(n1565), .Y(n1053) );
  OAI21X1 U401 ( .A(n2261), .B(n2285), .C(n1685), .Y(n1054) );
  OAI21X1 U403 ( .A(n2261), .B(n2284), .C(n1645), .Y(n1055) );
  OAI21X1 U405 ( .A(n2261), .B(n2283), .C(n1448), .Y(n1056) );
  OAI21X1 U407 ( .A(n2261), .B(n2282), .C(n304), .Y(n1057) );
  OAI21X1 U409 ( .A(n2261), .B(n2281), .C(n1523), .Y(n1058) );
  OAI21X1 U411 ( .A(n2261), .B(n2280), .C(n1486), .Y(n1059) );
  OAI21X1 U413 ( .A(n2261), .B(n2279), .C(n201), .Y(n1060) );
  OAI21X1 U415 ( .A(n2261), .B(n2278), .C(n171), .Y(n1061) );
  OAI21X1 U417 ( .A(n2261), .B(n2277), .C(n262), .Y(n1062) );
  OAI21X1 U419 ( .A(n2261), .B(n2276), .C(n231), .Y(n1063) );
  OAI21X1 U421 ( .A(n2261), .B(n2275), .C(n1606), .Y(n1064) );
  OAI21X1 U423 ( .A(n2261), .B(n2274), .C(n1564), .Y(n1065) );
  OAI21X1 U425 ( .A(n2261), .B(n2273), .C(n91), .Y(n1066) );
  OAI21X1 U427 ( .A(n2261), .B(n2272), .C(n45), .Y(n1067) );
  OAI21X1 U429 ( .A(n1462), .B(n1702), .C(reset), .Y(n492) );
  OAI21X1 U430 ( .A(n2260), .B(n2287), .C(n1563), .Y(n1068) );
  OAI21X1 U432 ( .A(n2260), .B(n2286), .C(n1605), .Y(n1069) );
  OAI21X1 U434 ( .A(n2260), .B(n2285), .C(n1644), .Y(n1070) );
  OAI21X1 U436 ( .A(n2260), .B(n2284), .C(n1684), .Y(n1071) );
  OAI21X1 U438 ( .A(n2260), .B(n2283), .C(n302), .Y(n1072) );
  OAI21X1 U440 ( .A(n2260), .B(n2282), .C(n1447), .Y(n1073) );
  OAI21X1 U442 ( .A(n2260), .B(n2281), .C(n1485), .Y(n1074) );
  OAI21X1 U444 ( .A(n2260), .B(n2280), .C(n1522), .Y(n1075) );
  OAI21X1 U446 ( .A(n2260), .B(n2279), .C(n170), .Y(n1076) );
  OAI21X1 U448 ( .A(n2260), .B(n2278), .C(n200), .Y(n1077) );
  OAI21X1 U450 ( .A(n2260), .B(n2277), .C(n230), .Y(n1078) );
  OAI21X1 U452 ( .A(n2260), .B(n2276), .C(n261), .Y(n1079) );
  OAI21X1 U454 ( .A(n2260), .B(n2275), .C(n1562), .Y(n1080) );
  OAI21X1 U456 ( .A(n2260), .B(n2274), .C(n1604), .Y(n1081) );
  OAI21X1 U458 ( .A(n2260), .B(n2273), .C(n44), .Y(n1082) );
  OAI21X1 U460 ( .A(n2260), .B(n2272), .C(n90), .Y(n1083) );
  OAI21X1 U462 ( .A(n1424), .B(n1702), .C(reset), .Y(n509) );
  OAI21X1 U463 ( .A(n2259), .B(n2287), .C(n1521), .Y(n1084) );
  OAI21X1 U465 ( .A(n2259), .B(n2286), .C(n1484), .Y(n1085) );
  OAI21X1 U467 ( .A(n2259), .B(n2285), .C(n1446), .Y(n1086) );
  OAI21X1 U469 ( .A(n2259), .B(n2284), .C(n300), .Y(n1087) );
  OAI21X1 U471 ( .A(n2259), .B(n2283), .C(n1683), .Y(n1088) );
  OAI21X1 U473 ( .A(n2259), .B(n2282), .C(n1643), .Y(n1089) );
  OAI21X1 U475 ( .A(n2259), .B(n2281), .C(n1603), .Y(n1090) );
  OAI21X1 U477 ( .A(n2259), .B(n2280), .C(n1561), .Y(n1091) );
  OAI21X1 U479 ( .A(n2259), .B(n2279), .C(n141), .Y(n1092) );
  OAI21X1 U481 ( .A(n2259), .B(n2278), .C(n115), .Y(n1093) );
  OAI21X1 U483 ( .A(n2259), .B(n2277), .C(n89), .Y(n1094) );
  OAI21X1 U485 ( .A(n2259), .B(n2276), .C(n43), .Y(n1095) );
  OAI21X1 U487 ( .A(n2259), .B(n2275), .C(n1520), .Y(n1096) );
  OAI21X1 U489 ( .A(n2259), .B(n2274), .C(n1483), .Y(n1097) );
  OAI21X1 U491 ( .A(n2259), .B(n2273), .C(n260), .Y(n1098) );
  OAI21X1 U493 ( .A(n2259), .B(n2272), .C(n229), .Y(n1099) );
  OAI21X1 U495 ( .A(n1423), .B(n1702), .C(reset), .Y(n526) );
  OAI21X1 U496 ( .A(n2258), .B(n2287), .C(n1482), .Y(n1100) );
  OAI21X1 U498 ( .A(n2258), .B(n2286), .C(n1519), .Y(n1101) );
  OAI21X1 U500 ( .A(n2258), .B(n2285), .C(n298), .Y(n1102) );
  OAI21X1 U502 ( .A(n2258), .B(n2284), .C(n1445), .Y(n1103) );
  OAI21X1 U504 ( .A(n2258), .B(n2283), .C(n1642), .Y(n1104) );
  OAI21X1 U506 ( .A(n2258), .B(n2282), .C(n1682), .Y(n1105) );
  OAI21X1 U508 ( .A(n2258), .B(n2281), .C(n1560), .Y(n1106) );
  OAI21X1 U510 ( .A(n2258), .B(n2280), .C(n1602), .Y(n1107) );
  OAI21X1 U512 ( .A(n2258), .B(n2279), .C(n114), .Y(n1108) );
  OAI21X1 U514 ( .A(n2258), .B(n2278), .C(n140), .Y(n1109) );
  OAI21X1 U516 ( .A(n2258), .B(n2277), .C(n42), .Y(n1110) );
  OAI21X1 U518 ( .A(n2258), .B(n2276), .C(n88), .Y(n1111) );
  OAI21X1 U520 ( .A(n2258), .B(n2275), .C(n1481), .Y(n1112) );
  OAI21X1 U522 ( .A(n2258), .B(n2274), .C(n1518), .Y(n1113) );
  OAI21X1 U524 ( .A(n2258), .B(n2273), .C(n228), .Y(n1114) );
  OAI21X1 U526 ( .A(n2258), .B(n2272), .C(n259), .Y(n1115) );
  OAI21X1 U528 ( .A(n1461), .B(n1702), .C(reset), .Y(n543) );
  OAI21X1 U529 ( .A(n2257), .B(n2287), .C(n1444), .Y(n1116) );
  OAI21X1 U531 ( .A(n2257), .B(n2286), .C(n296), .Y(n1117) );
  OAI21X1 U533 ( .A(n2257), .B(n2285), .C(n1517), .Y(n1118) );
  OAI21X1 U535 ( .A(n2257), .B(n2284), .C(n1480), .Y(n1119) );
  OAI21X1 U537 ( .A(n2257), .B(n2283), .C(n1601), .Y(n1120) );
  OAI21X1 U539 ( .A(n2257), .B(n2282), .C(n1559), .Y(n1121) );
  OAI21X1 U541 ( .A(n2257), .B(n2281), .C(n1681), .Y(n1122) );
  OAI21X1 U543 ( .A(n2257), .B(n2280), .C(n1641), .Y(n1123) );
  OAI21X1 U545 ( .A(n2257), .B(n2279), .C(n87), .Y(n1124) );
  OAI21X1 U547 ( .A(n2257), .B(n2278), .C(n41), .Y(n1125) );
  OAI21X1 U549 ( .A(n2257), .B(n2277), .C(n139), .Y(n1126) );
  OAI21X1 U551 ( .A(n2257), .B(n2276), .C(n113), .Y(n1127) );
  OAI21X1 U553 ( .A(n2257), .B(n2275), .C(n1443), .Y(n1128) );
  OAI21X1 U555 ( .A(n2257), .B(n2274), .C(n294), .Y(n1129) );
  OAI21X1 U557 ( .A(n2257), .B(n2273), .C(n199), .Y(n1130) );
  OAI21X1 U559 ( .A(n2257), .B(n2272), .C(n169), .Y(n1131) );
  OAI21X1 U561 ( .A(n1499), .B(n1702), .C(reset), .Y(n560) );
  OAI21X1 U562 ( .A(n2256), .B(n2287), .C(n292), .Y(n1132) );
  OAI21X1 U564 ( .A(n2256), .B(n2286), .C(n1442), .Y(n1133) );
  OAI21X1 U566 ( .A(n2256), .B(n2285), .C(n1479), .Y(n1134) );
  OAI21X1 U568 ( .A(n2256), .B(n2284), .C(n1516), .Y(n1135) );
  OAI21X1 U570 ( .A(n2256), .B(n2283), .C(n1558), .Y(n1136) );
  OAI21X1 U572 ( .A(n2256), .B(n2282), .C(n1600), .Y(n1137) );
  OAI21X1 U574 ( .A(n2256), .B(n2281), .C(n1640), .Y(n1138) );
  OAI21X1 U576 ( .A(n2256), .B(n2280), .C(n1680), .Y(n1139) );
  OAI21X1 U578 ( .A(n2256), .B(n2279), .C(n40), .Y(n1140) );
  OAI21X1 U580 ( .A(n2256), .B(n2278), .C(n86), .Y(n1141) );
  OAI21X1 U582 ( .A(n2256), .B(n2277), .C(n112), .Y(n1142) );
  OAI21X1 U584 ( .A(n2256), .B(n2276), .C(n138), .Y(n1143) );
  OAI21X1 U586 ( .A(n2256), .B(n2275), .C(n290), .Y(n1144) );
  OAI21X1 U588 ( .A(n2256), .B(n2274), .C(n1441), .Y(n1145) );
  OAI21X1 U590 ( .A(n2256), .B(n2273), .C(n168), .Y(n1146) );
  OAI21X1 U592 ( .A(n2256), .B(n2272), .C(n198), .Y(n1147) );
  OAI21X1 U594 ( .A(n1537), .B(n1702), .C(reset), .Y(n577) );
  NAND3X1 U595 ( .A(n852), .B(n2310), .C(wr_ptr[3]), .Y(n458) );
  OAI21X1 U596 ( .A(n2255), .B(n2287), .C(n258), .Y(n1148) );
  OAI21X1 U598 ( .A(n2255), .B(n2286), .C(n227), .Y(n1149) );
  OAI21X1 U600 ( .A(n2255), .B(n2285), .C(n197), .Y(n1150) );
  OAI21X1 U602 ( .A(n2255), .B(n2284), .C(n167), .Y(n1151) );
  OAI21X1 U604 ( .A(n2255), .B(n2283), .C(n137), .Y(n1152) );
  OAI21X1 U606 ( .A(n2255), .B(n2282), .C(n111), .Y(n1153) );
  OAI21X1 U608 ( .A(n2255), .B(n2281), .C(n85), .Y(n1154) );
  OAI21X1 U610 ( .A(n2255), .B(n2280), .C(n39), .Y(n1155) );
  OAI21X1 U612 ( .A(n2255), .B(n2279), .C(n1679), .Y(n1156) );
  OAI21X1 U614 ( .A(n2255), .B(n2278), .C(n1639), .Y(n1157) );
  OAI21X1 U616 ( .A(n2255), .B(n2277), .C(n1599), .Y(n1158) );
  OAI21X1 U618 ( .A(n2255), .B(n2276), .C(n1557), .Y(n1159) );
  OAI21X1 U620 ( .A(n2255), .B(n2275), .C(n257), .Y(n1160) );
  OAI21X1 U622 ( .A(n2255), .B(n2274), .C(n226), .Y(n1161) );
  OAI21X1 U624 ( .A(n2255), .B(n2273), .C(n1515), .Y(n1162) );
  OAI21X1 U626 ( .A(n2255), .B(n2272), .C(n1478), .Y(n1163) );
  OAI21X1 U628 ( .A(n1538), .B(n1661), .C(reset), .Y(n594) );
  OAI21X1 U629 ( .A(n2254), .B(n2287), .C(n225), .Y(n1164) );
  OAI21X1 U631 ( .A(n2254), .B(n2286), .C(n256), .Y(n1165) );
  OAI21X1 U633 ( .A(n2254), .B(n2285), .C(n166), .Y(n1166) );
  OAI21X1 U635 ( .A(n2254), .B(n2284), .C(n196), .Y(n1167) );
  OAI21X1 U637 ( .A(n2254), .B(n2283), .C(n110), .Y(n1168) );
  OAI21X1 U639 ( .A(n2254), .B(n2282), .C(n136), .Y(n1169) );
  OAI21X1 U641 ( .A(n2254), .B(n2281), .C(n38), .Y(n1170) );
  OAI21X1 U643 ( .A(n2254), .B(n2280), .C(n84), .Y(n1171) );
  OAI21X1 U645 ( .A(n2254), .B(n2279), .C(n1638), .Y(n1172) );
  OAI21X1 U647 ( .A(n2254), .B(n2278), .C(n1678), .Y(n1173) );
  OAI21X1 U649 ( .A(n2254), .B(n2277), .C(n1556), .Y(n1174) );
  OAI21X1 U651 ( .A(n2254), .B(n2276), .C(n1598), .Y(n1175) );
  OAI21X1 U653 ( .A(n2254), .B(n2275), .C(n224), .Y(n1176) );
  OAI21X1 U655 ( .A(n2254), .B(n2274), .C(n255), .Y(n1177) );
  OAI21X1 U657 ( .A(n2254), .B(n2273), .C(n1477), .Y(n1178) );
  OAI21X1 U659 ( .A(n2254), .B(n2272), .C(n1514), .Y(n1179) );
  OAI21X1 U661 ( .A(n1500), .B(n1661), .C(reset), .Y(n612) );
  OAI21X1 U662 ( .A(n2253), .B(n2287), .C(n195), .Y(n1180) );
  OAI21X1 U664 ( .A(n2253), .B(n2286), .C(n165), .Y(n1181) );
  OAI21X1 U666 ( .A(n2253), .B(n2285), .C(n254), .Y(n1182) );
  OAI21X1 U668 ( .A(n2253), .B(n2284), .C(n223), .Y(n1183) );
  OAI21X1 U670 ( .A(n2253), .B(n2283), .C(n83), .Y(n1184) );
  OAI21X1 U672 ( .A(n2253), .B(n2282), .C(n37), .Y(n1185) );
  OAI21X1 U674 ( .A(n2253), .B(n2281), .C(n135), .Y(n1186) );
  OAI21X1 U676 ( .A(n2253), .B(n2280), .C(n109), .Y(n1187) );
  OAI21X1 U678 ( .A(n2253), .B(n2279), .C(n1597), .Y(n1188) );
  OAI21X1 U680 ( .A(n2253), .B(n2278), .C(n1555), .Y(n1189) );
  OAI21X1 U682 ( .A(n2253), .B(n2277), .C(n1677), .Y(n1190) );
  OAI21X1 U684 ( .A(n2253), .B(n2276), .C(n1637), .Y(n1191) );
  OAI21X1 U686 ( .A(n2253), .B(n2275), .C(n194), .Y(n1192) );
  OAI21X1 U688 ( .A(n2253), .B(n2274), .C(n164), .Y(n1193) );
  OAI21X1 U690 ( .A(n2253), .B(n2273), .C(n1440), .Y(n1194) );
  OAI21X1 U692 ( .A(n2253), .B(n2272), .C(n288), .Y(n1195) );
  OAI21X1 U694 ( .A(n1462), .B(n1661), .C(reset), .Y(n629) );
  OAI21X1 U695 ( .A(n2252), .B(n2287), .C(n163), .Y(n1196) );
  OAI21X1 U697 ( .A(n2252), .B(n2286), .C(n193), .Y(n1197) );
  OAI21X1 U699 ( .A(n2252), .B(n2285), .C(n222), .Y(n1198) );
  OAI21X1 U701 ( .A(n2252), .B(n2284), .C(n253), .Y(n1199) );
  OAI21X1 U703 ( .A(n2252), .B(n2283), .C(n36), .Y(n1200) );
  OAI21X1 U705 ( .A(n2252), .B(n2282), .C(n82), .Y(n1201) );
  OAI21X1 U707 ( .A(n2252), .B(n2281), .C(n108), .Y(n1202) );
  OAI21X1 U709 ( .A(n2252), .B(n2280), .C(n134), .Y(n1203) );
  OAI21X1 U711 ( .A(n2252), .B(n2279), .C(n1554), .Y(n1204) );
  OAI21X1 U713 ( .A(n2252), .B(n2278), .C(n1596), .Y(n1205) );
  OAI21X1 U715 ( .A(n2252), .B(n2277), .C(n1636), .Y(n1206) );
  OAI21X1 U717 ( .A(n2252), .B(n2276), .C(n1676), .Y(n1207) );
  OAI21X1 U719 ( .A(n2252), .B(n2275), .C(n162), .Y(n1208) );
  OAI21X1 U721 ( .A(n2252), .B(n2274), .C(n192), .Y(n1209) );
  OAI21X1 U723 ( .A(n2252), .B(n2273), .C(n286), .Y(n1210) );
  OAI21X1 U725 ( .A(n2252), .B(n2272), .C(n1439), .Y(n1211) );
  OAI21X1 U727 ( .A(n1424), .B(n1661), .C(reset), .Y(n646) );
  OAI21X1 U728 ( .A(n2251), .B(n2287), .C(n1675), .Y(n1212) );
  OAI21X1 U730 ( .A(n2251), .B(n2286), .C(n1635), .Y(n1213) );
  OAI21X1 U732 ( .A(n2251), .B(n2285), .C(n1595), .Y(n1214) );
  OAI21X1 U734 ( .A(n2251), .B(n2284), .C(n1553), .Y(n1215) );
  OAI21X1 U736 ( .A(n2251), .B(n2283), .C(n1513), .Y(n1216) );
  OAI21X1 U738 ( .A(n2251), .B(n2282), .C(n1476), .Y(n1217) );
  OAI21X1 U740 ( .A(n2251), .B(n2281), .C(n1438), .Y(n1218) );
  OAI21X1 U742 ( .A(n2251), .B(n2280), .C(n284), .Y(n1219) );
  OAI21X1 U744 ( .A(n2251), .B(n2279), .C(n252), .Y(n1220) );
  OAI21X1 U746 ( .A(n2251), .B(n2278), .C(n221), .Y(n1221) );
  OAI21X1 U748 ( .A(n2251), .B(n2277), .C(n191), .Y(n1222) );
  OAI21X1 U750 ( .A(n2251), .B(n2276), .C(n161), .Y(n1223) );
  OAI21X1 U752 ( .A(n2251), .B(n2275), .C(n1674), .Y(n1224) );
  OAI21X1 U754 ( .A(n2251), .B(n2274), .C(n1634), .Y(n1225) );
  OAI21X1 U756 ( .A(n2251), .B(n2273), .C(n133), .Y(n1226) );
  OAI21X1 U758 ( .A(n2251), .B(n2272), .C(n107), .Y(n1227) );
  OAI21X1 U760 ( .A(n1423), .B(n1661), .C(reset), .Y(n663) );
  OAI21X1 U761 ( .A(n2250), .B(n2287), .C(n1633), .Y(n1228) );
  OAI21X1 U763 ( .A(n2250), .B(n2286), .C(n1673), .Y(n1229) );
  OAI21X1 U765 ( .A(n2250), .B(n2285), .C(n1552), .Y(n1230) );
  OAI21X1 U767 ( .A(n2250), .B(n2284), .C(n1594), .Y(n1231) );
  OAI21X1 U769 ( .A(n2250), .B(n2283), .C(n1475), .Y(n1232) );
  OAI21X1 U771 ( .A(n2250), .B(n2282), .C(n1512), .Y(n1233) );
  OAI21X1 U773 ( .A(n2250), .B(n2281), .C(n282), .Y(n1234) );
  OAI21X1 U775 ( .A(n2250), .B(n2280), .C(n1437), .Y(n1235) );
  OAI21X1 U777 ( .A(n2250), .B(n2279), .C(n220), .Y(n1236) );
  OAI21X1 U779 ( .A(n2250), .B(n2278), .C(n251), .Y(n1237) );
  OAI21X1 U781 ( .A(n2250), .B(n2277), .C(n160), .Y(n1238) );
  OAI21X1 U783 ( .A(n2250), .B(n2276), .C(n190), .Y(n1239) );
  OAI21X1 U785 ( .A(n2250), .B(n2275), .C(n1632), .Y(n1240) );
  OAI21X1 U787 ( .A(n2250), .B(n2274), .C(n1672), .Y(n1241) );
  OAI21X1 U789 ( .A(n2250), .B(n2273), .C(n106), .Y(n1242) );
  OAI21X1 U791 ( .A(n2250), .B(n2272), .C(n132), .Y(n1243) );
  OAI21X1 U793 ( .A(n1461), .B(n1661), .C(reset), .Y(n680) );
  OAI21X1 U794 ( .A(n2249), .B(n2287), .C(n1593), .Y(n1244) );
  OAI21X1 U796 ( .A(n2249), .B(n2286), .C(n1551), .Y(n1245) );
  OAI21X1 U798 ( .A(n2249), .B(n2285), .C(n1671), .Y(n1246) );
  OAI21X1 U800 ( .A(n2249), .B(n2284), .C(n1631), .Y(n1247) );
  OAI21X1 U802 ( .A(n2249), .B(n2283), .C(n1436), .Y(n1248) );
  OAI21X1 U804 ( .A(n2249), .B(n2282), .C(n280), .Y(n1249) );
  OAI21X1 U806 ( .A(n2249), .B(n2281), .C(n1511), .Y(n1250) );
  OAI21X1 U808 ( .A(n2249), .B(n2280), .C(n1474), .Y(n1251) );
  OAI21X1 U810 ( .A(n2249), .B(n2279), .C(n189), .Y(n1252) );
  OAI21X1 U812 ( .A(n2249), .B(n2278), .C(n159), .Y(n1253) );
  OAI21X1 U814 ( .A(n2249), .B(n2277), .C(n250), .Y(n1254) );
  OAI21X1 U816 ( .A(n2249), .B(n2276), .C(n219), .Y(n1255) );
  OAI21X1 U818 ( .A(n2249), .B(n2275), .C(n1592), .Y(n1256) );
  OAI21X1 U820 ( .A(n2249), .B(n2274), .C(n1550), .Y(n1257) );
  OAI21X1 U822 ( .A(n2249), .B(n2273), .C(n81), .Y(n1258) );
  OAI21X1 U824 ( .A(n2249), .B(n2272), .C(n35), .Y(n1259) );
  OAI21X1 U826 ( .A(n1499), .B(n1661), .C(reset), .Y(n697) );
  OAI21X1 U827 ( .A(n2248), .B(n2287), .C(n1549), .Y(n1260) );
  OAI21X1 U829 ( .A(n2248), .B(n2286), .C(n1591), .Y(n1261) );
  OAI21X1 U831 ( .A(n2248), .B(n2285), .C(n1630), .Y(n1262) );
  OAI21X1 U833 ( .A(n2248), .B(n2284), .C(n1670), .Y(n1263) );
  OAI21X1 U835 ( .A(n2248), .B(n2283), .C(n279), .Y(n1264) );
  OAI21X1 U837 ( .A(n2248), .B(n2282), .C(n1435), .Y(n1265) );
  OAI21X1 U839 ( .A(n2248), .B(n2281), .C(n1473), .Y(n1266) );
  OAI21X1 U841 ( .A(n2248), .B(n2280), .C(n1510), .Y(n1267) );
  OAI21X1 U843 ( .A(n2248), .B(n2279), .C(n158), .Y(n1268) );
  OAI21X1 U845 ( .A(n2248), .B(n2278), .C(n188), .Y(n1269) );
  OAI21X1 U847 ( .A(n2248), .B(n2277), .C(n218), .Y(n1270) );
  OAI21X1 U849 ( .A(n2248), .B(n2276), .C(n249), .Y(n1271) );
  OAI21X1 U851 ( .A(n2248), .B(n2275), .C(n1548), .Y(n1272) );
  OAI21X1 U853 ( .A(n2248), .B(n2274), .C(n1590), .Y(n1273) );
  OAI21X1 U855 ( .A(n2248), .B(n2273), .C(n34), .Y(n1274) );
  OAI21X1 U857 ( .A(n2248), .B(n2272), .C(n80), .Y(n1275) );
  OAI21X1 U859 ( .A(n1537), .B(n1661), .C(reset), .Y(n714) );
  NAND3X1 U860 ( .A(n852), .B(n2313), .C(wr_ptr[4]), .Y(n595) );
  OAI21X1 U861 ( .A(n2247), .B(n2287), .C(n1509), .Y(n1276) );
  OAI21X1 U863 ( .A(n2247), .B(n2286), .C(n1472), .Y(n1277) );
  OAI21X1 U865 ( .A(n2247), .B(n2285), .C(n1434), .Y(n1278) );
  OAI21X1 U867 ( .A(n2247), .B(n2284), .C(n278), .Y(n1279) );
  OAI21X1 U869 ( .A(n2247), .B(n2283), .C(n1669), .Y(n1280) );
  OAI21X1 U871 ( .A(n2247), .B(n2282), .C(n1629), .Y(n1281) );
  OAI21X1 U873 ( .A(n2247), .B(n2281), .C(n1589), .Y(n1282) );
  OAI21X1 U875 ( .A(n2247), .B(n2280), .C(n1547), .Y(n1283) );
  OAI21X1 U877 ( .A(n2247), .B(n2279), .C(n131), .Y(n1284) );
  OAI21X1 U879 ( .A(n2247), .B(n2278), .C(n105), .Y(n1285) );
  OAI21X1 U881 ( .A(n2247), .B(n2277), .C(n79), .Y(n1286) );
  OAI21X1 U883 ( .A(n2247), .B(n2276), .C(n33), .Y(n1287) );
  OAI21X1 U885 ( .A(n2247), .B(n2275), .C(n1508), .Y(n1288) );
  OAI21X1 U887 ( .A(n2247), .B(n2274), .C(n1471), .Y(n1289) );
  OAI21X1 U889 ( .A(n2247), .B(n2273), .C(n248), .Y(n1290) );
  OAI21X1 U891 ( .A(n2247), .B(n2272), .C(n217), .Y(n1291) );
  OAI21X1 U893 ( .A(n1538), .B(n1620), .C(reset), .Y(n731) );
  NAND3X1 U894 ( .A(n2311), .B(n2312), .C(n2309), .Y(n314) );
  OAI21X1 U895 ( .A(n2246), .B(n2287), .C(n1470), .Y(n1292) );
  OAI21X1 U897 ( .A(n2246), .B(n2286), .C(n1507), .Y(n1293) );
  OAI21X1 U899 ( .A(n2246), .B(n2285), .C(n277), .Y(n1294) );
  OAI21X1 U901 ( .A(n2246), .B(n2284), .C(n1433), .Y(n1295) );
  OAI21X1 U903 ( .A(n2246), .B(n2283), .C(n1628), .Y(n1296) );
  OAI21X1 U905 ( .A(n2246), .B(n2282), .C(n1668), .Y(n1297) );
  OAI21X1 U907 ( .A(n2246), .B(n2281), .C(n1546), .Y(n1298) );
  OAI21X1 U909 ( .A(n2246), .B(n2280), .C(n1588), .Y(n1299) );
  OAI21X1 U911 ( .A(n2246), .B(n2279), .C(n104), .Y(n1300) );
  OAI21X1 U913 ( .A(n2246), .B(n2278), .C(n130), .Y(n1301) );
  OAI21X1 U915 ( .A(n2246), .B(n2277), .C(n32), .Y(n1302) );
  OAI21X1 U917 ( .A(n2246), .B(n2276), .C(n78), .Y(n1303) );
  OAI21X1 U919 ( .A(n2246), .B(n2275), .C(n1469), .Y(n1304) );
  OAI21X1 U921 ( .A(n2246), .B(n2274), .C(n1506), .Y(n1305) );
  OAI21X1 U923 ( .A(n2246), .B(n2273), .C(n216), .Y(n1306) );
  OAI21X1 U925 ( .A(n2246), .B(n2272), .C(n247), .Y(n1307) );
  OAI21X1 U927 ( .A(n1500), .B(n1620), .C(reset), .Y(n749) );
  NAND3X1 U928 ( .A(n2311), .B(n2312), .C(wr_ptr[0]), .Y(n332) );
  OAI21X1 U929 ( .A(n2245), .B(n2287), .C(n1432), .Y(n1308) );
  OAI21X1 U931 ( .A(n2245), .B(n2286), .C(n276), .Y(n1309) );
  OAI21X1 U933 ( .A(n2245), .B(n2285), .C(n1505), .Y(n1310) );
  OAI21X1 U935 ( .A(n2245), .B(n2284), .C(n1468), .Y(n1311) );
  OAI21X1 U937 ( .A(n2245), .B(n2283), .C(n1587), .Y(n1312) );
  OAI21X1 U939 ( .A(n2245), .B(n2282), .C(n1545), .Y(n1313) );
  OAI21X1 U941 ( .A(n2245), .B(n2281), .C(n1667), .Y(n1314) );
  OAI21X1 U943 ( .A(n2245), .B(n2280), .C(n1627), .Y(n1315) );
  OAI21X1 U945 ( .A(n2245), .B(n2279), .C(n77), .Y(n1316) );
  OAI21X1 U947 ( .A(n2245), .B(n2278), .C(n31), .Y(n1317) );
  OAI21X1 U949 ( .A(n2245), .B(n2277), .C(n129), .Y(n1318) );
  OAI21X1 U951 ( .A(n2245), .B(n2276), .C(n103), .Y(n1319) );
  OAI21X1 U953 ( .A(n2245), .B(n2275), .C(n1431), .Y(n1320) );
  OAI21X1 U955 ( .A(n2245), .B(n2274), .C(n275), .Y(n1321) );
  OAI21X1 U957 ( .A(n2245), .B(n2273), .C(n187), .Y(n1322) );
  OAI21X1 U959 ( .A(n2245), .B(n2272), .C(n157), .Y(n1323) );
  OAI21X1 U961 ( .A(n1462), .B(n1620), .C(reset), .Y(n766) );
  NAND3X1 U962 ( .A(n2309), .B(n2312), .C(wr_ptr[1]), .Y(n350) );
  OAI21X1 U963 ( .A(n2244), .B(n2287), .C(n274), .Y(n1324) );
  OAI21X1 U965 ( .A(n2244), .B(n2286), .C(n1430), .Y(n1325) );
  OAI21X1 U967 ( .A(n2244), .B(n2285), .C(n1467), .Y(n1326) );
  OAI21X1 U969 ( .A(n2244), .B(n2284), .C(n1504), .Y(n1327) );
  OAI21X1 U971 ( .A(n2244), .B(n2283), .C(n1544), .Y(n1328) );
  OAI21X1 U973 ( .A(n2244), .B(n2282), .C(n1586), .Y(n1329) );
  OAI21X1 U975 ( .A(n2244), .B(n2281), .C(n1626), .Y(n1330) );
  OAI21X1 U977 ( .A(n2244), .B(n2280), .C(n1666), .Y(n1331) );
  OAI21X1 U979 ( .A(n2244), .B(n2279), .C(n30), .Y(n1332) );
  OAI21X1 U981 ( .A(n2244), .B(n2278), .C(n72), .Y(n1333) );
  OAI21X1 U983 ( .A(n2244), .B(n2277), .C(n102), .Y(n1334) );
  OAI21X1 U985 ( .A(n2244), .B(n2276), .C(n128), .Y(n1335) );
  OAI21X1 U987 ( .A(n2244), .B(n2275), .C(n273), .Y(n1336) );
  OAI21X1 U989 ( .A(n2244), .B(n2274), .C(n1429), .Y(n1337) );
  OAI21X1 U991 ( .A(n2244), .B(n2273), .C(n156), .Y(n1338) );
  OAI21X1 U993 ( .A(n2244), .B(n2272), .C(n186), .Y(n1339) );
  OAI21X1 U995 ( .A(n1424), .B(n1620), .C(reset), .Y(n783) );
  NAND3X1 U996 ( .A(wr_ptr[0]), .B(n2312), .C(wr_ptr[1]), .Y(n368) );
  OAI21X1 U997 ( .A(n2243), .B(n2287), .C(n246), .Y(n1340) );
  OAI21X1 U999 ( .A(n2243), .B(n2286), .C(n215), .Y(n1341) );
  OAI21X1 U1001 ( .A(n2243), .B(n2285), .C(n185), .Y(n1342) );
  OAI21X1 U1003 ( .A(n2243), .B(n2284), .C(n155), .Y(n1343) );
  OAI21X1 U1005 ( .A(n2243), .B(n2283), .C(n127), .Y(n1344) );
  OAI21X1 U1007 ( .A(n2243), .B(n2282), .C(n101), .Y(n1345) );
  OAI21X1 U1009 ( .A(n2243), .B(n2281), .C(n55), .Y(n1346) );
  OAI21X1 U1011 ( .A(n2243), .B(n2280), .C(n29), .Y(n1347) );
  OAI21X1 U1013 ( .A(n2243), .B(n2279), .C(n1665), .Y(n1348) );
  OAI21X1 U1015 ( .A(n2243), .B(n2278), .C(n1625), .Y(n1349) );
  OAI21X1 U1017 ( .A(n2243), .B(n2277), .C(n1585), .Y(n1350) );
  OAI21X1 U1019 ( .A(n2243), .B(n2276), .C(n1543), .Y(n1351) );
  OAI21X1 U1021 ( .A(n2243), .B(n2275), .C(n245), .Y(n1352) );
  OAI21X1 U1023 ( .A(n2243), .B(n2274), .C(n214), .Y(n1353) );
  OAI21X1 U1025 ( .A(n2243), .B(n2273), .C(n1503), .Y(n1354) );
  OAI21X1 U1027 ( .A(n2243), .B(n2272), .C(n1466), .Y(n1355) );
  OAI21X1 U1029 ( .A(n1423), .B(n1620), .C(reset), .Y(n800) );
  NAND3X1 U1030 ( .A(n2309), .B(n2311), .C(wr_ptr[2]), .Y(n386) );
  OAI21X1 U1031 ( .A(n2242), .B(n2287), .C(n213), .Y(n1356) );
  OAI21X1 U1033 ( .A(n2242), .B(n2286), .C(n244), .Y(n1357) );
  OAI21X1 U1035 ( .A(n2242), .B(n2285), .C(n154), .Y(n1358) );
  OAI21X1 U1037 ( .A(n2242), .B(n2284), .C(n184), .Y(n1359) );
  OAI21X1 U1039 ( .A(n2242), .B(n2283), .C(n100), .Y(n1360) );
  OAI21X1 U1041 ( .A(n2242), .B(n2282), .C(n126), .Y(n1361) );
  OAI21X1 U1043 ( .A(n2242), .B(n2281), .C(n28), .Y(n1362) );
  OAI21X1 U1045 ( .A(n2242), .B(n2280), .C(n54), .Y(n1363) );
  OAI21X1 U1047 ( .A(n2242), .B(n2279), .C(n1624), .Y(n1364) );
  OAI21X1 U1049 ( .A(n2242), .B(n2278), .C(n1664), .Y(n1365) );
  OAI21X1 U1051 ( .A(n2242), .B(n2277), .C(n1542), .Y(n1366) );
  OAI21X1 U1053 ( .A(n2242), .B(n2276), .C(n1584), .Y(n1367) );
  OAI21X1 U1055 ( .A(n2242), .B(n2275), .C(n212), .Y(n1368) );
  OAI21X1 U1057 ( .A(n2242), .B(n2274), .C(n243), .Y(n1369) );
  OAI21X1 U1059 ( .A(n2242), .B(n2273), .C(n1465), .Y(n1370) );
  OAI21X1 U1061 ( .A(n2242), .B(n2272), .C(n1502), .Y(n1371) );
  OAI21X1 U1063 ( .A(n1461), .B(n1620), .C(reset), .Y(n817) );
  NAND3X1 U1064 ( .A(wr_ptr[0]), .B(n2311), .C(wr_ptr[2]), .Y(n404) );
  OAI21X1 U1065 ( .A(n2241), .B(n2287), .C(n183), .Y(n1372) );
  OAI21X1 U1067 ( .A(n2241), .B(n2286), .C(n153), .Y(n1373) );
  OAI21X1 U1069 ( .A(n2241), .B(n2285), .C(n242), .Y(n1374) );
  OAI21X1 U1071 ( .A(n2241), .B(n2284), .C(n211), .Y(n1375) );
  OAI21X1 U1073 ( .A(n2241), .B(n2283), .C(n53), .Y(n1376) );
  OAI21X1 U1075 ( .A(n2241), .B(n2282), .C(n27), .Y(n1377) );
  OAI21X1 U1077 ( .A(n2241), .B(n2281), .C(n125), .Y(n1378) );
  OAI21X1 U1079 ( .A(n2241), .B(n2280), .C(n99), .Y(n1379) );
  OAI21X1 U1081 ( .A(n2241), .B(n2279), .C(n1583), .Y(n1380) );
  OAI21X1 U1083 ( .A(n2241), .B(n2278), .C(n1541), .Y(n1381) );
  OAI21X1 U1085 ( .A(n2241), .B(n2277), .C(n1663), .Y(n1382) );
  OAI21X1 U1087 ( .A(n2241), .B(n2276), .C(n1623), .Y(n1383) );
  OAI21X1 U1089 ( .A(n2241), .B(n2275), .C(n182), .Y(n1384) );
  OAI21X1 U1091 ( .A(n2241), .B(n2274), .C(n152), .Y(n1385) );
  OAI21X1 U1093 ( .A(n2241), .B(n2273), .C(n1428), .Y(n1386) );
  OAI21X1 U1095 ( .A(n2241), .B(n2272), .C(n272), .Y(n1387) );
  OAI21X1 U1097 ( .A(n1499), .B(n1620), .C(reset), .Y(n834) );
  NAND3X1 U1098 ( .A(wr_ptr[1]), .B(n2309), .C(wr_ptr[2]), .Y(n422) );
  OAI21X1 U1099 ( .A(n2240), .B(n2287), .C(n151), .Y(n1388) );
  OAI21X1 U1102 ( .A(n2240), .B(n2286), .C(n181), .Y(n1389) );
  OAI21X1 U1105 ( .A(n2240), .B(n2285), .C(n210), .Y(n1390) );
  OAI21X1 U1108 ( .A(n2240), .B(n2284), .C(n241), .Y(n1391) );
  OAI21X1 U1111 ( .A(n2240), .B(n2283), .C(n26), .Y(n1392) );
  OAI21X1 U1114 ( .A(n2240), .B(n2282), .C(n52), .Y(n1393) );
  OAI21X1 U1117 ( .A(n2240), .B(n2281), .C(n98), .Y(n1394) );
  OAI21X1 U1120 ( .A(n2240), .B(n2280), .C(n124), .Y(n1395) );
  OAI21X1 U1123 ( .A(n2240), .B(n2279), .C(n1540), .Y(n1396) );
  OAI21X1 U1126 ( .A(n2240), .B(n2278), .C(n1582), .Y(n1397) );
  OAI21X1 U1129 ( .A(n2240), .B(n2277), .C(n1622), .Y(n1398) );
  OAI21X1 U1132 ( .A(n2240), .B(n2276), .C(n1662), .Y(n1399) );
  OAI21X1 U1135 ( .A(n2240), .B(n2275), .C(n150), .Y(n1400) );
  OAI21X1 U1138 ( .A(n2240), .B(n2274), .C(n180), .Y(n1401) );
  OAI21X1 U1141 ( .A(n2240), .B(n2273), .C(n271), .Y(n1402) );
  OAI21X1 U1144 ( .A(n2240), .B(n2272), .C(n1427), .Y(n1403) );
  OAI21X1 U1147 ( .A(n1537), .B(n1620), .C(reset), .Y(n851) );
  NAND3X1 U1148 ( .A(wr_ptr[3]), .B(n852), .C(wr_ptr[4]), .Y(n732) );
  NAND3X1 U1149 ( .A(wr_ptr[1]), .B(wr_ptr[0]), .C(wr_ptr[2]), .Y(n440) );
  OAI21X1 U1150 ( .A(n2313), .B(n1660), .C(n1464), .Y(n1404) );
  OAI21X1 U1152 ( .A(n2312), .B(n1660), .C(n1581), .Y(n1405) );
  OAI21X1 U1154 ( .A(n2311), .B(n1660), .C(n240), .Y(n1406) );
  OAI21X1 U1156 ( .A(n2310), .B(n1660), .C(n1426), .Y(n1407) );
  OAI21X1 U1158 ( .A(n2288), .B(n1703), .C(n1621), .Y(n1408) );
  OAI21X1 U1160 ( .A(n2289), .B(n1703), .C(n1580), .Y(n1409) );
  OAI21X1 U1162 ( .A(n2290), .B(n1703), .C(n1501), .Y(n1410) );
  OAI21X1 U1164 ( .A(n2291), .B(n1703), .C(n1463), .Y(n1411) );
  OAI21X1 U1166 ( .A(n2292), .B(n1703), .C(n1425), .Y(n1412) );
  AOI22X1 U1168 ( .A(n56), .B(n861), .C(data_out[15]), .D(n859), .Y(n866) );
  AOI22X1 U1169 ( .A(n57), .B(n2239), .C(data_out[14]), .D(n859), .Y(n867) );
  AOI22X1 U1170 ( .A(n58), .B(n2238), .C(data_out[13]), .D(n859), .Y(n868) );
  AOI22X1 U1171 ( .A(n59), .B(n861), .C(data_out[12]), .D(n859), .Y(n869) );
  AOI22X1 U1172 ( .A(n60), .B(n2239), .C(data_out[11]), .D(n859), .Y(n870) );
  AOI22X1 U1173 ( .A(n61), .B(n2238), .C(data_out[10]), .D(n859), .Y(n871) );
  AOI22X1 U1174 ( .A(n62), .B(n861), .C(data_out[9]), .D(n859), .Y(n872) );
  AOI22X1 U1175 ( .A(n63), .B(n2239), .C(data_out[8]), .D(n859), .Y(n873) );
  AOI22X1 U1176 ( .A(n64), .B(n2238), .C(data_out[7]), .D(n859), .Y(n874) );
  AOI22X1 U1177 ( .A(n65), .B(n861), .C(data_out[6]), .D(n859), .Y(n875) );
  AOI22X1 U1178 ( .A(n66), .B(n2239), .C(data_out[5]), .D(n859), .Y(n876) );
  AOI22X1 U1179 ( .A(n67), .B(n2238), .C(data_out[4]), .D(n859), .Y(n877) );
  AOI22X1 U1180 ( .A(n68), .B(n861), .C(data_out[3]), .D(n859), .Y(n878) );
  AOI22X1 U1181 ( .A(n69), .B(n2239), .C(data_out[2]), .D(n859), .Y(n879) );
  AOI22X1 U1182 ( .A(n70), .B(n2238), .C(data_out[1]), .D(n859), .Y(n880) );
  AOI22X1 U1183 ( .A(n71), .B(n861), .C(data_out[0]), .D(n859), .Y(n881) );
  OAI21X1 U1186 ( .A(n2309), .B(n1660), .C(n1539), .Y(n1413) );
  NAND3X1 U1190 ( .A(n1701), .B(fillcount[5]), .C(n885), .Y(n2315) );
  NOR3X1 U1191 ( .A(fillcount[2]), .B(fillcount[4]), .C(fillcount[3]), .Y(n885) );
  NAND3X1 U1193 ( .A(n886), .B(n887), .C(n888), .Y(n2314) );
  NOR3X1 U1194 ( .A(n889), .B(n890), .C(n891), .Y(n888) );
  XNOR2X1 U1195 ( .A(n2312), .B(n14), .Y(n891) );
  XNOR2X1 U1196 ( .A(n2313), .B(n15), .Y(n890) );
  XNOR2X1 U1197 ( .A(n2309), .B(n12), .Y(n889) );
  XNOR2X1 U1198 ( .A(n13), .B(wr_ptr[1]), .Y(n887) );
  XNOR2X1 U1199 ( .A(n16), .B(wr_ptr[4]), .Y(n886) );
  HAX1 add_57_U1_1_1 ( .A(n13), .B(n12), .YC(add_57_carry[2]), .YS(n73) );
  HAX1 add_57_U1_1_2 ( .A(n14), .B(add_57_carry[2]), .YC(add_57_carry[3]), 
        .YS(n74) );
  HAX1 add_57_U1_1_3 ( .A(n15), .B(add_57_carry[3]), .YC(add_57_carry[4]), 
        .YS(n75) );
  HAX1 add_51_U1_1_1 ( .A(wr_ptr[1]), .B(wr_ptr[0]), .YC(add_51_carry[2]), 
        .YS(n20) );
  HAX1 add_51_U1_1_2 ( .A(wr_ptr[2]), .B(add_51_carry[2]), .YC(add_51_carry[3]), .YS(n21) );
  HAX1 add_51_U1_1_3 ( .A(wr_ptr[3]), .B(add_51_carry[3]), .YC(add_51_carry[4]), .YS(n22) );
  FAX1 sub_93_U2_1 ( .A(wr_ptr[1]), .B(n2290), .C(sub_93_carry[1]), .YC(
        sub_93_carry[2]), .YS(fillcount[1]) );
  FAX1 sub_93_U2_2 ( .A(wr_ptr[2]), .B(n2289), .C(sub_93_carry[2]), .YC(
        sub_93_carry[3]), .YS(fillcount[2]) );
  FAX1 sub_93_U2_3 ( .A(wr_ptr[3]), .B(n2288), .C(sub_93_carry[3]), .YC(
        sub_93_carry[4]), .YS(fillcount[3]) );
  FAX1 sub_93_U2_4 ( .A(wr_ptr[4]), .B(n2292), .C(sub_93_carry[4]), .YC(
        sub_93_carry[5]), .YS(fillcount[4]) );
  AND2X1 U3 ( .A(get), .B(empty_bar), .Y(n882) );
  AND2X1 U4 ( .A(reset), .B(n1536), .Y(n853) );
  AND2X1 U5 ( .A(reset), .B(n1704), .Y(n859) );
  BUFX2 U6 ( .A(n881), .Y(n1) );
  BUFX2 U7 ( .A(n880), .Y(n2) );
  BUFX2 U8 ( .A(n879), .Y(n3) );
  BUFX2 U9 ( .A(n878), .Y(n4) );
  BUFX2 U10 ( .A(n877), .Y(n5) );
  BUFX2 U11 ( .A(n876), .Y(n6) );
  BUFX2 U12 ( .A(n875), .Y(n7) );
  BUFX2 U13 ( .A(n874), .Y(n8) );
  BUFX2 U14 ( .A(n873), .Y(n9) );
  BUFX2 U15 ( .A(n872), .Y(n10) );
  BUFX2 U16 ( .A(n871), .Y(n11) );
  BUFX2 U17 ( .A(n870), .Y(n17) );
  BUFX2 U18 ( .A(n869), .Y(n18) );
  BUFX2 U19 ( .A(n868), .Y(n19) );
  BUFX2 U20 ( .A(n867), .Y(n24) );
  BUFX2 U21 ( .A(n866), .Y(n25) );
  AND2X1 U22 ( .A(mem[500]), .B(n2240), .Y(n839) );
  INVX1 U23 ( .A(n839), .Y(n26) );
  AND2X1 U24 ( .A(mem[485]), .B(n2241), .Y(n823) );
  INVX1 U25 ( .A(n823), .Y(n27) );
  AND2X1 U26 ( .A(mem[470]), .B(n2242), .Y(n807) );
  INVX1 U27 ( .A(n807), .Y(n28) );
  AND2X1 U28 ( .A(mem[455]), .B(n2243), .Y(n791) );
  INVX1 U29 ( .A(n791), .Y(n29) );
  AND2X1 U30 ( .A(mem[440]), .B(n2244), .Y(n775) );
  INVX1 U31 ( .A(n775), .Y(n30) );
  AND2X1 U32 ( .A(mem[425]), .B(n2245), .Y(n759) );
  INVX1 U33 ( .A(n759), .Y(n31) );
  AND2X1 U34 ( .A(mem[410]), .B(n2246), .Y(n743) );
  INVX1 U35 ( .A(n743), .Y(n32) );
  AND2X1 U36 ( .A(mem[395]), .B(n2247), .Y(n726) );
  INVX1 U37 ( .A(n726), .Y(n33) );
  AND2X1 U38 ( .A(mem[382]), .B(n2248), .Y(n712) );
  INVX1 U39 ( .A(n712), .Y(n34) );
  AND2X1 U40 ( .A(mem[367]), .B(n2249), .Y(n696) );
  INVX1 U41 ( .A(n696), .Y(n35) );
  AND2X1 U42 ( .A(mem[308]), .B(n2252), .Y(n634) );
  INVX1 U43 ( .A(n634), .Y(n36) );
  AND2X1 U44 ( .A(mem[293]), .B(n2253), .Y(n618) );
  INVX1 U45 ( .A(n618), .Y(n37) );
  AND2X1 U46 ( .A(mem[278]), .B(n2254), .Y(n602) );
  INVX1 U47 ( .A(n602), .Y(n38) );
  AND2X1 U48 ( .A(mem[263]), .B(n2255), .Y(n585) );
  INVX1 U49 ( .A(n585), .Y(n39) );
  AND2X1 U50 ( .A(mem[248]), .B(n2256), .Y(n569) );
  INVX1 U51 ( .A(n569), .Y(n40) );
  AND2X1 U52 ( .A(mem[233]), .B(n2257), .Y(n553) );
  INVX1 U53 ( .A(n553), .Y(n41) );
  AND2X1 U54 ( .A(mem[218]), .B(n2258), .Y(n537) );
  INVX1 U55 ( .A(n537), .Y(n42) );
  AND2X1 U56 ( .A(mem[203]), .B(n2259), .Y(n521) );
  INVX1 U57 ( .A(n521), .Y(n43) );
  AND2X1 U58 ( .A(mem[190]), .B(n2260), .Y(n507) );
  INVX1 U59 ( .A(n507), .Y(n44) );
  AND2X1 U60 ( .A(mem[175]), .B(n2261), .Y(n491) );
  INVX1 U61 ( .A(n491), .Y(n45) );
  AND2X1 U62 ( .A(mem[120]), .B(n2264), .Y(n431) );
  INVX1 U63 ( .A(n431), .Y(n46) );
  AND2X1 U64 ( .A(mem[105]), .B(n2265), .Y(n414) );
  INVX1 U65 ( .A(n414), .Y(n47) );
  AND2X1 U67 ( .A(mem[90]), .B(n2266), .Y(n397) );
  INVX1 U69 ( .A(n397), .Y(n48) );
  AND2X1 U71 ( .A(mem[75]), .B(n2267), .Y(n380) );
  INVX1 U73 ( .A(n380), .Y(n49) );
  AND2X1 U75 ( .A(mem[62]), .B(n2268), .Y(n365) );
  INVX1 U77 ( .A(n365), .Y(n50) );
  AND2X1 U79 ( .A(mem[47]), .B(n2269), .Y(n348) );
  INVX1 U81 ( .A(n348), .Y(n51) );
  AND2X1 U83 ( .A(mem[501]), .B(n2240), .Y(n840) );
  INVX1 U85 ( .A(n840), .Y(n52) );
  AND2X1 U87 ( .A(mem[484]), .B(n2241), .Y(n822) );
  INVX1 U89 ( .A(n822), .Y(n53) );
  AND2X1 U91 ( .A(mem[471]), .B(n2242), .Y(n808) );
  INVX1 U93 ( .A(n808), .Y(n54) );
  AND2X1 U95 ( .A(mem[454]), .B(n2243), .Y(n790) );
  INVX1 U97 ( .A(n790), .Y(n55) );
  AND2X1 U100 ( .A(mem[441]), .B(n2244), .Y(n776) );
  INVX1 U102 ( .A(n776), .Y(n72) );
  AND2X1 U104 ( .A(mem[424]), .B(n2245), .Y(n758) );
  INVX1 U106 ( .A(n758), .Y(n77) );
  AND2X1 U108 ( .A(mem[411]), .B(n2246), .Y(n744) );
  INVX1 U110 ( .A(n744), .Y(n78) );
  AND2X1 U112 ( .A(mem[394]), .B(n2247), .Y(n725) );
  INVX1 U114 ( .A(n725), .Y(n79) );
  AND2X1 U116 ( .A(mem[383]), .B(n2248), .Y(n713) );
  INVX1 U118 ( .A(n713), .Y(n80) );
  AND2X1 U120 ( .A(mem[366]), .B(n2249), .Y(n695) );
  INVX1 U122 ( .A(n695), .Y(n81) );
  AND2X1 U124 ( .A(mem[309]), .B(n2252), .Y(n635) );
  INVX1 U126 ( .A(n635), .Y(n82) );
  AND2X1 U128 ( .A(mem[292]), .B(n2253), .Y(n617) );
  INVX1 U130 ( .A(n617), .Y(n83) );
  AND2X1 U133 ( .A(mem[279]), .B(n2254), .Y(n603) );
  INVX1 U135 ( .A(n603), .Y(n84) );
  AND2X1 U137 ( .A(mem[262]), .B(n2255), .Y(n584) );
  INVX1 U139 ( .A(n584), .Y(n85) );
  AND2X1 U141 ( .A(mem[249]), .B(n2256), .Y(n570) );
  INVX1 U143 ( .A(n570), .Y(n86) );
  AND2X1 U145 ( .A(mem[232]), .B(n2257), .Y(n552) );
  INVX1 U147 ( .A(n552), .Y(n87) );
  AND2X1 U149 ( .A(mem[219]), .B(n2258), .Y(n538) );
  INVX1 U151 ( .A(n538), .Y(n88) );
  AND2X1 U153 ( .A(mem[202]), .B(n2259), .Y(n520) );
  INVX1 U155 ( .A(n520), .Y(n89) );
  AND2X1 U157 ( .A(mem[191]), .B(n2260), .Y(n508) );
  INVX1 U159 ( .A(n508), .Y(n90) );
  AND2X1 U161 ( .A(mem[174]), .B(n2261), .Y(n490) );
  INVX1 U163 ( .A(n490), .Y(n91) );
  AND2X1 U166 ( .A(mem[121]), .B(n2264), .Y(n432) );
  INVX1 U168 ( .A(n432), .Y(n92) );
  AND2X1 U170 ( .A(mem[104]), .B(n2265), .Y(n413) );
  INVX1 U172 ( .A(n413), .Y(n93) );
  AND2X1 U174 ( .A(mem[91]), .B(n2266), .Y(n398) );
  INVX1 U176 ( .A(n398), .Y(n94) );
  AND2X1 U178 ( .A(mem[74]), .B(n2267), .Y(n379) );
  INVX1 U180 ( .A(n379), .Y(n95) );
  AND2X1 U182 ( .A(mem[63]), .B(n2268), .Y(n366) );
  INVX1 U184 ( .A(n366), .Y(n96) );
  AND2X1 U186 ( .A(mem[46]), .B(n2269), .Y(n347) );
  INVX1 U188 ( .A(n347), .Y(n97) );
  AND2X1 U190 ( .A(mem[502]), .B(n2240), .Y(n841) );
  INVX1 U192 ( .A(n841), .Y(n98) );
  AND2X1 U194 ( .A(mem[487]), .B(n2241), .Y(n825) );
  INVX1 U196 ( .A(n825), .Y(n99) );
  AND2X1 U199 ( .A(mem[468]), .B(n2242), .Y(n805) );
  INVX1 U201 ( .A(n805), .Y(n100) );
  AND2X1 U203 ( .A(mem[453]), .B(n2243), .Y(n789) );
  INVX1 U205 ( .A(n789), .Y(n101) );
  AND2X1 U207 ( .A(mem[442]), .B(n2244), .Y(n777) );
  INVX1 U209 ( .A(n777), .Y(n102) );
  AND2X1 U211 ( .A(mem[427]), .B(n2245), .Y(n761) );
  INVX1 U213 ( .A(n761), .Y(n103) );
  AND2X1 U215 ( .A(mem[408]), .B(n2246), .Y(n741) );
  INVX1 U217 ( .A(n741), .Y(n104) );
  AND2X1 U219 ( .A(mem[393]), .B(n2247), .Y(n724) );
  INVX1 U221 ( .A(n724), .Y(n105) );
  AND2X1 U223 ( .A(mem[350]), .B(n2250), .Y(n678) );
  INVX1 U225 ( .A(n678), .Y(n106) );
  AND2X1 U227 ( .A(mem[335]), .B(n2251), .Y(n662) );
  INVX1 U229 ( .A(n662), .Y(n107) );
  AND2X1 U232 ( .A(mem[310]), .B(n2252), .Y(n636) );
  INVX1 U234 ( .A(n636), .Y(n108) );
  AND2X1 U236 ( .A(mem[295]), .B(n2253), .Y(n620) );
  INVX1 U238 ( .A(n620), .Y(n109) );
  AND2X1 U240 ( .A(mem[276]), .B(n2254), .Y(n600) );
  INVX1 U242 ( .A(n600), .Y(n110) );
  AND2X1 U244 ( .A(mem[261]), .B(n2255), .Y(n583) );
  INVX1 U246 ( .A(n583), .Y(n111) );
  AND2X1 U248 ( .A(mem[250]), .B(n2256), .Y(n571) );
  INVX1 U250 ( .A(n571), .Y(n112) );
  AND2X1 U252 ( .A(mem[235]), .B(n2257), .Y(n555) );
  INVX1 U254 ( .A(n555), .Y(n113) );
  AND2X1 U256 ( .A(mem[216]), .B(n2258), .Y(n535) );
  INVX1 U258 ( .A(n535), .Y(n114) );
  AND2X1 U260 ( .A(mem[201]), .B(n2259), .Y(n519) );
  INVX1 U262 ( .A(n519), .Y(n115) );
  AND2X1 U265 ( .A(mem[158]), .B(n2262), .Y(n473) );
  INVX1 U267 ( .A(n473), .Y(n116) );
  AND2X1 U269 ( .A(mem[143]), .B(n2263), .Y(n456) );
  INVX1 U271 ( .A(n456), .Y(n117) );
  AND2X1 U273 ( .A(mem[122]), .B(n2264), .Y(n433) );
  INVX1 U275 ( .A(n433), .Y(n118) );
  AND2X1 U277 ( .A(mem[107]), .B(n2265), .Y(n416) );
  INVX1 U279 ( .A(n416), .Y(n119) );
  AND2X1 U281 ( .A(mem[88]), .B(n2266), .Y(n395) );
  INVX1 U283 ( .A(n395), .Y(n120) );
  AND2X1 U285 ( .A(mem[73]), .B(n2267), .Y(n378) );
  INVX1 U287 ( .A(n378), .Y(n121) );
  AND2X1 U289 ( .A(mem[30]), .B(n2270), .Y(n329) );
  INVX1 U291 ( .A(n329), .Y(n122) );
  AND2X1 U293 ( .A(mem[15]), .B(n2271), .Y(n311) );
  INVX1 U295 ( .A(n311), .Y(n123) );
  AND2X1 U298 ( .A(mem[503]), .B(n2240), .Y(n842) );
  INVX1 U300 ( .A(n842), .Y(n124) );
  AND2X1 U302 ( .A(mem[486]), .B(n2241), .Y(n824) );
  INVX1 U304 ( .A(n824), .Y(n125) );
  AND2X1 U306 ( .A(mem[469]), .B(n2242), .Y(n806) );
  INVX1 U308 ( .A(n806), .Y(n126) );
  AND2X1 U310 ( .A(mem[452]), .B(n2243), .Y(n788) );
  INVX1 U312 ( .A(n788), .Y(n127) );
  AND2X1 U314 ( .A(mem[443]), .B(n2244), .Y(n778) );
  INVX1 U316 ( .A(n778), .Y(n128) );
  AND2X1 U318 ( .A(mem[426]), .B(n2245), .Y(n760) );
  INVX1 U320 ( .A(n760), .Y(n129) );
  AND2X1 U322 ( .A(mem[409]), .B(n2246), .Y(n742) );
  INVX1 U324 ( .A(n742), .Y(n130) );
  AND2X1 U326 ( .A(mem[392]), .B(n2247), .Y(n723) );
  INVX1 U328 ( .A(n723), .Y(n131) );
  AND2X1 U332 ( .A(mem[351]), .B(n2250), .Y(n679) );
  INVX1 U334 ( .A(n679), .Y(n132) );
  AND2X1 U336 ( .A(mem[334]), .B(n2251), .Y(n661) );
  INVX1 U338 ( .A(n661), .Y(n133) );
  AND2X1 U340 ( .A(mem[311]), .B(n2252), .Y(n637) );
  INVX1 U342 ( .A(n637), .Y(n134) );
  AND2X1 U344 ( .A(mem[294]), .B(n2253), .Y(n619) );
  INVX1 U346 ( .A(n619), .Y(n135) );
  AND2X1 U348 ( .A(mem[277]), .B(n2254), .Y(n601) );
  INVX1 U350 ( .A(n601), .Y(n136) );
  AND2X1 U352 ( .A(mem[260]), .B(n2255), .Y(n582) );
  INVX1 U354 ( .A(n582), .Y(n137) );
  AND2X1 U356 ( .A(mem[251]), .B(n2256), .Y(n572) );
  INVX1 U358 ( .A(n572), .Y(n138) );
  AND2X1 U360 ( .A(mem[234]), .B(n2257), .Y(n554) );
  INVX1 U362 ( .A(n554), .Y(n139) );
  AND2X1 U365 ( .A(mem[217]), .B(n2258), .Y(n536) );
  INVX1 U367 ( .A(n536), .Y(n140) );
  AND2X1 U369 ( .A(mem[200]), .B(n2259), .Y(n518) );
  INVX1 U371 ( .A(n518), .Y(n141) );
  AND2X1 U373 ( .A(mem[159]), .B(n2262), .Y(n474) );
  INVX1 U375 ( .A(n474), .Y(n142) );
  AND2X1 U377 ( .A(mem[142]), .B(n2263), .Y(n455) );
  INVX1 U379 ( .A(n455), .Y(n143) );
  AND2X1 U381 ( .A(mem[123]), .B(n2264), .Y(n434) );
  INVX1 U383 ( .A(n434), .Y(n144) );
  AND2X1 U385 ( .A(mem[106]), .B(n2265), .Y(n415) );
  INVX1 U387 ( .A(n415), .Y(n145) );
  AND2X1 U389 ( .A(mem[89]), .B(n2266), .Y(n396) );
  INVX1 U391 ( .A(n396), .Y(n146) );
  AND2X1 U393 ( .A(mem[72]), .B(n2267), .Y(n377) );
  INVX1 U395 ( .A(n377), .Y(n147) );
  AND2X1 U398 ( .A(mem[31]), .B(n2270), .Y(n330) );
  INVX1 U400 ( .A(n330), .Y(n148) );
  AND2X1 U402 ( .A(mem[14]), .B(n2271), .Y(n309) );
  INVX1 U404 ( .A(n309), .Y(n149) );
  AND2X1 U406 ( .A(mem[508]), .B(n2240), .Y(n847) );
  INVX1 U408 ( .A(n847), .Y(n150) );
  AND2X1 U410 ( .A(mem[496]), .B(n2240), .Y(n835) );
  INVX1 U412 ( .A(n835), .Y(n151) );
  AND2X1 U414 ( .A(mem[493]), .B(n2241), .Y(n831) );
  INVX1 U416 ( .A(n831), .Y(n152) );
  AND2X1 U418 ( .A(mem[481]), .B(n2241), .Y(n819) );
  INVX1 U420 ( .A(n819), .Y(n153) );
  AND2X1 U422 ( .A(mem[466]), .B(n2242), .Y(n803) );
  INVX1 U424 ( .A(n803), .Y(n154) );
  AND2X1 U426 ( .A(mem[451]), .B(n2243), .Y(n787) );
  INVX1 U428 ( .A(n787), .Y(n155) );
  AND2X1 U431 ( .A(mem[446]), .B(n2244), .Y(n781) );
  INVX1 U433 ( .A(n781), .Y(n156) );
  AND2X1 U435 ( .A(mem[431]), .B(n2245), .Y(n765) );
  INVX1 U437 ( .A(n765), .Y(n157) );
  AND2X1 U439 ( .A(mem[376]), .B(n2248), .Y(n706) );
  INVX1 U441 ( .A(n706), .Y(n158) );
  AND2X1 U443 ( .A(mem[361]), .B(n2249), .Y(n690) );
  INVX1 U445 ( .A(n690), .Y(n159) );
  AND2X1 U447 ( .A(mem[346]), .B(n2250), .Y(n674) );
  INVX1 U449 ( .A(n674), .Y(n160) );
  AND2X1 U451 ( .A(mem[331]), .B(n2251), .Y(n658) );
  INVX1 U453 ( .A(n658), .Y(n161) );
  AND2X1 U455 ( .A(mem[316]), .B(n2252), .Y(n642) );
  INVX1 U457 ( .A(n642), .Y(n162) );
  AND2X1 U459 ( .A(mem[304]), .B(n2252), .Y(n630) );
  INVX1 U461 ( .A(n630), .Y(n163) );
  AND2X1 U464 ( .A(mem[301]), .B(n2253), .Y(n626) );
  INVX1 U466 ( .A(n626), .Y(n164) );
  AND2X1 U468 ( .A(mem[289]), .B(n2253), .Y(n614) );
  INVX1 U470 ( .A(n614), .Y(n165) );
  AND2X1 U472 ( .A(mem[274]), .B(n2254), .Y(n598) );
  INVX1 U474 ( .A(n598), .Y(n166) );
  AND2X1 U476 ( .A(mem[259]), .B(n2255), .Y(n581) );
  INVX1 U478 ( .A(n581), .Y(n167) );
  AND2X1 U480 ( .A(mem[254]), .B(n2256), .Y(n575) );
  INVX1 U482 ( .A(n575), .Y(n168) );
  AND2X1 U484 ( .A(mem[239]), .B(n2257), .Y(n559) );
  INVX1 U486 ( .A(n559), .Y(n169) );
  AND2X1 U488 ( .A(mem[184]), .B(n2260), .Y(n501) );
  INVX1 U490 ( .A(n501), .Y(n170) );
  AND2X1 U492 ( .A(mem[169]), .B(n2261), .Y(n485) );
  INVX1 U494 ( .A(n485), .Y(n171) );
  AND2X1 U497 ( .A(mem[154]), .B(n2262), .Y(n469) );
  INVX1 U499 ( .A(n469), .Y(n172) );
  AND2X1 U501 ( .A(mem[139]), .B(n2263), .Y(n452) );
  INVX1 U503 ( .A(n452), .Y(n173) );
  AND2X1 U505 ( .A(mem[126]), .B(n2264), .Y(n437) );
  INVX1 U507 ( .A(n437), .Y(n174) );
  AND2X1 U509 ( .A(mem[111]), .B(n2265), .Y(n420) );
  INVX1 U511 ( .A(n420), .Y(n175) );
  AND2X1 U513 ( .A(mem[56]), .B(n2268), .Y(n359) );
  INVX1 U515 ( .A(n359), .Y(n176) );
  AND2X1 U517 ( .A(mem[41]), .B(n2269), .Y(n342) );
  INVX1 U519 ( .A(n342), .Y(n177) );
  AND2X1 U521 ( .A(mem[26]), .B(n2270), .Y(n325) );
  INVX1 U523 ( .A(n325), .Y(n178) );
  AND2X1 U525 ( .A(mem[11]), .B(n2271), .Y(n303) );
  INVX1 U527 ( .A(n303), .Y(n179) );
  AND2X1 U530 ( .A(mem[509]), .B(n2240), .Y(n848) );
  INVX1 U532 ( .A(n848), .Y(n180) );
  AND2X1 U534 ( .A(mem[497]), .B(n2240), .Y(n836) );
  INVX1 U536 ( .A(n836), .Y(n181) );
  AND2X1 U538 ( .A(mem[492]), .B(n2241), .Y(n830) );
  INVX1 U540 ( .A(n830), .Y(n182) );
  AND2X1 U542 ( .A(mem[480]), .B(n2241), .Y(n818) );
  INVX1 U544 ( .A(n818), .Y(n183) );
  AND2X1 U546 ( .A(mem[467]), .B(n2242), .Y(n804) );
  INVX1 U548 ( .A(n804), .Y(n184) );
  AND2X1 U550 ( .A(mem[450]), .B(n2243), .Y(n786) );
  INVX1 U552 ( .A(n786), .Y(n185) );
  AND2X1 U554 ( .A(mem[447]), .B(n2244), .Y(n782) );
  INVX1 U556 ( .A(n782), .Y(n186) );
  AND2X1 U558 ( .A(mem[430]), .B(n2245), .Y(n764) );
  INVX1 U560 ( .A(n764), .Y(n187) );
  AND2X1 U563 ( .A(mem[377]), .B(n2248), .Y(n707) );
  INVX1 U565 ( .A(n707), .Y(n188) );
  AND2X1 U567 ( .A(mem[360]), .B(n2249), .Y(n689) );
  INVX1 U569 ( .A(n689), .Y(n189) );
  AND2X1 U571 ( .A(mem[347]), .B(n2250), .Y(n675) );
  INVX1 U573 ( .A(n675), .Y(n190) );
  AND2X1 U575 ( .A(mem[330]), .B(n2251), .Y(n657) );
  INVX1 U577 ( .A(n657), .Y(n191) );
  AND2X1 U579 ( .A(mem[317]), .B(n2252), .Y(n643) );
  INVX1 U581 ( .A(n643), .Y(n192) );
  AND2X1 U583 ( .A(mem[305]), .B(n2252), .Y(n631) );
  INVX1 U585 ( .A(n631), .Y(n193) );
  AND2X1 U587 ( .A(mem[300]), .B(n2253), .Y(n625) );
  INVX1 U589 ( .A(n625), .Y(n194) );
  AND2X1 U591 ( .A(mem[288]), .B(n2253), .Y(n613) );
  INVX1 U593 ( .A(n613), .Y(n195) );
  AND2X1 U597 ( .A(mem[275]), .B(n2254), .Y(n599) );
  INVX1 U599 ( .A(n599), .Y(n196) );
  AND2X1 U601 ( .A(mem[258]), .B(n2255), .Y(n580) );
  INVX1 U603 ( .A(n580), .Y(n197) );
  AND2X1 U605 ( .A(mem[255]), .B(n2256), .Y(n576) );
  INVX1 U607 ( .A(n576), .Y(n198) );
  AND2X1 U609 ( .A(mem[238]), .B(n2257), .Y(n558) );
  INVX1 U611 ( .A(n558), .Y(n199) );
  AND2X1 U613 ( .A(mem[185]), .B(n2260), .Y(n502) );
  INVX1 U615 ( .A(n502), .Y(n200) );
  AND2X1 U617 ( .A(mem[168]), .B(n2261), .Y(n484) );
  INVX1 U619 ( .A(n484), .Y(n201) );
  AND2X1 U621 ( .A(mem[155]), .B(n2262), .Y(n470) );
  INVX1 U623 ( .A(n470), .Y(n202) );
  AND2X1 U625 ( .A(mem[138]), .B(n2263), .Y(n451) );
  INVX1 U627 ( .A(n451), .Y(n203) );
  AND2X1 U630 ( .A(mem[127]), .B(n2264), .Y(n438) );
  INVX1 U632 ( .A(n438), .Y(n204) );
  AND2X1 U634 ( .A(mem[110]), .B(n2265), .Y(n419) );
  INVX1 U636 ( .A(n419), .Y(n205) );
  AND2X1 U638 ( .A(mem[57]), .B(n2268), .Y(n360) );
  INVX1 U640 ( .A(n360), .Y(n206) );
  AND2X1 U642 ( .A(mem[40]), .B(n2269), .Y(n341) );
  INVX1 U644 ( .A(n341), .Y(n207) );
  AND2X1 U646 ( .A(mem[27]), .B(n2270), .Y(n326) );
  INVX1 U648 ( .A(n326), .Y(n208) );
  AND2X1 U650 ( .A(mem[10]), .B(n2271), .Y(n301) );
  INVX1 U652 ( .A(n301), .Y(n209) );
  AND2X1 U654 ( .A(mem[498]), .B(n2240), .Y(n837) );
  INVX1 U656 ( .A(n837), .Y(n210) );
  AND2X1 U658 ( .A(mem[483]), .B(n2241), .Y(n821) );
  INVX1 U660 ( .A(n821), .Y(n211) );
  AND2X1 U663 ( .A(mem[476]), .B(n2242), .Y(n813) );
  INVX1 U665 ( .A(n813), .Y(n212) );
  AND2X1 U667 ( .A(mem[464]), .B(n2242), .Y(n801) );
  INVX1 U669 ( .A(n801), .Y(n213) );
  AND2X1 U671 ( .A(mem[461]), .B(n2243), .Y(n797) );
  INVX1 U673 ( .A(n797), .Y(n214) );
  AND2X1 U675 ( .A(mem[449]), .B(n2243), .Y(n785) );
  INVX1 U677 ( .A(n785), .Y(n215) );
  AND2X1 U679 ( .A(mem[414]), .B(n2246), .Y(n747) );
  INVX1 U681 ( .A(n747), .Y(n216) );
  AND2X1 U683 ( .A(mem[399]), .B(n2247), .Y(n730) );
  INVX1 U685 ( .A(n730), .Y(n217) );
  AND2X1 U687 ( .A(mem[378]), .B(n2248), .Y(n708) );
  INVX1 U689 ( .A(n708), .Y(n218) );
  AND2X1 U691 ( .A(mem[363]), .B(n2249), .Y(n692) );
  INVX1 U693 ( .A(n692), .Y(n219) );
  AND2X1 U696 ( .A(mem[344]), .B(n2250), .Y(n672) );
  INVX1 U698 ( .A(n672), .Y(n220) );
  AND2X1 U700 ( .A(mem[329]), .B(n2251), .Y(n656) );
  INVX1 U702 ( .A(n656), .Y(n221) );
  AND2X1 U704 ( .A(mem[306]), .B(n2252), .Y(n632) );
  INVX1 U706 ( .A(n632), .Y(n222) );
  AND2X1 U708 ( .A(mem[291]), .B(n2253), .Y(n616) );
  INVX1 U710 ( .A(n616), .Y(n223) );
  AND2X1 U712 ( .A(mem[284]), .B(n2254), .Y(n608) );
  INVX1 U714 ( .A(n608), .Y(n224) );
  AND2X1 U716 ( .A(mem[272]), .B(n2254), .Y(n596) );
  INVX1 U718 ( .A(n596), .Y(n225) );
  AND2X1 U720 ( .A(mem[269]), .B(n2255), .Y(n591) );
  INVX1 U722 ( .A(n591), .Y(n226) );
  AND2X1 U724 ( .A(mem[257]), .B(n2255), .Y(n579) );
  INVX1 U726 ( .A(n579), .Y(n227) );
  AND2X1 U729 ( .A(mem[222]), .B(n2258), .Y(n541) );
  INVX1 U731 ( .A(n541), .Y(n228) );
  AND2X1 U733 ( .A(mem[207]), .B(n2259), .Y(n525) );
  INVX1 U735 ( .A(n525), .Y(n229) );
  AND2X1 U737 ( .A(mem[186]), .B(n2260), .Y(n503) );
  INVX1 U739 ( .A(n503), .Y(n230) );
  AND2X1 U741 ( .A(mem[171]), .B(n2261), .Y(n487) );
  INVX1 U743 ( .A(n487), .Y(n231) );
  AND2X1 U745 ( .A(mem[152]), .B(n2262), .Y(n467) );
  INVX1 U747 ( .A(n467), .Y(n232) );
  AND2X1 U749 ( .A(mem[137]), .B(n2263), .Y(n450) );
  INVX1 U751 ( .A(n450), .Y(n233) );
  AND2X1 U753 ( .A(mem[94]), .B(n2266), .Y(n401) );
  INVX1 U755 ( .A(n401), .Y(n234) );
  AND2X1 U757 ( .A(mem[79]), .B(n2267), .Y(n384) );
  INVX1 U759 ( .A(n384), .Y(n235) );
  AND2X1 U762 ( .A(mem[58]), .B(n2268), .Y(n361) );
  INVX1 U764 ( .A(n361), .Y(n236) );
  AND2X1 U766 ( .A(mem[43]), .B(n2269), .Y(n344) );
  INVX1 U768 ( .A(n344), .Y(n237) );
  AND2X1 U770 ( .A(mem[24]), .B(n2270), .Y(n323) );
  INVX1 U772 ( .A(n323), .Y(n238) );
  AND2X1 U774 ( .A(mem[9]), .B(n2271), .Y(n299) );
  INVX1 U776 ( .A(n299), .Y(n239) );
  AND2X1 U778 ( .A(n20), .B(n855), .Y(n857) );
  INVX1 U780 ( .A(n857), .Y(n240) );
  AND2X1 U782 ( .A(mem[499]), .B(n2240), .Y(n838) );
  INVX1 U784 ( .A(n838), .Y(n241) );
  AND2X1 U786 ( .A(mem[482]), .B(n2241), .Y(n820) );
  INVX1 U788 ( .A(n820), .Y(n242) );
  AND2X1 U790 ( .A(mem[477]), .B(n2242), .Y(n814) );
  INVX1 U792 ( .A(n814), .Y(n243) );
  AND2X1 U795 ( .A(mem[465]), .B(n2242), .Y(n802) );
  INVX1 U797 ( .A(n802), .Y(n244) );
  AND2X1 U799 ( .A(mem[460]), .B(n2243), .Y(n796) );
  INVX1 U801 ( .A(n796), .Y(n245) );
  AND2X1 U803 ( .A(mem[448]), .B(n2243), .Y(n784) );
  INVX1 U805 ( .A(n784), .Y(n246) );
  AND2X1 U807 ( .A(mem[415]), .B(n2246), .Y(n748) );
  INVX1 U809 ( .A(n748), .Y(n247) );
  AND2X1 U811 ( .A(mem[398]), .B(n2247), .Y(n729) );
  INVX1 U813 ( .A(n729), .Y(n248) );
  AND2X1 U815 ( .A(mem[379]), .B(n2248), .Y(n709) );
  INVX1 U817 ( .A(n709), .Y(n249) );
  AND2X1 U819 ( .A(mem[362]), .B(n2249), .Y(n691) );
  INVX1 U821 ( .A(n691), .Y(n250) );
  AND2X1 U823 ( .A(mem[345]), .B(n2250), .Y(n673) );
  INVX1 U825 ( .A(n673), .Y(n251) );
  AND2X1 U828 ( .A(mem[328]), .B(n2251), .Y(n655) );
  INVX1 U830 ( .A(n655), .Y(n252) );
  AND2X1 U832 ( .A(mem[307]), .B(n2252), .Y(n633) );
  INVX1 U834 ( .A(n633), .Y(n253) );
  AND2X1 U836 ( .A(mem[290]), .B(n2253), .Y(n615) );
  INVX1 U838 ( .A(n615), .Y(n254) );
  AND2X1 U840 ( .A(mem[285]), .B(n2254), .Y(n609) );
  INVX1 U842 ( .A(n609), .Y(n255) );
  AND2X1 U844 ( .A(mem[273]), .B(n2254), .Y(n597) );
  INVX1 U846 ( .A(n597), .Y(n256) );
  AND2X1 U848 ( .A(mem[268]), .B(n2255), .Y(n590) );
  INVX1 U850 ( .A(n590), .Y(n257) );
  AND2X1 U852 ( .A(mem[256]), .B(n2255), .Y(n578) );
  INVX1 U854 ( .A(n578), .Y(n258) );
  AND2X1 U856 ( .A(mem[223]), .B(n2258), .Y(n542) );
  INVX1 U858 ( .A(n542), .Y(n259) );
  AND2X1 U862 ( .A(mem[206]), .B(n2259), .Y(n524) );
  INVX1 U864 ( .A(n524), .Y(n260) );
  AND2X1 U866 ( .A(mem[187]), .B(n2260), .Y(n504) );
  INVX1 U868 ( .A(n504), .Y(n261) );
  AND2X1 U870 ( .A(mem[170]), .B(n2261), .Y(n486) );
  INVX1 U872 ( .A(n486), .Y(n262) );
  AND2X1 U874 ( .A(mem[153]), .B(n2262), .Y(n468) );
  INVX1 U876 ( .A(n468), .Y(n263) );
  AND2X1 U878 ( .A(mem[136]), .B(n2263), .Y(n449) );
  INVX1 U880 ( .A(n449), .Y(n264) );
  AND2X1 U882 ( .A(mem[95]), .B(n2266), .Y(n402) );
  INVX1 U884 ( .A(n402), .Y(n265) );
  AND2X1 U886 ( .A(mem[78]), .B(n2267), .Y(n383) );
  INVX1 U888 ( .A(n383), .Y(n266) );
  AND2X1 U890 ( .A(mem[59]), .B(n2268), .Y(n362) );
  INVX1 U892 ( .A(n362), .Y(n267) );
  AND2X1 U896 ( .A(mem[42]), .B(n2269), .Y(n343) );
  INVX1 U898 ( .A(n343), .Y(n268) );
  AND2X1 U900 ( .A(mem[25]), .B(n2270), .Y(n324) );
  INVX1 U902 ( .A(n324), .Y(n269) );
  AND2X1 U904 ( .A(mem[8]), .B(n2271), .Y(n297) );
  INVX1 U906 ( .A(n297), .Y(n270) );
  AND2X1 U908 ( .A(mem[510]), .B(n2240), .Y(n849) );
  INVX1 U910 ( .A(n849), .Y(n271) );
  AND2X1 U912 ( .A(mem[495]), .B(n2241), .Y(n833) );
  INVX1 U914 ( .A(n833), .Y(n272) );
  AND2X1 U916 ( .A(mem[444]), .B(n2244), .Y(n779) );
  INVX1 U918 ( .A(n779), .Y(n273) );
  AND2X1 U920 ( .A(mem[432]), .B(n2244), .Y(n767) );
  INVX1 U922 ( .A(n767), .Y(n274) );
  AND2X1 U924 ( .A(mem[429]), .B(n2245), .Y(n763) );
  INVX1 U926 ( .A(n763), .Y(n275) );
  AND2X1 U930 ( .A(mem[417]), .B(n2245), .Y(n751) );
  INVX1 U932 ( .A(n751), .Y(n276) );
  AND2X1 U934 ( .A(mem[402]), .B(n2246), .Y(n735) );
  INVX1 U936 ( .A(n735), .Y(n277) );
  AND2X1 U938 ( .A(mem[387]), .B(n2247), .Y(n718) );
  INVX1 U940 ( .A(n718), .Y(n278) );
  AND2X1 U942 ( .A(mem[372]), .B(n2248), .Y(n702) );
  INVX1 U944 ( .A(n702), .Y(n279) );
  AND2X1 U946 ( .A(mem[357]), .B(n2249), .Y(n686) );
  INVX1 U948 ( .A(n686), .Y(n280) );
  AND2X1 U950 ( .A(mem[342]), .B(n2250), .Y(n670) );
  INVX1 U952 ( .A(n670), .Y(n282) );
  AND2X1 U954 ( .A(mem[327]), .B(n2251), .Y(n654) );
  INVX1 U956 ( .A(n654), .Y(n284) );
  AND2X1 U958 ( .A(mem[318]), .B(n2252), .Y(n644) );
  INVX1 U960 ( .A(n644), .Y(n286) );
  AND2X1 U964 ( .A(mem[303]), .B(n2253), .Y(n628) );
  INVX1 U966 ( .A(n628), .Y(n288) );
  AND2X1 U968 ( .A(mem[252]), .B(n2256), .Y(n573) );
  INVX1 U970 ( .A(n573), .Y(n290) );
  AND2X1 U972 ( .A(mem[240]), .B(n2256), .Y(n561) );
  INVX1 U974 ( .A(n561), .Y(n292) );
  AND2X1 U976 ( .A(mem[237]), .B(n2257), .Y(n557) );
  INVX1 U978 ( .A(n557), .Y(n294) );
  AND2X1 U980 ( .A(mem[225]), .B(n2257), .Y(n545) );
  INVX1 U982 ( .A(n545), .Y(n296) );
  AND2X1 U984 ( .A(mem[210]), .B(n2258), .Y(n529) );
  INVX1 U986 ( .A(n529), .Y(n298) );
  AND2X1 U988 ( .A(mem[195]), .B(n2259), .Y(n513) );
  INVX1 U990 ( .A(n513), .Y(n300) );
  AND2X1 U992 ( .A(mem[180]), .B(n2260), .Y(n497) );
  INVX1 U994 ( .A(n497), .Y(n302) );
  AND2X1 U998 ( .A(mem[165]), .B(n2261), .Y(n481) );
  INVX1 U1000 ( .A(n481), .Y(n304) );
  AND2X1 U1002 ( .A(mem[150]), .B(n2262), .Y(n465) );
  INVX1 U1004 ( .A(n465), .Y(n306) );
  AND2X1 U1006 ( .A(mem[135]), .B(n2263), .Y(n448) );
  INVX1 U1008 ( .A(n448), .Y(n308) );
  AND2X1 U1010 ( .A(mem[124]), .B(n2264), .Y(n435) );
  INVX1 U1012 ( .A(n435), .Y(n310) );
  AND2X1 U1014 ( .A(mem[112]), .B(n2264), .Y(n423) );
  INVX1 U1016 ( .A(n423), .Y(n1414) );
  AND2X1 U1018 ( .A(mem[109]), .B(n2265), .Y(n418) );
  INVX1 U1020 ( .A(n418), .Y(n1415) );
  AND2X1 U1022 ( .A(mem[97]), .B(n2265), .Y(n406) );
  INVX1 U1024 ( .A(n406), .Y(n1416) );
  AND2X1 U1026 ( .A(mem[82]), .B(n2266), .Y(n389) );
  INVX1 U1028 ( .A(n389), .Y(n1417) );
  AND2X1 U1032 ( .A(mem[67]), .B(n2267), .Y(n372) );
  INVX1 U1034 ( .A(n372), .Y(n1418) );
  AND2X1 U1036 ( .A(mem[52]), .B(n2268), .Y(n355) );
  INVX1 U1038 ( .A(n355), .Y(n1419) );
  AND2X1 U1040 ( .A(mem[37]), .B(n2269), .Y(n338) );
  INVX1 U1042 ( .A(n338), .Y(n1420) );
  AND2X1 U1044 ( .A(mem[22]), .B(n2270), .Y(n321) );
  INVX1 U1046 ( .A(n321), .Y(n1421) );
  AND2X1 U1048 ( .A(mem[7]), .B(n2271), .Y(n295) );
  INVX1 U1050 ( .A(n295), .Y(n1422) );
  BUFX2 U1052 ( .A(n386), .Y(n1423) );
  BUFX2 U1054 ( .A(n368), .Y(n1424) );
  AND2X1 U1056 ( .A(n76), .B(n2238), .Y(n865) );
  INVX1 U1058 ( .A(n865), .Y(n1425) );
  AND2X1 U1060 ( .A(n23), .B(n855), .Y(n858) );
  INVX1 U1062 ( .A(n858), .Y(n1426) );
  AND2X1 U1066 ( .A(mem[511]), .B(n2240), .Y(n850) );
  INVX1 U1068 ( .A(n850), .Y(n1427) );
  AND2X1 U1070 ( .A(mem[494]), .B(n2241), .Y(n832) );
  INVX1 U1072 ( .A(n832), .Y(n1428) );
  AND2X1 U1074 ( .A(mem[445]), .B(n2244), .Y(n780) );
  INVX1 U1076 ( .A(n780), .Y(n1429) );
  AND2X1 U1078 ( .A(mem[433]), .B(n2244), .Y(n768) );
  INVX1 U1080 ( .A(n768), .Y(n1430) );
  AND2X1 U1082 ( .A(mem[428]), .B(n2245), .Y(n762) );
  INVX1 U1084 ( .A(n762), .Y(n1431) );
  AND2X1 U1086 ( .A(mem[416]), .B(n2245), .Y(n750) );
  INVX1 U1088 ( .A(n750), .Y(n1432) );
  AND2X1 U1090 ( .A(mem[403]), .B(n2246), .Y(n736) );
  INVX1 U1092 ( .A(n736), .Y(n1433) );
  AND2X1 U1094 ( .A(mem[386]), .B(n2247), .Y(n717) );
  INVX1 U1096 ( .A(n717), .Y(n1434) );
  AND2X1 U1100 ( .A(mem[373]), .B(n2248), .Y(n703) );
  INVX1 U1101 ( .A(n703), .Y(n1435) );
  AND2X1 U1103 ( .A(mem[356]), .B(n2249), .Y(n685) );
  INVX1 U1104 ( .A(n685), .Y(n1436) );
  AND2X1 U1106 ( .A(mem[343]), .B(n2250), .Y(n671) );
  INVX1 U1107 ( .A(n671), .Y(n1437) );
  AND2X1 U1109 ( .A(mem[326]), .B(n2251), .Y(n653) );
  INVX1 U1110 ( .A(n653), .Y(n1438) );
  AND2X1 U1112 ( .A(mem[319]), .B(n2252), .Y(n645) );
  INVX1 U1113 ( .A(n645), .Y(n1439) );
  AND2X1 U1115 ( .A(mem[302]), .B(n2253), .Y(n627) );
  INVX1 U1116 ( .A(n627), .Y(n1440) );
  AND2X1 U1118 ( .A(mem[253]), .B(n2256), .Y(n574) );
  INVX1 U1119 ( .A(n574), .Y(n1441) );
  AND2X1 U1121 ( .A(mem[241]), .B(n2256), .Y(n562) );
  INVX1 U1122 ( .A(n562), .Y(n1442) );
  AND2X1 U1124 ( .A(mem[236]), .B(n2257), .Y(n556) );
  INVX1 U1125 ( .A(n556), .Y(n1443) );
  AND2X1 U1127 ( .A(mem[224]), .B(n2257), .Y(n544) );
  INVX1 U1128 ( .A(n544), .Y(n1444) );
  AND2X1 U1130 ( .A(mem[211]), .B(n2258), .Y(n530) );
  INVX1 U1131 ( .A(n530), .Y(n1445) );
  AND2X1 U1133 ( .A(mem[194]), .B(n2259), .Y(n512) );
  INVX1 U1134 ( .A(n512), .Y(n1446) );
  AND2X1 U1136 ( .A(mem[181]), .B(n2260), .Y(n498) );
  INVX1 U1137 ( .A(n498), .Y(n1447) );
  AND2X1 U1139 ( .A(mem[164]), .B(n2261), .Y(n480) );
  INVX1 U1140 ( .A(n480), .Y(n1448) );
  AND2X1 U1142 ( .A(mem[151]), .B(n2262), .Y(n466) );
  INVX1 U1143 ( .A(n466), .Y(n1449) );
  AND2X1 U1145 ( .A(mem[134]), .B(n2263), .Y(n447) );
  INVX1 U1146 ( .A(n447), .Y(n1450) );
  AND2X1 U1151 ( .A(mem[125]), .B(n2264), .Y(n436) );
  INVX1 U1153 ( .A(n436), .Y(n1451) );
  AND2X1 U1155 ( .A(mem[113]), .B(n2264), .Y(n424) );
  INVX1 U1157 ( .A(n424), .Y(n1452) );
  AND2X1 U1159 ( .A(mem[108]), .B(n2265), .Y(n417) );
  INVX1 U1161 ( .A(n417), .Y(n1453) );
  AND2X1 U1163 ( .A(mem[96]), .B(n2265), .Y(n405) );
  INVX1 U1165 ( .A(n405), .Y(n1454) );
  AND2X1 U1167 ( .A(mem[83]), .B(n2266), .Y(n390) );
  INVX1 U1184 ( .A(n390), .Y(n1455) );
  AND2X1 U1185 ( .A(mem[66]), .B(n2267), .Y(n371) );
  INVX1 U1187 ( .A(n371), .Y(n1456) );
  AND2X1 U1188 ( .A(mem[53]), .B(n2268), .Y(n356) );
  INVX1 U1189 ( .A(n356), .Y(n1457) );
  AND2X1 U1192 ( .A(mem[36]), .B(n2269), .Y(n337) );
  INVX1 U1200 ( .A(n337), .Y(n1458) );
  AND2X1 U1201 ( .A(mem[23]), .B(n2270), .Y(n322) );
  INVX1 U1202 ( .A(n322), .Y(n1459) );
  AND2X1 U1203 ( .A(mem[6]), .B(n2271), .Y(n293) );
  INVX1 U1204 ( .A(n293), .Y(n1460) );
  BUFX2 U1205 ( .A(n404), .Y(n1461) );
  BUFX2 U1206 ( .A(n350), .Y(n1462) );
  AND2X1 U1207 ( .A(n2291), .B(n2239), .Y(n864) );
  INVX1 U1208 ( .A(n864), .Y(n1463) );
  AND2X1 U1209 ( .A(n22), .B(n855), .Y(n854) );
  INVX1 U1210 ( .A(n854), .Y(n1464) );
  AND2X1 U1211 ( .A(mem[478]), .B(n2242), .Y(n815) );
  INVX1 U1212 ( .A(n815), .Y(n1465) );
  AND2X1 U1213 ( .A(mem[463]), .B(n2243), .Y(n799) );
  INVX1 U1214 ( .A(n799), .Y(n1466) );
  AND2X1 U1215 ( .A(mem[434]), .B(n2244), .Y(n769) );
  INVX1 U1216 ( .A(n769), .Y(n1467) );
  AND2X1 U1217 ( .A(mem[419]), .B(n2245), .Y(n753) );
  INVX1 U1218 ( .A(n753), .Y(n1468) );
  AND2X1 U1219 ( .A(mem[412]), .B(n2246), .Y(n745) );
  INVX1 U1220 ( .A(n745), .Y(n1469) );
  AND2X1 U1221 ( .A(mem[400]), .B(n2246), .Y(n733) );
  INVX1 U1222 ( .A(n733), .Y(n1470) );
  AND2X1 U1223 ( .A(mem[397]), .B(n2247), .Y(n728) );
  INVX1 U1224 ( .A(n728), .Y(n1471) );
  AND2X1 U1225 ( .A(mem[385]), .B(n2247), .Y(n716) );
  INVX1 U1226 ( .A(n716), .Y(n1472) );
  AND2X1 U1227 ( .A(mem[374]), .B(n2248), .Y(n704) );
  INVX1 U1228 ( .A(n704), .Y(n1473) );
  AND2X1 U1229 ( .A(mem[359]), .B(n2249), .Y(n688) );
  INVX1 U1230 ( .A(n688), .Y(n1474) );
  AND2X1 U1231 ( .A(mem[340]), .B(n2250), .Y(n668) );
  INVX1 U1232 ( .A(n668), .Y(n1475) );
  AND2X1 U1233 ( .A(mem[325]), .B(n2251), .Y(n652) );
  INVX1 U1234 ( .A(n652), .Y(n1476) );
  AND2X1 U1235 ( .A(mem[286]), .B(n2254), .Y(n610) );
  INVX1 U1236 ( .A(n610), .Y(n1477) );
  AND2X1 U1237 ( .A(mem[271]), .B(n2255), .Y(n593) );
  INVX1 U1238 ( .A(n593), .Y(n1478) );
  AND2X1 U1239 ( .A(mem[242]), .B(n2256), .Y(n563) );
  INVX1 U1240 ( .A(n563), .Y(n1479) );
  AND2X1 U1241 ( .A(mem[227]), .B(n2257), .Y(n547) );
  INVX1 U1242 ( .A(n547), .Y(n1480) );
  AND2X1 U1243 ( .A(mem[220]), .B(n2258), .Y(n539) );
  INVX1 U1244 ( .A(n539), .Y(n1481) );
  AND2X1 U1245 ( .A(mem[208]), .B(n2258), .Y(n527) );
  INVX1 U1246 ( .A(n527), .Y(n1482) );
  AND2X1 U1247 ( .A(mem[205]), .B(n2259), .Y(n523) );
  INVX1 U1248 ( .A(n523), .Y(n1483) );
  AND2X1 U1249 ( .A(mem[193]), .B(n2259), .Y(n511) );
  INVX1 U1250 ( .A(n511), .Y(n1484) );
  AND2X1 U1251 ( .A(mem[182]), .B(n2260), .Y(n499) );
  INVX1 U1252 ( .A(n499), .Y(n1485) );
  AND2X1 U1253 ( .A(mem[167]), .B(n2261), .Y(n483) );
  INVX1 U1254 ( .A(n483), .Y(n1486) );
  AND2X1 U1255 ( .A(mem[148]), .B(n2262), .Y(n463) );
  INVX1 U1256 ( .A(n463), .Y(n1487) );
  AND2X1 U1257 ( .A(mem[133]), .B(n2263), .Y(n446) );
  INVX1 U1258 ( .A(n446), .Y(n1488) );
  AND2X1 U1259 ( .A(mem[114]), .B(n2264), .Y(n425) );
  INVX1 U1260 ( .A(n425), .Y(n1489) );
  AND2X1 U1261 ( .A(mem[99]), .B(n2265), .Y(n408) );
  INVX1 U1262 ( .A(n408), .Y(n1490) );
  AND2X1 U1263 ( .A(mem[92]), .B(n2266), .Y(n399) );
  INVX1 U1264 ( .A(n399), .Y(n1491) );
  AND2X1 U1265 ( .A(mem[80]), .B(n2266), .Y(n387) );
  INVX1 U1266 ( .A(n387), .Y(n1492) );
  AND2X1 U1267 ( .A(mem[77]), .B(n2267), .Y(n382) );
  INVX1 U1268 ( .A(n382), .Y(n1493) );
  AND2X1 U1269 ( .A(mem[65]), .B(n2267), .Y(n370) );
  INVX1 U1270 ( .A(n370), .Y(n1494) );
  AND2X1 U1271 ( .A(mem[54]), .B(n2268), .Y(n357) );
  INVX1 U1272 ( .A(n357), .Y(n1495) );
  AND2X1 U1273 ( .A(mem[39]), .B(n2269), .Y(n340) );
  INVX1 U1274 ( .A(n340), .Y(n1496) );
  AND2X1 U1275 ( .A(mem[20]), .B(n2270), .Y(n319) );
  INVX1 U1276 ( .A(n319), .Y(n1497) );
  AND2X1 U1277 ( .A(mem[5]), .B(n2271), .Y(n291) );
  INVX1 U1278 ( .A(n291), .Y(n1498) );
  BUFX2 U1279 ( .A(n422), .Y(n1499) );
  BUFX2 U1280 ( .A(n332), .Y(n1500) );
  AND2X1 U1281 ( .A(n73), .B(n861), .Y(n863) );
  INVX1 U1282 ( .A(n863), .Y(n1501) );
  AND2X1 U1283 ( .A(reset), .B(n1703), .Y(n861) );
  AND2X1 U1284 ( .A(mem[479]), .B(n2242), .Y(n816) );
  INVX1 U1285 ( .A(n816), .Y(n1502) );
  AND2X1 U1286 ( .A(mem[462]), .B(n2243), .Y(n798) );
  INVX1 U1287 ( .A(n798), .Y(n1503) );
  AND2X1 U1288 ( .A(mem[435]), .B(n2244), .Y(n770) );
  INVX1 U1289 ( .A(n770), .Y(n1504) );
  AND2X1 U1290 ( .A(mem[418]), .B(n2245), .Y(n752) );
  INVX1 U1291 ( .A(n752), .Y(n1505) );
  AND2X1 U1292 ( .A(mem[413]), .B(n2246), .Y(n746) );
  INVX1 U1293 ( .A(n746), .Y(n1506) );
  AND2X1 U1294 ( .A(mem[401]), .B(n2246), .Y(n734) );
  INVX1 U1295 ( .A(n734), .Y(n1507) );
  AND2X1 U1296 ( .A(mem[396]), .B(n2247), .Y(n727) );
  INVX1 U1297 ( .A(n727), .Y(n1508) );
  AND2X1 U1298 ( .A(mem[384]), .B(n2247), .Y(n715) );
  INVX1 U1299 ( .A(n715), .Y(n1509) );
  AND2X1 U1300 ( .A(mem[375]), .B(n2248), .Y(n705) );
  INVX1 U1301 ( .A(n705), .Y(n1510) );
  AND2X1 U1302 ( .A(mem[358]), .B(n2249), .Y(n687) );
  INVX1 U1303 ( .A(n687), .Y(n1511) );
  AND2X1 U1304 ( .A(mem[341]), .B(n2250), .Y(n669) );
  INVX1 U1305 ( .A(n669), .Y(n1512) );
  AND2X1 U1306 ( .A(mem[324]), .B(n2251), .Y(n651) );
  INVX1 U1307 ( .A(n651), .Y(n1513) );
  AND2X1 U1308 ( .A(mem[287]), .B(n2254), .Y(n611) );
  INVX1 U1309 ( .A(n611), .Y(n1514) );
  AND2X1 U1310 ( .A(mem[270]), .B(n2255), .Y(n592) );
  INVX1 U1311 ( .A(n592), .Y(n1515) );
  AND2X1 U1312 ( .A(mem[243]), .B(n2256), .Y(n564) );
  INVX1 U1313 ( .A(n564), .Y(n1516) );
  AND2X1 U1314 ( .A(mem[226]), .B(n2257), .Y(n546) );
  INVX1 U1315 ( .A(n546), .Y(n1517) );
  AND2X1 U1316 ( .A(mem[221]), .B(n2258), .Y(n540) );
  INVX1 U1317 ( .A(n540), .Y(n1518) );
  AND2X1 U1318 ( .A(mem[209]), .B(n2258), .Y(n528) );
  INVX1 U1319 ( .A(n528), .Y(n1519) );
  AND2X1 U1320 ( .A(mem[204]), .B(n2259), .Y(n522) );
  INVX1 U1321 ( .A(n522), .Y(n1520) );
  AND2X1 U1322 ( .A(mem[192]), .B(n2259), .Y(n510) );
  INVX1 U1323 ( .A(n510), .Y(n1521) );
  AND2X1 U1324 ( .A(mem[183]), .B(n2260), .Y(n500) );
  INVX1 U1325 ( .A(n500), .Y(n1522) );
  AND2X1 U1326 ( .A(mem[166]), .B(n2261), .Y(n482) );
  INVX1 U1327 ( .A(n482), .Y(n1523) );
  AND2X1 U1328 ( .A(mem[149]), .B(n2262), .Y(n464) );
  INVX1 U1329 ( .A(n464), .Y(n1524) );
  AND2X1 U1330 ( .A(mem[132]), .B(n2263), .Y(n445) );
  INVX1 U1331 ( .A(n445), .Y(n1525) );
  AND2X1 U1332 ( .A(mem[115]), .B(n2264), .Y(n426) );
  INVX1 U1333 ( .A(n426), .Y(n1526) );
  AND2X1 U1334 ( .A(mem[98]), .B(n2265), .Y(n407) );
  INVX1 U1335 ( .A(n407), .Y(n1527) );
  AND2X1 U1336 ( .A(mem[93]), .B(n2266), .Y(n400) );
  INVX1 U1337 ( .A(n400), .Y(n1528) );
  AND2X1 U1338 ( .A(mem[81]), .B(n2266), .Y(n388) );
  INVX1 U1339 ( .A(n388), .Y(n1529) );
  AND2X1 U1340 ( .A(mem[76]), .B(n2267), .Y(n381) );
  INVX1 U1341 ( .A(n381), .Y(n1530) );
  AND2X1 U1342 ( .A(mem[64]), .B(n2267), .Y(n369) );
  INVX1 U1343 ( .A(n369), .Y(n1531) );
  AND2X1 U1344 ( .A(mem[55]), .B(n2268), .Y(n358) );
  INVX1 U1345 ( .A(n358), .Y(n1532) );
  AND2X1 U1346 ( .A(mem[38]), .B(n2269), .Y(n339) );
  INVX1 U1347 ( .A(n339), .Y(n1533) );
  AND2X1 U1348 ( .A(mem[21]), .B(n2270), .Y(n320) );
  INVX1 U1349 ( .A(n320), .Y(n1534) );
  AND2X1 U1350 ( .A(mem[4]), .B(n2271), .Y(n289) );
  INVX1 U1351 ( .A(n289), .Y(n1535) );
  AND2X1 U1352 ( .A(put), .B(full_bar), .Y(n852) );
  INVX1 U1353 ( .A(n852), .Y(n1536) );
  BUFX2 U1354 ( .A(n440), .Y(n1537) );
  BUFX2 U1355 ( .A(n314), .Y(n1538) );
  AND2X1 U1356 ( .A(n2309), .B(n855), .Y(n883) );
  INVX1 U1357 ( .A(n883), .Y(n1539) );
  AND2X1 U1358 ( .A(mem[504]), .B(n2240), .Y(n843) );
  INVX1 U1359 ( .A(n843), .Y(n1540) );
  AND2X1 U1360 ( .A(mem[489]), .B(n2241), .Y(n827) );
  INVX1 U1361 ( .A(n827), .Y(n1541) );
  AND2X1 U1362 ( .A(mem[474]), .B(n2242), .Y(n811) );
  INVX1 U1363 ( .A(n811), .Y(n1542) );
  AND2X1 U1364 ( .A(mem[459]), .B(n2243), .Y(n795) );
  INVX1 U1365 ( .A(n795), .Y(n1543) );
  AND2X1 U1366 ( .A(mem[436]), .B(n2244), .Y(n771) );
  INVX1 U1367 ( .A(n771), .Y(n1544) );
  AND2X1 U1368 ( .A(mem[421]), .B(n2245), .Y(n755) );
  INVX1 U1369 ( .A(n755), .Y(n1545) );
  AND2X1 U1370 ( .A(mem[406]), .B(n2246), .Y(n739) );
  INVX1 U1371 ( .A(n739), .Y(n1546) );
  AND2X1 U1372 ( .A(mem[391]), .B(n2247), .Y(n722) );
  INVX1 U1373 ( .A(n722), .Y(n1547) );
  AND2X1 U1374 ( .A(mem[380]), .B(n2248), .Y(n710) );
  INVX1 U1375 ( .A(n710), .Y(n1548) );
  AND2X1 U1376 ( .A(mem[368]), .B(n2248), .Y(n698) );
  INVX1 U1377 ( .A(n698), .Y(n1549) );
  AND2X1 U1378 ( .A(mem[365]), .B(n2249), .Y(n694) );
  INVX1 U1379 ( .A(n694), .Y(n1550) );
  AND2X1 U1380 ( .A(mem[353]), .B(n2249), .Y(n682) );
  INVX1 U1381 ( .A(n682), .Y(n1551) );
  AND2X1 U1382 ( .A(mem[338]), .B(n2250), .Y(n666) );
  INVX1 U1383 ( .A(n666), .Y(n1552) );
  AND2X1 U1384 ( .A(mem[323]), .B(n2251), .Y(n650) );
  INVX1 U1385 ( .A(n650), .Y(n1553) );
  AND2X1 U1386 ( .A(mem[312]), .B(n2252), .Y(n638) );
  INVX1 U1387 ( .A(n638), .Y(n1554) );
  AND2X1 U1388 ( .A(mem[297]), .B(n2253), .Y(n622) );
  INVX1 U1389 ( .A(n622), .Y(n1555) );
  AND2X1 U1390 ( .A(mem[282]), .B(n2254), .Y(n606) );
  INVX1 U1391 ( .A(n606), .Y(n1556) );
  AND2X1 U1392 ( .A(mem[267]), .B(n2255), .Y(n589) );
  INVX1 U1393 ( .A(n589), .Y(n1557) );
  AND2X1 U1394 ( .A(mem[244]), .B(n2256), .Y(n565) );
  INVX1 U1395 ( .A(n565), .Y(n1558) );
  AND2X1 U1396 ( .A(mem[229]), .B(n2257), .Y(n549) );
  INVX1 U1397 ( .A(n549), .Y(n1559) );
  AND2X1 U1398 ( .A(mem[214]), .B(n2258), .Y(n533) );
  INVX1 U1399 ( .A(n533), .Y(n1560) );
  AND2X1 U1400 ( .A(mem[199]), .B(n2259), .Y(n517) );
  INVX1 U1401 ( .A(n517), .Y(n1561) );
  AND2X1 U1402 ( .A(mem[188]), .B(n2260), .Y(n505) );
  INVX1 U1403 ( .A(n505), .Y(n1562) );
  AND2X1 U1404 ( .A(mem[176]), .B(n2260), .Y(n493) );
  INVX1 U1405 ( .A(n493), .Y(n1563) );
  AND2X1 U1406 ( .A(mem[173]), .B(n2261), .Y(n489) );
  INVX1 U1407 ( .A(n489), .Y(n1564) );
  AND2X1 U1408 ( .A(mem[161]), .B(n2261), .Y(n477) );
  INVX1 U1409 ( .A(n477), .Y(n1565) );
  AND2X1 U1410 ( .A(mem[146]), .B(n2262), .Y(n461) );
  INVX1 U1411 ( .A(n461), .Y(n1566) );
  AND2X1 U1412 ( .A(mem[131]), .B(n2263), .Y(n444) );
  INVX1 U1413 ( .A(n444), .Y(n1567) );
  AND2X1 U1414 ( .A(mem[116]), .B(n2264), .Y(n427) );
  INVX1 U1415 ( .A(n427), .Y(n1568) );
  AND2X1 U1416 ( .A(mem[101]), .B(n2265), .Y(n410) );
  INVX1 U1417 ( .A(n410), .Y(n1569) );
  AND2X1 U1418 ( .A(mem[86]), .B(n2266), .Y(n393) );
  INVX1 U1419 ( .A(n393), .Y(n1570) );
  AND2X1 U1420 ( .A(mem[71]), .B(n2267), .Y(n376) );
  INVX1 U1421 ( .A(n376), .Y(n1571) );
  AND2X1 U1422 ( .A(mem[60]), .B(n2268), .Y(n363) );
  INVX1 U1423 ( .A(n363), .Y(n1572) );
  AND2X1 U1424 ( .A(mem[48]), .B(n2268), .Y(n351) );
  INVX1 U1425 ( .A(n351), .Y(n1573) );
  AND2X1 U1426 ( .A(mem[45]), .B(n2269), .Y(n346) );
  INVX1 U1427 ( .A(n346), .Y(n1574) );
  AND2X1 U1428 ( .A(mem[33]), .B(n2269), .Y(n334) );
  INVX1 U1429 ( .A(n334), .Y(n1575) );
  AND2X1 U1430 ( .A(mem[18]), .B(n2270), .Y(n317) );
  INVX1 U1431 ( .A(n317), .Y(n1576) );
  AND2X1 U1432 ( .A(mem[3]), .B(n2271), .Y(n287) );
  INVX1 U1433 ( .A(n287), .Y(n1577) );
  BUFX2 U1434 ( .A(n2314), .Y(empty_bar) );
  BUFX2 U1435 ( .A(n313), .Y(n1579) );
  AND2X1 U1436 ( .A(n74), .B(n2238), .Y(n862) );
  INVX1 U1437 ( .A(n862), .Y(n1580) );
  AND2X1 U1438 ( .A(reset), .B(n1703), .Y(n2238) );
  AND2X1 U1439 ( .A(n21), .B(n855), .Y(n856) );
  INVX1 U1440 ( .A(n856), .Y(n1581) );
  AND2X1 U1441 ( .A(reset), .B(n1660), .Y(n855) );
  AND2X1 U1442 ( .A(mem[505]), .B(n2240), .Y(n844) );
  INVX1 U1443 ( .A(n844), .Y(n1582) );
  AND2X1 U1444 ( .A(mem[488]), .B(n2241), .Y(n826) );
  INVX1 U1445 ( .A(n826), .Y(n1583) );
  AND2X1 U1446 ( .A(mem[475]), .B(n2242), .Y(n812) );
  INVX1 U1447 ( .A(n812), .Y(n1584) );
  AND2X1 U1448 ( .A(mem[458]), .B(n2243), .Y(n794) );
  INVX1 U1449 ( .A(n794), .Y(n1585) );
  AND2X1 U1450 ( .A(mem[437]), .B(n2244), .Y(n772) );
  INVX1 U1451 ( .A(n772), .Y(n1586) );
  AND2X1 U1452 ( .A(mem[420]), .B(n2245), .Y(n754) );
  INVX1 U1453 ( .A(n754), .Y(n1587) );
  AND2X1 U1454 ( .A(mem[407]), .B(n2246), .Y(n740) );
  INVX1 U1455 ( .A(n740), .Y(n1588) );
  AND2X1 U1456 ( .A(mem[390]), .B(n2247), .Y(n721) );
  INVX1 U1457 ( .A(n721), .Y(n1589) );
  AND2X1 U1458 ( .A(mem[381]), .B(n2248), .Y(n711) );
  INVX1 U1459 ( .A(n711), .Y(n1590) );
  AND2X1 U1460 ( .A(mem[369]), .B(n2248), .Y(n699) );
  INVX1 U1461 ( .A(n699), .Y(n1591) );
  AND2X1 U1462 ( .A(mem[364]), .B(n2249), .Y(n693) );
  INVX1 U1463 ( .A(n693), .Y(n1592) );
  AND2X1 U1464 ( .A(mem[352]), .B(n2249), .Y(n681) );
  INVX1 U1465 ( .A(n681), .Y(n1593) );
  AND2X1 U1466 ( .A(mem[339]), .B(n2250), .Y(n667) );
  INVX1 U1467 ( .A(n667), .Y(n1594) );
  AND2X1 U1468 ( .A(mem[322]), .B(n2251), .Y(n649) );
  INVX1 U1469 ( .A(n649), .Y(n1595) );
  AND2X1 U1470 ( .A(mem[313]), .B(n2252), .Y(n639) );
  INVX1 U1471 ( .A(n639), .Y(n1596) );
  AND2X1 U1472 ( .A(mem[296]), .B(n2253), .Y(n621) );
  INVX1 U1473 ( .A(n621), .Y(n1597) );
  AND2X1 U1474 ( .A(mem[283]), .B(n2254), .Y(n607) );
  INVX1 U1475 ( .A(n607), .Y(n1598) );
  AND2X1 U1476 ( .A(mem[266]), .B(n2255), .Y(n588) );
  INVX1 U1477 ( .A(n588), .Y(n1599) );
  AND2X1 U1478 ( .A(mem[245]), .B(n2256), .Y(n566) );
  INVX1 U1479 ( .A(n566), .Y(n1600) );
  AND2X1 U1480 ( .A(mem[228]), .B(n2257), .Y(n548) );
  INVX1 U1481 ( .A(n548), .Y(n1601) );
  AND2X1 U1482 ( .A(mem[215]), .B(n2258), .Y(n534) );
  INVX1 U1483 ( .A(n534), .Y(n1602) );
  AND2X1 U1484 ( .A(mem[198]), .B(n2259), .Y(n516) );
  INVX1 U1485 ( .A(n516), .Y(n1603) );
  AND2X1 U1486 ( .A(mem[189]), .B(n2260), .Y(n506) );
  INVX1 U1487 ( .A(n506), .Y(n1604) );
  AND2X1 U1488 ( .A(mem[177]), .B(n2260), .Y(n494) );
  INVX1 U1489 ( .A(n494), .Y(n1605) );
  AND2X1 U1490 ( .A(mem[172]), .B(n2261), .Y(n488) );
  INVX1 U1491 ( .A(n488), .Y(n1606) );
  AND2X1 U1492 ( .A(mem[160]), .B(n2261), .Y(n476) );
  INVX1 U1493 ( .A(n476), .Y(n1607) );
  AND2X1 U1494 ( .A(mem[147]), .B(n2262), .Y(n462) );
  INVX1 U1495 ( .A(n462), .Y(n1608) );
  AND2X1 U1496 ( .A(mem[130]), .B(n2263), .Y(n443) );
  INVX1 U1497 ( .A(n443), .Y(n1609) );
  AND2X1 U1498 ( .A(mem[117]), .B(n2264), .Y(n428) );
  INVX1 U1499 ( .A(n428), .Y(n1610) );
  AND2X1 U1500 ( .A(mem[100]), .B(n2265), .Y(n409) );
  INVX1 U1501 ( .A(n409), .Y(n1611) );
  AND2X1 U1502 ( .A(mem[87]), .B(n2266), .Y(n394) );
  INVX1 U1503 ( .A(n394), .Y(n1612) );
  AND2X1 U1504 ( .A(mem[70]), .B(n2267), .Y(n375) );
  INVX1 U1505 ( .A(n375), .Y(n1613) );
  AND2X1 U1506 ( .A(mem[61]), .B(n2268), .Y(n364) );
  INVX1 U1507 ( .A(n364), .Y(n1614) );
  AND2X1 U1508 ( .A(mem[49]), .B(n2268), .Y(n352) );
  INVX1 U1509 ( .A(n352), .Y(n1615) );
  AND2X1 U1510 ( .A(mem[44]), .B(n2269), .Y(n345) );
  INVX1 U1511 ( .A(n345), .Y(n1616) );
  AND2X1 U1512 ( .A(mem[32]), .B(n2269), .Y(n333) );
  INVX1 U1513 ( .A(n333), .Y(n1617) );
  AND2X1 U1514 ( .A(mem[19]), .B(n2270), .Y(n318) );
  INVX1 U1515 ( .A(n318), .Y(n1618) );
  AND2X1 U1516 ( .A(mem[2]), .B(n2271), .Y(n285) );
  INVX1 U1517 ( .A(n285), .Y(n1619) );
  BUFX2 U1518 ( .A(n732), .Y(n1620) );
  AND2X1 U1519 ( .A(n75), .B(n2239), .Y(n860) );
  INVX1 U1520 ( .A(n860), .Y(n1621) );
  AND2X1 U1521 ( .A(reset), .B(n1703), .Y(n2239) );
  AND2X1 U1522 ( .A(mem[506]), .B(n2240), .Y(n845) );
  INVX1 U1523 ( .A(n845), .Y(n1622) );
  AND2X1 U1524 ( .A(mem[491]), .B(n2241), .Y(n829) );
  INVX1 U1525 ( .A(n829), .Y(n1623) );
  AND2X1 U1526 ( .A(mem[472]), .B(n2242), .Y(n809) );
  INVX1 U1527 ( .A(n809), .Y(n1624) );
  AND2X1 U1528 ( .A(mem[457]), .B(n2243), .Y(n793) );
  INVX1 U1529 ( .A(n793), .Y(n1625) );
  AND2X1 U1530 ( .A(mem[438]), .B(n2244), .Y(n773) );
  INVX1 U1531 ( .A(n773), .Y(n1626) );
  AND2X1 U1532 ( .A(mem[423]), .B(n2245), .Y(n757) );
  INVX1 U1533 ( .A(n757), .Y(n1627) );
  AND2X1 U1534 ( .A(mem[404]), .B(n2246), .Y(n737) );
  INVX1 U1535 ( .A(n737), .Y(n1628) );
  AND2X1 U1536 ( .A(mem[389]), .B(n2247), .Y(n720) );
  INVX1 U1537 ( .A(n720), .Y(n1629) );
  AND2X1 U1538 ( .A(mem[370]), .B(n2248), .Y(n700) );
  INVX1 U1539 ( .A(n700), .Y(n1630) );
  AND2X1 U1540 ( .A(mem[355]), .B(n2249), .Y(n684) );
  INVX1 U1541 ( .A(n684), .Y(n1631) );
  AND2X1 U1542 ( .A(mem[348]), .B(n2250), .Y(n676) );
  INVX1 U1543 ( .A(n676), .Y(n1632) );
  AND2X1 U1544 ( .A(mem[336]), .B(n2250), .Y(n664) );
  INVX1 U1545 ( .A(n664), .Y(n1633) );
  AND2X1 U1546 ( .A(mem[333]), .B(n2251), .Y(n660) );
  INVX1 U1547 ( .A(n660), .Y(n1634) );
  AND2X1 U1548 ( .A(mem[321]), .B(n2251), .Y(n648) );
  INVX1 U1549 ( .A(n648), .Y(n1635) );
  AND2X1 U1550 ( .A(mem[314]), .B(n2252), .Y(n640) );
  INVX1 U1551 ( .A(n640), .Y(n1636) );
  AND2X1 U1552 ( .A(mem[299]), .B(n2253), .Y(n624) );
  INVX1 U1553 ( .A(n624), .Y(n1637) );
  AND2X1 U1554 ( .A(mem[280]), .B(n2254), .Y(n604) );
  INVX1 U1555 ( .A(n604), .Y(n1638) );
  AND2X1 U1556 ( .A(mem[265]), .B(n2255), .Y(n587) );
  INVX1 U1557 ( .A(n587), .Y(n1639) );
  AND2X1 U1558 ( .A(mem[246]), .B(n2256), .Y(n567) );
  INVX1 U1559 ( .A(n567), .Y(n1640) );
  AND2X1 U1560 ( .A(mem[231]), .B(n2257), .Y(n551) );
  INVX1 U1561 ( .A(n551), .Y(n1641) );
  AND2X1 U1562 ( .A(mem[212]), .B(n2258), .Y(n531) );
  INVX1 U1563 ( .A(n531), .Y(n1642) );
  AND2X1 U1564 ( .A(mem[197]), .B(n2259), .Y(n515) );
  INVX1 U1565 ( .A(n515), .Y(n1643) );
  AND2X1 U1566 ( .A(mem[178]), .B(n2260), .Y(n495) );
  INVX1 U1567 ( .A(n495), .Y(n1644) );
  AND2X1 U1568 ( .A(mem[163]), .B(n2261), .Y(n479) );
  INVX1 U1569 ( .A(n479), .Y(n1645) );
  AND2X1 U1570 ( .A(mem[156]), .B(n2262), .Y(n471) );
  INVX1 U1571 ( .A(n471), .Y(n1646) );
  AND2X1 U1572 ( .A(mem[144]), .B(n2262), .Y(n459) );
  INVX1 U1573 ( .A(n459), .Y(n1647) );
  AND2X1 U1574 ( .A(mem[141]), .B(n2263), .Y(n454) );
  INVX1 U1575 ( .A(n454), .Y(n1648) );
  AND2X1 U1576 ( .A(mem[129]), .B(n2263), .Y(n442) );
  INVX1 U1577 ( .A(n442), .Y(n1649) );
  AND2X1 U1578 ( .A(mem[118]), .B(n2264), .Y(n429) );
  INVX1 U1579 ( .A(n429), .Y(n1650) );
  AND2X1 U1580 ( .A(mem[103]), .B(n2265), .Y(n412) );
  INVX1 U1581 ( .A(n412), .Y(n1651) );
  AND2X1 U1582 ( .A(mem[84]), .B(n2266), .Y(n391) );
  INVX1 U1583 ( .A(n391), .Y(n1652) );
  AND2X1 U1584 ( .A(mem[69]), .B(n2267), .Y(n374) );
  INVX1 U1585 ( .A(n374), .Y(n1653) );
  AND2X1 U1586 ( .A(mem[50]), .B(n2268), .Y(n353) );
  INVX1 U1587 ( .A(n353), .Y(n1654) );
  AND2X1 U1588 ( .A(mem[35]), .B(n2269), .Y(n336) );
  INVX1 U1589 ( .A(n336), .Y(n1655) );
  AND2X1 U1590 ( .A(mem[28]), .B(n2270), .Y(n327) );
  INVX1 U1591 ( .A(n327), .Y(n1656) );
  AND2X1 U1592 ( .A(mem[16]), .B(n2270), .Y(n315) );
  INVX1 U1593 ( .A(n315), .Y(n1657) );
  AND2X1 U1594 ( .A(mem[13]), .B(n2271), .Y(n307) );
  INVX1 U1595 ( .A(n307), .Y(n1658) );
  AND2X1 U1596 ( .A(mem[1]), .B(n2271), .Y(n283) );
  INVX1 U1597 ( .A(n283), .Y(n1659) );
  INVX1 U1598 ( .A(n853), .Y(n1660) );
  BUFX2 U1599 ( .A(n595), .Y(n1661) );
  AND2X1 U1600 ( .A(mem[507]), .B(n2240), .Y(n846) );
  INVX1 U1601 ( .A(n846), .Y(n1662) );
  AND2X1 U1602 ( .A(mem[490]), .B(n2241), .Y(n828) );
  INVX1 U1603 ( .A(n828), .Y(n1663) );
  AND2X1 U1604 ( .A(mem[473]), .B(n2242), .Y(n810) );
  INVX1 U1605 ( .A(n810), .Y(n1664) );
  AND2X1 U1606 ( .A(mem[456]), .B(n2243), .Y(n792) );
  INVX1 U1607 ( .A(n792), .Y(n1665) );
  AND2X1 U1608 ( .A(mem[439]), .B(n2244), .Y(n774) );
  INVX1 U1609 ( .A(n774), .Y(n1666) );
  AND2X1 U1610 ( .A(mem[422]), .B(n2245), .Y(n756) );
  INVX1 U1611 ( .A(n756), .Y(n1667) );
  AND2X1 U1612 ( .A(mem[405]), .B(n2246), .Y(n738) );
  INVX1 U1613 ( .A(n738), .Y(n1668) );
  AND2X1 U1614 ( .A(mem[388]), .B(n2247), .Y(n719) );
  INVX1 U1615 ( .A(n719), .Y(n1669) );
  AND2X1 U1616 ( .A(mem[371]), .B(n2248), .Y(n701) );
  INVX1 U1617 ( .A(n701), .Y(n1670) );
  AND2X1 U1618 ( .A(mem[354]), .B(n2249), .Y(n683) );
  INVX1 U1619 ( .A(n683), .Y(n1671) );
  AND2X1 U1620 ( .A(mem[349]), .B(n2250), .Y(n677) );
  INVX1 U1621 ( .A(n677), .Y(n1672) );
  AND2X1 U1622 ( .A(mem[337]), .B(n2250), .Y(n665) );
  INVX1 U1623 ( .A(n665), .Y(n1673) );
  AND2X1 U1624 ( .A(mem[332]), .B(n2251), .Y(n659) );
  INVX1 U1625 ( .A(n659), .Y(n1674) );
  AND2X1 U1626 ( .A(mem[320]), .B(n2251), .Y(n647) );
  INVX1 U1627 ( .A(n647), .Y(n1675) );
  AND2X1 U1628 ( .A(mem[315]), .B(n2252), .Y(n641) );
  INVX1 U1629 ( .A(n641), .Y(n1676) );
  AND2X1 U1630 ( .A(mem[298]), .B(n2253), .Y(n623) );
  INVX1 U1631 ( .A(n623), .Y(n1677) );
  AND2X1 U1632 ( .A(mem[281]), .B(n2254), .Y(n605) );
  INVX1 U1633 ( .A(n605), .Y(n1678) );
  AND2X1 U1634 ( .A(mem[264]), .B(n2255), .Y(n586) );
  INVX1 U1635 ( .A(n586), .Y(n1679) );
  AND2X1 U1636 ( .A(mem[247]), .B(n2256), .Y(n568) );
  INVX1 U1637 ( .A(n568), .Y(n1680) );
  AND2X1 U1638 ( .A(mem[230]), .B(n2257), .Y(n550) );
  INVX1 U1639 ( .A(n550), .Y(n1681) );
  AND2X1 U1640 ( .A(mem[213]), .B(n2258), .Y(n532) );
  INVX1 U1641 ( .A(n532), .Y(n1682) );
  AND2X1 U1642 ( .A(mem[196]), .B(n2259), .Y(n514) );
  INVX1 U1643 ( .A(n514), .Y(n1683) );
  AND2X1 U1644 ( .A(mem[179]), .B(n2260), .Y(n496) );
  INVX1 U1645 ( .A(n496), .Y(n1684) );
  AND2X1 U1646 ( .A(mem[162]), .B(n2261), .Y(n478) );
  INVX1 U1647 ( .A(n478), .Y(n1685) );
  AND2X1 U1648 ( .A(mem[157]), .B(n2262), .Y(n472) );
  INVX1 U1649 ( .A(n472), .Y(n1686) );
  AND2X1 U1650 ( .A(mem[145]), .B(n2262), .Y(n460) );
  INVX1 U1651 ( .A(n460), .Y(n1687) );
  AND2X1 U1652 ( .A(mem[140]), .B(n2263), .Y(n453) );
  INVX1 U1653 ( .A(n453), .Y(n1688) );
  AND2X1 U1654 ( .A(mem[128]), .B(n2263), .Y(n441) );
  INVX1 U1655 ( .A(n441), .Y(n1689) );
  AND2X1 U1656 ( .A(mem[119]), .B(n2264), .Y(n430) );
  INVX1 U1657 ( .A(n430), .Y(n1690) );
  AND2X1 U1658 ( .A(mem[102]), .B(n2265), .Y(n411) );
  INVX1 U1659 ( .A(n411), .Y(n1691) );
  AND2X1 U1660 ( .A(mem[85]), .B(n2266), .Y(n392) );
  INVX1 U1661 ( .A(n392), .Y(n1692) );
  AND2X1 U1662 ( .A(mem[68]), .B(n2267), .Y(n373) );
  INVX1 U1663 ( .A(n373), .Y(n1693) );
  AND2X1 U1664 ( .A(mem[51]), .B(n2268), .Y(n354) );
  INVX1 U1665 ( .A(n354), .Y(n1694) );
  AND2X1 U1666 ( .A(mem[34]), .B(n2269), .Y(n335) );
  INVX1 U1667 ( .A(n335), .Y(n1695) );
  AND2X1 U1668 ( .A(mem[29]), .B(n2270), .Y(n328) );
  INVX1 U1669 ( .A(n328), .Y(n1696) );
  AND2X1 U1670 ( .A(mem[17]), .B(n2270), .Y(n316) );
  INVX1 U1671 ( .A(n316), .Y(n1697) );
  AND2X1 U1672 ( .A(mem[12]), .B(n2271), .Y(n305) );
  INVX1 U1673 ( .A(n305), .Y(n1698) );
  AND2X1 U1674 ( .A(mem[0]), .B(n2271), .Y(n281) );
  INVX1 U1675 ( .A(n281), .Y(n1699) );
  BUFX2 U1676 ( .A(n2315), .Y(full_bar) );
  OR2X1 U1677 ( .A(fillcount[1]), .B(fillcount[0]), .Y(n884) );
  INVX1 U1678 ( .A(n884), .Y(n1701) );
  BUFX2 U1679 ( .A(n458), .Y(n1702) );
  INVX1 U1680 ( .A(n859), .Y(n1703) );
  INVX1 U1681 ( .A(n882), .Y(n1704) );
  INVX1 U1682 ( .A(n2291), .Y(n2217) );
  INVX1 U1683 ( .A(n2291), .Y(n2218) );
  INVX1 U1684 ( .A(n2291), .Y(n2219) );
  INVX1 U1685 ( .A(n2291), .Y(n2220) );
  INVX1 U1686 ( .A(n2291), .Y(n2221) );
  INVX1 U1687 ( .A(n2291), .Y(n2222) );
  INVX1 U1688 ( .A(n2291), .Y(n2223) );
  INVX1 U1689 ( .A(n2291), .Y(n2224) );
  INVX1 U1690 ( .A(n2291), .Y(n2225) );
  INVX1 U1691 ( .A(n2291), .Y(n2226) );
  INVX1 U1692 ( .A(n2291), .Y(n2227) );
  INVX1 U1693 ( .A(n2291), .Y(n2228) );
  INVX1 U1694 ( .A(n2291), .Y(n2229) );
  INVX1 U1695 ( .A(n2291), .Y(n2230) );
  INVX1 U1696 ( .A(n2291), .Y(n2231) );
  INVX1 U1697 ( .A(n2291), .Y(n2232) );
  INVX1 U1698 ( .A(n2290), .Y(n2236) );
  INVX1 U1699 ( .A(n2290), .Y(n2237) );
  INVX1 U1700 ( .A(n2291), .Y(n2233) );
  INVX1 U1701 ( .A(n2291), .Y(n2234) );
  INVX1 U1702 ( .A(n2291), .Y(n2235) );
  INVX1 U1703 ( .A(n312), .Y(n2271) );
  INVX1 U1704 ( .A(n663), .Y(n2251) );
  INVX1 U1705 ( .A(n680), .Y(n2250) );
  INVX1 U1706 ( .A(n697), .Y(n2249) );
  INVX1 U1707 ( .A(n714), .Y(n2248) );
  INVX1 U1708 ( .A(n731), .Y(n2247) );
  INVX1 U1709 ( .A(n749), .Y(n2246) );
  INVX1 U1710 ( .A(n766), .Y(n2245) );
  INVX1 U1711 ( .A(n783), .Y(n2244) );
  INVX1 U1712 ( .A(n800), .Y(n2243) );
  INVX1 U1713 ( .A(n817), .Y(n2242) );
  INVX1 U1714 ( .A(n834), .Y(n2241) );
  INVX1 U1715 ( .A(n331), .Y(n2270) );
  INVX1 U1716 ( .A(n349), .Y(n2269) );
  INVX1 U1717 ( .A(n367), .Y(n2268) );
  INVX1 U1718 ( .A(n385), .Y(n2267) );
  INVX1 U1719 ( .A(n403), .Y(n2266) );
  INVX1 U1720 ( .A(n421), .Y(n2265) );
  INVX1 U1721 ( .A(n439), .Y(n2264) );
  INVX1 U1722 ( .A(n457), .Y(n2263) );
  INVX1 U1723 ( .A(n475), .Y(n2262) );
  INVX1 U1724 ( .A(n492), .Y(n2261) );
  INVX1 U1725 ( .A(n509), .Y(n2260) );
  INVX1 U1726 ( .A(n526), .Y(n2259) );
  INVX1 U1727 ( .A(n543), .Y(n2258) );
  INVX1 U1728 ( .A(n560), .Y(n2257) );
  INVX1 U1729 ( .A(n577), .Y(n2256) );
  INVX1 U1730 ( .A(n594), .Y(n2255) );
  INVX1 U1731 ( .A(n612), .Y(n2254) );
  INVX1 U1732 ( .A(n629), .Y(n2253) );
  INVX1 U1733 ( .A(n646), .Y(n2252) );
  INVX1 U1734 ( .A(n851), .Y(n2240) );
  INVX1 U1735 ( .A(sub_93_carry[5]), .Y(fillcount[5]) );
  INVX1 U1736 ( .A(n1705), .Y(n2282) );
  INVX1 U1737 ( .A(n1706), .Y(n2281) );
  INVX1 U1738 ( .A(n1707), .Y(n2280) );
  INVX1 U1739 ( .A(n1708), .Y(n2279) );
  INVX1 U1740 ( .A(n1709), .Y(n2278) );
  INVX1 U1741 ( .A(n1710), .Y(n2277) );
  INVX1 U1742 ( .A(n1711), .Y(n2276) );
  INVX1 U1743 ( .A(n1712), .Y(n2275) );
  INVX1 U1744 ( .A(n1713), .Y(n2274) );
  INVX1 U1745 ( .A(n1714), .Y(n2273) );
  INVX1 U1746 ( .A(n1715), .Y(n2272) );
  INVX1 U1747 ( .A(n1716), .Y(n2287) );
  INVX1 U1748 ( .A(n1717), .Y(n2286) );
  INVX1 U1749 ( .A(n1718), .Y(n2285) );
  INVX1 U1750 ( .A(n1719), .Y(n2284) );
  INVX1 U1751 ( .A(n1720), .Y(n2283) );
  INVX1 U1752 ( .A(n16), .Y(n2292) );
  INVX1 U1753 ( .A(n12), .Y(n2291) );
  INVX1 U1754 ( .A(wr_ptr[2]), .Y(n2312) );
  INVX1 U1755 ( .A(wr_ptr[0]), .Y(n2309) );
  INVX1 U1756 ( .A(n1), .Y(n2293) );
  INVX1 U1757 ( .A(n2201), .Y(n71) );
  INVX1 U1758 ( .A(n2), .Y(n2294) );
  INVX1 U1759 ( .A(n2202), .Y(n70) );
  INVX1 U1760 ( .A(n3), .Y(n2295) );
  INVX1 U1761 ( .A(n2203), .Y(n69) );
  INVX1 U1762 ( .A(n4), .Y(n2296) );
  INVX1 U1763 ( .A(n2204), .Y(n68) );
  INVX1 U1764 ( .A(n5), .Y(n2297) );
  INVX1 U1765 ( .A(n2205), .Y(n67) );
  INVX1 U1766 ( .A(n6), .Y(n2298) );
  INVX1 U1767 ( .A(n2206), .Y(n66) );
  INVX1 U1768 ( .A(n7), .Y(n2299) );
  INVX1 U1769 ( .A(n2207), .Y(n65) );
  INVX1 U1770 ( .A(n8), .Y(n2300) );
  INVX1 U1771 ( .A(n2208), .Y(n64) );
  INVX1 U1772 ( .A(n9), .Y(n2301) );
  INVX1 U1773 ( .A(n2209), .Y(n63) );
  INVX1 U1774 ( .A(n10), .Y(n2302) );
  INVX1 U1775 ( .A(n2210), .Y(n62) );
  INVX1 U1776 ( .A(n11), .Y(n2303) );
  INVX1 U1777 ( .A(n2211), .Y(n61) );
  INVX1 U1778 ( .A(n17), .Y(n2304) );
  INVX1 U1779 ( .A(n2212), .Y(n60) );
  INVX1 U1780 ( .A(n18), .Y(n2305) );
  INVX1 U1781 ( .A(n2213), .Y(n59) );
  INVX1 U1782 ( .A(n19), .Y(n2306) );
  INVX1 U1783 ( .A(n2214), .Y(n58) );
  INVX1 U1784 ( .A(n24), .Y(n2307) );
  INVX1 U1785 ( .A(n2215), .Y(n57) );
  INVX1 U1786 ( .A(n25), .Y(n2308) );
  INVX1 U1787 ( .A(n2216), .Y(n56) );
  INVX1 U1788 ( .A(wr_ptr[1]), .Y(n2311) );
  INVX1 U1789 ( .A(wr_ptr[3]), .Y(n2313) );
  INVX1 U1790 ( .A(wr_ptr[4]), .Y(n2310) );
  AND2X1 U1791 ( .A(data_in[5]), .B(reset), .Y(n1705) );
  AND2X1 U1792 ( .A(data_in[6]), .B(reset), .Y(n1706) );
  AND2X1 U1793 ( .A(data_in[7]), .B(reset), .Y(n1707) );
  AND2X1 U1794 ( .A(data_in[8]), .B(reset), .Y(n1708) );
  AND2X1 U1795 ( .A(data_in[9]), .B(reset), .Y(n1709) );
  AND2X1 U1796 ( .A(data_in[10]), .B(reset), .Y(n1710) );
  AND2X1 U1797 ( .A(data_in[11]), .B(reset), .Y(n1711) );
  AND2X1 U1798 ( .A(data_in[12]), .B(reset), .Y(n1712) );
  AND2X1 U1799 ( .A(data_in[13]), .B(reset), .Y(n1713) );
  AND2X1 U1800 ( .A(data_in[14]), .B(reset), .Y(n1714) );
  AND2X1 U1801 ( .A(data_in[15]), .B(reset), .Y(n1715) );
  AND2X1 U1802 ( .A(data_in[0]), .B(reset), .Y(n1716) );
  AND2X1 U1803 ( .A(data_in[1]), .B(reset), .Y(n1717) );
  AND2X1 U1804 ( .A(data_in[2]), .B(reset), .Y(n1718) );
  AND2X1 U1805 ( .A(data_in[3]), .B(reset), .Y(n1719) );
  AND2X1 U1806 ( .A(data_in[4]), .B(reset), .Y(n1720) );
  INVX1 U1807 ( .A(n13), .Y(n2290) );
  INVX1 U1808 ( .A(n14), .Y(n2289) );
  INVX1 U1809 ( .A(n15), .Y(n2288) );
  MUX2X1 U1810 ( .B(n1722), .A(n1723), .S(n13), .Y(n1721) );
  MUX2X1 U1811 ( .B(n1725), .A(n1726), .S(n2237), .Y(n1724) );
  MUX2X1 U1812 ( .B(n1728), .A(n1729), .S(n2236), .Y(n1727) );
  MUX2X1 U1813 ( .B(n1731), .A(n1732), .S(n13), .Y(n1730) );
  MUX2X1 U1814 ( .B(n1734), .A(n1735), .S(n15), .Y(n1733) );
  MUX2X1 U1815 ( .B(n1737), .A(n1738), .S(n13), .Y(n1736) );
  MUX2X1 U1816 ( .B(n1740), .A(n1741), .S(n2236), .Y(n1739) );
  MUX2X1 U1817 ( .B(n1743), .A(n1744), .S(n2237), .Y(n1742) );
  MUX2X1 U1818 ( .B(n1746), .A(n1747), .S(n13), .Y(n1745) );
  MUX2X1 U1819 ( .B(n1749), .A(n1750), .S(n15), .Y(n1748) );
  MUX2X1 U1820 ( .B(n1752), .A(n1753), .S(n2236), .Y(n1751) );
  MUX2X1 U1821 ( .B(n1755), .A(n1756), .S(n2236), .Y(n1754) );
  MUX2X1 U1822 ( .B(n1758), .A(n1759), .S(n2236), .Y(n1757) );
  MUX2X1 U1823 ( .B(n1761), .A(n1762), .S(n2236), .Y(n1760) );
  MUX2X1 U1824 ( .B(n1764), .A(n1765), .S(n15), .Y(n1763) );
  MUX2X1 U1825 ( .B(n1767), .A(n1768), .S(n2236), .Y(n1766) );
  MUX2X1 U1826 ( .B(n1770), .A(n1771), .S(n2236), .Y(n1769) );
  MUX2X1 U1827 ( .B(n1773), .A(n1774), .S(n2236), .Y(n1772) );
  MUX2X1 U1828 ( .B(n1776), .A(n1777), .S(n2236), .Y(n1775) );
  MUX2X1 U1829 ( .B(n1779), .A(n1780), .S(n15), .Y(n1778) );
  MUX2X1 U1830 ( .B(n1782), .A(n1783), .S(n2236), .Y(n1781) );
  MUX2X1 U1831 ( .B(n1785), .A(n1786), .S(n2236), .Y(n1784) );
  MUX2X1 U1832 ( .B(n1788), .A(n1789), .S(n2236), .Y(n1787) );
  MUX2X1 U1833 ( .B(n1791), .A(n1792), .S(n2236), .Y(n1790) );
  MUX2X1 U1834 ( .B(n1794), .A(n1795), .S(n15), .Y(n1793) );
  MUX2X1 U1835 ( .B(n1797), .A(n1798), .S(n2236), .Y(n1796) );
  MUX2X1 U1836 ( .B(n1800), .A(n1801), .S(n2236), .Y(n1799) );
  MUX2X1 U1837 ( .B(n1803), .A(n1804), .S(n2236), .Y(n1802) );
  MUX2X1 U1838 ( .B(n1806), .A(n1807), .S(n2237), .Y(n1805) );
  MUX2X1 U1839 ( .B(n1809), .A(n1810), .S(n15), .Y(n1808) );
  MUX2X1 U1840 ( .B(n1812), .A(n1813), .S(n2237), .Y(n1811) );
  MUX2X1 U1841 ( .B(n1815), .A(n1816), .S(n13), .Y(n1814) );
  MUX2X1 U1842 ( .B(n1818), .A(n1819), .S(n2236), .Y(n1817) );
  MUX2X1 U1843 ( .B(n1821), .A(n1822), .S(n2236), .Y(n1820) );
  MUX2X1 U1844 ( .B(n1824), .A(n1825), .S(n15), .Y(n1823) );
  MUX2X1 U1845 ( .B(n1827), .A(n1828), .S(n13), .Y(n1826) );
  MUX2X1 U1846 ( .B(n1830), .A(n1831), .S(n2237), .Y(n1829) );
  MUX2X1 U1847 ( .B(n1833), .A(n1834), .S(n13), .Y(n1832) );
  MUX2X1 U1848 ( .B(n1836), .A(n1837), .S(n13), .Y(n1835) );
  MUX2X1 U1849 ( .B(n1839), .A(n1840), .S(n15), .Y(n1838) );
  MUX2X1 U1850 ( .B(n1842), .A(n1843), .S(n2237), .Y(n1841) );
  MUX2X1 U1851 ( .B(n1845), .A(n1846), .S(n2237), .Y(n1844) );
  MUX2X1 U1852 ( .B(n1848), .A(n1849), .S(n2237), .Y(n1847) );
  MUX2X1 U1853 ( .B(n1851), .A(n1852), .S(n2237), .Y(n1850) );
  MUX2X1 U1854 ( .B(n1854), .A(n1855), .S(n15), .Y(n1853) );
  MUX2X1 U1855 ( .B(n1857), .A(n1858), .S(n2237), .Y(n1856) );
  MUX2X1 U1856 ( .B(n1860), .A(n1861), .S(n2237), .Y(n1859) );
  MUX2X1 U1857 ( .B(n1863), .A(n1864), .S(n2237), .Y(n1862) );
  MUX2X1 U1858 ( .B(n1866), .A(n1867), .S(n2237), .Y(n1865) );
  MUX2X1 U1859 ( .B(n1869), .A(n1870), .S(n15), .Y(n1868) );
  MUX2X1 U1860 ( .B(n1872), .A(n1873), .S(n2237), .Y(n1871) );
  MUX2X1 U1861 ( .B(n1875), .A(n1876), .S(n2237), .Y(n1874) );
  MUX2X1 U1862 ( .B(n1878), .A(n1879), .S(n2237), .Y(n1877) );
  MUX2X1 U1863 ( .B(n1881), .A(n1882), .S(n2237), .Y(n1880) );
  MUX2X1 U1864 ( .B(n1884), .A(n1885), .S(n15), .Y(n1883) );
  MUX2X1 U1865 ( .B(n1887), .A(n1888), .S(n13), .Y(n1886) );
  MUX2X1 U1866 ( .B(n1890), .A(n1891), .S(n13), .Y(n1889) );
  MUX2X1 U1867 ( .B(n1893), .A(n1894), .S(n13), .Y(n1892) );
  MUX2X1 U1868 ( .B(n1896), .A(n1897), .S(n13), .Y(n1895) );
  MUX2X1 U1869 ( .B(n1899), .A(n1900), .S(n15), .Y(n1898) );
  MUX2X1 U1870 ( .B(n1902), .A(n1903), .S(n13), .Y(n1901) );
  MUX2X1 U1871 ( .B(n1905), .A(n1906), .S(n13), .Y(n1904) );
  MUX2X1 U1872 ( .B(n1908), .A(n1909), .S(n13), .Y(n1907) );
  MUX2X1 U1873 ( .B(n1911), .A(n1912), .S(n13), .Y(n1910) );
  MUX2X1 U1874 ( .B(n1914), .A(n1915), .S(n15), .Y(n1913) );
  MUX2X1 U1875 ( .B(n1917), .A(n1918), .S(n13), .Y(n1916) );
  MUX2X1 U1876 ( .B(n1920), .A(n1921), .S(n13), .Y(n1919) );
  MUX2X1 U1877 ( .B(n1923), .A(n1924), .S(n13), .Y(n1922) );
  MUX2X1 U1878 ( .B(n1926), .A(n1927), .S(n13), .Y(n1925) );
  MUX2X1 U1879 ( .B(n1929), .A(n1930), .S(n15), .Y(n1928) );
  MUX2X1 U1880 ( .B(n1932), .A(n1933), .S(n2236), .Y(n1931) );
  MUX2X1 U1881 ( .B(n1935), .A(n1936), .S(n2237), .Y(n1934) );
  MUX2X1 U1882 ( .B(n1938), .A(n1939), .S(n13), .Y(n1937) );
  MUX2X1 U1883 ( .B(n1941), .A(n1942), .S(n13), .Y(n1940) );
  MUX2X1 U1884 ( .B(n1944), .A(n1945), .S(n15), .Y(n1943) );
  MUX2X1 U1885 ( .B(n1947), .A(n1948), .S(n2237), .Y(n1946) );
  MUX2X1 U1886 ( .B(n1950), .A(n1951), .S(n2237), .Y(n1949) );
  MUX2X1 U1887 ( .B(n1953), .A(n1954), .S(n13), .Y(n1952) );
  MUX2X1 U1888 ( .B(n1956), .A(n1957), .S(n2237), .Y(n1955) );
  MUX2X1 U1889 ( .B(n1959), .A(n1960), .S(n15), .Y(n1958) );
  MUX2X1 U1890 ( .B(n1962), .A(n1963), .S(n13), .Y(n1961) );
  MUX2X1 U1891 ( .B(n1965), .A(n1966), .S(n13), .Y(n1964) );
  MUX2X1 U1892 ( .B(n1968), .A(n1969), .S(n2236), .Y(n1967) );
  MUX2X1 U1893 ( .B(n1971), .A(n1972), .S(n2237), .Y(n1970) );
  MUX2X1 U1894 ( .B(n1974), .A(n1975), .S(n15), .Y(n1973) );
  MUX2X1 U1895 ( .B(n1977), .A(n1978), .S(n13), .Y(n1976) );
  MUX2X1 U1896 ( .B(n1980), .A(n1981), .S(n13), .Y(n1979) );
  MUX2X1 U1897 ( .B(n1983), .A(n1984), .S(n13), .Y(n1982) );
  MUX2X1 U1898 ( .B(n1986), .A(n1987), .S(n13), .Y(n1985) );
  MUX2X1 U1899 ( .B(n1989), .A(n1990), .S(n15), .Y(n1988) );
  MUX2X1 U1900 ( .B(n1992), .A(n1993), .S(n13), .Y(n1991) );
  MUX2X1 U1901 ( .B(n1995), .A(n1996), .S(n13), .Y(n1994) );
  MUX2X1 U1902 ( .B(n1998), .A(n1999), .S(n13), .Y(n1997) );
  MUX2X1 U1903 ( .B(n2001), .A(n2002), .S(n13), .Y(n2000) );
  MUX2X1 U1904 ( .B(n2004), .A(n2005), .S(n15), .Y(n2003) );
  MUX2X1 U1905 ( .B(n2007), .A(n2008), .S(n13), .Y(n2006) );
  MUX2X1 U1906 ( .B(n2010), .A(n2011), .S(n2236), .Y(n2009) );
  MUX2X1 U1907 ( .B(n2013), .A(n2014), .S(n13), .Y(n2012) );
  MUX2X1 U1908 ( .B(n2016), .A(n2017), .S(n13), .Y(n2015) );
  MUX2X1 U1909 ( .B(n2019), .A(n2020), .S(n15), .Y(n2018) );
  MUX2X1 U1910 ( .B(n2022), .A(n2023), .S(n13), .Y(n2021) );
  MUX2X1 U1911 ( .B(n2025), .A(n2026), .S(n2237), .Y(n2024) );
  MUX2X1 U1912 ( .B(n2028), .A(n2029), .S(n13), .Y(n2027) );
  MUX2X1 U1913 ( .B(n2031), .A(n2032), .S(n13), .Y(n2030) );
  MUX2X1 U1914 ( .B(n2034), .A(n2035), .S(n15), .Y(n2033) );
  MUX2X1 U1915 ( .B(n2037), .A(n2038), .S(n13), .Y(n2036) );
  MUX2X1 U1916 ( .B(n2040), .A(n2041), .S(n2237), .Y(n2039) );
  MUX2X1 U1917 ( .B(n2043), .A(n2044), .S(n13), .Y(n2042) );
  MUX2X1 U1918 ( .B(n2046), .A(n2047), .S(n13), .Y(n2045) );
  MUX2X1 U1919 ( .B(n2049), .A(n2050), .S(n15), .Y(n2048) );
  MUX2X1 U1920 ( .B(n2052), .A(n2053), .S(n13), .Y(n2051) );
  MUX2X1 U1921 ( .B(n2055), .A(n2056), .S(n13), .Y(n2054) );
  MUX2X1 U1922 ( .B(n2058), .A(n2059), .S(n2236), .Y(n2057) );
  MUX2X1 U1923 ( .B(n2061), .A(n2062), .S(n2236), .Y(n2060) );
  MUX2X1 U1924 ( .B(n2064), .A(n2065), .S(n15), .Y(n2063) );
  MUX2X1 U1925 ( .B(n2067), .A(n2068), .S(n2236), .Y(n2066) );
  MUX2X1 U1926 ( .B(n2070), .A(n2071), .S(n13), .Y(n2069) );
  MUX2X1 U1927 ( .B(n2073), .A(n2074), .S(n2236), .Y(n2072) );
  MUX2X1 U1928 ( .B(n2076), .A(n2077), .S(n2236), .Y(n2075) );
  MUX2X1 U1929 ( .B(n2079), .A(n2080), .S(n15), .Y(n2078) );
  MUX2X1 U1930 ( .B(n2082), .A(n2083), .S(n13), .Y(n2081) );
  MUX2X1 U1931 ( .B(n2085), .A(n2086), .S(n2237), .Y(n2084) );
  MUX2X1 U1932 ( .B(n2088), .A(n2089), .S(n2237), .Y(n2087) );
  MUX2X1 U1933 ( .B(n2091), .A(n2092), .S(n2236), .Y(n2090) );
  MUX2X1 U1934 ( .B(n2094), .A(n2095), .S(n15), .Y(n2093) );
  MUX2X1 U1935 ( .B(n2097), .A(n2098), .S(n2236), .Y(n2096) );
  MUX2X1 U1936 ( .B(n2100), .A(n2101), .S(n13), .Y(n2099) );
  MUX2X1 U1937 ( .B(n2103), .A(n2104), .S(n13), .Y(n2102) );
  MUX2X1 U1938 ( .B(n2106), .A(n2107), .S(n13), .Y(n2105) );
  MUX2X1 U1939 ( .B(n2109), .A(n2110), .S(n15), .Y(n2108) );
  MUX2X1 U1940 ( .B(n2112), .A(n2113), .S(n13), .Y(n2111) );
  MUX2X1 U1941 ( .B(n2115), .A(n2116), .S(n2236), .Y(n2114) );
  MUX2X1 U1942 ( .B(n2118), .A(n2119), .S(n2237), .Y(n2117) );
  MUX2X1 U1943 ( .B(n2121), .A(n2122), .S(n2236), .Y(n2120) );
  MUX2X1 U1944 ( .B(n2124), .A(n2125), .S(n15), .Y(n2123) );
  MUX2X1 U1945 ( .B(n2127), .A(n2128), .S(n2236), .Y(n2126) );
  MUX2X1 U1946 ( .B(n2130), .A(n2131), .S(n2237), .Y(n2129) );
  MUX2X1 U1947 ( .B(n2133), .A(n2134), .S(n13), .Y(n2132) );
  MUX2X1 U1948 ( .B(n2136), .A(n2137), .S(n13), .Y(n2135) );
  MUX2X1 U1949 ( .B(n2139), .A(n2140), .S(n15), .Y(n2138) );
  MUX2X1 U1950 ( .B(n2142), .A(n2143), .S(n2237), .Y(n2141) );
  MUX2X1 U1951 ( .B(n2145), .A(n2146), .S(n13), .Y(n2144) );
  MUX2X1 U1952 ( .B(n2148), .A(n2149), .S(n2237), .Y(n2147) );
  MUX2X1 U1953 ( .B(n2151), .A(n2152), .S(n2237), .Y(n2150) );
  MUX2X1 U1954 ( .B(n2154), .A(n2155), .S(n15), .Y(n2153) );
  MUX2X1 U1955 ( .B(n2157), .A(n2158), .S(n13), .Y(n2156) );
  MUX2X1 U1956 ( .B(n2160), .A(n2161), .S(n13), .Y(n2159) );
  MUX2X1 U1957 ( .B(n2163), .A(n2164), .S(n13), .Y(n2162) );
  MUX2X1 U1958 ( .B(n2166), .A(n2167), .S(n2236), .Y(n2165) );
  MUX2X1 U1959 ( .B(n2169), .A(n2170), .S(n15), .Y(n2168) );
  MUX2X1 U1960 ( .B(n2172), .A(n2173), .S(n2237), .Y(n2171) );
  MUX2X1 U1961 ( .B(n2175), .A(n2176), .S(n13), .Y(n2174) );
  MUX2X1 U1962 ( .B(n2178), .A(n2179), .S(n2236), .Y(n2177) );
  MUX2X1 U1963 ( .B(n2181), .A(n2182), .S(n13), .Y(n2180) );
  MUX2X1 U1964 ( .B(n2184), .A(n2185), .S(n15), .Y(n2183) );
  MUX2X1 U1965 ( .B(n2187), .A(n2188), .S(n13), .Y(n2186) );
  MUX2X1 U1966 ( .B(n2190), .A(n2191), .S(n13), .Y(n2189) );
  MUX2X1 U1967 ( .B(n2193), .A(n2194), .S(n2237), .Y(n2192) );
  MUX2X1 U1968 ( .B(n2196), .A(n2197), .S(n2237), .Y(n2195) );
  MUX2X1 U1969 ( .B(n2199), .A(n2200), .S(n15), .Y(n2198) );
  MUX2X1 U1970 ( .B(mem[480]), .A(mem[496]), .S(n2220), .Y(n1723) );
  MUX2X1 U1971 ( .B(mem[448]), .A(mem[464]), .S(n2229), .Y(n1722) );
  MUX2X1 U1972 ( .B(mem[416]), .A(mem[432]), .S(n2227), .Y(n1726) );
  MUX2X1 U1973 ( .B(mem[384]), .A(mem[400]), .S(n2231), .Y(n1725) );
  MUX2X1 U1974 ( .B(n1724), .A(n1721), .S(n14), .Y(n1735) );
  MUX2X1 U1975 ( .B(mem[352]), .A(mem[368]), .S(n2217), .Y(n1729) );
  MUX2X1 U1976 ( .B(mem[320]), .A(mem[336]), .S(n2217), .Y(n1728) );
  MUX2X1 U1977 ( .B(mem[288]), .A(mem[304]), .S(n2217), .Y(n1732) );
  MUX2X1 U1978 ( .B(mem[256]), .A(mem[272]), .S(n2217), .Y(n1731) );
  MUX2X1 U1979 ( .B(n1730), .A(n1727), .S(n14), .Y(n1734) );
  MUX2X1 U1980 ( .B(mem[224]), .A(mem[240]), .S(n2217), .Y(n1738) );
  MUX2X1 U1981 ( .B(mem[192]), .A(mem[208]), .S(n2217), .Y(n1737) );
  MUX2X1 U1982 ( .B(mem[160]), .A(mem[176]), .S(n2217), .Y(n1741) );
  MUX2X1 U1983 ( .B(mem[128]), .A(mem[144]), .S(n2217), .Y(n1740) );
  MUX2X1 U1984 ( .B(n1739), .A(n1736), .S(n14), .Y(n1750) );
  MUX2X1 U1985 ( .B(mem[96]), .A(mem[112]), .S(n2217), .Y(n1744) );
  MUX2X1 U1986 ( .B(mem[64]), .A(mem[80]), .S(n2217), .Y(n1743) );
  MUX2X1 U1987 ( .B(mem[32]), .A(mem[48]), .S(n2217), .Y(n1747) );
  MUX2X1 U1988 ( .B(mem[0]), .A(mem[16]), .S(n2217), .Y(n1746) );
  MUX2X1 U1989 ( .B(n1745), .A(n1742), .S(n14), .Y(n1749) );
  MUX2X1 U1990 ( .B(n1748), .A(n1733), .S(n16), .Y(n2201) );
  MUX2X1 U1991 ( .B(mem[481]), .A(mem[497]), .S(n2218), .Y(n1753) );
  MUX2X1 U1992 ( .B(mem[449]), .A(mem[465]), .S(n2218), .Y(n1752) );
  MUX2X1 U1993 ( .B(mem[417]), .A(mem[433]), .S(n2218), .Y(n1756) );
  MUX2X1 U1994 ( .B(mem[385]), .A(mem[401]), .S(n2218), .Y(n1755) );
  MUX2X1 U1995 ( .B(n1754), .A(n1751), .S(n14), .Y(n1765) );
  MUX2X1 U1996 ( .B(mem[353]), .A(mem[369]), .S(n2218), .Y(n1759) );
  MUX2X1 U1997 ( .B(mem[321]), .A(mem[337]), .S(n2218), .Y(n1758) );
  MUX2X1 U1998 ( .B(mem[289]), .A(mem[305]), .S(n2218), .Y(n1762) );
  MUX2X1 U1999 ( .B(mem[257]), .A(mem[273]), .S(n2218), .Y(n1761) );
  MUX2X1 U2000 ( .B(n1760), .A(n1757), .S(n14), .Y(n1764) );
  MUX2X1 U2001 ( .B(mem[225]), .A(mem[241]), .S(n2218), .Y(n1768) );
  MUX2X1 U2002 ( .B(mem[193]), .A(mem[209]), .S(n2218), .Y(n1767) );
  MUX2X1 U2003 ( .B(mem[161]), .A(mem[177]), .S(n2218), .Y(n1771) );
  MUX2X1 U2004 ( .B(mem[129]), .A(mem[145]), .S(n2218), .Y(n1770) );
  MUX2X1 U2005 ( .B(n1769), .A(n1766), .S(n14), .Y(n1780) );
  MUX2X1 U2006 ( .B(mem[97]), .A(mem[113]), .S(n2219), .Y(n1774) );
  MUX2X1 U2007 ( .B(mem[65]), .A(mem[81]), .S(n2219), .Y(n1773) );
  MUX2X1 U2008 ( .B(mem[33]), .A(mem[49]), .S(n2219), .Y(n1777) );
  MUX2X1 U2009 ( .B(mem[1]), .A(mem[17]), .S(n2219), .Y(n1776) );
  MUX2X1 U2010 ( .B(n1775), .A(n1772), .S(n14), .Y(n1779) );
  MUX2X1 U2011 ( .B(n1778), .A(n1763), .S(n16), .Y(n2202) );
  MUX2X1 U2012 ( .B(mem[482]), .A(mem[498]), .S(n2219), .Y(n1783) );
  MUX2X1 U2013 ( .B(mem[450]), .A(mem[466]), .S(n2219), .Y(n1782) );
  MUX2X1 U2014 ( .B(mem[418]), .A(mem[434]), .S(n2219), .Y(n1786) );
  MUX2X1 U2015 ( .B(mem[386]), .A(mem[402]), .S(n2219), .Y(n1785) );
  MUX2X1 U2016 ( .B(n1784), .A(n1781), .S(n14), .Y(n1795) );
  MUX2X1 U2017 ( .B(mem[354]), .A(mem[370]), .S(n2219), .Y(n1789) );
  MUX2X1 U2018 ( .B(mem[322]), .A(mem[338]), .S(n2219), .Y(n1788) );
  MUX2X1 U2019 ( .B(mem[290]), .A(mem[306]), .S(n2219), .Y(n1792) );
  MUX2X1 U2020 ( .B(mem[258]), .A(mem[274]), .S(n2219), .Y(n1791) );
  MUX2X1 U2021 ( .B(n1790), .A(n1787), .S(n14), .Y(n1794) );
  MUX2X1 U2022 ( .B(mem[226]), .A(mem[242]), .S(n2220), .Y(n1798) );
  MUX2X1 U2023 ( .B(mem[194]), .A(mem[210]), .S(n2220), .Y(n1797) );
  MUX2X1 U2024 ( .B(mem[162]), .A(mem[178]), .S(n2220), .Y(n1801) );
  MUX2X1 U2025 ( .B(mem[130]), .A(mem[146]), .S(n2220), .Y(n1800) );
  MUX2X1 U2026 ( .B(n1799), .A(n1796), .S(n14), .Y(n1810) );
  MUX2X1 U2027 ( .B(mem[98]), .A(mem[114]), .S(n2220), .Y(n1804) );
  MUX2X1 U2028 ( .B(mem[66]), .A(mem[82]), .S(n2220), .Y(n1803) );
  MUX2X1 U2029 ( .B(mem[34]), .A(mem[50]), .S(n2220), .Y(n1807) );
  MUX2X1 U2030 ( .B(mem[2]), .A(mem[18]), .S(n2220), .Y(n1806) );
  MUX2X1 U2031 ( .B(n1805), .A(n1802), .S(n14), .Y(n1809) );
  MUX2X1 U2032 ( .B(n1808), .A(n1793), .S(n16), .Y(n2203) );
  MUX2X1 U2033 ( .B(mem[483]), .A(mem[499]), .S(n2220), .Y(n1813) );
  MUX2X1 U2034 ( .B(mem[451]), .A(mem[467]), .S(n2220), .Y(n1812) );
  MUX2X1 U2035 ( .B(mem[419]), .A(mem[435]), .S(n2220), .Y(n1816) );
  MUX2X1 U2036 ( .B(mem[387]), .A(mem[403]), .S(n2220), .Y(n1815) );
  MUX2X1 U2037 ( .B(n1814), .A(n1811), .S(n14), .Y(n1825) );
  MUX2X1 U2038 ( .B(mem[355]), .A(mem[371]), .S(n2221), .Y(n1819) );
  MUX2X1 U2039 ( .B(mem[323]), .A(mem[339]), .S(n2221), .Y(n1818) );
  MUX2X1 U2040 ( .B(mem[291]), .A(mem[307]), .S(n2221), .Y(n1822) );
  MUX2X1 U2041 ( .B(mem[259]), .A(mem[275]), .S(n2221), .Y(n1821) );
  MUX2X1 U2042 ( .B(n1820), .A(n1817), .S(n14), .Y(n1824) );
  MUX2X1 U2043 ( .B(mem[227]), .A(mem[243]), .S(n2221), .Y(n1828) );
  MUX2X1 U2044 ( .B(mem[195]), .A(mem[211]), .S(n2221), .Y(n1827) );
  MUX2X1 U2045 ( .B(mem[163]), .A(mem[179]), .S(n2221), .Y(n1831) );
  MUX2X1 U2046 ( .B(mem[131]), .A(mem[147]), .S(n2221), .Y(n1830) );
  MUX2X1 U2047 ( .B(n1829), .A(n1826), .S(n14), .Y(n1840) );
  MUX2X1 U2048 ( .B(mem[99]), .A(mem[115]), .S(n2221), .Y(n1834) );
  MUX2X1 U2049 ( .B(mem[67]), .A(mem[83]), .S(n2221), .Y(n1833) );
  MUX2X1 U2050 ( .B(mem[35]), .A(mem[51]), .S(n2221), .Y(n1837) );
  MUX2X1 U2051 ( .B(mem[3]), .A(mem[19]), .S(n2221), .Y(n1836) );
  MUX2X1 U2052 ( .B(n1835), .A(n1832), .S(n14), .Y(n1839) );
  MUX2X1 U2053 ( .B(n1838), .A(n1823), .S(n16), .Y(n2204) );
  MUX2X1 U2054 ( .B(mem[484]), .A(mem[500]), .S(n2222), .Y(n1843) );
  MUX2X1 U2055 ( .B(mem[452]), .A(mem[468]), .S(n2222), .Y(n1842) );
  MUX2X1 U2056 ( .B(mem[420]), .A(mem[436]), .S(n2222), .Y(n1846) );
  MUX2X1 U2057 ( .B(mem[388]), .A(mem[404]), .S(n2222), .Y(n1845) );
  MUX2X1 U2058 ( .B(n1844), .A(n1841), .S(n14), .Y(n1855) );
  MUX2X1 U2059 ( .B(mem[356]), .A(mem[372]), .S(n2222), .Y(n1849) );
  MUX2X1 U2060 ( .B(mem[324]), .A(mem[340]), .S(n2222), .Y(n1848) );
  MUX2X1 U2061 ( .B(mem[292]), .A(mem[308]), .S(n2222), .Y(n1852) );
  MUX2X1 U2062 ( .B(mem[260]), .A(mem[276]), .S(n2222), .Y(n1851) );
  MUX2X1 U2063 ( .B(n1850), .A(n1847), .S(n14), .Y(n1854) );
  MUX2X1 U2064 ( .B(mem[228]), .A(mem[244]), .S(n2222), .Y(n1858) );
  MUX2X1 U2065 ( .B(mem[196]), .A(mem[212]), .S(n2222), .Y(n1857) );
  MUX2X1 U2066 ( .B(mem[164]), .A(mem[180]), .S(n2222), .Y(n1861) );
  MUX2X1 U2067 ( .B(mem[132]), .A(mem[148]), .S(n2222), .Y(n1860) );
  MUX2X1 U2068 ( .B(n1859), .A(n1856), .S(n14), .Y(n1870) );
  MUX2X1 U2069 ( .B(mem[100]), .A(mem[116]), .S(n2223), .Y(n1864) );
  MUX2X1 U2070 ( .B(mem[68]), .A(mem[84]), .S(n2223), .Y(n1863) );
  MUX2X1 U2071 ( .B(mem[36]), .A(mem[52]), .S(n2223), .Y(n1867) );
  MUX2X1 U2072 ( .B(mem[4]), .A(mem[20]), .S(n2223), .Y(n1866) );
  MUX2X1 U2073 ( .B(n1865), .A(n1862), .S(n14), .Y(n1869) );
  MUX2X1 U2074 ( .B(n1868), .A(n1853), .S(n16), .Y(n2205) );
  MUX2X1 U2075 ( .B(mem[485]), .A(mem[501]), .S(n2223), .Y(n1873) );
  MUX2X1 U2076 ( .B(mem[453]), .A(mem[469]), .S(n2223), .Y(n1872) );
  MUX2X1 U2077 ( .B(mem[421]), .A(mem[437]), .S(n2223), .Y(n1876) );
  MUX2X1 U2078 ( .B(mem[389]), .A(mem[405]), .S(n2223), .Y(n1875) );
  MUX2X1 U2079 ( .B(n1874), .A(n1871), .S(n14), .Y(n1885) );
  MUX2X1 U2080 ( .B(mem[357]), .A(mem[373]), .S(n2223), .Y(n1879) );
  MUX2X1 U2081 ( .B(mem[325]), .A(mem[341]), .S(n2223), .Y(n1878) );
  MUX2X1 U2082 ( .B(mem[293]), .A(mem[309]), .S(n2223), .Y(n1882) );
  MUX2X1 U2083 ( .B(mem[261]), .A(mem[277]), .S(n2223), .Y(n1881) );
  MUX2X1 U2084 ( .B(n1880), .A(n1877), .S(n14), .Y(n1884) );
  MUX2X1 U2085 ( .B(mem[229]), .A(mem[245]), .S(n2224), .Y(n1888) );
  MUX2X1 U2086 ( .B(mem[197]), .A(mem[213]), .S(n2224), .Y(n1887) );
  MUX2X1 U2087 ( .B(mem[165]), .A(mem[181]), .S(n2224), .Y(n1891) );
  MUX2X1 U2088 ( .B(mem[133]), .A(mem[149]), .S(n2224), .Y(n1890) );
  MUX2X1 U2089 ( .B(n1889), .A(n1886), .S(n14), .Y(n1900) );
  MUX2X1 U2090 ( .B(mem[101]), .A(mem[117]), .S(n2224), .Y(n1894) );
  MUX2X1 U2091 ( .B(mem[69]), .A(mem[85]), .S(n2224), .Y(n1893) );
  MUX2X1 U2092 ( .B(mem[37]), .A(mem[53]), .S(n2224), .Y(n1897) );
  MUX2X1 U2093 ( .B(mem[5]), .A(mem[21]), .S(n2224), .Y(n1896) );
  MUX2X1 U2094 ( .B(n1895), .A(n1892), .S(n14), .Y(n1899) );
  MUX2X1 U2095 ( .B(n1898), .A(n1883), .S(n16), .Y(n2206) );
  MUX2X1 U2096 ( .B(mem[486]), .A(mem[502]), .S(n2224), .Y(n1903) );
  MUX2X1 U2097 ( .B(mem[454]), .A(mem[470]), .S(n2224), .Y(n1902) );
  MUX2X1 U2098 ( .B(mem[422]), .A(mem[438]), .S(n2224), .Y(n1906) );
  MUX2X1 U2099 ( .B(mem[390]), .A(mem[406]), .S(n2224), .Y(n1905) );
  MUX2X1 U2100 ( .B(n1904), .A(n1901), .S(n14), .Y(n1915) );
  MUX2X1 U2101 ( .B(mem[358]), .A(mem[374]), .S(n2225), .Y(n1909) );
  MUX2X1 U2102 ( .B(mem[326]), .A(mem[342]), .S(n2225), .Y(n1908) );
  MUX2X1 U2103 ( .B(mem[294]), .A(mem[310]), .S(n2225), .Y(n1912) );
  MUX2X1 U2104 ( .B(mem[262]), .A(mem[278]), .S(n2225), .Y(n1911) );
  MUX2X1 U2105 ( .B(n1910), .A(n1907), .S(n14), .Y(n1914) );
  MUX2X1 U2106 ( .B(mem[230]), .A(mem[246]), .S(n2225), .Y(n1918) );
  MUX2X1 U2107 ( .B(mem[198]), .A(mem[214]), .S(n2225), .Y(n1917) );
  MUX2X1 U2108 ( .B(mem[166]), .A(mem[182]), .S(n2225), .Y(n1921) );
  MUX2X1 U2109 ( .B(mem[134]), .A(mem[150]), .S(n2225), .Y(n1920) );
  MUX2X1 U2110 ( .B(n1919), .A(n1916), .S(n14), .Y(n1930) );
  MUX2X1 U2111 ( .B(mem[102]), .A(mem[118]), .S(n2225), .Y(n1924) );
  MUX2X1 U2112 ( .B(mem[70]), .A(mem[86]), .S(n2225), .Y(n1923) );
  MUX2X1 U2113 ( .B(mem[38]), .A(mem[54]), .S(n2225), .Y(n1927) );
  MUX2X1 U2114 ( .B(mem[6]), .A(mem[22]), .S(n2225), .Y(n1926) );
  MUX2X1 U2115 ( .B(n1925), .A(n1922), .S(n14), .Y(n1929) );
  MUX2X1 U2116 ( .B(n1928), .A(n1913), .S(n16), .Y(n2207) );
  MUX2X1 U2117 ( .B(mem[487]), .A(mem[503]), .S(n2226), .Y(n1933) );
  MUX2X1 U2118 ( .B(mem[455]), .A(mem[471]), .S(n2226), .Y(n1932) );
  MUX2X1 U2119 ( .B(mem[423]), .A(mem[439]), .S(n2226), .Y(n1936) );
  MUX2X1 U2120 ( .B(mem[391]), .A(mem[407]), .S(n2226), .Y(n1935) );
  MUX2X1 U2121 ( .B(n1934), .A(n1931), .S(n14), .Y(n1945) );
  MUX2X1 U2122 ( .B(mem[359]), .A(mem[375]), .S(n2226), .Y(n1939) );
  MUX2X1 U2123 ( .B(mem[327]), .A(mem[343]), .S(n2226), .Y(n1938) );
  MUX2X1 U2124 ( .B(mem[295]), .A(mem[311]), .S(n2226), .Y(n1942) );
  MUX2X1 U2125 ( .B(mem[263]), .A(mem[279]), .S(n2226), .Y(n1941) );
  MUX2X1 U2126 ( .B(n1940), .A(n1937), .S(n14), .Y(n1944) );
  MUX2X1 U2127 ( .B(mem[231]), .A(mem[247]), .S(n2226), .Y(n1948) );
  MUX2X1 U2128 ( .B(mem[199]), .A(mem[215]), .S(n2226), .Y(n1947) );
  MUX2X1 U2129 ( .B(mem[167]), .A(mem[183]), .S(n2226), .Y(n1951) );
  MUX2X1 U2130 ( .B(mem[135]), .A(mem[151]), .S(n2226), .Y(n1950) );
  MUX2X1 U2131 ( .B(n1949), .A(n1946), .S(n14), .Y(n1960) );
  MUX2X1 U2132 ( .B(mem[103]), .A(mem[119]), .S(n2227), .Y(n1954) );
  MUX2X1 U2133 ( .B(mem[71]), .A(mem[87]), .S(n2227), .Y(n1953) );
  MUX2X1 U2134 ( .B(mem[39]), .A(mem[55]), .S(n2227), .Y(n1957) );
  MUX2X1 U2135 ( .B(mem[7]), .A(mem[23]), .S(n2227), .Y(n1956) );
  MUX2X1 U2136 ( .B(n1955), .A(n1952), .S(n14), .Y(n1959) );
  MUX2X1 U2137 ( .B(n1958), .A(n1943), .S(n16), .Y(n2208) );
  MUX2X1 U2138 ( .B(mem[488]), .A(mem[504]), .S(n2227), .Y(n1963) );
  MUX2X1 U2139 ( .B(mem[456]), .A(mem[472]), .S(n2227), .Y(n1962) );
  MUX2X1 U2140 ( .B(mem[424]), .A(mem[440]), .S(n2227), .Y(n1966) );
  MUX2X1 U2141 ( .B(mem[392]), .A(mem[408]), .S(n2227), .Y(n1965) );
  MUX2X1 U2142 ( .B(n1964), .A(n1961), .S(n14), .Y(n1975) );
  MUX2X1 U2143 ( .B(mem[360]), .A(mem[376]), .S(n2227), .Y(n1969) );
  MUX2X1 U2144 ( .B(mem[328]), .A(mem[344]), .S(n2227), .Y(n1968) );
  MUX2X1 U2145 ( .B(mem[296]), .A(mem[312]), .S(n2227), .Y(n1972) );
  MUX2X1 U2146 ( .B(mem[264]), .A(mem[280]), .S(n2227), .Y(n1971) );
  MUX2X1 U2147 ( .B(n1970), .A(n1967), .S(n14), .Y(n1974) );
  MUX2X1 U2148 ( .B(mem[232]), .A(mem[248]), .S(n2228), .Y(n1978) );
  MUX2X1 U2149 ( .B(mem[200]), .A(mem[216]), .S(n2228), .Y(n1977) );
  MUX2X1 U2150 ( .B(mem[168]), .A(mem[184]), .S(n2228), .Y(n1981) );
  MUX2X1 U2151 ( .B(mem[136]), .A(mem[152]), .S(n2228), .Y(n1980) );
  MUX2X1 U2152 ( .B(n1979), .A(n1976), .S(n14), .Y(n1990) );
  MUX2X1 U2153 ( .B(mem[104]), .A(mem[120]), .S(n2228), .Y(n1984) );
  MUX2X1 U2154 ( .B(mem[72]), .A(mem[88]), .S(n2228), .Y(n1983) );
  MUX2X1 U2155 ( .B(mem[40]), .A(mem[56]), .S(n2228), .Y(n1987) );
  MUX2X1 U2156 ( .B(mem[8]), .A(mem[24]), .S(n2228), .Y(n1986) );
  MUX2X1 U2157 ( .B(n1985), .A(n1982), .S(n14), .Y(n1989) );
  MUX2X1 U2158 ( .B(n1988), .A(n1973), .S(n16), .Y(n2209) );
  MUX2X1 U2159 ( .B(mem[489]), .A(mem[505]), .S(n2228), .Y(n1993) );
  MUX2X1 U2160 ( .B(mem[457]), .A(mem[473]), .S(n2228), .Y(n1992) );
  MUX2X1 U2161 ( .B(mem[425]), .A(mem[441]), .S(n2228), .Y(n1996) );
  MUX2X1 U2162 ( .B(mem[393]), .A(mem[409]), .S(n2228), .Y(n1995) );
  MUX2X1 U2163 ( .B(n1994), .A(n1991), .S(n14), .Y(n2005) );
  MUX2X1 U2164 ( .B(mem[361]), .A(mem[377]), .S(n2229), .Y(n1999) );
  MUX2X1 U2165 ( .B(mem[329]), .A(mem[345]), .S(n2229), .Y(n1998) );
  MUX2X1 U2166 ( .B(mem[297]), .A(mem[313]), .S(n2229), .Y(n2002) );
  MUX2X1 U2167 ( .B(mem[265]), .A(mem[281]), .S(n2229), .Y(n2001) );
  MUX2X1 U2168 ( .B(n2000), .A(n1997), .S(n14), .Y(n2004) );
  MUX2X1 U2169 ( .B(mem[233]), .A(mem[249]), .S(n2229), .Y(n2008) );
  MUX2X1 U2170 ( .B(mem[201]), .A(mem[217]), .S(n2229), .Y(n2007) );
  MUX2X1 U2171 ( .B(mem[169]), .A(mem[185]), .S(n2229), .Y(n2011) );
  MUX2X1 U2172 ( .B(mem[137]), .A(mem[153]), .S(n2229), .Y(n2010) );
  MUX2X1 U2173 ( .B(n2009), .A(n2006), .S(n14), .Y(n2020) );
  MUX2X1 U2174 ( .B(mem[105]), .A(mem[121]), .S(n2229), .Y(n2014) );
  MUX2X1 U2175 ( .B(mem[73]), .A(mem[89]), .S(n2229), .Y(n2013) );
  MUX2X1 U2176 ( .B(mem[41]), .A(mem[57]), .S(n2229), .Y(n2017) );
  MUX2X1 U2177 ( .B(mem[9]), .A(mem[25]), .S(n2229), .Y(n2016) );
  MUX2X1 U2178 ( .B(n2015), .A(n2012), .S(n14), .Y(n2019) );
  MUX2X1 U2179 ( .B(n2018), .A(n2003), .S(n16), .Y(n2210) );
  MUX2X1 U2180 ( .B(mem[490]), .A(mem[506]), .S(n2230), .Y(n2023) );
  MUX2X1 U2181 ( .B(mem[458]), .A(mem[474]), .S(n2223), .Y(n2022) );
  MUX2X1 U2182 ( .B(mem[426]), .A(mem[442]), .S(n2227), .Y(n2026) );
  MUX2X1 U2183 ( .B(mem[394]), .A(mem[410]), .S(n2219), .Y(n2025) );
  MUX2X1 U2184 ( .B(n2024), .A(n2021), .S(n14), .Y(n2035) );
  MUX2X1 U2185 ( .B(mem[362]), .A(mem[378]), .S(n2224), .Y(n2029) );
  MUX2X1 U2186 ( .B(mem[330]), .A(mem[346]), .S(n2231), .Y(n2028) );
  MUX2X1 U2187 ( .B(mem[298]), .A(mem[314]), .S(n2228), .Y(n2032) );
  MUX2X1 U2188 ( .B(mem[266]), .A(mem[282]), .S(n2222), .Y(n2031) );
  MUX2X1 U2189 ( .B(n2030), .A(n2027), .S(n14), .Y(n2034) );
  MUX2X1 U2190 ( .B(mem[234]), .A(mem[250]), .S(n2224), .Y(n2038) );
  MUX2X1 U2191 ( .B(mem[202]), .A(mem[218]), .S(n2234), .Y(n2037) );
  MUX2X1 U2192 ( .B(mem[170]), .A(mem[186]), .S(n2228), .Y(n2041) );
  MUX2X1 U2193 ( .B(mem[138]), .A(mem[154]), .S(n2222), .Y(n2040) );
  MUX2X1 U2194 ( .B(n2039), .A(n2036), .S(n14), .Y(n2050) );
  MUX2X1 U2195 ( .B(mem[106]), .A(mem[122]), .S(n2230), .Y(n2044) );
  MUX2X1 U2196 ( .B(mem[74]), .A(mem[90]), .S(n2230), .Y(n2043) );
  MUX2X1 U2197 ( .B(mem[42]), .A(mem[58]), .S(n2230), .Y(n2047) );
  MUX2X1 U2198 ( .B(mem[10]), .A(mem[26]), .S(n2230), .Y(n2046) );
  MUX2X1 U2199 ( .B(n2045), .A(n2042), .S(n14), .Y(n2049) );
  MUX2X1 U2200 ( .B(n2048), .A(n2033), .S(n16), .Y(n2211) );
  MUX2X1 U2201 ( .B(mem[491]), .A(mem[507]), .S(n2230), .Y(n2053) );
  MUX2X1 U2202 ( .B(mem[459]), .A(mem[475]), .S(n2230), .Y(n2052) );
  MUX2X1 U2203 ( .B(mem[427]), .A(mem[443]), .S(n2230), .Y(n2056) );
  MUX2X1 U2204 ( .B(mem[395]), .A(mem[411]), .S(n2230), .Y(n2055) );
  MUX2X1 U2205 ( .B(n2054), .A(n2051), .S(n14), .Y(n2065) );
  MUX2X1 U2206 ( .B(mem[363]), .A(mem[379]), .S(n2230), .Y(n2059) );
  MUX2X1 U2207 ( .B(mem[331]), .A(mem[347]), .S(n2230), .Y(n2058) );
  MUX2X1 U2208 ( .B(mem[299]), .A(mem[315]), .S(n2230), .Y(n2062) );
  MUX2X1 U2209 ( .B(mem[267]), .A(mem[283]), .S(n2230), .Y(n2061) );
  MUX2X1 U2210 ( .B(n2060), .A(n2057), .S(n14), .Y(n2064) );
  MUX2X1 U2211 ( .B(mem[235]), .A(mem[251]), .S(n2231), .Y(n2068) );
  MUX2X1 U2212 ( .B(mem[203]), .A(mem[219]), .S(n2231), .Y(n2067) );
  MUX2X1 U2213 ( .B(mem[171]), .A(mem[187]), .S(n2231), .Y(n2071) );
  MUX2X1 U2214 ( .B(mem[139]), .A(mem[155]), .S(n2231), .Y(n2070) );
  MUX2X1 U2215 ( .B(n2069), .A(n2066), .S(n14), .Y(n2080) );
  MUX2X1 U2216 ( .B(mem[107]), .A(mem[123]), .S(n2231), .Y(n2074) );
  MUX2X1 U2217 ( .B(mem[75]), .A(mem[91]), .S(n2231), .Y(n2073) );
  MUX2X1 U2218 ( .B(mem[43]), .A(mem[59]), .S(n2231), .Y(n2077) );
  MUX2X1 U2219 ( .B(mem[11]), .A(mem[27]), .S(n2231), .Y(n2076) );
  MUX2X1 U2220 ( .B(n2075), .A(n2072), .S(n14), .Y(n2079) );
  MUX2X1 U2221 ( .B(n2078), .A(n2063), .S(n16), .Y(n2212) );
  MUX2X1 U2222 ( .B(mem[492]), .A(mem[508]), .S(n2231), .Y(n2083) );
  MUX2X1 U2223 ( .B(mem[460]), .A(mem[476]), .S(n2231), .Y(n2082) );
  MUX2X1 U2224 ( .B(mem[428]), .A(mem[444]), .S(n2231), .Y(n2086) );
  MUX2X1 U2225 ( .B(mem[396]), .A(mem[412]), .S(n2231), .Y(n2085) );
  MUX2X1 U2226 ( .B(n2084), .A(n2081), .S(n14), .Y(n2095) );
  MUX2X1 U2227 ( .B(mem[364]), .A(mem[380]), .S(n2232), .Y(n2089) );
  MUX2X1 U2228 ( .B(mem[332]), .A(mem[348]), .S(n2232), .Y(n2088) );
  MUX2X1 U2229 ( .B(mem[300]), .A(mem[316]), .S(n2232), .Y(n2092) );
  MUX2X1 U2230 ( .B(mem[268]), .A(mem[284]), .S(n2232), .Y(n2091) );
  MUX2X1 U2231 ( .B(n2090), .A(n2087), .S(n14), .Y(n2094) );
  MUX2X1 U2232 ( .B(mem[236]), .A(mem[252]), .S(n2232), .Y(n2098) );
  MUX2X1 U2233 ( .B(mem[204]), .A(mem[220]), .S(n2232), .Y(n2097) );
  MUX2X1 U2234 ( .B(mem[172]), .A(mem[188]), .S(n2232), .Y(n2101) );
  MUX2X1 U2235 ( .B(mem[140]), .A(mem[156]), .S(n2232), .Y(n2100) );
  MUX2X1 U2236 ( .B(n2099), .A(n2096), .S(n14), .Y(n2110) );
  MUX2X1 U2237 ( .B(mem[108]), .A(mem[124]), .S(n2232), .Y(n2104) );
  MUX2X1 U2238 ( .B(mem[76]), .A(mem[92]), .S(n2232), .Y(n2103) );
  MUX2X1 U2239 ( .B(mem[44]), .A(mem[60]), .S(n2232), .Y(n2107) );
  MUX2X1 U2240 ( .B(mem[12]), .A(mem[28]), .S(n2232), .Y(n2106) );
  MUX2X1 U2241 ( .B(n2105), .A(n2102), .S(n14), .Y(n2109) );
  MUX2X1 U2242 ( .B(n2108), .A(n2093), .S(n16), .Y(n2213) );
  MUX2X1 U2243 ( .B(mem[493]), .A(mem[509]), .S(n2233), .Y(n2113) );
  MUX2X1 U2244 ( .B(mem[461]), .A(mem[477]), .S(n2233), .Y(n2112) );
  MUX2X1 U2245 ( .B(mem[429]), .A(mem[445]), .S(n2233), .Y(n2116) );
  MUX2X1 U2246 ( .B(mem[397]), .A(mem[413]), .S(n2233), .Y(n2115) );
  MUX2X1 U2247 ( .B(n2114), .A(n2111), .S(n14), .Y(n2125) );
  MUX2X1 U2248 ( .B(mem[365]), .A(mem[381]), .S(n2233), .Y(n2119) );
  MUX2X1 U2249 ( .B(mem[333]), .A(mem[349]), .S(n2233), .Y(n2118) );
  MUX2X1 U2250 ( .B(mem[301]), .A(mem[317]), .S(n2233), .Y(n2122) );
  MUX2X1 U2251 ( .B(mem[269]), .A(mem[285]), .S(n2233), .Y(n2121) );
  MUX2X1 U2252 ( .B(n2120), .A(n2117), .S(n14), .Y(n2124) );
  MUX2X1 U2253 ( .B(mem[237]), .A(mem[253]), .S(n2233), .Y(n2128) );
  MUX2X1 U2254 ( .B(mem[205]), .A(mem[221]), .S(n2233), .Y(n2127) );
  MUX2X1 U2255 ( .B(mem[173]), .A(mem[189]), .S(n2233), .Y(n2131) );
  MUX2X1 U2256 ( .B(mem[141]), .A(mem[157]), .S(n2233), .Y(n2130) );
  MUX2X1 U2257 ( .B(n2129), .A(n2126), .S(n14), .Y(n2140) );
  MUX2X1 U2258 ( .B(mem[109]), .A(mem[125]), .S(n2234), .Y(n2134) );
  MUX2X1 U2259 ( .B(mem[77]), .A(mem[93]), .S(n2234), .Y(n2133) );
  MUX2X1 U2260 ( .B(mem[45]), .A(mem[61]), .S(n2234), .Y(n2137) );
  MUX2X1 U2261 ( .B(mem[13]), .A(mem[29]), .S(n2234), .Y(n2136) );
  MUX2X1 U2262 ( .B(n2135), .A(n2132), .S(n14), .Y(n2139) );
  MUX2X1 U2263 ( .B(n2138), .A(n2123), .S(n16), .Y(n2214) );
  MUX2X1 U2264 ( .B(mem[494]), .A(mem[510]), .S(n2234), .Y(n2143) );
  MUX2X1 U2265 ( .B(mem[462]), .A(mem[478]), .S(n2234), .Y(n2142) );
  MUX2X1 U2266 ( .B(mem[430]), .A(mem[446]), .S(n2234), .Y(n2146) );
  MUX2X1 U2267 ( .B(mem[398]), .A(mem[414]), .S(n2234), .Y(n2145) );
  MUX2X1 U2268 ( .B(n2144), .A(n2141), .S(n14), .Y(n2155) );
  MUX2X1 U2269 ( .B(mem[366]), .A(mem[382]), .S(n2234), .Y(n2149) );
  MUX2X1 U2270 ( .B(mem[334]), .A(mem[350]), .S(n2234), .Y(n2148) );
  MUX2X1 U2271 ( .B(mem[302]), .A(mem[318]), .S(n2234), .Y(n2152) );
  MUX2X1 U2272 ( .B(mem[270]), .A(mem[286]), .S(n2234), .Y(n2151) );
  MUX2X1 U2273 ( .B(n2150), .A(n2147), .S(n14), .Y(n2154) );
  MUX2X1 U2274 ( .B(mem[238]), .A(mem[254]), .S(n2235), .Y(n2158) );
  MUX2X1 U2275 ( .B(mem[206]), .A(mem[222]), .S(n2235), .Y(n2157) );
  MUX2X1 U2276 ( .B(mem[174]), .A(mem[190]), .S(n2235), .Y(n2161) );
  MUX2X1 U2277 ( .B(mem[142]), .A(mem[158]), .S(n2235), .Y(n2160) );
  MUX2X1 U2278 ( .B(n2159), .A(n2156), .S(n14), .Y(n2170) );
  MUX2X1 U2279 ( .B(mem[110]), .A(mem[126]), .S(n2235), .Y(n2164) );
  MUX2X1 U2280 ( .B(mem[78]), .A(mem[94]), .S(n2235), .Y(n2163) );
  MUX2X1 U2281 ( .B(mem[46]), .A(mem[62]), .S(n2235), .Y(n2167) );
  MUX2X1 U2282 ( .B(mem[14]), .A(mem[30]), .S(n2235), .Y(n2166) );
  MUX2X1 U2283 ( .B(n2165), .A(n2162), .S(n14), .Y(n2169) );
  MUX2X1 U2284 ( .B(n2168), .A(n2153), .S(n16), .Y(n2215) );
  MUX2X1 U2285 ( .B(mem[495]), .A(mem[511]), .S(n2235), .Y(n2173) );
  MUX2X1 U2286 ( .B(mem[463]), .A(mem[479]), .S(n2235), .Y(n2172) );
  MUX2X1 U2287 ( .B(mem[431]), .A(mem[447]), .S(n2235), .Y(n2176) );
  MUX2X1 U2288 ( .B(mem[399]), .A(mem[415]), .S(n2235), .Y(n2175) );
  MUX2X1 U2289 ( .B(n2174), .A(n2171), .S(n14), .Y(n2185) );
  MUX2X1 U2290 ( .B(mem[367]), .A(mem[383]), .S(n2233), .Y(n2179) );
  MUX2X1 U2291 ( .B(mem[335]), .A(mem[351]), .S(n2232), .Y(n2178) );
  MUX2X1 U2292 ( .B(mem[303]), .A(mem[319]), .S(n2235), .Y(n2182) );
  MUX2X1 U2293 ( .B(mem[271]), .A(mem[287]), .S(n2218), .Y(n2181) );
  MUX2X1 U2294 ( .B(n2180), .A(n2177), .S(n14), .Y(n2184) );
  MUX2X1 U2295 ( .B(mem[239]), .A(mem[255]), .S(n2223), .Y(n2188) );
  MUX2X1 U2296 ( .B(mem[207]), .A(mem[223]), .S(n2226), .Y(n2187) );
  MUX2X1 U2297 ( .B(mem[175]), .A(mem[191]), .S(n2221), .Y(n2191) );
  MUX2X1 U2298 ( .B(mem[143]), .A(mem[159]), .S(n2219), .Y(n2190) );
  MUX2X1 U2299 ( .B(n2189), .A(n2186), .S(n14), .Y(n2200) );
  MUX2X1 U2300 ( .B(mem[111]), .A(mem[127]), .S(n2225), .Y(n2194) );
  MUX2X1 U2301 ( .B(mem[79]), .A(mem[95]), .S(n2217), .Y(n2193) );
  MUX2X1 U2302 ( .B(mem[47]), .A(mem[63]), .S(n2234), .Y(n2197) );
  MUX2X1 U2303 ( .B(mem[15]), .A(mem[31]), .S(n2230), .Y(n2196) );
  MUX2X1 U2304 ( .B(n2195), .A(n2192), .S(n14), .Y(n2199) );
  MUX2X1 U2305 ( .B(n2198), .A(n2183), .S(n16), .Y(n2216) );
  OR2X1 U2306 ( .A(n2291), .B(wr_ptr[0]), .Y(sub_93_carry[1]) );
  XNOR2X1 U2307 ( .A(wr_ptr[0]), .B(n2291), .Y(fillcount[0]) );
  XOR2X1 U2308 ( .A(add_51_carry[4]), .B(wr_ptr[4]), .Y(n23) );
  XOR2X1 U2309 ( .A(add_57_carry[4]), .B(n16), .Y(n76) );
endmodule


module FIFO_DEPTH_P25_WIDTH33 ( clk, reset, data_in, put, get, data_out, 
        empty_bar, full_bar, fillcount );
  input [32:0] data_in;
  output [32:0] data_out;
  output [5:0] fillcount;
  input clk, reset, put, get;
  output empty_bar, full_bar;
  wire   n12, n13, n14, n15, n16, n4624, n4625, n20, n21, n22, n23, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n90, n91, n92, n93, n349, n351, n353, n355, n357, n359,
         n361, n363, n365, n367, n369, n371, n373, n375, n377, n379, n381,
         n383, n385, n387, n389, n391, n393, n395, n397, n399, n401, n403,
         n405, n407, n409, n411, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n17, n18, n19,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n89, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n350, n352, n354, n356, n358, n360,
         n362, n364, n366, n368, n370, n372, n374, n376, n378, n380, n382,
         n384, n386, n388, n390, n392, n394, n396, n398, n400, n402, n404,
         n406, n408, n410, n412, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
         n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623;
  wire   [4:0] wr_ptr;
  wire   [1055:0] mem;
  wire   [4:2] add_57_carry;
  wire   [4:2] add_51_carry;
  wire   [5:1] sub_93_carry;

  DFFPOSX1 wr_ptr_reg_0_ ( .D(n2603), .CLK(clk), .Q(wr_ptr[0]) );
  DFFPOSX1 rd_ptr_reg_4_ ( .D(n2602), .CLK(clk), .Q(n16) );
  DFFPOSX1 rd_ptr_reg_0_ ( .D(n2601), .CLK(clk), .Q(n12) );
  DFFPOSX1 rd_ptr_reg_1_ ( .D(n2600), .CLK(clk), .Q(n13) );
  DFFPOSX1 rd_ptr_reg_2_ ( .D(n2599), .CLK(clk), .Q(n14) );
  DFFPOSX1 rd_ptr_reg_3_ ( .D(n2598), .CLK(clk), .Q(n15) );
  DFFPOSX1 wr_ptr_reg_4_ ( .D(n2597), .CLK(clk), .Q(wr_ptr[4]) );
  DFFPOSX1 wr_ptr_reg_1_ ( .D(n2596), .CLK(clk), .Q(wr_ptr[1]) );
  DFFPOSX1 wr_ptr_reg_2_ ( .D(n2595), .CLK(clk), .Q(wr_ptr[2]) );
  DFFPOSX1 wr_ptr_reg_3_ ( .D(n2594), .CLK(clk), .Q(wr_ptr[3]) );
  DFFPOSX1 data_out_reg_32_ ( .D(n4618), .CLK(clk), .Q(data_out[32]) );
  DFFPOSX1 data_out_reg_31_ ( .D(n4617), .CLK(clk), .Q(data_out[31]) );
  DFFPOSX1 data_out_reg_30_ ( .D(n4616), .CLK(clk), .Q(data_out[30]) );
  DFFPOSX1 data_out_reg_29_ ( .D(n4615), .CLK(clk), .Q(data_out[29]) );
  DFFPOSX1 data_out_reg_28_ ( .D(n4614), .CLK(clk), .Q(data_out[28]) );
  DFFPOSX1 data_out_reg_27_ ( .D(n4613), .CLK(clk), .Q(data_out[27]) );
  DFFPOSX1 data_out_reg_26_ ( .D(n4612), .CLK(clk), .Q(data_out[26]) );
  DFFPOSX1 data_out_reg_25_ ( .D(n4611), .CLK(clk), .Q(data_out[25]) );
  DFFPOSX1 data_out_reg_24_ ( .D(n4610), .CLK(clk), .Q(data_out[24]) );
  DFFPOSX1 data_out_reg_23_ ( .D(n4609), .CLK(clk), .Q(data_out[23]) );
  DFFPOSX1 data_out_reg_22_ ( .D(n4608), .CLK(clk), .Q(data_out[22]) );
  DFFPOSX1 data_out_reg_21_ ( .D(n4607), .CLK(clk), .Q(data_out[21]) );
  DFFPOSX1 data_out_reg_20_ ( .D(n4606), .CLK(clk), .Q(data_out[20]) );
  DFFPOSX1 data_out_reg_19_ ( .D(n4605), .CLK(clk), .Q(data_out[19]) );
  DFFPOSX1 data_out_reg_18_ ( .D(n4604), .CLK(clk), .Q(data_out[18]) );
  DFFPOSX1 data_out_reg_17_ ( .D(n4603), .CLK(clk), .Q(data_out[17]) );
  DFFPOSX1 data_out_reg_16_ ( .D(n4602), .CLK(clk), .Q(data_out[16]) );
  DFFPOSX1 data_out_reg_15_ ( .D(n4601), .CLK(clk), .Q(data_out[15]) );
  DFFPOSX1 data_out_reg_14_ ( .D(n4600), .CLK(clk), .Q(data_out[14]) );
  DFFPOSX1 data_out_reg_13_ ( .D(n4599), .CLK(clk), .Q(data_out[13]) );
  DFFPOSX1 data_out_reg_12_ ( .D(n4598), .CLK(clk), .Q(data_out[12]) );
  DFFPOSX1 data_out_reg_11_ ( .D(n4597), .CLK(clk), .Q(data_out[11]) );
  DFFPOSX1 data_out_reg_10_ ( .D(n4596), .CLK(clk), .Q(data_out[10]) );
  DFFPOSX1 data_out_reg_9_ ( .D(n4595), .CLK(clk), .Q(data_out[9]) );
  DFFPOSX1 data_out_reg_8_ ( .D(n4594), .CLK(clk), .Q(data_out[8]) );
  DFFPOSX1 data_out_reg_7_ ( .D(n4593), .CLK(clk), .Q(data_out[7]) );
  DFFPOSX1 data_out_reg_6_ ( .D(n4592), .CLK(clk), .Q(data_out[6]) );
  DFFPOSX1 data_out_reg_5_ ( .D(n4591), .CLK(clk), .Q(data_out[5]) );
  DFFPOSX1 data_out_reg_4_ ( .D(n4590), .CLK(clk), .Q(data_out[4]) );
  DFFPOSX1 data_out_reg_3_ ( .D(n4589), .CLK(clk), .Q(data_out[3]) );
  DFFPOSX1 data_out_reg_2_ ( .D(n4588), .CLK(clk), .Q(data_out[2]) );
  DFFPOSX1 data_out_reg_1_ ( .D(n4587), .CLK(clk), .Q(data_out[1]) );
  DFFPOSX1 data_out_reg_0_ ( .D(n4586), .CLK(clk), .Q(data_out[0]) );
  DFFPOSX1 mem_reg_31__32_ ( .D(n2593), .CLK(clk), .Q(mem[1055]) );
  DFFPOSX1 mem_reg_31__31_ ( .D(n2592), .CLK(clk), .Q(mem[1054]) );
  DFFPOSX1 mem_reg_31__30_ ( .D(n2591), .CLK(clk), .Q(mem[1053]) );
  DFFPOSX1 mem_reg_31__29_ ( .D(n2590), .CLK(clk), .Q(mem[1052]) );
  DFFPOSX1 mem_reg_31__28_ ( .D(n2589), .CLK(clk), .Q(mem[1051]) );
  DFFPOSX1 mem_reg_31__27_ ( .D(n2588), .CLK(clk), .Q(mem[1050]) );
  DFFPOSX1 mem_reg_31__26_ ( .D(n2587), .CLK(clk), .Q(mem[1049]) );
  DFFPOSX1 mem_reg_31__25_ ( .D(n2586), .CLK(clk), .Q(mem[1048]) );
  DFFPOSX1 mem_reg_31__24_ ( .D(n2585), .CLK(clk), .Q(mem[1047]) );
  DFFPOSX1 mem_reg_31__23_ ( .D(n2584), .CLK(clk), .Q(mem[1046]) );
  DFFPOSX1 mem_reg_31__22_ ( .D(n2583), .CLK(clk), .Q(mem[1045]) );
  DFFPOSX1 mem_reg_31__21_ ( .D(n2582), .CLK(clk), .Q(mem[1044]) );
  DFFPOSX1 mem_reg_31__20_ ( .D(n2581), .CLK(clk), .Q(mem[1043]) );
  DFFPOSX1 mem_reg_31__19_ ( .D(n2580), .CLK(clk), .Q(mem[1042]) );
  DFFPOSX1 mem_reg_31__18_ ( .D(n2579), .CLK(clk), .Q(mem[1041]) );
  DFFPOSX1 mem_reg_31__17_ ( .D(n2578), .CLK(clk), .Q(mem[1040]) );
  DFFPOSX1 mem_reg_31__16_ ( .D(n2577), .CLK(clk), .Q(mem[1039]) );
  DFFPOSX1 mem_reg_31__15_ ( .D(n2576), .CLK(clk), .Q(mem[1038]) );
  DFFPOSX1 mem_reg_31__14_ ( .D(n2575), .CLK(clk), .Q(mem[1037]) );
  DFFPOSX1 mem_reg_31__13_ ( .D(n2574), .CLK(clk), .Q(mem[1036]) );
  DFFPOSX1 mem_reg_31__12_ ( .D(n2573), .CLK(clk), .Q(mem[1035]) );
  DFFPOSX1 mem_reg_31__11_ ( .D(n2572), .CLK(clk), .Q(mem[1034]) );
  DFFPOSX1 mem_reg_31__10_ ( .D(n2571), .CLK(clk), .Q(mem[1033]) );
  DFFPOSX1 mem_reg_31__9_ ( .D(n2570), .CLK(clk), .Q(mem[1032]) );
  DFFPOSX1 mem_reg_31__8_ ( .D(n2569), .CLK(clk), .Q(mem[1031]) );
  DFFPOSX1 mem_reg_31__7_ ( .D(n2568), .CLK(clk), .Q(mem[1030]) );
  DFFPOSX1 mem_reg_31__6_ ( .D(n2567), .CLK(clk), .Q(mem[1029]) );
  DFFPOSX1 mem_reg_31__5_ ( .D(n2566), .CLK(clk), .Q(mem[1028]) );
  DFFPOSX1 mem_reg_31__4_ ( .D(n2565), .CLK(clk), .Q(mem[1027]) );
  DFFPOSX1 mem_reg_31__3_ ( .D(n2564), .CLK(clk), .Q(mem[1026]) );
  DFFPOSX1 mem_reg_31__2_ ( .D(n2563), .CLK(clk), .Q(mem[1025]) );
  DFFPOSX1 mem_reg_31__1_ ( .D(n2562), .CLK(clk), .Q(mem[1024]) );
  DFFPOSX1 mem_reg_31__0_ ( .D(n2561), .CLK(clk), .Q(mem[1023]) );
  DFFPOSX1 mem_reg_30__32_ ( .D(n2560), .CLK(clk), .Q(mem[1022]) );
  DFFPOSX1 mem_reg_30__31_ ( .D(n2559), .CLK(clk), .Q(mem[1021]) );
  DFFPOSX1 mem_reg_30__30_ ( .D(n2558), .CLK(clk), .Q(mem[1020]) );
  DFFPOSX1 mem_reg_30__29_ ( .D(n2557), .CLK(clk), .Q(mem[1019]) );
  DFFPOSX1 mem_reg_30__28_ ( .D(n2556), .CLK(clk), .Q(mem[1018]) );
  DFFPOSX1 mem_reg_30__27_ ( .D(n2555), .CLK(clk), .Q(mem[1017]) );
  DFFPOSX1 mem_reg_30__26_ ( .D(n2554), .CLK(clk), .Q(mem[1016]) );
  DFFPOSX1 mem_reg_30__25_ ( .D(n2553), .CLK(clk), .Q(mem[1015]) );
  DFFPOSX1 mem_reg_30__24_ ( .D(n2552), .CLK(clk), .Q(mem[1014]) );
  DFFPOSX1 mem_reg_30__23_ ( .D(n2551), .CLK(clk), .Q(mem[1013]) );
  DFFPOSX1 mem_reg_30__22_ ( .D(n2550), .CLK(clk), .Q(mem[1012]) );
  DFFPOSX1 mem_reg_30__21_ ( .D(n2549), .CLK(clk), .Q(mem[1011]) );
  DFFPOSX1 mem_reg_30__20_ ( .D(n2548), .CLK(clk), .Q(mem[1010]) );
  DFFPOSX1 mem_reg_30__19_ ( .D(n2547), .CLK(clk), .Q(mem[1009]) );
  DFFPOSX1 mem_reg_30__18_ ( .D(n2546), .CLK(clk), .Q(mem[1008]) );
  DFFPOSX1 mem_reg_30__17_ ( .D(n2545), .CLK(clk), .Q(mem[1007]) );
  DFFPOSX1 mem_reg_30__16_ ( .D(n2544), .CLK(clk), .Q(mem[1006]) );
  DFFPOSX1 mem_reg_30__15_ ( .D(n2543), .CLK(clk), .Q(mem[1005]) );
  DFFPOSX1 mem_reg_30__14_ ( .D(n2542), .CLK(clk), .Q(mem[1004]) );
  DFFPOSX1 mem_reg_30__13_ ( .D(n2541), .CLK(clk), .Q(mem[1003]) );
  DFFPOSX1 mem_reg_30__12_ ( .D(n2540), .CLK(clk), .Q(mem[1002]) );
  DFFPOSX1 mem_reg_30__11_ ( .D(n2539), .CLK(clk), .Q(mem[1001]) );
  DFFPOSX1 mem_reg_30__10_ ( .D(n2538), .CLK(clk), .Q(mem[1000]) );
  DFFPOSX1 mem_reg_30__9_ ( .D(n2537), .CLK(clk), .Q(mem[999]) );
  DFFPOSX1 mem_reg_30__8_ ( .D(n2536), .CLK(clk), .Q(mem[998]) );
  DFFPOSX1 mem_reg_30__7_ ( .D(n2535), .CLK(clk), .Q(mem[997]) );
  DFFPOSX1 mem_reg_30__6_ ( .D(n2534), .CLK(clk), .Q(mem[996]) );
  DFFPOSX1 mem_reg_30__5_ ( .D(n2533), .CLK(clk), .Q(mem[995]) );
  DFFPOSX1 mem_reg_30__4_ ( .D(n2532), .CLK(clk), .Q(mem[994]) );
  DFFPOSX1 mem_reg_30__3_ ( .D(n2531), .CLK(clk), .Q(mem[993]) );
  DFFPOSX1 mem_reg_30__2_ ( .D(n2530), .CLK(clk), .Q(mem[992]) );
  DFFPOSX1 mem_reg_30__1_ ( .D(n2529), .CLK(clk), .Q(mem[991]) );
  DFFPOSX1 mem_reg_30__0_ ( .D(n2528), .CLK(clk), .Q(mem[990]) );
  DFFPOSX1 mem_reg_29__32_ ( .D(n2527), .CLK(clk), .Q(mem[989]) );
  DFFPOSX1 mem_reg_29__31_ ( .D(n2526), .CLK(clk), .Q(mem[988]) );
  DFFPOSX1 mem_reg_29__30_ ( .D(n2525), .CLK(clk), .Q(mem[987]) );
  DFFPOSX1 mem_reg_29__29_ ( .D(n2524), .CLK(clk), .Q(mem[986]) );
  DFFPOSX1 mem_reg_29__28_ ( .D(n2523), .CLK(clk), .Q(mem[985]) );
  DFFPOSX1 mem_reg_29__27_ ( .D(n2522), .CLK(clk), .Q(mem[984]) );
  DFFPOSX1 mem_reg_29__26_ ( .D(n2521), .CLK(clk), .Q(mem[983]) );
  DFFPOSX1 mem_reg_29__25_ ( .D(n2520), .CLK(clk), .Q(mem[982]) );
  DFFPOSX1 mem_reg_29__24_ ( .D(n2519), .CLK(clk), .Q(mem[981]) );
  DFFPOSX1 mem_reg_29__23_ ( .D(n2518), .CLK(clk), .Q(mem[980]) );
  DFFPOSX1 mem_reg_29__22_ ( .D(n2517), .CLK(clk), .Q(mem[979]) );
  DFFPOSX1 mem_reg_29__21_ ( .D(n2516), .CLK(clk), .Q(mem[978]) );
  DFFPOSX1 mem_reg_29__20_ ( .D(n2515), .CLK(clk), .Q(mem[977]) );
  DFFPOSX1 mem_reg_29__19_ ( .D(n2514), .CLK(clk), .Q(mem[976]) );
  DFFPOSX1 mem_reg_29__18_ ( .D(n2513), .CLK(clk), .Q(mem[975]) );
  DFFPOSX1 mem_reg_29__17_ ( .D(n2512), .CLK(clk), .Q(mem[974]) );
  DFFPOSX1 mem_reg_29__16_ ( .D(n2511), .CLK(clk), .Q(mem[973]) );
  DFFPOSX1 mem_reg_29__15_ ( .D(n2510), .CLK(clk), .Q(mem[972]) );
  DFFPOSX1 mem_reg_29__14_ ( .D(n2509), .CLK(clk), .Q(mem[971]) );
  DFFPOSX1 mem_reg_29__13_ ( .D(n2508), .CLK(clk), .Q(mem[970]) );
  DFFPOSX1 mem_reg_29__12_ ( .D(n2507), .CLK(clk), .Q(mem[969]) );
  DFFPOSX1 mem_reg_29__11_ ( .D(n2506), .CLK(clk), .Q(mem[968]) );
  DFFPOSX1 mem_reg_29__10_ ( .D(n2505), .CLK(clk), .Q(mem[967]) );
  DFFPOSX1 mem_reg_29__9_ ( .D(n2504), .CLK(clk), .Q(mem[966]) );
  DFFPOSX1 mem_reg_29__8_ ( .D(n2503), .CLK(clk), .Q(mem[965]) );
  DFFPOSX1 mem_reg_29__7_ ( .D(n2502), .CLK(clk), .Q(mem[964]) );
  DFFPOSX1 mem_reg_29__6_ ( .D(n2501), .CLK(clk), .Q(mem[963]) );
  DFFPOSX1 mem_reg_29__5_ ( .D(n2500), .CLK(clk), .Q(mem[962]) );
  DFFPOSX1 mem_reg_29__4_ ( .D(n2499), .CLK(clk), .Q(mem[961]) );
  DFFPOSX1 mem_reg_29__3_ ( .D(n2498), .CLK(clk), .Q(mem[960]) );
  DFFPOSX1 mem_reg_29__2_ ( .D(n2497), .CLK(clk), .Q(mem[959]) );
  DFFPOSX1 mem_reg_29__1_ ( .D(n2496), .CLK(clk), .Q(mem[958]) );
  DFFPOSX1 mem_reg_29__0_ ( .D(n2495), .CLK(clk), .Q(mem[957]) );
  DFFPOSX1 mem_reg_28__32_ ( .D(n2494), .CLK(clk), .Q(mem[956]) );
  DFFPOSX1 mem_reg_28__31_ ( .D(n2493), .CLK(clk), .Q(mem[955]) );
  DFFPOSX1 mem_reg_28__30_ ( .D(n2492), .CLK(clk), .Q(mem[954]) );
  DFFPOSX1 mem_reg_28__29_ ( .D(n2491), .CLK(clk), .Q(mem[953]) );
  DFFPOSX1 mem_reg_28__28_ ( .D(n2490), .CLK(clk), .Q(mem[952]) );
  DFFPOSX1 mem_reg_28__27_ ( .D(n2489), .CLK(clk), .Q(mem[951]) );
  DFFPOSX1 mem_reg_28__26_ ( .D(n2488), .CLK(clk), .Q(mem[950]) );
  DFFPOSX1 mem_reg_28__25_ ( .D(n2487), .CLK(clk), .Q(mem[949]) );
  DFFPOSX1 mem_reg_28__24_ ( .D(n2486), .CLK(clk), .Q(mem[948]) );
  DFFPOSX1 mem_reg_28__23_ ( .D(n2485), .CLK(clk), .Q(mem[947]) );
  DFFPOSX1 mem_reg_28__22_ ( .D(n2484), .CLK(clk), .Q(mem[946]) );
  DFFPOSX1 mem_reg_28__21_ ( .D(n2483), .CLK(clk), .Q(mem[945]) );
  DFFPOSX1 mem_reg_28__20_ ( .D(n2482), .CLK(clk), .Q(mem[944]) );
  DFFPOSX1 mem_reg_28__19_ ( .D(n2481), .CLK(clk), .Q(mem[943]) );
  DFFPOSX1 mem_reg_28__18_ ( .D(n2480), .CLK(clk), .Q(mem[942]) );
  DFFPOSX1 mem_reg_28__17_ ( .D(n2479), .CLK(clk), .Q(mem[941]) );
  DFFPOSX1 mem_reg_28__16_ ( .D(n2478), .CLK(clk), .Q(mem[940]) );
  DFFPOSX1 mem_reg_28__15_ ( .D(n2477), .CLK(clk), .Q(mem[939]) );
  DFFPOSX1 mem_reg_28__14_ ( .D(n2476), .CLK(clk), .Q(mem[938]) );
  DFFPOSX1 mem_reg_28__13_ ( .D(n2475), .CLK(clk), .Q(mem[937]) );
  DFFPOSX1 mem_reg_28__12_ ( .D(n2474), .CLK(clk), .Q(mem[936]) );
  DFFPOSX1 mem_reg_28__11_ ( .D(n2473), .CLK(clk), .Q(mem[935]) );
  DFFPOSX1 mem_reg_28__10_ ( .D(n2472), .CLK(clk), .Q(mem[934]) );
  DFFPOSX1 mem_reg_28__9_ ( .D(n2471), .CLK(clk), .Q(mem[933]) );
  DFFPOSX1 mem_reg_28__8_ ( .D(n2470), .CLK(clk), .Q(mem[932]) );
  DFFPOSX1 mem_reg_28__7_ ( .D(n2469), .CLK(clk), .Q(mem[931]) );
  DFFPOSX1 mem_reg_28__6_ ( .D(n2468), .CLK(clk), .Q(mem[930]) );
  DFFPOSX1 mem_reg_28__5_ ( .D(n2467), .CLK(clk), .Q(mem[929]) );
  DFFPOSX1 mem_reg_28__4_ ( .D(n2466), .CLK(clk), .Q(mem[928]) );
  DFFPOSX1 mem_reg_28__3_ ( .D(n2465), .CLK(clk), .Q(mem[927]) );
  DFFPOSX1 mem_reg_28__2_ ( .D(n2464), .CLK(clk), .Q(mem[926]) );
  DFFPOSX1 mem_reg_28__1_ ( .D(n2463), .CLK(clk), .Q(mem[925]) );
  DFFPOSX1 mem_reg_28__0_ ( .D(n2462), .CLK(clk), .Q(mem[924]) );
  DFFPOSX1 mem_reg_27__32_ ( .D(n2461), .CLK(clk), .Q(mem[923]) );
  DFFPOSX1 mem_reg_27__31_ ( .D(n2460), .CLK(clk), .Q(mem[922]) );
  DFFPOSX1 mem_reg_27__30_ ( .D(n2459), .CLK(clk), .Q(mem[921]) );
  DFFPOSX1 mem_reg_27__29_ ( .D(n2458), .CLK(clk), .Q(mem[920]) );
  DFFPOSX1 mem_reg_27__28_ ( .D(n2457), .CLK(clk), .Q(mem[919]) );
  DFFPOSX1 mem_reg_27__27_ ( .D(n2456), .CLK(clk), .Q(mem[918]) );
  DFFPOSX1 mem_reg_27__26_ ( .D(n2455), .CLK(clk), .Q(mem[917]) );
  DFFPOSX1 mem_reg_27__25_ ( .D(n2454), .CLK(clk), .Q(mem[916]) );
  DFFPOSX1 mem_reg_27__24_ ( .D(n2453), .CLK(clk), .Q(mem[915]) );
  DFFPOSX1 mem_reg_27__23_ ( .D(n2452), .CLK(clk), .Q(mem[914]) );
  DFFPOSX1 mem_reg_27__22_ ( .D(n2451), .CLK(clk), .Q(mem[913]) );
  DFFPOSX1 mem_reg_27__21_ ( .D(n2450), .CLK(clk), .Q(mem[912]) );
  DFFPOSX1 mem_reg_27__20_ ( .D(n2449), .CLK(clk), .Q(mem[911]) );
  DFFPOSX1 mem_reg_27__19_ ( .D(n2448), .CLK(clk), .Q(mem[910]) );
  DFFPOSX1 mem_reg_27__18_ ( .D(n2447), .CLK(clk), .Q(mem[909]) );
  DFFPOSX1 mem_reg_27__17_ ( .D(n2446), .CLK(clk), .Q(mem[908]) );
  DFFPOSX1 mem_reg_27__16_ ( .D(n2445), .CLK(clk), .Q(mem[907]) );
  DFFPOSX1 mem_reg_27__15_ ( .D(n2444), .CLK(clk), .Q(mem[906]) );
  DFFPOSX1 mem_reg_27__14_ ( .D(n2443), .CLK(clk), .Q(mem[905]) );
  DFFPOSX1 mem_reg_27__13_ ( .D(n2442), .CLK(clk), .Q(mem[904]) );
  DFFPOSX1 mem_reg_27__12_ ( .D(n2441), .CLK(clk), .Q(mem[903]) );
  DFFPOSX1 mem_reg_27__11_ ( .D(n2440), .CLK(clk), .Q(mem[902]) );
  DFFPOSX1 mem_reg_27__10_ ( .D(n2439), .CLK(clk), .Q(mem[901]) );
  DFFPOSX1 mem_reg_27__9_ ( .D(n2438), .CLK(clk), .Q(mem[900]) );
  DFFPOSX1 mem_reg_27__8_ ( .D(n2437), .CLK(clk), .Q(mem[899]) );
  DFFPOSX1 mem_reg_27__7_ ( .D(n2436), .CLK(clk), .Q(mem[898]) );
  DFFPOSX1 mem_reg_27__6_ ( .D(n2435), .CLK(clk), .Q(mem[897]) );
  DFFPOSX1 mem_reg_27__5_ ( .D(n2434), .CLK(clk), .Q(mem[896]) );
  DFFPOSX1 mem_reg_27__4_ ( .D(n2433), .CLK(clk), .Q(mem[895]) );
  DFFPOSX1 mem_reg_27__3_ ( .D(n2432), .CLK(clk), .Q(mem[894]) );
  DFFPOSX1 mem_reg_27__2_ ( .D(n2431), .CLK(clk), .Q(mem[893]) );
  DFFPOSX1 mem_reg_27__1_ ( .D(n2430), .CLK(clk), .Q(mem[892]) );
  DFFPOSX1 mem_reg_27__0_ ( .D(n2429), .CLK(clk), .Q(mem[891]) );
  DFFPOSX1 mem_reg_26__32_ ( .D(n2428), .CLK(clk), .Q(mem[890]) );
  DFFPOSX1 mem_reg_26__31_ ( .D(n2427), .CLK(clk), .Q(mem[889]) );
  DFFPOSX1 mem_reg_26__30_ ( .D(n2426), .CLK(clk), .Q(mem[888]) );
  DFFPOSX1 mem_reg_26__29_ ( .D(n2425), .CLK(clk), .Q(mem[887]) );
  DFFPOSX1 mem_reg_26__28_ ( .D(n2424), .CLK(clk), .Q(mem[886]) );
  DFFPOSX1 mem_reg_26__27_ ( .D(n2423), .CLK(clk), .Q(mem[885]) );
  DFFPOSX1 mem_reg_26__26_ ( .D(n2422), .CLK(clk), .Q(mem[884]) );
  DFFPOSX1 mem_reg_26__25_ ( .D(n2421), .CLK(clk), .Q(mem[883]) );
  DFFPOSX1 mem_reg_26__24_ ( .D(n2420), .CLK(clk), .Q(mem[882]) );
  DFFPOSX1 mem_reg_26__23_ ( .D(n2419), .CLK(clk), .Q(mem[881]) );
  DFFPOSX1 mem_reg_26__22_ ( .D(n2418), .CLK(clk), .Q(mem[880]) );
  DFFPOSX1 mem_reg_26__21_ ( .D(n2417), .CLK(clk), .Q(mem[879]) );
  DFFPOSX1 mem_reg_26__20_ ( .D(n2416), .CLK(clk), .Q(mem[878]) );
  DFFPOSX1 mem_reg_26__19_ ( .D(n2415), .CLK(clk), .Q(mem[877]) );
  DFFPOSX1 mem_reg_26__18_ ( .D(n2414), .CLK(clk), .Q(mem[876]) );
  DFFPOSX1 mem_reg_26__17_ ( .D(n2413), .CLK(clk), .Q(mem[875]) );
  DFFPOSX1 mem_reg_26__16_ ( .D(n2412), .CLK(clk), .Q(mem[874]) );
  DFFPOSX1 mem_reg_26__15_ ( .D(n2411), .CLK(clk), .Q(mem[873]) );
  DFFPOSX1 mem_reg_26__14_ ( .D(n2410), .CLK(clk), .Q(mem[872]) );
  DFFPOSX1 mem_reg_26__13_ ( .D(n2409), .CLK(clk), .Q(mem[871]) );
  DFFPOSX1 mem_reg_26__12_ ( .D(n2408), .CLK(clk), .Q(mem[870]) );
  DFFPOSX1 mem_reg_26__11_ ( .D(n2407), .CLK(clk), .Q(mem[869]) );
  DFFPOSX1 mem_reg_26__10_ ( .D(n2406), .CLK(clk), .Q(mem[868]) );
  DFFPOSX1 mem_reg_26__9_ ( .D(n2405), .CLK(clk), .Q(mem[867]) );
  DFFPOSX1 mem_reg_26__8_ ( .D(n2404), .CLK(clk), .Q(mem[866]) );
  DFFPOSX1 mem_reg_26__7_ ( .D(n2403), .CLK(clk), .Q(mem[865]) );
  DFFPOSX1 mem_reg_26__6_ ( .D(n2402), .CLK(clk), .Q(mem[864]) );
  DFFPOSX1 mem_reg_26__5_ ( .D(n2401), .CLK(clk), .Q(mem[863]) );
  DFFPOSX1 mem_reg_26__4_ ( .D(n2400), .CLK(clk), .Q(mem[862]) );
  DFFPOSX1 mem_reg_26__3_ ( .D(n2399), .CLK(clk), .Q(mem[861]) );
  DFFPOSX1 mem_reg_26__2_ ( .D(n2398), .CLK(clk), .Q(mem[860]) );
  DFFPOSX1 mem_reg_26__1_ ( .D(n2397), .CLK(clk), .Q(mem[859]) );
  DFFPOSX1 mem_reg_26__0_ ( .D(n2396), .CLK(clk), .Q(mem[858]) );
  DFFPOSX1 mem_reg_25__32_ ( .D(n2395), .CLK(clk), .Q(mem[857]) );
  DFFPOSX1 mem_reg_25__31_ ( .D(n2394), .CLK(clk), .Q(mem[856]) );
  DFFPOSX1 mem_reg_25__30_ ( .D(n2393), .CLK(clk), .Q(mem[855]) );
  DFFPOSX1 mem_reg_25__29_ ( .D(n2392), .CLK(clk), .Q(mem[854]) );
  DFFPOSX1 mem_reg_25__28_ ( .D(n2391), .CLK(clk), .Q(mem[853]) );
  DFFPOSX1 mem_reg_25__27_ ( .D(n2390), .CLK(clk), .Q(mem[852]) );
  DFFPOSX1 mem_reg_25__26_ ( .D(n2389), .CLK(clk), .Q(mem[851]) );
  DFFPOSX1 mem_reg_25__25_ ( .D(n2388), .CLK(clk), .Q(mem[850]) );
  DFFPOSX1 mem_reg_25__24_ ( .D(n2387), .CLK(clk), .Q(mem[849]) );
  DFFPOSX1 mem_reg_25__23_ ( .D(n2386), .CLK(clk), .Q(mem[848]) );
  DFFPOSX1 mem_reg_25__22_ ( .D(n2385), .CLK(clk), .Q(mem[847]) );
  DFFPOSX1 mem_reg_25__21_ ( .D(n2384), .CLK(clk), .Q(mem[846]) );
  DFFPOSX1 mem_reg_25__20_ ( .D(n2383), .CLK(clk), .Q(mem[845]) );
  DFFPOSX1 mem_reg_25__19_ ( .D(n2382), .CLK(clk), .Q(mem[844]) );
  DFFPOSX1 mem_reg_25__18_ ( .D(n2381), .CLK(clk), .Q(mem[843]) );
  DFFPOSX1 mem_reg_25__17_ ( .D(n2380), .CLK(clk), .Q(mem[842]) );
  DFFPOSX1 mem_reg_25__16_ ( .D(n2379), .CLK(clk), .Q(mem[841]) );
  DFFPOSX1 mem_reg_25__15_ ( .D(n2378), .CLK(clk), .Q(mem[840]) );
  DFFPOSX1 mem_reg_25__14_ ( .D(n2377), .CLK(clk), .Q(mem[839]) );
  DFFPOSX1 mem_reg_25__13_ ( .D(n2376), .CLK(clk), .Q(mem[838]) );
  DFFPOSX1 mem_reg_25__12_ ( .D(n2375), .CLK(clk), .Q(mem[837]) );
  DFFPOSX1 mem_reg_25__11_ ( .D(n2374), .CLK(clk), .Q(mem[836]) );
  DFFPOSX1 mem_reg_25__10_ ( .D(n2373), .CLK(clk), .Q(mem[835]) );
  DFFPOSX1 mem_reg_25__9_ ( .D(n2372), .CLK(clk), .Q(mem[834]) );
  DFFPOSX1 mem_reg_25__8_ ( .D(n2371), .CLK(clk), .Q(mem[833]) );
  DFFPOSX1 mem_reg_25__7_ ( .D(n2370), .CLK(clk), .Q(mem[832]) );
  DFFPOSX1 mem_reg_25__6_ ( .D(n2369), .CLK(clk), .Q(mem[831]) );
  DFFPOSX1 mem_reg_25__5_ ( .D(n2368), .CLK(clk), .Q(mem[830]) );
  DFFPOSX1 mem_reg_25__4_ ( .D(n2367), .CLK(clk), .Q(mem[829]) );
  DFFPOSX1 mem_reg_25__3_ ( .D(n2366), .CLK(clk), .Q(mem[828]) );
  DFFPOSX1 mem_reg_25__2_ ( .D(n2365), .CLK(clk), .Q(mem[827]) );
  DFFPOSX1 mem_reg_25__1_ ( .D(n2364), .CLK(clk), .Q(mem[826]) );
  DFFPOSX1 mem_reg_25__0_ ( .D(n2363), .CLK(clk), .Q(mem[825]) );
  DFFPOSX1 mem_reg_24__32_ ( .D(n2362), .CLK(clk), .Q(mem[824]) );
  DFFPOSX1 mem_reg_24__31_ ( .D(n2361), .CLK(clk), .Q(mem[823]) );
  DFFPOSX1 mem_reg_24__30_ ( .D(n2360), .CLK(clk), .Q(mem[822]) );
  DFFPOSX1 mem_reg_24__29_ ( .D(n2359), .CLK(clk), .Q(mem[821]) );
  DFFPOSX1 mem_reg_24__28_ ( .D(n2358), .CLK(clk), .Q(mem[820]) );
  DFFPOSX1 mem_reg_24__27_ ( .D(n2357), .CLK(clk), .Q(mem[819]) );
  DFFPOSX1 mem_reg_24__26_ ( .D(n2356), .CLK(clk), .Q(mem[818]) );
  DFFPOSX1 mem_reg_24__25_ ( .D(n2355), .CLK(clk), .Q(mem[817]) );
  DFFPOSX1 mem_reg_24__24_ ( .D(n2354), .CLK(clk), .Q(mem[816]) );
  DFFPOSX1 mem_reg_24__23_ ( .D(n2353), .CLK(clk), .Q(mem[815]) );
  DFFPOSX1 mem_reg_24__22_ ( .D(n2352), .CLK(clk), .Q(mem[814]) );
  DFFPOSX1 mem_reg_24__21_ ( .D(n2351), .CLK(clk), .Q(mem[813]) );
  DFFPOSX1 mem_reg_24__20_ ( .D(n2350), .CLK(clk), .Q(mem[812]) );
  DFFPOSX1 mem_reg_24__19_ ( .D(n2349), .CLK(clk), .Q(mem[811]) );
  DFFPOSX1 mem_reg_24__18_ ( .D(n2348), .CLK(clk), .Q(mem[810]) );
  DFFPOSX1 mem_reg_24__17_ ( .D(n2347), .CLK(clk), .Q(mem[809]) );
  DFFPOSX1 mem_reg_24__16_ ( .D(n2346), .CLK(clk), .Q(mem[808]) );
  DFFPOSX1 mem_reg_24__15_ ( .D(n2345), .CLK(clk), .Q(mem[807]) );
  DFFPOSX1 mem_reg_24__14_ ( .D(n2344), .CLK(clk), .Q(mem[806]) );
  DFFPOSX1 mem_reg_24__13_ ( .D(n2343), .CLK(clk), .Q(mem[805]) );
  DFFPOSX1 mem_reg_24__12_ ( .D(n2342), .CLK(clk), .Q(mem[804]) );
  DFFPOSX1 mem_reg_24__11_ ( .D(n2341), .CLK(clk), .Q(mem[803]) );
  DFFPOSX1 mem_reg_24__10_ ( .D(n2340), .CLK(clk), .Q(mem[802]) );
  DFFPOSX1 mem_reg_24__9_ ( .D(n2339), .CLK(clk), .Q(mem[801]) );
  DFFPOSX1 mem_reg_24__8_ ( .D(n2338), .CLK(clk), .Q(mem[800]) );
  DFFPOSX1 mem_reg_24__7_ ( .D(n2337), .CLK(clk), .Q(mem[799]) );
  DFFPOSX1 mem_reg_24__6_ ( .D(n2336), .CLK(clk), .Q(mem[798]) );
  DFFPOSX1 mem_reg_24__5_ ( .D(n2335), .CLK(clk), .Q(mem[797]) );
  DFFPOSX1 mem_reg_24__4_ ( .D(n2334), .CLK(clk), .Q(mem[796]) );
  DFFPOSX1 mem_reg_24__3_ ( .D(n2333), .CLK(clk), .Q(mem[795]) );
  DFFPOSX1 mem_reg_24__2_ ( .D(n2332), .CLK(clk), .Q(mem[794]) );
  DFFPOSX1 mem_reg_24__1_ ( .D(n2331), .CLK(clk), .Q(mem[793]) );
  DFFPOSX1 mem_reg_24__0_ ( .D(n2330), .CLK(clk), .Q(mem[792]) );
  DFFPOSX1 mem_reg_23__32_ ( .D(n2329), .CLK(clk), .Q(mem[791]) );
  DFFPOSX1 mem_reg_23__31_ ( .D(n2328), .CLK(clk), .Q(mem[790]) );
  DFFPOSX1 mem_reg_23__30_ ( .D(n2327), .CLK(clk), .Q(mem[789]) );
  DFFPOSX1 mem_reg_23__29_ ( .D(n2326), .CLK(clk), .Q(mem[788]) );
  DFFPOSX1 mem_reg_23__28_ ( .D(n2325), .CLK(clk), .Q(mem[787]) );
  DFFPOSX1 mem_reg_23__27_ ( .D(n2324), .CLK(clk), .Q(mem[786]) );
  DFFPOSX1 mem_reg_23__26_ ( .D(n2323), .CLK(clk), .Q(mem[785]) );
  DFFPOSX1 mem_reg_23__25_ ( .D(n2322), .CLK(clk), .Q(mem[784]) );
  DFFPOSX1 mem_reg_23__24_ ( .D(n2321), .CLK(clk), .Q(mem[783]) );
  DFFPOSX1 mem_reg_23__23_ ( .D(n2320), .CLK(clk), .Q(mem[782]) );
  DFFPOSX1 mem_reg_23__22_ ( .D(n2319), .CLK(clk), .Q(mem[781]) );
  DFFPOSX1 mem_reg_23__21_ ( .D(n2318), .CLK(clk), .Q(mem[780]) );
  DFFPOSX1 mem_reg_23__20_ ( .D(n2317), .CLK(clk), .Q(mem[779]) );
  DFFPOSX1 mem_reg_23__19_ ( .D(n2316), .CLK(clk), .Q(mem[778]) );
  DFFPOSX1 mem_reg_23__18_ ( .D(n2315), .CLK(clk), .Q(mem[777]) );
  DFFPOSX1 mem_reg_23__17_ ( .D(n2314), .CLK(clk), .Q(mem[776]) );
  DFFPOSX1 mem_reg_23__16_ ( .D(n2313), .CLK(clk), .Q(mem[775]) );
  DFFPOSX1 mem_reg_23__15_ ( .D(n2312), .CLK(clk), .Q(mem[774]) );
  DFFPOSX1 mem_reg_23__14_ ( .D(n2311), .CLK(clk), .Q(mem[773]) );
  DFFPOSX1 mem_reg_23__13_ ( .D(n2310), .CLK(clk), .Q(mem[772]) );
  DFFPOSX1 mem_reg_23__12_ ( .D(n2309), .CLK(clk), .Q(mem[771]) );
  DFFPOSX1 mem_reg_23__11_ ( .D(n2308), .CLK(clk), .Q(mem[770]) );
  DFFPOSX1 mem_reg_23__10_ ( .D(n2307), .CLK(clk), .Q(mem[769]) );
  DFFPOSX1 mem_reg_23__9_ ( .D(n2306), .CLK(clk), .Q(mem[768]) );
  DFFPOSX1 mem_reg_23__8_ ( .D(n2305), .CLK(clk), .Q(mem[767]) );
  DFFPOSX1 mem_reg_23__7_ ( .D(n2304), .CLK(clk), .Q(mem[766]) );
  DFFPOSX1 mem_reg_23__6_ ( .D(n2303), .CLK(clk), .Q(mem[765]) );
  DFFPOSX1 mem_reg_23__5_ ( .D(n2302), .CLK(clk), .Q(mem[764]) );
  DFFPOSX1 mem_reg_23__4_ ( .D(n2301), .CLK(clk), .Q(mem[763]) );
  DFFPOSX1 mem_reg_23__3_ ( .D(n2300), .CLK(clk), .Q(mem[762]) );
  DFFPOSX1 mem_reg_23__2_ ( .D(n2299), .CLK(clk), .Q(mem[761]) );
  DFFPOSX1 mem_reg_23__1_ ( .D(n2298), .CLK(clk), .Q(mem[760]) );
  DFFPOSX1 mem_reg_23__0_ ( .D(n2297), .CLK(clk), .Q(mem[759]) );
  DFFPOSX1 mem_reg_22__32_ ( .D(n2296), .CLK(clk), .Q(mem[758]) );
  DFFPOSX1 mem_reg_22__31_ ( .D(n2295), .CLK(clk), .Q(mem[757]) );
  DFFPOSX1 mem_reg_22__30_ ( .D(n2294), .CLK(clk), .Q(mem[756]) );
  DFFPOSX1 mem_reg_22__29_ ( .D(n2293), .CLK(clk), .Q(mem[755]) );
  DFFPOSX1 mem_reg_22__28_ ( .D(n2292), .CLK(clk), .Q(mem[754]) );
  DFFPOSX1 mem_reg_22__27_ ( .D(n2291), .CLK(clk), .Q(mem[753]) );
  DFFPOSX1 mem_reg_22__26_ ( .D(n2290), .CLK(clk), .Q(mem[752]) );
  DFFPOSX1 mem_reg_22__25_ ( .D(n2289), .CLK(clk), .Q(mem[751]) );
  DFFPOSX1 mem_reg_22__24_ ( .D(n2288), .CLK(clk), .Q(mem[750]) );
  DFFPOSX1 mem_reg_22__23_ ( .D(n2287), .CLK(clk), .Q(mem[749]) );
  DFFPOSX1 mem_reg_22__22_ ( .D(n2286), .CLK(clk), .Q(mem[748]) );
  DFFPOSX1 mem_reg_22__21_ ( .D(n2285), .CLK(clk), .Q(mem[747]) );
  DFFPOSX1 mem_reg_22__20_ ( .D(n2284), .CLK(clk), .Q(mem[746]) );
  DFFPOSX1 mem_reg_22__19_ ( .D(n2283), .CLK(clk), .Q(mem[745]) );
  DFFPOSX1 mem_reg_22__18_ ( .D(n2282), .CLK(clk), .Q(mem[744]) );
  DFFPOSX1 mem_reg_22__17_ ( .D(n2281), .CLK(clk), .Q(mem[743]) );
  DFFPOSX1 mem_reg_22__16_ ( .D(n2280), .CLK(clk), .Q(mem[742]) );
  DFFPOSX1 mem_reg_22__15_ ( .D(n2279), .CLK(clk), .Q(mem[741]) );
  DFFPOSX1 mem_reg_22__14_ ( .D(n2278), .CLK(clk), .Q(mem[740]) );
  DFFPOSX1 mem_reg_22__13_ ( .D(n2277), .CLK(clk), .Q(mem[739]) );
  DFFPOSX1 mem_reg_22__12_ ( .D(n2276), .CLK(clk), .Q(mem[738]) );
  DFFPOSX1 mem_reg_22__11_ ( .D(n2275), .CLK(clk), .Q(mem[737]) );
  DFFPOSX1 mem_reg_22__10_ ( .D(n2274), .CLK(clk), .Q(mem[736]) );
  DFFPOSX1 mem_reg_22__9_ ( .D(n2273), .CLK(clk), .Q(mem[735]) );
  DFFPOSX1 mem_reg_22__8_ ( .D(n2272), .CLK(clk), .Q(mem[734]) );
  DFFPOSX1 mem_reg_22__7_ ( .D(n2271), .CLK(clk), .Q(mem[733]) );
  DFFPOSX1 mem_reg_22__6_ ( .D(n2270), .CLK(clk), .Q(mem[732]) );
  DFFPOSX1 mem_reg_22__5_ ( .D(n2269), .CLK(clk), .Q(mem[731]) );
  DFFPOSX1 mem_reg_22__4_ ( .D(n2268), .CLK(clk), .Q(mem[730]) );
  DFFPOSX1 mem_reg_22__3_ ( .D(n2267), .CLK(clk), .Q(mem[729]) );
  DFFPOSX1 mem_reg_22__2_ ( .D(n2266), .CLK(clk), .Q(mem[728]) );
  DFFPOSX1 mem_reg_22__1_ ( .D(n2265), .CLK(clk), .Q(mem[727]) );
  DFFPOSX1 mem_reg_22__0_ ( .D(n2264), .CLK(clk), .Q(mem[726]) );
  DFFPOSX1 mem_reg_21__32_ ( .D(n2263), .CLK(clk), .Q(mem[725]) );
  DFFPOSX1 mem_reg_21__31_ ( .D(n2262), .CLK(clk), .Q(mem[724]) );
  DFFPOSX1 mem_reg_21__30_ ( .D(n2261), .CLK(clk), .Q(mem[723]) );
  DFFPOSX1 mem_reg_21__29_ ( .D(n2260), .CLK(clk), .Q(mem[722]) );
  DFFPOSX1 mem_reg_21__28_ ( .D(n2259), .CLK(clk), .Q(mem[721]) );
  DFFPOSX1 mem_reg_21__27_ ( .D(n2258), .CLK(clk), .Q(mem[720]) );
  DFFPOSX1 mem_reg_21__26_ ( .D(n2257), .CLK(clk), .Q(mem[719]) );
  DFFPOSX1 mem_reg_21__25_ ( .D(n2256), .CLK(clk), .Q(mem[718]) );
  DFFPOSX1 mem_reg_21__24_ ( .D(n2255), .CLK(clk), .Q(mem[717]) );
  DFFPOSX1 mem_reg_21__23_ ( .D(n2254), .CLK(clk), .Q(mem[716]) );
  DFFPOSX1 mem_reg_21__22_ ( .D(n2253), .CLK(clk), .Q(mem[715]) );
  DFFPOSX1 mem_reg_21__21_ ( .D(n2252), .CLK(clk), .Q(mem[714]) );
  DFFPOSX1 mem_reg_21__20_ ( .D(n2251), .CLK(clk), .Q(mem[713]) );
  DFFPOSX1 mem_reg_21__19_ ( .D(n2250), .CLK(clk), .Q(mem[712]) );
  DFFPOSX1 mem_reg_21__18_ ( .D(n2249), .CLK(clk), .Q(mem[711]) );
  DFFPOSX1 mem_reg_21__17_ ( .D(n2248), .CLK(clk), .Q(mem[710]) );
  DFFPOSX1 mem_reg_21__16_ ( .D(n2247), .CLK(clk), .Q(mem[709]) );
  DFFPOSX1 mem_reg_21__15_ ( .D(n2246), .CLK(clk), .Q(mem[708]) );
  DFFPOSX1 mem_reg_21__14_ ( .D(n2245), .CLK(clk), .Q(mem[707]) );
  DFFPOSX1 mem_reg_21__13_ ( .D(n2244), .CLK(clk), .Q(mem[706]) );
  DFFPOSX1 mem_reg_21__12_ ( .D(n2243), .CLK(clk), .Q(mem[705]) );
  DFFPOSX1 mem_reg_21__11_ ( .D(n2242), .CLK(clk), .Q(mem[704]) );
  DFFPOSX1 mem_reg_21__10_ ( .D(n2241), .CLK(clk), .Q(mem[703]) );
  DFFPOSX1 mem_reg_21__9_ ( .D(n2240), .CLK(clk), .Q(mem[702]) );
  DFFPOSX1 mem_reg_21__8_ ( .D(n2239), .CLK(clk), .Q(mem[701]) );
  DFFPOSX1 mem_reg_21__7_ ( .D(n2238), .CLK(clk), .Q(mem[700]) );
  DFFPOSX1 mem_reg_21__6_ ( .D(n2237), .CLK(clk), .Q(mem[699]) );
  DFFPOSX1 mem_reg_21__5_ ( .D(n2236), .CLK(clk), .Q(mem[698]) );
  DFFPOSX1 mem_reg_21__4_ ( .D(n2235), .CLK(clk), .Q(mem[697]) );
  DFFPOSX1 mem_reg_21__3_ ( .D(n2234), .CLK(clk), .Q(mem[696]) );
  DFFPOSX1 mem_reg_21__2_ ( .D(n2233), .CLK(clk), .Q(mem[695]) );
  DFFPOSX1 mem_reg_21__1_ ( .D(n2232), .CLK(clk), .Q(mem[694]) );
  DFFPOSX1 mem_reg_21__0_ ( .D(n2231), .CLK(clk), .Q(mem[693]) );
  DFFPOSX1 mem_reg_20__32_ ( .D(n2230), .CLK(clk), .Q(mem[692]) );
  DFFPOSX1 mem_reg_20__31_ ( .D(n2229), .CLK(clk), .Q(mem[691]) );
  DFFPOSX1 mem_reg_20__30_ ( .D(n2228), .CLK(clk), .Q(mem[690]) );
  DFFPOSX1 mem_reg_20__29_ ( .D(n2227), .CLK(clk), .Q(mem[689]) );
  DFFPOSX1 mem_reg_20__28_ ( .D(n2226), .CLK(clk), .Q(mem[688]) );
  DFFPOSX1 mem_reg_20__27_ ( .D(n2225), .CLK(clk), .Q(mem[687]) );
  DFFPOSX1 mem_reg_20__26_ ( .D(n2224), .CLK(clk), .Q(mem[686]) );
  DFFPOSX1 mem_reg_20__25_ ( .D(n2223), .CLK(clk), .Q(mem[685]) );
  DFFPOSX1 mem_reg_20__24_ ( .D(n2222), .CLK(clk), .Q(mem[684]) );
  DFFPOSX1 mem_reg_20__23_ ( .D(n2221), .CLK(clk), .Q(mem[683]) );
  DFFPOSX1 mem_reg_20__22_ ( .D(n2220), .CLK(clk), .Q(mem[682]) );
  DFFPOSX1 mem_reg_20__21_ ( .D(n2219), .CLK(clk), .Q(mem[681]) );
  DFFPOSX1 mem_reg_20__20_ ( .D(n2218), .CLK(clk), .Q(mem[680]) );
  DFFPOSX1 mem_reg_20__19_ ( .D(n2217), .CLK(clk), .Q(mem[679]) );
  DFFPOSX1 mem_reg_20__18_ ( .D(n2216), .CLK(clk), .Q(mem[678]) );
  DFFPOSX1 mem_reg_20__17_ ( .D(n2215), .CLK(clk), .Q(mem[677]) );
  DFFPOSX1 mem_reg_20__16_ ( .D(n2214), .CLK(clk), .Q(mem[676]) );
  DFFPOSX1 mem_reg_20__15_ ( .D(n2213), .CLK(clk), .Q(mem[675]) );
  DFFPOSX1 mem_reg_20__14_ ( .D(n2212), .CLK(clk), .Q(mem[674]) );
  DFFPOSX1 mem_reg_20__13_ ( .D(n2211), .CLK(clk), .Q(mem[673]) );
  DFFPOSX1 mem_reg_20__12_ ( .D(n2210), .CLK(clk), .Q(mem[672]) );
  DFFPOSX1 mem_reg_20__11_ ( .D(n2209), .CLK(clk), .Q(mem[671]) );
  DFFPOSX1 mem_reg_20__10_ ( .D(n2208), .CLK(clk), .Q(mem[670]) );
  DFFPOSX1 mem_reg_20__9_ ( .D(n2207), .CLK(clk), .Q(mem[669]) );
  DFFPOSX1 mem_reg_20__8_ ( .D(n2206), .CLK(clk), .Q(mem[668]) );
  DFFPOSX1 mem_reg_20__7_ ( .D(n2205), .CLK(clk), .Q(mem[667]) );
  DFFPOSX1 mem_reg_20__6_ ( .D(n2204), .CLK(clk), .Q(mem[666]) );
  DFFPOSX1 mem_reg_20__5_ ( .D(n2203), .CLK(clk), .Q(mem[665]) );
  DFFPOSX1 mem_reg_20__4_ ( .D(n2202), .CLK(clk), .Q(mem[664]) );
  DFFPOSX1 mem_reg_20__3_ ( .D(n2201), .CLK(clk), .Q(mem[663]) );
  DFFPOSX1 mem_reg_20__2_ ( .D(n2200), .CLK(clk), .Q(mem[662]) );
  DFFPOSX1 mem_reg_20__1_ ( .D(n2199), .CLK(clk), .Q(mem[661]) );
  DFFPOSX1 mem_reg_20__0_ ( .D(n2198), .CLK(clk), .Q(mem[660]) );
  DFFPOSX1 mem_reg_19__32_ ( .D(n2197), .CLK(clk), .Q(mem[659]) );
  DFFPOSX1 mem_reg_19__31_ ( .D(n2196), .CLK(clk), .Q(mem[658]) );
  DFFPOSX1 mem_reg_19__30_ ( .D(n2195), .CLK(clk), .Q(mem[657]) );
  DFFPOSX1 mem_reg_19__29_ ( .D(n2194), .CLK(clk), .Q(mem[656]) );
  DFFPOSX1 mem_reg_19__28_ ( .D(n2193), .CLK(clk), .Q(mem[655]) );
  DFFPOSX1 mem_reg_19__27_ ( .D(n2192), .CLK(clk), .Q(mem[654]) );
  DFFPOSX1 mem_reg_19__26_ ( .D(n2191), .CLK(clk), .Q(mem[653]) );
  DFFPOSX1 mem_reg_19__25_ ( .D(n2190), .CLK(clk), .Q(mem[652]) );
  DFFPOSX1 mem_reg_19__24_ ( .D(n2189), .CLK(clk), .Q(mem[651]) );
  DFFPOSX1 mem_reg_19__23_ ( .D(n2188), .CLK(clk), .Q(mem[650]) );
  DFFPOSX1 mem_reg_19__22_ ( .D(n2187), .CLK(clk), .Q(mem[649]) );
  DFFPOSX1 mem_reg_19__21_ ( .D(n2186), .CLK(clk), .Q(mem[648]) );
  DFFPOSX1 mem_reg_19__20_ ( .D(n2185), .CLK(clk), .Q(mem[647]) );
  DFFPOSX1 mem_reg_19__19_ ( .D(n2184), .CLK(clk), .Q(mem[646]) );
  DFFPOSX1 mem_reg_19__18_ ( .D(n2183), .CLK(clk), .Q(mem[645]) );
  DFFPOSX1 mem_reg_19__17_ ( .D(n2182), .CLK(clk), .Q(mem[644]) );
  DFFPOSX1 mem_reg_19__16_ ( .D(n2181), .CLK(clk), .Q(mem[643]) );
  DFFPOSX1 mem_reg_19__15_ ( .D(n2180), .CLK(clk), .Q(mem[642]) );
  DFFPOSX1 mem_reg_19__14_ ( .D(n2179), .CLK(clk), .Q(mem[641]) );
  DFFPOSX1 mem_reg_19__13_ ( .D(n2178), .CLK(clk), .Q(mem[640]) );
  DFFPOSX1 mem_reg_19__12_ ( .D(n2177), .CLK(clk), .Q(mem[639]) );
  DFFPOSX1 mem_reg_19__11_ ( .D(n2176), .CLK(clk), .Q(mem[638]) );
  DFFPOSX1 mem_reg_19__10_ ( .D(n2175), .CLK(clk), .Q(mem[637]) );
  DFFPOSX1 mem_reg_19__9_ ( .D(n2174), .CLK(clk), .Q(mem[636]) );
  DFFPOSX1 mem_reg_19__8_ ( .D(n2173), .CLK(clk), .Q(mem[635]) );
  DFFPOSX1 mem_reg_19__7_ ( .D(n2172), .CLK(clk), .Q(mem[634]) );
  DFFPOSX1 mem_reg_19__6_ ( .D(n2171), .CLK(clk), .Q(mem[633]) );
  DFFPOSX1 mem_reg_19__5_ ( .D(n2170), .CLK(clk), .Q(mem[632]) );
  DFFPOSX1 mem_reg_19__4_ ( .D(n2169), .CLK(clk), .Q(mem[631]) );
  DFFPOSX1 mem_reg_19__3_ ( .D(n2168), .CLK(clk), .Q(mem[630]) );
  DFFPOSX1 mem_reg_19__2_ ( .D(n2167), .CLK(clk), .Q(mem[629]) );
  DFFPOSX1 mem_reg_19__1_ ( .D(n2166), .CLK(clk), .Q(mem[628]) );
  DFFPOSX1 mem_reg_19__0_ ( .D(n2165), .CLK(clk), .Q(mem[627]) );
  DFFPOSX1 mem_reg_18__32_ ( .D(n2164), .CLK(clk), .Q(mem[626]) );
  DFFPOSX1 mem_reg_18__31_ ( .D(n2163), .CLK(clk), .Q(mem[625]) );
  DFFPOSX1 mem_reg_18__30_ ( .D(n2162), .CLK(clk), .Q(mem[624]) );
  DFFPOSX1 mem_reg_18__29_ ( .D(n2161), .CLK(clk), .Q(mem[623]) );
  DFFPOSX1 mem_reg_18__28_ ( .D(n2160), .CLK(clk), .Q(mem[622]) );
  DFFPOSX1 mem_reg_18__27_ ( .D(n2159), .CLK(clk), .Q(mem[621]) );
  DFFPOSX1 mem_reg_18__26_ ( .D(n2158), .CLK(clk), .Q(mem[620]) );
  DFFPOSX1 mem_reg_18__25_ ( .D(n2157), .CLK(clk), .Q(mem[619]) );
  DFFPOSX1 mem_reg_18__24_ ( .D(n2156), .CLK(clk), .Q(mem[618]) );
  DFFPOSX1 mem_reg_18__23_ ( .D(n2155), .CLK(clk), .Q(mem[617]) );
  DFFPOSX1 mem_reg_18__22_ ( .D(n2154), .CLK(clk), .Q(mem[616]) );
  DFFPOSX1 mem_reg_18__21_ ( .D(n2153), .CLK(clk), .Q(mem[615]) );
  DFFPOSX1 mem_reg_18__20_ ( .D(n2152), .CLK(clk), .Q(mem[614]) );
  DFFPOSX1 mem_reg_18__19_ ( .D(n2151), .CLK(clk), .Q(mem[613]) );
  DFFPOSX1 mem_reg_18__18_ ( .D(n2150), .CLK(clk), .Q(mem[612]) );
  DFFPOSX1 mem_reg_18__17_ ( .D(n2149), .CLK(clk), .Q(mem[611]) );
  DFFPOSX1 mem_reg_18__16_ ( .D(n2148), .CLK(clk), .Q(mem[610]) );
  DFFPOSX1 mem_reg_18__15_ ( .D(n2147), .CLK(clk), .Q(mem[609]) );
  DFFPOSX1 mem_reg_18__14_ ( .D(n2146), .CLK(clk), .Q(mem[608]) );
  DFFPOSX1 mem_reg_18__13_ ( .D(n2145), .CLK(clk), .Q(mem[607]) );
  DFFPOSX1 mem_reg_18__12_ ( .D(n2144), .CLK(clk), .Q(mem[606]) );
  DFFPOSX1 mem_reg_18__11_ ( .D(n2143), .CLK(clk), .Q(mem[605]) );
  DFFPOSX1 mem_reg_18__10_ ( .D(n2142), .CLK(clk), .Q(mem[604]) );
  DFFPOSX1 mem_reg_18__9_ ( .D(n2141), .CLK(clk), .Q(mem[603]) );
  DFFPOSX1 mem_reg_18__8_ ( .D(n2140), .CLK(clk), .Q(mem[602]) );
  DFFPOSX1 mem_reg_18__7_ ( .D(n2139), .CLK(clk), .Q(mem[601]) );
  DFFPOSX1 mem_reg_18__6_ ( .D(n2138), .CLK(clk), .Q(mem[600]) );
  DFFPOSX1 mem_reg_18__5_ ( .D(n2137), .CLK(clk), .Q(mem[599]) );
  DFFPOSX1 mem_reg_18__4_ ( .D(n2136), .CLK(clk), .Q(mem[598]) );
  DFFPOSX1 mem_reg_18__3_ ( .D(n2135), .CLK(clk), .Q(mem[597]) );
  DFFPOSX1 mem_reg_18__2_ ( .D(n2134), .CLK(clk), .Q(mem[596]) );
  DFFPOSX1 mem_reg_18__1_ ( .D(n2133), .CLK(clk), .Q(mem[595]) );
  DFFPOSX1 mem_reg_18__0_ ( .D(n2132), .CLK(clk), .Q(mem[594]) );
  DFFPOSX1 mem_reg_17__32_ ( .D(n2131), .CLK(clk), .Q(mem[593]) );
  DFFPOSX1 mem_reg_17__31_ ( .D(n2130), .CLK(clk), .Q(mem[592]) );
  DFFPOSX1 mem_reg_17__30_ ( .D(n2129), .CLK(clk), .Q(mem[591]) );
  DFFPOSX1 mem_reg_17__29_ ( .D(n2128), .CLK(clk), .Q(mem[590]) );
  DFFPOSX1 mem_reg_17__28_ ( .D(n2127), .CLK(clk), .Q(mem[589]) );
  DFFPOSX1 mem_reg_17__27_ ( .D(n2126), .CLK(clk), .Q(mem[588]) );
  DFFPOSX1 mem_reg_17__26_ ( .D(n2125), .CLK(clk), .Q(mem[587]) );
  DFFPOSX1 mem_reg_17__25_ ( .D(n2124), .CLK(clk), .Q(mem[586]) );
  DFFPOSX1 mem_reg_17__24_ ( .D(n2123), .CLK(clk), .Q(mem[585]) );
  DFFPOSX1 mem_reg_17__23_ ( .D(n2122), .CLK(clk), .Q(mem[584]) );
  DFFPOSX1 mem_reg_17__22_ ( .D(n2121), .CLK(clk), .Q(mem[583]) );
  DFFPOSX1 mem_reg_17__21_ ( .D(n2120), .CLK(clk), .Q(mem[582]) );
  DFFPOSX1 mem_reg_17__20_ ( .D(n2119), .CLK(clk), .Q(mem[581]) );
  DFFPOSX1 mem_reg_17__19_ ( .D(n2118), .CLK(clk), .Q(mem[580]) );
  DFFPOSX1 mem_reg_17__18_ ( .D(n2117), .CLK(clk), .Q(mem[579]) );
  DFFPOSX1 mem_reg_17__17_ ( .D(n2116), .CLK(clk), .Q(mem[578]) );
  DFFPOSX1 mem_reg_17__16_ ( .D(n2115), .CLK(clk), .Q(mem[577]) );
  DFFPOSX1 mem_reg_17__15_ ( .D(n2114), .CLK(clk), .Q(mem[576]) );
  DFFPOSX1 mem_reg_17__14_ ( .D(n2113), .CLK(clk), .Q(mem[575]) );
  DFFPOSX1 mem_reg_17__13_ ( .D(n2112), .CLK(clk), .Q(mem[574]) );
  DFFPOSX1 mem_reg_17__12_ ( .D(n2111), .CLK(clk), .Q(mem[573]) );
  DFFPOSX1 mem_reg_17__11_ ( .D(n2110), .CLK(clk), .Q(mem[572]) );
  DFFPOSX1 mem_reg_17__10_ ( .D(n2109), .CLK(clk), .Q(mem[571]) );
  DFFPOSX1 mem_reg_17__9_ ( .D(n2108), .CLK(clk), .Q(mem[570]) );
  DFFPOSX1 mem_reg_17__8_ ( .D(n2107), .CLK(clk), .Q(mem[569]) );
  DFFPOSX1 mem_reg_17__7_ ( .D(n2106), .CLK(clk), .Q(mem[568]) );
  DFFPOSX1 mem_reg_17__6_ ( .D(n2105), .CLK(clk), .Q(mem[567]) );
  DFFPOSX1 mem_reg_17__5_ ( .D(n2104), .CLK(clk), .Q(mem[566]) );
  DFFPOSX1 mem_reg_17__4_ ( .D(n2103), .CLK(clk), .Q(mem[565]) );
  DFFPOSX1 mem_reg_17__3_ ( .D(n2102), .CLK(clk), .Q(mem[564]) );
  DFFPOSX1 mem_reg_17__2_ ( .D(n2101), .CLK(clk), .Q(mem[563]) );
  DFFPOSX1 mem_reg_17__1_ ( .D(n2100), .CLK(clk), .Q(mem[562]) );
  DFFPOSX1 mem_reg_17__0_ ( .D(n2099), .CLK(clk), .Q(mem[561]) );
  DFFPOSX1 mem_reg_16__32_ ( .D(n2098), .CLK(clk), .Q(mem[560]) );
  DFFPOSX1 mem_reg_16__31_ ( .D(n2097), .CLK(clk), .Q(mem[559]) );
  DFFPOSX1 mem_reg_16__30_ ( .D(n2096), .CLK(clk), .Q(mem[558]) );
  DFFPOSX1 mem_reg_16__29_ ( .D(n2095), .CLK(clk), .Q(mem[557]) );
  DFFPOSX1 mem_reg_16__28_ ( .D(n2094), .CLK(clk), .Q(mem[556]) );
  DFFPOSX1 mem_reg_16__27_ ( .D(n2093), .CLK(clk), .Q(mem[555]) );
  DFFPOSX1 mem_reg_16__26_ ( .D(n2092), .CLK(clk), .Q(mem[554]) );
  DFFPOSX1 mem_reg_16__25_ ( .D(n2091), .CLK(clk), .Q(mem[553]) );
  DFFPOSX1 mem_reg_16__24_ ( .D(n2090), .CLK(clk), .Q(mem[552]) );
  DFFPOSX1 mem_reg_16__23_ ( .D(n2089), .CLK(clk), .Q(mem[551]) );
  DFFPOSX1 mem_reg_16__22_ ( .D(n2088), .CLK(clk), .Q(mem[550]) );
  DFFPOSX1 mem_reg_16__21_ ( .D(n2087), .CLK(clk), .Q(mem[549]) );
  DFFPOSX1 mem_reg_16__20_ ( .D(n2086), .CLK(clk), .Q(mem[548]) );
  DFFPOSX1 mem_reg_16__19_ ( .D(n2085), .CLK(clk), .Q(mem[547]) );
  DFFPOSX1 mem_reg_16__18_ ( .D(n2084), .CLK(clk), .Q(mem[546]) );
  DFFPOSX1 mem_reg_16__17_ ( .D(n2083), .CLK(clk), .Q(mem[545]) );
  DFFPOSX1 mem_reg_16__16_ ( .D(n2082), .CLK(clk), .Q(mem[544]) );
  DFFPOSX1 mem_reg_16__15_ ( .D(n2081), .CLK(clk), .Q(mem[543]) );
  DFFPOSX1 mem_reg_16__14_ ( .D(n2080), .CLK(clk), .Q(mem[542]) );
  DFFPOSX1 mem_reg_16__13_ ( .D(n2079), .CLK(clk), .Q(mem[541]) );
  DFFPOSX1 mem_reg_16__12_ ( .D(n2078), .CLK(clk), .Q(mem[540]) );
  DFFPOSX1 mem_reg_16__11_ ( .D(n2077), .CLK(clk), .Q(mem[539]) );
  DFFPOSX1 mem_reg_16__10_ ( .D(n2076), .CLK(clk), .Q(mem[538]) );
  DFFPOSX1 mem_reg_16__9_ ( .D(n2075), .CLK(clk), .Q(mem[537]) );
  DFFPOSX1 mem_reg_16__8_ ( .D(n2074), .CLK(clk), .Q(mem[536]) );
  DFFPOSX1 mem_reg_16__7_ ( .D(n2073), .CLK(clk), .Q(mem[535]) );
  DFFPOSX1 mem_reg_16__6_ ( .D(n2072), .CLK(clk), .Q(mem[534]) );
  DFFPOSX1 mem_reg_16__5_ ( .D(n2071), .CLK(clk), .Q(mem[533]) );
  DFFPOSX1 mem_reg_16__4_ ( .D(n2070), .CLK(clk), .Q(mem[532]) );
  DFFPOSX1 mem_reg_16__3_ ( .D(n2069), .CLK(clk), .Q(mem[531]) );
  DFFPOSX1 mem_reg_16__2_ ( .D(n2068), .CLK(clk), .Q(mem[530]) );
  DFFPOSX1 mem_reg_16__1_ ( .D(n2067), .CLK(clk), .Q(mem[529]) );
  DFFPOSX1 mem_reg_16__0_ ( .D(n2066), .CLK(clk), .Q(mem[528]) );
  DFFPOSX1 mem_reg_15__32_ ( .D(n2065), .CLK(clk), .Q(mem[527]) );
  DFFPOSX1 mem_reg_15__31_ ( .D(n2064), .CLK(clk), .Q(mem[526]) );
  DFFPOSX1 mem_reg_15__30_ ( .D(n2063), .CLK(clk), .Q(mem[525]) );
  DFFPOSX1 mem_reg_15__29_ ( .D(n2062), .CLK(clk), .Q(mem[524]) );
  DFFPOSX1 mem_reg_15__28_ ( .D(n2061), .CLK(clk), .Q(mem[523]) );
  DFFPOSX1 mem_reg_15__27_ ( .D(n2060), .CLK(clk), .Q(mem[522]) );
  DFFPOSX1 mem_reg_15__26_ ( .D(n2059), .CLK(clk), .Q(mem[521]) );
  DFFPOSX1 mem_reg_15__25_ ( .D(n2058), .CLK(clk), .Q(mem[520]) );
  DFFPOSX1 mem_reg_15__24_ ( .D(n2057), .CLK(clk), .Q(mem[519]) );
  DFFPOSX1 mem_reg_15__23_ ( .D(n2056), .CLK(clk), .Q(mem[518]) );
  DFFPOSX1 mem_reg_15__22_ ( .D(n2055), .CLK(clk), .Q(mem[517]) );
  DFFPOSX1 mem_reg_15__21_ ( .D(n2054), .CLK(clk), .Q(mem[516]) );
  DFFPOSX1 mem_reg_15__20_ ( .D(n2053), .CLK(clk), .Q(mem[515]) );
  DFFPOSX1 mem_reg_15__19_ ( .D(n2052), .CLK(clk), .Q(mem[514]) );
  DFFPOSX1 mem_reg_15__18_ ( .D(n2051), .CLK(clk), .Q(mem[513]) );
  DFFPOSX1 mem_reg_15__17_ ( .D(n2050), .CLK(clk), .Q(mem[512]) );
  DFFPOSX1 mem_reg_15__16_ ( .D(n2049), .CLK(clk), .Q(mem[511]) );
  DFFPOSX1 mem_reg_15__15_ ( .D(n2048), .CLK(clk), .Q(mem[510]) );
  DFFPOSX1 mem_reg_15__14_ ( .D(n2047), .CLK(clk), .Q(mem[509]) );
  DFFPOSX1 mem_reg_15__13_ ( .D(n2046), .CLK(clk), .Q(mem[508]) );
  DFFPOSX1 mem_reg_15__12_ ( .D(n2045), .CLK(clk), .Q(mem[507]) );
  DFFPOSX1 mem_reg_15__11_ ( .D(n2044), .CLK(clk), .Q(mem[506]) );
  DFFPOSX1 mem_reg_15__10_ ( .D(n2043), .CLK(clk), .Q(mem[505]) );
  DFFPOSX1 mem_reg_15__9_ ( .D(n2042), .CLK(clk), .Q(mem[504]) );
  DFFPOSX1 mem_reg_15__8_ ( .D(n2041), .CLK(clk), .Q(mem[503]) );
  DFFPOSX1 mem_reg_15__7_ ( .D(n2040), .CLK(clk), .Q(mem[502]) );
  DFFPOSX1 mem_reg_15__6_ ( .D(n2039), .CLK(clk), .Q(mem[501]) );
  DFFPOSX1 mem_reg_15__5_ ( .D(n2038), .CLK(clk), .Q(mem[500]) );
  DFFPOSX1 mem_reg_15__4_ ( .D(n2037), .CLK(clk), .Q(mem[499]) );
  DFFPOSX1 mem_reg_15__3_ ( .D(n2036), .CLK(clk), .Q(mem[498]) );
  DFFPOSX1 mem_reg_15__2_ ( .D(n2035), .CLK(clk), .Q(mem[497]) );
  DFFPOSX1 mem_reg_15__1_ ( .D(n2034), .CLK(clk), .Q(mem[496]) );
  DFFPOSX1 mem_reg_15__0_ ( .D(n2033), .CLK(clk), .Q(mem[495]) );
  DFFPOSX1 mem_reg_14__32_ ( .D(n2032), .CLK(clk), .Q(mem[494]) );
  DFFPOSX1 mem_reg_14__31_ ( .D(n2031), .CLK(clk), .Q(mem[493]) );
  DFFPOSX1 mem_reg_14__30_ ( .D(n2030), .CLK(clk), .Q(mem[492]) );
  DFFPOSX1 mem_reg_14__29_ ( .D(n2029), .CLK(clk), .Q(mem[491]) );
  DFFPOSX1 mem_reg_14__28_ ( .D(n2028), .CLK(clk), .Q(mem[490]) );
  DFFPOSX1 mem_reg_14__27_ ( .D(n2027), .CLK(clk), .Q(mem[489]) );
  DFFPOSX1 mem_reg_14__26_ ( .D(n2026), .CLK(clk), .Q(mem[488]) );
  DFFPOSX1 mem_reg_14__25_ ( .D(n2025), .CLK(clk), .Q(mem[487]) );
  DFFPOSX1 mem_reg_14__24_ ( .D(n2024), .CLK(clk), .Q(mem[486]) );
  DFFPOSX1 mem_reg_14__23_ ( .D(n2023), .CLK(clk), .Q(mem[485]) );
  DFFPOSX1 mem_reg_14__22_ ( .D(n2022), .CLK(clk), .Q(mem[484]) );
  DFFPOSX1 mem_reg_14__21_ ( .D(n2021), .CLK(clk), .Q(mem[483]) );
  DFFPOSX1 mem_reg_14__20_ ( .D(n2020), .CLK(clk), .Q(mem[482]) );
  DFFPOSX1 mem_reg_14__19_ ( .D(n2019), .CLK(clk), .Q(mem[481]) );
  DFFPOSX1 mem_reg_14__18_ ( .D(n2018), .CLK(clk), .Q(mem[480]) );
  DFFPOSX1 mem_reg_14__17_ ( .D(n2017), .CLK(clk), .Q(mem[479]) );
  DFFPOSX1 mem_reg_14__16_ ( .D(n2016), .CLK(clk), .Q(mem[478]) );
  DFFPOSX1 mem_reg_14__15_ ( .D(n2015), .CLK(clk), .Q(mem[477]) );
  DFFPOSX1 mem_reg_14__14_ ( .D(n2014), .CLK(clk), .Q(mem[476]) );
  DFFPOSX1 mem_reg_14__13_ ( .D(n2013), .CLK(clk), .Q(mem[475]) );
  DFFPOSX1 mem_reg_14__12_ ( .D(n2012), .CLK(clk), .Q(mem[474]) );
  DFFPOSX1 mem_reg_14__11_ ( .D(n2011), .CLK(clk), .Q(mem[473]) );
  DFFPOSX1 mem_reg_14__10_ ( .D(n2010), .CLK(clk), .Q(mem[472]) );
  DFFPOSX1 mem_reg_14__9_ ( .D(n2009), .CLK(clk), .Q(mem[471]) );
  DFFPOSX1 mem_reg_14__8_ ( .D(n2008), .CLK(clk), .Q(mem[470]) );
  DFFPOSX1 mem_reg_14__7_ ( .D(n2007), .CLK(clk), .Q(mem[469]) );
  DFFPOSX1 mem_reg_14__6_ ( .D(n2006), .CLK(clk), .Q(mem[468]) );
  DFFPOSX1 mem_reg_14__5_ ( .D(n2005), .CLK(clk), .Q(mem[467]) );
  DFFPOSX1 mem_reg_14__4_ ( .D(n2004), .CLK(clk), .Q(mem[466]) );
  DFFPOSX1 mem_reg_14__3_ ( .D(n2003), .CLK(clk), .Q(mem[465]) );
  DFFPOSX1 mem_reg_14__2_ ( .D(n2002), .CLK(clk), .Q(mem[464]) );
  DFFPOSX1 mem_reg_14__1_ ( .D(n2001), .CLK(clk), .Q(mem[463]) );
  DFFPOSX1 mem_reg_14__0_ ( .D(n2000), .CLK(clk), .Q(mem[462]) );
  DFFPOSX1 mem_reg_13__32_ ( .D(n1999), .CLK(clk), .Q(mem[461]) );
  DFFPOSX1 mem_reg_13__31_ ( .D(n1998), .CLK(clk), .Q(mem[460]) );
  DFFPOSX1 mem_reg_13__30_ ( .D(n1997), .CLK(clk), .Q(mem[459]) );
  DFFPOSX1 mem_reg_13__29_ ( .D(n1996), .CLK(clk), .Q(mem[458]) );
  DFFPOSX1 mem_reg_13__28_ ( .D(n1995), .CLK(clk), .Q(mem[457]) );
  DFFPOSX1 mem_reg_13__27_ ( .D(n1994), .CLK(clk), .Q(mem[456]) );
  DFFPOSX1 mem_reg_13__26_ ( .D(n1993), .CLK(clk), .Q(mem[455]) );
  DFFPOSX1 mem_reg_13__25_ ( .D(n1992), .CLK(clk), .Q(mem[454]) );
  DFFPOSX1 mem_reg_13__24_ ( .D(n1991), .CLK(clk), .Q(mem[453]) );
  DFFPOSX1 mem_reg_13__23_ ( .D(n1990), .CLK(clk), .Q(mem[452]) );
  DFFPOSX1 mem_reg_13__22_ ( .D(n1989), .CLK(clk), .Q(mem[451]) );
  DFFPOSX1 mem_reg_13__21_ ( .D(n1988), .CLK(clk), .Q(mem[450]) );
  DFFPOSX1 mem_reg_13__20_ ( .D(n1987), .CLK(clk), .Q(mem[449]) );
  DFFPOSX1 mem_reg_13__19_ ( .D(n1986), .CLK(clk), .Q(mem[448]) );
  DFFPOSX1 mem_reg_13__18_ ( .D(n1985), .CLK(clk), .Q(mem[447]) );
  DFFPOSX1 mem_reg_13__17_ ( .D(n1984), .CLK(clk), .Q(mem[446]) );
  DFFPOSX1 mem_reg_13__16_ ( .D(n1983), .CLK(clk), .Q(mem[445]) );
  DFFPOSX1 mem_reg_13__15_ ( .D(n1982), .CLK(clk), .Q(mem[444]) );
  DFFPOSX1 mem_reg_13__14_ ( .D(n1981), .CLK(clk), .Q(mem[443]) );
  DFFPOSX1 mem_reg_13__13_ ( .D(n1980), .CLK(clk), .Q(mem[442]) );
  DFFPOSX1 mem_reg_13__12_ ( .D(n1979), .CLK(clk), .Q(mem[441]) );
  DFFPOSX1 mem_reg_13__11_ ( .D(n1978), .CLK(clk), .Q(mem[440]) );
  DFFPOSX1 mem_reg_13__10_ ( .D(n1977), .CLK(clk), .Q(mem[439]) );
  DFFPOSX1 mem_reg_13__9_ ( .D(n1976), .CLK(clk), .Q(mem[438]) );
  DFFPOSX1 mem_reg_13__8_ ( .D(n1975), .CLK(clk), .Q(mem[437]) );
  DFFPOSX1 mem_reg_13__7_ ( .D(n1974), .CLK(clk), .Q(mem[436]) );
  DFFPOSX1 mem_reg_13__6_ ( .D(n1973), .CLK(clk), .Q(mem[435]) );
  DFFPOSX1 mem_reg_13__5_ ( .D(n1972), .CLK(clk), .Q(mem[434]) );
  DFFPOSX1 mem_reg_13__4_ ( .D(n1971), .CLK(clk), .Q(mem[433]) );
  DFFPOSX1 mem_reg_13__3_ ( .D(n1970), .CLK(clk), .Q(mem[432]) );
  DFFPOSX1 mem_reg_13__2_ ( .D(n1969), .CLK(clk), .Q(mem[431]) );
  DFFPOSX1 mem_reg_13__1_ ( .D(n1968), .CLK(clk), .Q(mem[430]) );
  DFFPOSX1 mem_reg_13__0_ ( .D(n1967), .CLK(clk), .Q(mem[429]) );
  DFFPOSX1 mem_reg_12__32_ ( .D(n1966), .CLK(clk), .Q(mem[428]) );
  DFFPOSX1 mem_reg_12__31_ ( .D(n1965), .CLK(clk), .Q(mem[427]) );
  DFFPOSX1 mem_reg_12__30_ ( .D(n1964), .CLK(clk), .Q(mem[426]) );
  DFFPOSX1 mem_reg_12__29_ ( .D(n1963), .CLK(clk), .Q(mem[425]) );
  DFFPOSX1 mem_reg_12__28_ ( .D(n1962), .CLK(clk), .Q(mem[424]) );
  DFFPOSX1 mem_reg_12__27_ ( .D(n1961), .CLK(clk), .Q(mem[423]) );
  DFFPOSX1 mem_reg_12__26_ ( .D(n1960), .CLK(clk), .Q(mem[422]) );
  DFFPOSX1 mem_reg_12__25_ ( .D(n1959), .CLK(clk), .Q(mem[421]) );
  DFFPOSX1 mem_reg_12__24_ ( .D(n1958), .CLK(clk), .Q(mem[420]) );
  DFFPOSX1 mem_reg_12__23_ ( .D(n1957), .CLK(clk), .Q(mem[419]) );
  DFFPOSX1 mem_reg_12__22_ ( .D(n1956), .CLK(clk), .Q(mem[418]) );
  DFFPOSX1 mem_reg_12__21_ ( .D(n1955), .CLK(clk), .Q(mem[417]) );
  DFFPOSX1 mem_reg_12__20_ ( .D(n1954), .CLK(clk), .Q(mem[416]) );
  DFFPOSX1 mem_reg_12__19_ ( .D(n1953), .CLK(clk), .Q(mem[415]) );
  DFFPOSX1 mem_reg_12__18_ ( .D(n1952), .CLK(clk), .Q(mem[414]) );
  DFFPOSX1 mem_reg_12__17_ ( .D(n1951), .CLK(clk), .Q(mem[413]) );
  DFFPOSX1 mem_reg_12__16_ ( .D(n1950), .CLK(clk), .Q(mem[412]) );
  DFFPOSX1 mem_reg_12__15_ ( .D(n1949), .CLK(clk), .Q(mem[411]) );
  DFFPOSX1 mem_reg_12__14_ ( .D(n1948), .CLK(clk), .Q(mem[410]) );
  DFFPOSX1 mem_reg_12__13_ ( .D(n1947), .CLK(clk), .Q(mem[409]) );
  DFFPOSX1 mem_reg_12__12_ ( .D(n1946), .CLK(clk), .Q(mem[408]) );
  DFFPOSX1 mem_reg_12__11_ ( .D(n1945), .CLK(clk), .Q(mem[407]) );
  DFFPOSX1 mem_reg_12__10_ ( .D(n1944), .CLK(clk), .Q(mem[406]) );
  DFFPOSX1 mem_reg_12__9_ ( .D(n1943), .CLK(clk), .Q(mem[405]) );
  DFFPOSX1 mem_reg_12__8_ ( .D(n1942), .CLK(clk), .Q(mem[404]) );
  DFFPOSX1 mem_reg_12__7_ ( .D(n1941), .CLK(clk), .Q(mem[403]) );
  DFFPOSX1 mem_reg_12__6_ ( .D(n1940), .CLK(clk), .Q(mem[402]) );
  DFFPOSX1 mem_reg_12__5_ ( .D(n1939), .CLK(clk), .Q(mem[401]) );
  DFFPOSX1 mem_reg_12__4_ ( .D(n1938), .CLK(clk), .Q(mem[400]) );
  DFFPOSX1 mem_reg_12__3_ ( .D(n1937), .CLK(clk), .Q(mem[399]) );
  DFFPOSX1 mem_reg_12__2_ ( .D(n1936), .CLK(clk), .Q(mem[398]) );
  DFFPOSX1 mem_reg_12__1_ ( .D(n1935), .CLK(clk), .Q(mem[397]) );
  DFFPOSX1 mem_reg_12__0_ ( .D(n1934), .CLK(clk), .Q(mem[396]) );
  DFFPOSX1 mem_reg_11__32_ ( .D(n1933), .CLK(clk), .Q(mem[395]) );
  DFFPOSX1 mem_reg_11__31_ ( .D(n1932), .CLK(clk), .Q(mem[394]) );
  DFFPOSX1 mem_reg_11__30_ ( .D(n1931), .CLK(clk), .Q(mem[393]) );
  DFFPOSX1 mem_reg_11__29_ ( .D(n1930), .CLK(clk), .Q(mem[392]) );
  DFFPOSX1 mem_reg_11__28_ ( .D(n1929), .CLK(clk), .Q(mem[391]) );
  DFFPOSX1 mem_reg_11__27_ ( .D(n1928), .CLK(clk), .Q(mem[390]) );
  DFFPOSX1 mem_reg_11__26_ ( .D(n1927), .CLK(clk), .Q(mem[389]) );
  DFFPOSX1 mem_reg_11__25_ ( .D(n1926), .CLK(clk), .Q(mem[388]) );
  DFFPOSX1 mem_reg_11__24_ ( .D(n1925), .CLK(clk), .Q(mem[387]) );
  DFFPOSX1 mem_reg_11__23_ ( .D(n1924), .CLK(clk), .Q(mem[386]) );
  DFFPOSX1 mem_reg_11__22_ ( .D(n1923), .CLK(clk), .Q(mem[385]) );
  DFFPOSX1 mem_reg_11__21_ ( .D(n1922), .CLK(clk), .Q(mem[384]) );
  DFFPOSX1 mem_reg_11__20_ ( .D(n1921), .CLK(clk), .Q(mem[383]) );
  DFFPOSX1 mem_reg_11__19_ ( .D(n1920), .CLK(clk), .Q(mem[382]) );
  DFFPOSX1 mem_reg_11__18_ ( .D(n1919), .CLK(clk), .Q(mem[381]) );
  DFFPOSX1 mem_reg_11__17_ ( .D(n1918), .CLK(clk), .Q(mem[380]) );
  DFFPOSX1 mem_reg_11__16_ ( .D(n1917), .CLK(clk), .Q(mem[379]) );
  DFFPOSX1 mem_reg_11__15_ ( .D(n1916), .CLK(clk), .Q(mem[378]) );
  DFFPOSX1 mem_reg_11__14_ ( .D(n1915), .CLK(clk), .Q(mem[377]) );
  DFFPOSX1 mem_reg_11__13_ ( .D(n1914), .CLK(clk), .Q(mem[376]) );
  DFFPOSX1 mem_reg_11__12_ ( .D(n1913), .CLK(clk), .Q(mem[375]) );
  DFFPOSX1 mem_reg_11__11_ ( .D(n1912), .CLK(clk), .Q(mem[374]) );
  DFFPOSX1 mem_reg_11__10_ ( .D(n1911), .CLK(clk), .Q(mem[373]) );
  DFFPOSX1 mem_reg_11__9_ ( .D(n1910), .CLK(clk), .Q(mem[372]) );
  DFFPOSX1 mem_reg_11__8_ ( .D(n1909), .CLK(clk), .Q(mem[371]) );
  DFFPOSX1 mem_reg_11__7_ ( .D(n1908), .CLK(clk), .Q(mem[370]) );
  DFFPOSX1 mem_reg_11__6_ ( .D(n1907), .CLK(clk), .Q(mem[369]) );
  DFFPOSX1 mem_reg_11__5_ ( .D(n1906), .CLK(clk), .Q(mem[368]) );
  DFFPOSX1 mem_reg_11__4_ ( .D(n1905), .CLK(clk), .Q(mem[367]) );
  DFFPOSX1 mem_reg_11__3_ ( .D(n1904), .CLK(clk), .Q(mem[366]) );
  DFFPOSX1 mem_reg_11__2_ ( .D(n1903), .CLK(clk), .Q(mem[365]) );
  DFFPOSX1 mem_reg_11__1_ ( .D(n1902), .CLK(clk), .Q(mem[364]) );
  DFFPOSX1 mem_reg_11__0_ ( .D(n1901), .CLK(clk), .Q(mem[363]) );
  DFFPOSX1 mem_reg_10__32_ ( .D(n1900), .CLK(clk), .Q(mem[362]) );
  DFFPOSX1 mem_reg_10__31_ ( .D(n1899), .CLK(clk), .Q(mem[361]) );
  DFFPOSX1 mem_reg_10__30_ ( .D(n1898), .CLK(clk), .Q(mem[360]) );
  DFFPOSX1 mem_reg_10__29_ ( .D(n1897), .CLK(clk), .Q(mem[359]) );
  DFFPOSX1 mem_reg_10__28_ ( .D(n1896), .CLK(clk), .Q(mem[358]) );
  DFFPOSX1 mem_reg_10__27_ ( .D(n1895), .CLK(clk), .Q(mem[357]) );
  DFFPOSX1 mem_reg_10__26_ ( .D(n1894), .CLK(clk), .Q(mem[356]) );
  DFFPOSX1 mem_reg_10__25_ ( .D(n1893), .CLK(clk), .Q(mem[355]) );
  DFFPOSX1 mem_reg_10__24_ ( .D(n1892), .CLK(clk), .Q(mem[354]) );
  DFFPOSX1 mem_reg_10__23_ ( .D(n1891), .CLK(clk), .Q(mem[353]) );
  DFFPOSX1 mem_reg_10__22_ ( .D(n1890), .CLK(clk), .Q(mem[352]) );
  DFFPOSX1 mem_reg_10__21_ ( .D(n1889), .CLK(clk), .Q(mem[351]) );
  DFFPOSX1 mem_reg_10__20_ ( .D(n1888), .CLK(clk), .Q(mem[350]) );
  DFFPOSX1 mem_reg_10__19_ ( .D(n1887), .CLK(clk), .Q(mem[349]) );
  DFFPOSX1 mem_reg_10__18_ ( .D(n1886), .CLK(clk), .Q(mem[348]) );
  DFFPOSX1 mem_reg_10__17_ ( .D(n1885), .CLK(clk), .Q(mem[347]) );
  DFFPOSX1 mem_reg_10__16_ ( .D(n1884), .CLK(clk), .Q(mem[346]) );
  DFFPOSX1 mem_reg_10__15_ ( .D(n1883), .CLK(clk), .Q(mem[345]) );
  DFFPOSX1 mem_reg_10__14_ ( .D(n1882), .CLK(clk), .Q(mem[344]) );
  DFFPOSX1 mem_reg_10__13_ ( .D(n1881), .CLK(clk), .Q(mem[343]) );
  DFFPOSX1 mem_reg_10__12_ ( .D(n1880), .CLK(clk), .Q(mem[342]) );
  DFFPOSX1 mem_reg_10__11_ ( .D(n1879), .CLK(clk), .Q(mem[341]) );
  DFFPOSX1 mem_reg_10__10_ ( .D(n1878), .CLK(clk), .Q(mem[340]) );
  DFFPOSX1 mem_reg_10__9_ ( .D(n1877), .CLK(clk), .Q(mem[339]) );
  DFFPOSX1 mem_reg_10__8_ ( .D(n1876), .CLK(clk), .Q(mem[338]) );
  DFFPOSX1 mem_reg_10__7_ ( .D(n1875), .CLK(clk), .Q(mem[337]) );
  DFFPOSX1 mem_reg_10__6_ ( .D(n1874), .CLK(clk), .Q(mem[336]) );
  DFFPOSX1 mem_reg_10__5_ ( .D(n1873), .CLK(clk), .Q(mem[335]) );
  DFFPOSX1 mem_reg_10__4_ ( .D(n1872), .CLK(clk), .Q(mem[334]) );
  DFFPOSX1 mem_reg_10__3_ ( .D(n1871), .CLK(clk), .Q(mem[333]) );
  DFFPOSX1 mem_reg_10__2_ ( .D(n1870), .CLK(clk), .Q(mem[332]) );
  DFFPOSX1 mem_reg_10__1_ ( .D(n1869), .CLK(clk), .Q(mem[331]) );
  DFFPOSX1 mem_reg_10__0_ ( .D(n1868), .CLK(clk), .Q(mem[330]) );
  DFFPOSX1 mem_reg_9__32_ ( .D(n1867), .CLK(clk), .Q(mem[329]) );
  DFFPOSX1 mem_reg_9__31_ ( .D(n1866), .CLK(clk), .Q(mem[328]) );
  DFFPOSX1 mem_reg_9__30_ ( .D(n1865), .CLK(clk), .Q(mem[327]) );
  DFFPOSX1 mem_reg_9__29_ ( .D(n1864), .CLK(clk), .Q(mem[326]) );
  DFFPOSX1 mem_reg_9__28_ ( .D(n1863), .CLK(clk), .Q(mem[325]) );
  DFFPOSX1 mem_reg_9__27_ ( .D(n1862), .CLK(clk), .Q(mem[324]) );
  DFFPOSX1 mem_reg_9__26_ ( .D(n1861), .CLK(clk), .Q(mem[323]) );
  DFFPOSX1 mem_reg_9__25_ ( .D(n1860), .CLK(clk), .Q(mem[322]) );
  DFFPOSX1 mem_reg_9__24_ ( .D(n1859), .CLK(clk), .Q(mem[321]) );
  DFFPOSX1 mem_reg_9__23_ ( .D(n1858), .CLK(clk), .Q(mem[320]) );
  DFFPOSX1 mem_reg_9__22_ ( .D(n1857), .CLK(clk), .Q(mem[319]) );
  DFFPOSX1 mem_reg_9__21_ ( .D(n1856), .CLK(clk), .Q(mem[318]) );
  DFFPOSX1 mem_reg_9__20_ ( .D(n1855), .CLK(clk), .Q(mem[317]) );
  DFFPOSX1 mem_reg_9__19_ ( .D(n1854), .CLK(clk), .Q(mem[316]) );
  DFFPOSX1 mem_reg_9__18_ ( .D(n1853), .CLK(clk), .Q(mem[315]) );
  DFFPOSX1 mem_reg_9__17_ ( .D(n1852), .CLK(clk), .Q(mem[314]) );
  DFFPOSX1 mem_reg_9__16_ ( .D(n1851), .CLK(clk), .Q(mem[313]) );
  DFFPOSX1 mem_reg_9__15_ ( .D(n1850), .CLK(clk), .Q(mem[312]) );
  DFFPOSX1 mem_reg_9__14_ ( .D(n1849), .CLK(clk), .Q(mem[311]) );
  DFFPOSX1 mem_reg_9__13_ ( .D(n1848), .CLK(clk), .Q(mem[310]) );
  DFFPOSX1 mem_reg_9__12_ ( .D(n1847), .CLK(clk), .Q(mem[309]) );
  DFFPOSX1 mem_reg_9__11_ ( .D(n1846), .CLK(clk), .Q(mem[308]) );
  DFFPOSX1 mem_reg_9__10_ ( .D(n1845), .CLK(clk), .Q(mem[307]) );
  DFFPOSX1 mem_reg_9__9_ ( .D(n1844), .CLK(clk), .Q(mem[306]) );
  DFFPOSX1 mem_reg_9__8_ ( .D(n1843), .CLK(clk), .Q(mem[305]) );
  DFFPOSX1 mem_reg_9__7_ ( .D(n1842), .CLK(clk), .Q(mem[304]) );
  DFFPOSX1 mem_reg_9__6_ ( .D(n1841), .CLK(clk), .Q(mem[303]) );
  DFFPOSX1 mem_reg_9__5_ ( .D(n1840), .CLK(clk), .Q(mem[302]) );
  DFFPOSX1 mem_reg_9__4_ ( .D(n1839), .CLK(clk), .Q(mem[301]) );
  DFFPOSX1 mem_reg_9__3_ ( .D(n1838), .CLK(clk), .Q(mem[300]) );
  DFFPOSX1 mem_reg_9__2_ ( .D(n1837), .CLK(clk), .Q(mem[299]) );
  DFFPOSX1 mem_reg_9__1_ ( .D(n1836), .CLK(clk), .Q(mem[298]) );
  DFFPOSX1 mem_reg_9__0_ ( .D(n1835), .CLK(clk), .Q(mem[297]) );
  DFFPOSX1 mem_reg_8__32_ ( .D(n1834), .CLK(clk), .Q(mem[296]) );
  DFFPOSX1 mem_reg_8__31_ ( .D(n1833), .CLK(clk), .Q(mem[295]) );
  DFFPOSX1 mem_reg_8__30_ ( .D(n1832), .CLK(clk), .Q(mem[294]) );
  DFFPOSX1 mem_reg_8__29_ ( .D(n1831), .CLK(clk), .Q(mem[293]) );
  DFFPOSX1 mem_reg_8__28_ ( .D(n1830), .CLK(clk), .Q(mem[292]) );
  DFFPOSX1 mem_reg_8__27_ ( .D(n1829), .CLK(clk), .Q(mem[291]) );
  DFFPOSX1 mem_reg_8__26_ ( .D(n1828), .CLK(clk), .Q(mem[290]) );
  DFFPOSX1 mem_reg_8__25_ ( .D(n1827), .CLK(clk), .Q(mem[289]) );
  DFFPOSX1 mem_reg_8__24_ ( .D(n1826), .CLK(clk), .Q(mem[288]) );
  DFFPOSX1 mem_reg_8__23_ ( .D(n1825), .CLK(clk), .Q(mem[287]) );
  DFFPOSX1 mem_reg_8__22_ ( .D(n1824), .CLK(clk), .Q(mem[286]) );
  DFFPOSX1 mem_reg_8__21_ ( .D(n1823), .CLK(clk), .Q(mem[285]) );
  DFFPOSX1 mem_reg_8__20_ ( .D(n1822), .CLK(clk), .Q(mem[284]) );
  DFFPOSX1 mem_reg_8__19_ ( .D(n1821), .CLK(clk), .Q(mem[283]) );
  DFFPOSX1 mem_reg_8__18_ ( .D(n1820), .CLK(clk), .Q(mem[282]) );
  DFFPOSX1 mem_reg_8__17_ ( .D(n1819), .CLK(clk), .Q(mem[281]) );
  DFFPOSX1 mem_reg_8__16_ ( .D(n1818), .CLK(clk), .Q(mem[280]) );
  DFFPOSX1 mem_reg_8__15_ ( .D(n1817), .CLK(clk), .Q(mem[279]) );
  DFFPOSX1 mem_reg_8__14_ ( .D(n1816), .CLK(clk), .Q(mem[278]) );
  DFFPOSX1 mem_reg_8__13_ ( .D(n1815), .CLK(clk), .Q(mem[277]) );
  DFFPOSX1 mem_reg_8__12_ ( .D(n1814), .CLK(clk), .Q(mem[276]) );
  DFFPOSX1 mem_reg_8__11_ ( .D(n1813), .CLK(clk), .Q(mem[275]) );
  DFFPOSX1 mem_reg_8__10_ ( .D(n1812), .CLK(clk), .Q(mem[274]) );
  DFFPOSX1 mem_reg_8__9_ ( .D(n1811), .CLK(clk), .Q(mem[273]) );
  DFFPOSX1 mem_reg_8__8_ ( .D(n1810), .CLK(clk), .Q(mem[272]) );
  DFFPOSX1 mem_reg_8__7_ ( .D(n1809), .CLK(clk), .Q(mem[271]) );
  DFFPOSX1 mem_reg_8__6_ ( .D(n1808), .CLK(clk), .Q(mem[270]) );
  DFFPOSX1 mem_reg_8__5_ ( .D(n1807), .CLK(clk), .Q(mem[269]) );
  DFFPOSX1 mem_reg_8__4_ ( .D(n1806), .CLK(clk), .Q(mem[268]) );
  DFFPOSX1 mem_reg_8__3_ ( .D(n1805), .CLK(clk), .Q(mem[267]) );
  DFFPOSX1 mem_reg_8__2_ ( .D(n1804), .CLK(clk), .Q(mem[266]) );
  DFFPOSX1 mem_reg_8__1_ ( .D(n1803), .CLK(clk), .Q(mem[265]) );
  DFFPOSX1 mem_reg_8__0_ ( .D(n1802), .CLK(clk), .Q(mem[264]) );
  DFFPOSX1 mem_reg_7__32_ ( .D(n1801), .CLK(clk), .Q(mem[263]) );
  DFFPOSX1 mem_reg_7__31_ ( .D(n1800), .CLK(clk), .Q(mem[262]) );
  DFFPOSX1 mem_reg_7__30_ ( .D(n1799), .CLK(clk), .Q(mem[261]) );
  DFFPOSX1 mem_reg_7__29_ ( .D(n1798), .CLK(clk), .Q(mem[260]) );
  DFFPOSX1 mem_reg_7__28_ ( .D(n1797), .CLK(clk), .Q(mem[259]) );
  DFFPOSX1 mem_reg_7__27_ ( .D(n1796), .CLK(clk), .Q(mem[258]) );
  DFFPOSX1 mem_reg_7__26_ ( .D(n1795), .CLK(clk), .Q(mem[257]) );
  DFFPOSX1 mem_reg_7__25_ ( .D(n1794), .CLK(clk), .Q(mem[256]) );
  DFFPOSX1 mem_reg_7__24_ ( .D(n1793), .CLK(clk), .Q(mem[255]) );
  DFFPOSX1 mem_reg_7__23_ ( .D(n1792), .CLK(clk), .Q(mem[254]) );
  DFFPOSX1 mem_reg_7__22_ ( .D(n1791), .CLK(clk), .Q(mem[253]) );
  DFFPOSX1 mem_reg_7__21_ ( .D(n1790), .CLK(clk), .Q(mem[252]) );
  DFFPOSX1 mem_reg_7__20_ ( .D(n1789), .CLK(clk), .Q(mem[251]) );
  DFFPOSX1 mem_reg_7__19_ ( .D(n1788), .CLK(clk), .Q(mem[250]) );
  DFFPOSX1 mem_reg_7__18_ ( .D(n1787), .CLK(clk), .Q(mem[249]) );
  DFFPOSX1 mem_reg_7__17_ ( .D(n1786), .CLK(clk), .Q(mem[248]) );
  DFFPOSX1 mem_reg_7__16_ ( .D(n1785), .CLK(clk), .Q(mem[247]) );
  DFFPOSX1 mem_reg_7__15_ ( .D(n1784), .CLK(clk), .Q(mem[246]) );
  DFFPOSX1 mem_reg_7__14_ ( .D(n1783), .CLK(clk), .Q(mem[245]) );
  DFFPOSX1 mem_reg_7__13_ ( .D(n1782), .CLK(clk), .Q(mem[244]) );
  DFFPOSX1 mem_reg_7__12_ ( .D(n1781), .CLK(clk), .Q(mem[243]) );
  DFFPOSX1 mem_reg_7__11_ ( .D(n1780), .CLK(clk), .Q(mem[242]) );
  DFFPOSX1 mem_reg_7__10_ ( .D(n1779), .CLK(clk), .Q(mem[241]) );
  DFFPOSX1 mem_reg_7__9_ ( .D(n1778), .CLK(clk), .Q(mem[240]) );
  DFFPOSX1 mem_reg_7__8_ ( .D(n1777), .CLK(clk), .Q(mem[239]) );
  DFFPOSX1 mem_reg_7__7_ ( .D(n1776), .CLK(clk), .Q(mem[238]) );
  DFFPOSX1 mem_reg_7__6_ ( .D(n1775), .CLK(clk), .Q(mem[237]) );
  DFFPOSX1 mem_reg_7__5_ ( .D(n1774), .CLK(clk), .Q(mem[236]) );
  DFFPOSX1 mem_reg_7__4_ ( .D(n1773), .CLK(clk), .Q(mem[235]) );
  DFFPOSX1 mem_reg_7__3_ ( .D(n1772), .CLK(clk), .Q(mem[234]) );
  DFFPOSX1 mem_reg_7__2_ ( .D(n1771), .CLK(clk), .Q(mem[233]) );
  DFFPOSX1 mem_reg_7__1_ ( .D(n1770), .CLK(clk), .Q(mem[232]) );
  DFFPOSX1 mem_reg_7__0_ ( .D(n1769), .CLK(clk), .Q(mem[231]) );
  DFFPOSX1 mem_reg_6__32_ ( .D(n1768), .CLK(clk), .Q(mem[230]) );
  DFFPOSX1 mem_reg_6__31_ ( .D(n1767), .CLK(clk), .Q(mem[229]) );
  DFFPOSX1 mem_reg_6__30_ ( .D(n1766), .CLK(clk), .Q(mem[228]) );
  DFFPOSX1 mem_reg_6__29_ ( .D(n1765), .CLK(clk), .Q(mem[227]) );
  DFFPOSX1 mem_reg_6__28_ ( .D(n1764), .CLK(clk), .Q(mem[226]) );
  DFFPOSX1 mem_reg_6__27_ ( .D(n1763), .CLK(clk), .Q(mem[225]) );
  DFFPOSX1 mem_reg_6__26_ ( .D(n1762), .CLK(clk), .Q(mem[224]) );
  DFFPOSX1 mem_reg_6__25_ ( .D(n1761), .CLK(clk), .Q(mem[223]) );
  DFFPOSX1 mem_reg_6__24_ ( .D(n1760), .CLK(clk), .Q(mem[222]) );
  DFFPOSX1 mem_reg_6__23_ ( .D(n1759), .CLK(clk), .Q(mem[221]) );
  DFFPOSX1 mem_reg_6__22_ ( .D(n1758), .CLK(clk), .Q(mem[220]) );
  DFFPOSX1 mem_reg_6__21_ ( .D(n1757), .CLK(clk), .Q(mem[219]) );
  DFFPOSX1 mem_reg_6__20_ ( .D(n1756), .CLK(clk), .Q(mem[218]) );
  DFFPOSX1 mem_reg_6__19_ ( .D(n1755), .CLK(clk), .Q(mem[217]) );
  DFFPOSX1 mem_reg_6__18_ ( .D(n1754), .CLK(clk), .Q(mem[216]) );
  DFFPOSX1 mem_reg_6__17_ ( .D(n1753), .CLK(clk), .Q(mem[215]) );
  DFFPOSX1 mem_reg_6__16_ ( .D(n1752), .CLK(clk), .Q(mem[214]) );
  DFFPOSX1 mem_reg_6__15_ ( .D(n1751), .CLK(clk), .Q(mem[213]) );
  DFFPOSX1 mem_reg_6__14_ ( .D(n1750), .CLK(clk), .Q(mem[212]) );
  DFFPOSX1 mem_reg_6__13_ ( .D(n1749), .CLK(clk), .Q(mem[211]) );
  DFFPOSX1 mem_reg_6__12_ ( .D(n1748), .CLK(clk), .Q(mem[210]) );
  DFFPOSX1 mem_reg_6__11_ ( .D(n1747), .CLK(clk), .Q(mem[209]) );
  DFFPOSX1 mem_reg_6__10_ ( .D(n1746), .CLK(clk), .Q(mem[208]) );
  DFFPOSX1 mem_reg_6__9_ ( .D(n1745), .CLK(clk), .Q(mem[207]) );
  DFFPOSX1 mem_reg_6__8_ ( .D(n1744), .CLK(clk), .Q(mem[206]) );
  DFFPOSX1 mem_reg_6__7_ ( .D(n1743), .CLK(clk), .Q(mem[205]) );
  DFFPOSX1 mem_reg_6__6_ ( .D(n1742), .CLK(clk), .Q(mem[204]) );
  DFFPOSX1 mem_reg_6__5_ ( .D(n1741), .CLK(clk), .Q(mem[203]) );
  DFFPOSX1 mem_reg_6__4_ ( .D(n1740), .CLK(clk), .Q(mem[202]) );
  DFFPOSX1 mem_reg_6__3_ ( .D(n1739), .CLK(clk), .Q(mem[201]) );
  DFFPOSX1 mem_reg_6__2_ ( .D(n1738), .CLK(clk), .Q(mem[200]) );
  DFFPOSX1 mem_reg_6__1_ ( .D(n1737), .CLK(clk), .Q(mem[199]) );
  DFFPOSX1 mem_reg_6__0_ ( .D(n1736), .CLK(clk), .Q(mem[198]) );
  DFFPOSX1 mem_reg_5__32_ ( .D(n1735), .CLK(clk), .Q(mem[197]) );
  DFFPOSX1 mem_reg_5__31_ ( .D(n1734), .CLK(clk), .Q(mem[196]) );
  DFFPOSX1 mem_reg_5__30_ ( .D(n1733), .CLK(clk), .Q(mem[195]) );
  DFFPOSX1 mem_reg_5__29_ ( .D(n1732), .CLK(clk), .Q(mem[194]) );
  DFFPOSX1 mem_reg_5__28_ ( .D(n1731), .CLK(clk), .Q(mem[193]) );
  DFFPOSX1 mem_reg_5__27_ ( .D(n1730), .CLK(clk), .Q(mem[192]) );
  DFFPOSX1 mem_reg_5__26_ ( .D(n1729), .CLK(clk), .Q(mem[191]) );
  DFFPOSX1 mem_reg_5__25_ ( .D(n1728), .CLK(clk), .Q(mem[190]) );
  DFFPOSX1 mem_reg_5__24_ ( .D(n1727), .CLK(clk), .Q(mem[189]) );
  DFFPOSX1 mem_reg_5__23_ ( .D(n1726), .CLK(clk), .Q(mem[188]) );
  DFFPOSX1 mem_reg_5__22_ ( .D(n1725), .CLK(clk), .Q(mem[187]) );
  DFFPOSX1 mem_reg_5__21_ ( .D(n1724), .CLK(clk), .Q(mem[186]) );
  DFFPOSX1 mem_reg_5__20_ ( .D(n1723), .CLK(clk), .Q(mem[185]) );
  DFFPOSX1 mem_reg_5__19_ ( .D(n1722), .CLK(clk), .Q(mem[184]) );
  DFFPOSX1 mem_reg_5__18_ ( .D(n1721), .CLK(clk), .Q(mem[183]) );
  DFFPOSX1 mem_reg_5__17_ ( .D(n1720), .CLK(clk), .Q(mem[182]) );
  DFFPOSX1 mem_reg_5__16_ ( .D(n1719), .CLK(clk), .Q(mem[181]) );
  DFFPOSX1 mem_reg_5__15_ ( .D(n1718), .CLK(clk), .Q(mem[180]) );
  DFFPOSX1 mem_reg_5__14_ ( .D(n1717), .CLK(clk), .Q(mem[179]) );
  DFFPOSX1 mem_reg_5__13_ ( .D(n1716), .CLK(clk), .Q(mem[178]) );
  DFFPOSX1 mem_reg_5__12_ ( .D(n1715), .CLK(clk), .Q(mem[177]) );
  DFFPOSX1 mem_reg_5__11_ ( .D(n1714), .CLK(clk), .Q(mem[176]) );
  DFFPOSX1 mem_reg_5__10_ ( .D(n1713), .CLK(clk), .Q(mem[175]) );
  DFFPOSX1 mem_reg_5__9_ ( .D(n1712), .CLK(clk), .Q(mem[174]) );
  DFFPOSX1 mem_reg_5__8_ ( .D(n1711), .CLK(clk), .Q(mem[173]) );
  DFFPOSX1 mem_reg_5__7_ ( .D(n1710), .CLK(clk), .Q(mem[172]) );
  DFFPOSX1 mem_reg_5__6_ ( .D(n1709), .CLK(clk), .Q(mem[171]) );
  DFFPOSX1 mem_reg_5__5_ ( .D(n1708), .CLK(clk), .Q(mem[170]) );
  DFFPOSX1 mem_reg_5__4_ ( .D(n1707), .CLK(clk), .Q(mem[169]) );
  DFFPOSX1 mem_reg_5__3_ ( .D(n1706), .CLK(clk), .Q(mem[168]) );
  DFFPOSX1 mem_reg_5__2_ ( .D(n1705), .CLK(clk), .Q(mem[167]) );
  DFFPOSX1 mem_reg_5__1_ ( .D(n1704), .CLK(clk), .Q(mem[166]) );
  DFFPOSX1 mem_reg_5__0_ ( .D(n1703), .CLK(clk), .Q(mem[165]) );
  DFFPOSX1 mem_reg_4__32_ ( .D(n1702), .CLK(clk), .Q(mem[164]) );
  DFFPOSX1 mem_reg_4__31_ ( .D(n1701), .CLK(clk), .Q(mem[163]) );
  DFFPOSX1 mem_reg_4__30_ ( .D(n1700), .CLK(clk), .Q(mem[162]) );
  DFFPOSX1 mem_reg_4__29_ ( .D(n1699), .CLK(clk), .Q(mem[161]) );
  DFFPOSX1 mem_reg_4__28_ ( .D(n1698), .CLK(clk), .Q(mem[160]) );
  DFFPOSX1 mem_reg_4__27_ ( .D(n1697), .CLK(clk), .Q(mem[159]) );
  DFFPOSX1 mem_reg_4__26_ ( .D(n1696), .CLK(clk), .Q(mem[158]) );
  DFFPOSX1 mem_reg_4__25_ ( .D(n1695), .CLK(clk), .Q(mem[157]) );
  DFFPOSX1 mem_reg_4__24_ ( .D(n1694), .CLK(clk), .Q(mem[156]) );
  DFFPOSX1 mem_reg_4__23_ ( .D(n1693), .CLK(clk), .Q(mem[155]) );
  DFFPOSX1 mem_reg_4__22_ ( .D(n1692), .CLK(clk), .Q(mem[154]) );
  DFFPOSX1 mem_reg_4__21_ ( .D(n1691), .CLK(clk), .Q(mem[153]) );
  DFFPOSX1 mem_reg_4__20_ ( .D(n1690), .CLK(clk), .Q(mem[152]) );
  DFFPOSX1 mem_reg_4__19_ ( .D(n1689), .CLK(clk), .Q(mem[151]) );
  DFFPOSX1 mem_reg_4__18_ ( .D(n1688), .CLK(clk), .Q(mem[150]) );
  DFFPOSX1 mem_reg_4__17_ ( .D(n1687), .CLK(clk), .Q(mem[149]) );
  DFFPOSX1 mem_reg_4__16_ ( .D(n1686), .CLK(clk), .Q(mem[148]) );
  DFFPOSX1 mem_reg_4__15_ ( .D(n1685), .CLK(clk), .Q(mem[147]) );
  DFFPOSX1 mem_reg_4__14_ ( .D(n1684), .CLK(clk), .Q(mem[146]) );
  DFFPOSX1 mem_reg_4__13_ ( .D(n1683), .CLK(clk), .Q(mem[145]) );
  DFFPOSX1 mem_reg_4__12_ ( .D(n1682), .CLK(clk), .Q(mem[144]) );
  DFFPOSX1 mem_reg_4__11_ ( .D(n1681), .CLK(clk), .Q(mem[143]) );
  DFFPOSX1 mem_reg_4__10_ ( .D(n1680), .CLK(clk), .Q(mem[142]) );
  DFFPOSX1 mem_reg_4__9_ ( .D(n1679), .CLK(clk), .Q(mem[141]) );
  DFFPOSX1 mem_reg_4__8_ ( .D(n1678), .CLK(clk), .Q(mem[140]) );
  DFFPOSX1 mem_reg_4__7_ ( .D(n1677), .CLK(clk), .Q(mem[139]) );
  DFFPOSX1 mem_reg_4__6_ ( .D(n1676), .CLK(clk), .Q(mem[138]) );
  DFFPOSX1 mem_reg_4__5_ ( .D(n1675), .CLK(clk), .Q(mem[137]) );
  DFFPOSX1 mem_reg_4__4_ ( .D(n1674), .CLK(clk), .Q(mem[136]) );
  DFFPOSX1 mem_reg_4__3_ ( .D(n1673), .CLK(clk), .Q(mem[135]) );
  DFFPOSX1 mem_reg_4__2_ ( .D(n1672), .CLK(clk), .Q(mem[134]) );
  DFFPOSX1 mem_reg_4__1_ ( .D(n1671), .CLK(clk), .Q(mem[133]) );
  DFFPOSX1 mem_reg_4__0_ ( .D(n1670), .CLK(clk), .Q(mem[132]) );
  DFFPOSX1 mem_reg_3__32_ ( .D(n1669), .CLK(clk), .Q(mem[131]) );
  DFFPOSX1 mem_reg_3__31_ ( .D(n1668), .CLK(clk), .Q(mem[130]) );
  DFFPOSX1 mem_reg_3__30_ ( .D(n1667), .CLK(clk), .Q(mem[129]) );
  DFFPOSX1 mem_reg_3__29_ ( .D(n1666), .CLK(clk), .Q(mem[128]) );
  DFFPOSX1 mem_reg_3__28_ ( .D(n1665), .CLK(clk), .Q(mem[127]) );
  DFFPOSX1 mem_reg_3__27_ ( .D(n1664), .CLK(clk), .Q(mem[126]) );
  DFFPOSX1 mem_reg_3__26_ ( .D(n1663), .CLK(clk), .Q(mem[125]) );
  DFFPOSX1 mem_reg_3__25_ ( .D(n1662), .CLK(clk), .Q(mem[124]) );
  DFFPOSX1 mem_reg_3__24_ ( .D(n1661), .CLK(clk), .Q(mem[123]) );
  DFFPOSX1 mem_reg_3__23_ ( .D(n1660), .CLK(clk), .Q(mem[122]) );
  DFFPOSX1 mem_reg_3__22_ ( .D(n1659), .CLK(clk), .Q(mem[121]) );
  DFFPOSX1 mem_reg_3__21_ ( .D(n1658), .CLK(clk), .Q(mem[120]) );
  DFFPOSX1 mem_reg_3__20_ ( .D(n1657), .CLK(clk), .Q(mem[119]) );
  DFFPOSX1 mem_reg_3__19_ ( .D(n1656), .CLK(clk), .Q(mem[118]) );
  DFFPOSX1 mem_reg_3__18_ ( .D(n1655), .CLK(clk), .Q(mem[117]) );
  DFFPOSX1 mem_reg_3__17_ ( .D(n1654), .CLK(clk), .Q(mem[116]) );
  DFFPOSX1 mem_reg_3__16_ ( .D(n1653), .CLK(clk), .Q(mem[115]) );
  DFFPOSX1 mem_reg_3__15_ ( .D(n1652), .CLK(clk), .Q(mem[114]) );
  DFFPOSX1 mem_reg_3__14_ ( .D(n1651), .CLK(clk), .Q(mem[113]) );
  DFFPOSX1 mem_reg_3__13_ ( .D(n1650), .CLK(clk), .Q(mem[112]) );
  DFFPOSX1 mem_reg_3__12_ ( .D(n1649), .CLK(clk), .Q(mem[111]) );
  DFFPOSX1 mem_reg_3__11_ ( .D(n1648), .CLK(clk), .Q(mem[110]) );
  DFFPOSX1 mem_reg_3__10_ ( .D(n1647), .CLK(clk), .Q(mem[109]) );
  DFFPOSX1 mem_reg_3__9_ ( .D(n1646), .CLK(clk), .Q(mem[108]) );
  DFFPOSX1 mem_reg_3__8_ ( .D(n1645), .CLK(clk), .Q(mem[107]) );
  DFFPOSX1 mem_reg_3__7_ ( .D(n1644), .CLK(clk), .Q(mem[106]) );
  DFFPOSX1 mem_reg_3__6_ ( .D(n1643), .CLK(clk), .Q(mem[105]) );
  DFFPOSX1 mem_reg_3__5_ ( .D(n1642), .CLK(clk), .Q(mem[104]) );
  DFFPOSX1 mem_reg_3__4_ ( .D(n1641), .CLK(clk), .Q(mem[103]) );
  DFFPOSX1 mem_reg_3__3_ ( .D(n1640), .CLK(clk), .Q(mem[102]) );
  DFFPOSX1 mem_reg_3__2_ ( .D(n1639), .CLK(clk), .Q(mem[101]) );
  DFFPOSX1 mem_reg_3__1_ ( .D(n1638), .CLK(clk), .Q(mem[100]) );
  DFFPOSX1 mem_reg_3__0_ ( .D(n1637), .CLK(clk), .Q(mem[99]) );
  DFFPOSX1 mem_reg_2__32_ ( .D(n1636), .CLK(clk), .Q(mem[98]) );
  DFFPOSX1 mem_reg_2__31_ ( .D(n1635), .CLK(clk), .Q(mem[97]) );
  DFFPOSX1 mem_reg_2__30_ ( .D(n1634), .CLK(clk), .Q(mem[96]) );
  DFFPOSX1 mem_reg_2__29_ ( .D(n1633), .CLK(clk), .Q(mem[95]) );
  DFFPOSX1 mem_reg_2__28_ ( .D(n1632), .CLK(clk), .Q(mem[94]) );
  DFFPOSX1 mem_reg_2__27_ ( .D(n1631), .CLK(clk), .Q(mem[93]) );
  DFFPOSX1 mem_reg_2__26_ ( .D(n1630), .CLK(clk), .Q(mem[92]) );
  DFFPOSX1 mem_reg_2__25_ ( .D(n1629), .CLK(clk), .Q(mem[91]) );
  DFFPOSX1 mem_reg_2__24_ ( .D(n1628), .CLK(clk), .Q(mem[90]) );
  DFFPOSX1 mem_reg_2__23_ ( .D(n1627), .CLK(clk), .Q(mem[89]) );
  DFFPOSX1 mem_reg_2__22_ ( .D(n1626), .CLK(clk), .Q(mem[88]) );
  DFFPOSX1 mem_reg_2__21_ ( .D(n1625), .CLK(clk), .Q(mem[87]) );
  DFFPOSX1 mem_reg_2__20_ ( .D(n1624), .CLK(clk), .Q(mem[86]) );
  DFFPOSX1 mem_reg_2__19_ ( .D(n1623), .CLK(clk), .Q(mem[85]) );
  DFFPOSX1 mem_reg_2__18_ ( .D(n1622), .CLK(clk), .Q(mem[84]) );
  DFFPOSX1 mem_reg_2__17_ ( .D(n1621), .CLK(clk), .Q(mem[83]) );
  DFFPOSX1 mem_reg_2__16_ ( .D(n1620), .CLK(clk), .Q(mem[82]) );
  DFFPOSX1 mem_reg_2__15_ ( .D(n1619), .CLK(clk), .Q(mem[81]) );
  DFFPOSX1 mem_reg_2__14_ ( .D(n1618), .CLK(clk), .Q(mem[80]) );
  DFFPOSX1 mem_reg_2__13_ ( .D(n1617), .CLK(clk), .Q(mem[79]) );
  DFFPOSX1 mem_reg_2__12_ ( .D(n1616), .CLK(clk), .Q(mem[78]) );
  DFFPOSX1 mem_reg_2__11_ ( .D(n1615), .CLK(clk), .Q(mem[77]) );
  DFFPOSX1 mem_reg_2__10_ ( .D(n1614), .CLK(clk), .Q(mem[76]) );
  DFFPOSX1 mem_reg_2__9_ ( .D(n1613), .CLK(clk), .Q(mem[75]) );
  DFFPOSX1 mem_reg_2__8_ ( .D(n1612), .CLK(clk), .Q(mem[74]) );
  DFFPOSX1 mem_reg_2__7_ ( .D(n1611), .CLK(clk), .Q(mem[73]) );
  DFFPOSX1 mem_reg_2__6_ ( .D(n1610), .CLK(clk), .Q(mem[72]) );
  DFFPOSX1 mem_reg_2__5_ ( .D(n1609), .CLK(clk), .Q(mem[71]) );
  DFFPOSX1 mem_reg_2__4_ ( .D(n1608), .CLK(clk), .Q(mem[70]) );
  DFFPOSX1 mem_reg_2__3_ ( .D(n1607), .CLK(clk), .Q(mem[69]) );
  DFFPOSX1 mem_reg_2__2_ ( .D(n1606), .CLK(clk), .Q(mem[68]) );
  DFFPOSX1 mem_reg_2__1_ ( .D(n1605), .CLK(clk), .Q(mem[67]) );
  DFFPOSX1 mem_reg_2__0_ ( .D(n1604), .CLK(clk), .Q(mem[66]) );
  DFFPOSX1 mem_reg_1__32_ ( .D(n1603), .CLK(clk), .Q(mem[65]) );
  DFFPOSX1 mem_reg_1__31_ ( .D(n1602), .CLK(clk), .Q(mem[64]) );
  DFFPOSX1 mem_reg_1__30_ ( .D(n1601), .CLK(clk), .Q(mem[63]) );
  DFFPOSX1 mem_reg_1__29_ ( .D(n1600), .CLK(clk), .Q(mem[62]) );
  DFFPOSX1 mem_reg_1__28_ ( .D(n1599), .CLK(clk), .Q(mem[61]) );
  DFFPOSX1 mem_reg_1__27_ ( .D(n1598), .CLK(clk), .Q(mem[60]) );
  DFFPOSX1 mem_reg_1__26_ ( .D(n1597), .CLK(clk), .Q(mem[59]) );
  DFFPOSX1 mem_reg_1__25_ ( .D(n1596), .CLK(clk), .Q(mem[58]) );
  DFFPOSX1 mem_reg_1__24_ ( .D(n1595), .CLK(clk), .Q(mem[57]) );
  DFFPOSX1 mem_reg_1__23_ ( .D(n1594), .CLK(clk), .Q(mem[56]) );
  DFFPOSX1 mem_reg_1__22_ ( .D(n1593), .CLK(clk), .Q(mem[55]) );
  DFFPOSX1 mem_reg_1__21_ ( .D(n1592), .CLK(clk), .Q(mem[54]) );
  DFFPOSX1 mem_reg_1__20_ ( .D(n1591), .CLK(clk), .Q(mem[53]) );
  DFFPOSX1 mem_reg_1__19_ ( .D(n1590), .CLK(clk), .Q(mem[52]) );
  DFFPOSX1 mem_reg_1__18_ ( .D(n1589), .CLK(clk), .Q(mem[51]) );
  DFFPOSX1 mem_reg_1__17_ ( .D(n1588), .CLK(clk), .Q(mem[50]) );
  DFFPOSX1 mem_reg_1__16_ ( .D(n1587), .CLK(clk), .Q(mem[49]) );
  DFFPOSX1 mem_reg_1__15_ ( .D(n1586), .CLK(clk), .Q(mem[48]) );
  DFFPOSX1 mem_reg_1__14_ ( .D(n1585), .CLK(clk), .Q(mem[47]) );
  DFFPOSX1 mem_reg_1__13_ ( .D(n1584), .CLK(clk), .Q(mem[46]) );
  DFFPOSX1 mem_reg_1__12_ ( .D(n1583), .CLK(clk), .Q(mem[45]) );
  DFFPOSX1 mem_reg_1__11_ ( .D(n1582), .CLK(clk), .Q(mem[44]) );
  DFFPOSX1 mem_reg_1__10_ ( .D(n1581), .CLK(clk), .Q(mem[43]) );
  DFFPOSX1 mem_reg_1__9_ ( .D(n1580), .CLK(clk), .Q(mem[42]) );
  DFFPOSX1 mem_reg_1__8_ ( .D(n1579), .CLK(clk), .Q(mem[41]) );
  DFFPOSX1 mem_reg_1__7_ ( .D(n1578), .CLK(clk), .Q(mem[40]) );
  DFFPOSX1 mem_reg_1__6_ ( .D(n1577), .CLK(clk), .Q(mem[39]) );
  DFFPOSX1 mem_reg_1__5_ ( .D(n1576), .CLK(clk), .Q(mem[38]) );
  DFFPOSX1 mem_reg_1__4_ ( .D(n1575), .CLK(clk), .Q(mem[37]) );
  DFFPOSX1 mem_reg_1__3_ ( .D(n1574), .CLK(clk), .Q(mem[36]) );
  DFFPOSX1 mem_reg_1__2_ ( .D(n1573), .CLK(clk), .Q(mem[35]) );
  DFFPOSX1 mem_reg_1__1_ ( .D(n1572), .CLK(clk), .Q(mem[34]) );
  DFFPOSX1 mem_reg_1__0_ ( .D(n1571), .CLK(clk), .Q(mem[33]) );
  DFFPOSX1 mem_reg_0__32_ ( .D(n1570), .CLK(clk), .Q(mem[32]) );
  DFFPOSX1 mem_reg_0__31_ ( .D(n1569), .CLK(clk), .Q(mem[31]) );
  DFFPOSX1 mem_reg_0__30_ ( .D(n1568), .CLK(clk), .Q(mem[30]) );
  DFFPOSX1 mem_reg_0__29_ ( .D(n1567), .CLK(clk), .Q(mem[29]) );
  DFFPOSX1 mem_reg_0__28_ ( .D(n1566), .CLK(clk), .Q(mem[28]) );
  DFFPOSX1 mem_reg_0__27_ ( .D(n1565), .CLK(clk), .Q(mem[27]) );
  DFFPOSX1 mem_reg_0__26_ ( .D(n1564), .CLK(clk), .Q(mem[26]) );
  DFFPOSX1 mem_reg_0__25_ ( .D(n1563), .CLK(clk), .Q(mem[25]) );
  DFFPOSX1 mem_reg_0__24_ ( .D(n1562), .CLK(clk), .Q(mem[24]) );
  DFFPOSX1 mem_reg_0__23_ ( .D(n1561), .CLK(clk), .Q(mem[23]) );
  DFFPOSX1 mem_reg_0__22_ ( .D(n1560), .CLK(clk), .Q(mem[22]) );
  DFFPOSX1 mem_reg_0__21_ ( .D(n1559), .CLK(clk), .Q(mem[21]) );
  DFFPOSX1 mem_reg_0__20_ ( .D(n1558), .CLK(clk), .Q(mem[20]) );
  DFFPOSX1 mem_reg_0__19_ ( .D(n1557), .CLK(clk), .Q(mem[19]) );
  DFFPOSX1 mem_reg_0__18_ ( .D(n1556), .CLK(clk), .Q(mem[18]) );
  DFFPOSX1 mem_reg_0__17_ ( .D(n1555), .CLK(clk), .Q(mem[17]) );
  DFFPOSX1 mem_reg_0__16_ ( .D(n1554), .CLK(clk), .Q(mem[16]) );
  DFFPOSX1 mem_reg_0__15_ ( .D(n1553), .CLK(clk), .Q(mem[15]) );
  DFFPOSX1 mem_reg_0__14_ ( .D(n1552), .CLK(clk), .Q(mem[14]) );
  DFFPOSX1 mem_reg_0__13_ ( .D(n1551), .CLK(clk), .Q(mem[13]) );
  DFFPOSX1 mem_reg_0__12_ ( .D(n1550), .CLK(clk), .Q(mem[12]) );
  DFFPOSX1 mem_reg_0__11_ ( .D(n1549), .CLK(clk), .Q(mem[11]) );
  DFFPOSX1 mem_reg_0__10_ ( .D(n1548), .CLK(clk), .Q(mem[10]) );
  DFFPOSX1 mem_reg_0__9_ ( .D(n1547), .CLK(clk), .Q(mem[9]) );
  DFFPOSX1 mem_reg_0__8_ ( .D(n1546), .CLK(clk), .Q(mem[8]) );
  DFFPOSX1 mem_reg_0__7_ ( .D(n1545), .CLK(clk), .Q(mem[7]) );
  DFFPOSX1 mem_reg_0__6_ ( .D(n1544), .CLK(clk), .Q(mem[6]) );
  DFFPOSX1 mem_reg_0__5_ ( .D(n1543), .CLK(clk), .Q(mem[5]) );
  DFFPOSX1 mem_reg_0__4_ ( .D(n1542), .CLK(clk), .Q(mem[4]) );
  DFFPOSX1 mem_reg_0__3_ ( .D(n1541), .CLK(clk), .Q(mem[3]) );
  DFFPOSX1 mem_reg_0__2_ ( .D(n1540), .CLK(clk), .Q(mem[2]) );
  DFFPOSX1 mem_reg_0__1_ ( .D(n1539), .CLK(clk), .Q(mem[1]) );
  DFFPOSX1 mem_reg_0__0_ ( .D(n1538), .CLK(clk), .Q(mem[0]) );
  OAI21X1 U83 ( .A(n4548), .B(n4581), .C(n3383), .Y(n1538) );
  OAI21X1 U85 ( .A(n4548), .B(n4580), .C(n3317), .Y(n1539) );
  OAI21X1 U87 ( .A(n4548), .B(n4579), .C(n3251), .Y(n1540) );
  OAI21X1 U89 ( .A(n4548), .B(n4578), .C(n3184), .Y(n1541) );
  OAI21X1 U91 ( .A(n4548), .B(n4577), .C(n3183), .Y(n1542) );
  OAI21X1 U93 ( .A(n4548), .B(n4576), .C(n3382), .Y(n1543) );
  OAI21X1 U95 ( .A(n4548), .B(n4575), .C(n3316), .Y(n1544) );
  OAI21X1 U97 ( .A(n4548), .B(n4574), .C(n3113), .Y(n1545) );
  OAI21X1 U99 ( .A(n4548), .B(n4573), .C(n3250), .Y(n1546) );
  OAI21X1 U101 ( .A(n4548), .B(n4572), .C(n3046), .Y(n1547) );
  OAI21X1 U103 ( .A(n4548), .B(n4571), .C(n2978), .Y(n1548) );
  OAI21X1 U105 ( .A(n4548), .B(n4570), .C(n2911), .Y(n1549) );
  OAI21X1 U107 ( .A(n4548), .B(n4569), .C(n2847), .Y(n1550) );
  OAI21X1 U109 ( .A(n4548), .B(n4568), .C(n2782), .Y(n1551) );
  OAI21X1 U111 ( .A(n4548), .B(n4567), .C(n2718), .Y(n1552) );
  OAI21X1 U113 ( .A(n4548), .B(n4566), .C(n2654), .Y(n1553) );
  OAI21X1 U115 ( .A(n4548), .B(n4565), .C(n386), .Y(n1554) );
  OAI21X1 U117 ( .A(n4548), .B(n4564), .C(n303), .Y(n1555) );
  OAI21X1 U119 ( .A(n4548), .B(n4563), .C(n239), .Y(n1556) );
  OAI21X1 U121 ( .A(n4548), .B(n4562), .C(n175), .Y(n1557) );
  OAI21X1 U123 ( .A(n4548), .B(n4561), .C(n3112), .Y(n1558) );
  OAI21X1 U125 ( .A(n4548), .B(n4560), .C(n3045), .Y(n1559) );
  OAI21X1 U127 ( .A(n4548), .B(n4559), .C(n2977), .Y(n1560) );
  OAI21X1 U129 ( .A(n4548), .B(n4558), .C(n2910), .Y(n1561) );
  OAI21X1 U131 ( .A(n4548), .B(n4557), .C(n2846), .Y(n1562) );
  OAI21X1 U133 ( .A(n4548), .B(n4556), .C(n2781), .Y(n1563) );
  OAI21X1 U135 ( .A(n4548), .B(n4555), .C(n2717), .Y(n1564) );
  OAI21X1 U137 ( .A(n4548), .B(n4554), .C(n2653), .Y(n1565) );
  OAI21X1 U139 ( .A(n4548), .B(n4553), .C(n384), .Y(n1566) );
  OAI21X1 U141 ( .A(n4548), .B(n4552), .C(n302), .Y(n1567) );
  OAI21X1 U143 ( .A(n4548), .B(n4551), .C(n238), .Y(n1568) );
  OAI21X1 U145 ( .A(n4548), .B(n4550), .C(n174), .Y(n1569) );
  OAI21X1 U147 ( .A(n4548), .B(n4549), .C(n111), .Y(n1570) );
  OAI21X1 U149 ( .A(n3185), .B(n3118), .C(reset), .Y(n414) );
  OAI21X1 U150 ( .A(n4547), .B(n4581), .C(n3315), .Y(n1571) );
  OAI21X1 U152 ( .A(n4547), .B(n4580), .C(n3381), .Y(n1572) );
  OAI21X1 U154 ( .A(n4547), .B(n4579), .C(n3182), .Y(n1573) );
  OAI21X1 U156 ( .A(n4547), .B(n4578), .C(n3249), .Y(n1574) );
  OAI21X1 U158 ( .A(n4547), .B(n4577), .C(n3248), .Y(n1575) );
  OAI21X1 U160 ( .A(n4547), .B(n4576), .C(n3314), .Y(n1576) );
  OAI21X1 U162 ( .A(n4547), .B(n4575), .C(n3380), .Y(n1577) );
  OAI21X1 U164 ( .A(n4547), .B(n4574), .C(n3044), .Y(n1578) );
  OAI21X1 U166 ( .A(n4547), .B(n4573), .C(n3181), .Y(n1579) );
  OAI21X1 U168 ( .A(n4547), .B(n4572), .C(n3111), .Y(n1580) );
  OAI21X1 U170 ( .A(n4547), .B(n4571), .C(n2909), .Y(n1581) );
  OAI21X1 U172 ( .A(n4547), .B(n4570), .C(n2976), .Y(n1582) );
  OAI21X1 U174 ( .A(n4547), .B(n4569), .C(n2780), .Y(n1583) );
  OAI21X1 U176 ( .A(n4547), .B(n4568), .C(n2845), .Y(n1584) );
  OAI21X1 U178 ( .A(n4547), .B(n4567), .C(n2652), .Y(n1585) );
  OAI21X1 U180 ( .A(n4547), .B(n4566), .C(n2716), .Y(n1586) );
  OAI21X1 U182 ( .A(n4547), .B(n4565), .C(n301), .Y(n1587) );
  OAI21X1 U184 ( .A(n4547), .B(n4564), .C(n382), .Y(n1588) );
  OAI21X1 U186 ( .A(n4547), .B(n4563), .C(n173), .Y(n1589) );
  OAI21X1 U188 ( .A(n4547), .B(n4562), .C(n237), .Y(n1590) );
  OAI21X1 U190 ( .A(n4547), .B(n4561), .C(n3043), .Y(n1591) );
  OAI21X1 U192 ( .A(n4547), .B(n4560), .C(n3110), .Y(n1592) );
  OAI21X1 U194 ( .A(n4547), .B(n4559), .C(n2908), .Y(n1593) );
  OAI21X1 U196 ( .A(n4547), .B(n4558), .C(n2975), .Y(n1594) );
  OAI21X1 U198 ( .A(n4547), .B(n4557), .C(n2779), .Y(n1595) );
  OAI21X1 U200 ( .A(n4547), .B(n4556), .C(n2844), .Y(n1596) );
  OAI21X1 U202 ( .A(n4547), .B(n4555), .C(n2651), .Y(n1597) );
  OAI21X1 U204 ( .A(n4547), .B(n4554), .C(n2715), .Y(n1598) );
  OAI21X1 U206 ( .A(n4547), .B(n4553), .C(n300), .Y(n1599) );
  OAI21X1 U208 ( .A(n4547), .B(n4552), .C(n380), .Y(n1600) );
  OAI21X1 U210 ( .A(n4547), .B(n4551), .C(n172), .Y(n1601) );
  OAI21X1 U212 ( .A(n4547), .B(n4550), .C(n236), .Y(n1602) );
  OAI21X1 U214 ( .A(n4547), .B(n4549), .C(n110), .Y(n1603) );
  OAI21X1 U216 ( .A(n3185), .B(n3048), .C(reset), .Y(n450) );
  OAI21X1 U217 ( .A(n4546), .B(n4581), .C(n3247), .Y(n1604) );
  OAI21X1 U219 ( .A(n4546), .B(n4580), .C(n3180), .Y(n1605) );
  OAI21X1 U221 ( .A(n4546), .B(n4579), .C(n3379), .Y(n1606) );
  OAI21X1 U223 ( .A(n4546), .B(n4578), .C(n3313), .Y(n1607) );
  OAI21X1 U225 ( .A(n4546), .B(n4577), .C(n3312), .Y(n1608) );
  OAI21X1 U227 ( .A(n4546), .B(n4576), .C(n3246), .Y(n1609) );
  OAI21X1 U229 ( .A(n4546), .B(n4575), .C(n3179), .Y(n1610) );
  OAI21X1 U231 ( .A(n4546), .B(n4574), .C(n2974), .Y(n1611) );
  OAI21X1 U233 ( .A(n4546), .B(n4573), .C(n3378), .Y(n1612) );
  OAI21X1 U235 ( .A(n4546), .B(n4572), .C(n2907), .Y(n1613) );
  OAI21X1 U237 ( .A(n4546), .B(n4571), .C(n3109), .Y(n1614) );
  OAI21X1 U239 ( .A(n4546), .B(n4570), .C(n3042), .Y(n1615) );
  OAI21X1 U241 ( .A(n4546), .B(n4569), .C(n2714), .Y(n1616) );
  OAI21X1 U243 ( .A(n4546), .B(n4568), .C(n2650), .Y(n1617) );
  OAI21X1 U245 ( .A(n4546), .B(n4567), .C(n2843), .Y(n1618) );
  OAI21X1 U247 ( .A(n4546), .B(n4566), .C(n2778), .Y(n1619) );
  OAI21X1 U249 ( .A(n4546), .B(n4565), .C(n235), .Y(n1620) );
  OAI21X1 U251 ( .A(n4546), .B(n4564), .C(n171), .Y(n1621) );
  OAI21X1 U253 ( .A(n4546), .B(n4563), .C(n378), .Y(n1622) );
  OAI21X1 U255 ( .A(n4546), .B(n4562), .C(n299), .Y(n1623) );
  OAI21X1 U257 ( .A(n4546), .B(n4561), .C(n2973), .Y(n1624) );
  OAI21X1 U259 ( .A(n4546), .B(n4560), .C(n2906), .Y(n1625) );
  OAI21X1 U261 ( .A(n4546), .B(n4559), .C(n3108), .Y(n1626) );
  OAI21X1 U263 ( .A(n4546), .B(n4558), .C(n3041), .Y(n1627) );
  OAI21X1 U265 ( .A(n4546), .B(n4557), .C(n2713), .Y(n1628) );
  OAI21X1 U267 ( .A(n4546), .B(n4556), .C(n2649), .Y(n1629) );
  OAI21X1 U269 ( .A(n4546), .B(n4555), .C(n2842), .Y(n1630) );
  OAI21X1 U271 ( .A(n4546), .B(n4554), .C(n2777), .Y(n1631) );
  OAI21X1 U273 ( .A(n4546), .B(n4553), .C(n234), .Y(n1632) );
  OAI21X1 U275 ( .A(n4546), .B(n4552), .C(n170), .Y(n1633) );
  OAI21X1 U277 ( .A(n4546), .B(n4551), .C(n376), .Y(n1634) );
  OAI21X1 U279 ( .A(n4546), .B(n4550), .C(n298), .Y(n1635) );
  OAI21X1 U281 ( .A(n4546), .B(n4549), .C(n109), .Y(n1636) );
  OAI21X1 U283 ( .A(n3185), .B(n2980), .C(reset), .Y(n485) );
  OAI21X1 U284 ( .A(n4545), .B(n4581), .C(n3178), .Y(n1637) );
  OAI21X1 U286 ( .A(n4545), .B(n4580), .C(n3245), .Y(n1638) );
  OAI21X1 U288 ( .A(n4545), .B(n4579), .C(n3311), .Y(n1639) );
  OAI21X1 U290 ( .A(n4545), .B(n4578), .C(n3377), .Y(n1640) );
  OAI21X1 U292 ( .A(n4545), .B(n4577), .C(n3376), .Y(n1641) );
  OAI21X1 U294 ( .A(n4545), .B(n4576), .C(n3177), .Y(n1642) );
  OAI21X1 U296 ( .A(n4545), .B(n4575), .C(n3244), .Y(n1643) );
  OAI21X1 U298 ( .A(n4545), .B(n4574), .C(n2905), .Y(n1644) );
  OAI21X1 U300 ( .A(n4545), .B(n4573), .C(n3310), .Y(n1645) );
  OAI21X1 U302 ( .A(n4545), .B(n4572), .C(n2972), .Y(n1646) );
  OAI21X1 U304 ( .A(n4545), .B(n4571), .C(n3040), .Y(n1647) );
  OAI21X1 U306 ( .A(n4545), .B(n4570), .C(n3107), .Y(n1648) );
  OAI21X1 U308 ( .A(n4545), .B(n4569), .C(n2648), .Y(n1649) );
  OAI21X1 U310 ( .A(n4545), .B(n4568), .C(n2712), .Y(n1650) );
  OAI21X1 U312 ( .A(n4545), .B(n4567), .C(n2776), .Y(n1651) );
  OAI21X1 U314 ( .A(n4545), .B(n4566), .C(n2841), .Y(n1652) );
  OAI21X1 U316 ( .A(n4545), .B(n4565), .C(n169), .Y(n1653) );
  OAI21X1 U318 ( .A(n4545), .B(n4564), .C(n233), .Y(n1654) );
  OAI21X1 U320 ( .A(n4545), .B(n4563), .C(n297), .Y(n1655) );
  OAI21X1 U322 ( .A(n4545), .B(n4562), .C(n374), .Y(n1656) );
  OAI21X1 U324 ( .A(n4545), .B(n4561), .C(n2904), .Y(n1657) );
  OAI21X1 U326 ( .A(n4545), .B(n4560), .C(n2971), .Y(n1658) );
  OAI21X1 U328 ( .A(n4545), .B(n4559), .C(n3039), .Y(n1659) );
  OAI21X1 U330 ( .A(n4545), .B(n4558), .C(n3106), .Y(n1660) );
  OAI21X1 U332 ( .A(n4545), .B(n4557), .C(n2647), .Y(n1661) );
  OAI21X1 U334 ( .A(n4545), .B(n4556), .C(n2711), .Y(n1662) );
  OAI21X1 U336 ( .A(n4545), .B(n4555), .C(n2775), .Y(n1663) );
  OAI21X1 U338 ( .A(n4545), .B(n4554), .C(n2840), .Y(n1664) );
  OAI21X1 U340 ( .A(n4545), .B(n4553), .C(n168), .Y(n1665) );
  OAI21X1 U342 ( .A(n4545), .B(n4552), .C(n232), .Y(n1666) );
  OAI21X1 U344 ( .A(n4545), .B(n4551), .C(n296), .Y(n1667) );
  OAI21X1 U346 ( .A(n4545), .B(n4550), .C(n372), .Y(n1668) );
  OAI21X1 U348 ( .A(n4545), .B(n4549), .C(n108), .Y(n1669) );
  OAI21X1 U350 ( .A(n3185), .B(n2913), .C(reset), .Y(n520) );
  OAI21X1 U351 ( .A(n4544), .B(n4581), .C(n3105), .Y(n1670) );
  OAI21X1 U353 ( .A(n4544), .B(n4580), .C(n3038), .Y(n1671) );
  OAI21X1 U355 ( .A(n4544), .B(n4579), .C(n2970), .Y(n1672) );
  OAI21X1 U357 ( .A(n4544), .B(n4578), .C(n2903), .Y(n1673) );
  OAI21X1 U359 ( .A(n4544), .B(n4577), .C(n2902), .Y(n1674) );
  OAI21X1 U361 ( .A(n4544), .B(n4576), .C(n3104), .Y(n1675) );
  OAI21X1 U363 ( .A(n4544), .B(n4575), .C(n3037), .Y(n1676) );
  OAI21X1 U365 ( .A(n4544), .B(n4574), .C(n3375), .Y(n1677) );
  OAI21X1 U367 ( .A(n4544), .B(n4573), .C(n2969), .Y(n1678) );
  OAI21X1 U369 ( .A(n4544), .B(n4572), .C(n3309), .Y(n1679) );
  OAI21X1 U371 ( .A(n4544), .B(n4571), .C(n3243), .Y(n1680) );
  OAI21X1 U373 ( .A(n4544), .B(n4570), .C(n3176), .Y(n1681) );
  OAI21X1 U375 ( .A(n4544), .B(n4569), .C(n370), .Y(n1682) );
  OAI21X1 U377 ( .A(n4544), .B(n4568), .C(n295), .Y(n1683) );
  OAI21X1 U379 ( .A(n4544), .B(n4567), .C(n231), .Y(n1684) );
  OAI21X1 U381 ( .A(n4544), .B(n4566), .C(n167), .Y(n1685) );
  OAI21X1 U383 ( .A(n4544), .B(n4565), .C(n2839), .Y(n1686) );
  OAI21X1 U385 ( .A(n4544), .B(n4564), .C(n2774), .Y(n1687) );
  OAI21X1 U387 ( .A(n4544), .B(n4563), .C(n2710), .Y(n1688) );
  OAI21X1 U389 ( .A(n4544), .B(n4562), .C(n2646), .Y(n1689) );
  OAI21X1 U391 ( .A(n4544), .B(n4561), .C(n3374), .Y(n1690) );
  OAI21X1 U393 ( .A(n4544), .B(n4560), .C(n3308), .Y(n1691) );
  OAI21X1 U395 ( .A(n4544), .B(n4559), .C(n3242), .Y(n1692) );
  OAI21X1 U397 ( .A(n4544), .B(n4558), .C(n3175), .Y(n1693) );
  OAI21X1 U399 ( .A(n4544), .B(n4557), .C(n368), .Y(n1694) );
  OAI21X1 U401 ( .A(n4544), .B(n4556), .C(n294), .Y(n1695) );
  OAI21X1 U403 ( .A(n4544), .B(n4555), .C(n230), .Y(n1696) );
  OAI21X1 U405 ( .A(n4544), .B(n4554), .C(n166), .Y(n1697) );
  OAI21X1 U407 ( .A(n4544), .B(n4553), .C(n2838), .Y(n1698) );
  OAI21X1 U409 ( .A(n4544), .B(n4552), .C(n2773), .Y(n1699) );
  OAI21X1 U411 ( .A(n4544), .B(n4551), .C(n2709), .Y(n1700) );
  OAI21X1 U413 ( .A(n4544), .B(n4550), .C(n2645), .Y(n1701) );
  OAI21X1 U415 ( .A(n4544), .B(n4549), .C(n107), .Y(n1702) );
  OAI21X1 U417 ( .A(n3185), .B(n2912), .C(reset), .Y(n555) );
  OAI21X1 U418 ( .A(n4543), .B(n4581), .C(n3036), .Y(n1703) );
  OAI21X1 U420 ( .A(n4543), .B(n4580), .C(n3103), .Y(n1704) );
  OAI21X1 U422 ( .A(n4543), .B(n4579), .C(n2901), .Y(n1705) );
  OAI21X1 U424 ( .A(n4543), .B(n4578), .C(n2968), .Y(n1706) );
  OAI21X1 U426 ( .A(n4543), .B(n4577), .C(n2967), .Y(n1707) );
  OAI21X1 U428 ( .A(n4543), .B(n4576), .C(n3035), .Y(n1708) );
  OAI21X1 U430 ( .A(n4543), .B(n4575), .C(n3102), .Y(n1709) );
  OAI21X1 U432 ( .A(n4543), .B(n4574), .C(n3307), .Y(n1710) );
  OAI21X1 U434 ( .A(n4543), .B(n4573), .C(n2900), .Y(n1711) );
  OAI21X1 U436 ( .A(n4543), .B(n4572), .C(n3373), .Y(n1712) );
  OAI21X1 U438 ( .A(n4543), .B(n4571), .C(n3174), .Y(n1713) );
  OAI21X1 U440 ( .A(n4543), .B(n4570), .C(n3241), .Y(n1714) );
  OAI21X1 U442 ( .A(n4543), .B(n4569), .C(n293), .Y(n1715) );
  OAI21X1 U444 ( .A(n4543), .B(n4568), .C(n366), .Y(n1716) );
  OAI21X1 U446 ( .A(n4543), .B(n4567), .C(n165), .Y(n1717) );
  OAI21X1 U448 ( .A(n4543), .B(n4566), .C(n229), .Y(n1718) );
  OAI21X1 U450 ( .A(n4543), .B(n4565), .C(n2772), .Y(n1719) );
  OAI21X1 U452 ( .A(n4543), .B(n4564), .C(n2837), .Y(n1720) );
  OAI21X1 U454 ( .A(n4543), .B(n4563), .C(n2644), .Y(n1721) );
  OAI21X1 U456 ( .A(n4543), .B(n4562), .C(n2708), .Y(n1722) );
  OAI21X1 U458 ( .A(n4543), .B(n4561), .C(n3306), .Y(n1723) );
  OAI21X1 U460 ( .A(n4543), .B(n4560), .C(n3372), .Y(n1724) );
  OAI21X1 U462 ( .A(n4543), .B(n4559), .C(n3173), .Y(n1725) );
  OAI21X1 U464 ( .A(n4543), .B(n4558), .C(n3240), .Y(n1726) );
  OAI21X1 U466 ( .A(n4543), .B(n4557), .C(n292), .Y(n1727) );
  OAI21X1 U468 ( .A(n4543), .B(n4556), .C(n364), .Y(n1728) );
  OAI21X1 U470 ( .A(n4543), .B(n4555), .C(n164), .Y(n1729) );
  OAI21X1 U472 ( .A(n4543), .B(n4554), .C(n228), .Y(n1730) );
  OAI21X1 U474 ( .A(n4543), .B(n4553), .C(n2771), .Y(n1731) );
  OAI21X1 U476 ( .A(n4543), .B(n4552), .C(n2836), .Y(n1732) );
  OAI21X1 U478 ( .A(n4543), .B(n4551), .C(n2643), .Y(n1733) );
  OAI21X1 U480 ( .A(n4543), .B(n4550), .C(n2707), .Y(n1734) );
  OAI21X1 U482 ( .A(n4543), .B(n4549), .C(n106), .Y(n1735) );
  OAI21X1 U484 ( .A(n3185), .B(n2979), .C(reset), .Y(n590) );
  OAI21X1 U485 ( .A(n4542), .B(n4581), .C(n2966), .Y(n1736) );
  OAI21X1 U487 ( .A(n4542), .B(n4580), .C(n2899), .Y(n1737) );
  OAI21X1 U489 ( .A(n4542), .B(n4579), .C(n3101), .Y(n1738) );
  OAI21X1 U491 ( .A(n4542), .B(n4578), .C(n3034), .Y(n1739) );
  OAI21X1 U493 ( .A(n4542), .B(n4577), .C(n3033), .Y(n1740) );
  OAI21X1 U495 ( .A(n4542), .B(n4576), .C(n2965), .Y(n1741) );
  OAI21X1 U497 ( .A(n4542), .B(n4575), .C(n2898), .Y(n1742) );
  OAI21X1 U499 ( .A(n4542), .B(n4574), .C(n3239), .Y(n1743) );
  OAI21X1 U501 ( .A(n4542), .B(n4573), .C(n3100), .Y(n1744) );
  OAI21X1 U503 ( .A(n4542), .B(n4572), .C(n3172), .Y(n1745) );
  OAI21X1 U505 ( .A(n4542), .B(n4571), .C(n3371), .Y(n1746) );
  OAI21X1 U507 ( .A(n4542), .B(n4570), .C(n3305), .Y(n1747) );
  OAI21X1 U509 ( .A(n4542), .B(n4569), .C(n227), .Y(n1748) );
  OAI21X1 U511 ( .A(n4542), .B(n4568), .C(n163), .Y(n1749) );
  OAI21X1 U513 ( .A(n4542), .B(n4567), .C(n362), .Y(n1750) );
  OAI21X1 U515 ( .A(n4542), .B(n4566), .C(n291), .Y(n1751) );
  OAI21X1 U517 ( .A(n4542), .B(n4565), .C(n2706), .Y(n1752) );
  OAI21X1 U519 ( .A(n4542), .B(n4564), .C(n2642), .Y(n1753) );
  OAI21X1 U521 ( .A(n4542), .B(n4563), .C(n2835), .Y(n1754) );
  OAI21X1 U523 ( .A(n4542), .B(n4562), .C(n2770), .Y(n1755) );
  OAI21X1 U525 ( .A(n4542), .B(n4561), .C(n3238), .Y(n1756) );
  OAI21X1 U527 ( .A(n4542), .B(n4560), .C(n3171), .Y(n1757) );
  OAI21X1 U529 ( .A(n4542), .B(n4559), .C(n3370), .Y(n1758) );
  OAI21X1 U531 ( .A(n4542), .B(n4558), .C(n3304), .Y(n1759) );
  OAI21X1 U533 ( .A(n4542), .B(n4557), .C(n226), .Y(n1760) );
  OAI21X1 U535 ( .A(n4542), .B(n4556), .C(n162), .Y(n1761) );
  OAI21X1 U537 ( .A(n4542), .B(n4555), .C(n360), .Y(n1762) );
  OAI21X1 U539 ( .A(n4542), .B(n4554), .C(n290), .Y(n1763) );
  OAI21X1 U541 ( .A(n4542), .B(n4553), .C(n2705), .Y(n1764) );
  OAI21X1 U543 ( .A(n4542), .B(n4552), .C(n2641), .Y(n1765) );
  OAI21X1 U545 ( .A(n4542), .B(n4551), .C(n2834), .Y(n1766) );
  OAI21X1 U547 ( .A(n4542), .B(n4550), .C(n2769), .Y(n1767) );
  OAI21X1 U549 ( .A(n4542), .B(n4549), .C(n105), .Y(n1768) );
  OAI21X1 U551 ( .A(n3185), .B(n3047), .C(reset), .Y(n625) );
  OAI21X1 U552 ( .A(n4541), .B(n4581), .C(n2897), .Y(n1769) );
  OAI21X1 U554 ( .A(n4541), .B(n4580), .C(n2964), .Y(n1770) );
  OAI21X1 U556 ( .A(n4541), .B(n4579), .C(n3032), .Y(n1771) );
  OAI21X1 U558 ( .A(n4541), .B(n4578), .C(n3099), .Y(n1772) );
  OAI21X1 U560 ( .A(n4541), .B(n4577), .C(n3098), .Y(n1773) );
  OAI21X1 U562 ( .A(n4541), .B(n4576), .C(n2896), .Y(n1774) );
  OAI21X1 U564 ( .A(n4541), .B(n4575), .C(n2963), .Y(n1775) );
  OAI21X1 U566 ( .A(n4541), .B(n4574), .C(n3170), .Y(n1776) );
  OAI21X1 U568 ( .A(n4541), .B(n4573), .C(n3031), .Y(n1777) );
  OAI21X1 U570 ( .A(n4541), .B(n4572), .C(n3237), .Y(n1778) );
  OAI21X1 U572 ( .A(n4541), .B(n4571), .C(n3303), .Y(n1779) );
  OAI21X1 U574 ( .A(n4541), .B(n4570), .C(n3369), .Y(n1780) );
  OAI21X1 U576 ( .A(n4541), .B(n4569), .C(n161), .Y(n1781) );
  OAI21X1 U578 ( .A(n4541), .B(n4568), .C(n225), .Y(n1782) );
  OAI21X1 U580 ( .A(n4541), .B(n4567), .C(n289), .Y(n1783) );
  OAI21X1 U582 ( .A(n4541), .B(n4566), .C(n358), .Y(n1784) );
  OAI21X1 U584 ( .A(n4541), .B(n4565), .C(n2640), .Y(n1785) );
  OAI21X1 U586 ( .A(n4541), .B(n4564), .C(n2704), .Y(n1786) );
  OAI21X1 U588 ( .A(n4541), .B(n4563), .C(n2768), .Y(n1787) );
  OAI21X1 U590 ( .A(n4541), .B(n4562), .C(n2833), .Y(n1788) );
  OAI21X1 U592 ( .A(n4541), .B(n4561), .C(n3169), .Y(n1789) );
  OAI21X1 U594 ( .A(n4541), .B(n4560), .C(n3236), .Y(n1790) );
  OAI21X1 U596 ( .A(n4541), .B(n4559), .C(n3302), .Y(n1791) );
  OAI21X1 U598 ( .A(n4541), .B(n4558), .C(n3368), .Y(n1792) );
  OAI21X1 U600 ( .A(n4541), .B(n4557), .C(n160), .Y(n1793) );
  OAI21X1 U602 ( .A(n4541), .B(n4556), .C(n224), .Y(n1794) );
  OAI21X1 U604 ( .A(n4541), .B(n4555), .C(n288), .Y(n1795) );
  OAI21X1 U606 ( .A(n4541), .B(n4554), .C(n356), .Y(n1796) );
  OAI21X1 U608 ( .A(n4541), .B(n4553), .C(n2639), .Y(n1797) );
  OAI21X1 U610 ( .A(n4541), .B(n4552), .C(n2703), .Y(n1798) );
  OAI21X1 U612 ( .A(n4541), .B(n4551), .C(n2767), .Y(n1799) );
  OAI21X1 U614 ( .A(n4541), .B(n4550), .C(n2832), .Y(n1800) );
  OAI21X1 U616 ( .A(n4541), .B(n4549), .C(n104), .Y(n1801) );
  OAI21X1 U618 ( .A(n3185), .B(n3117), .C(reset), .Y(n660) );
  NAND3X1 U619 ( .A(n4623), .B(n4620), .C(n1481), .Y(n415) );
  OAI21X1 U620 ( .A(n4540), .B(n4581), .C(n3367), .Y(n1802) );
  OAI21X1 U622 ( .A(n4540), .B(n4580), .C(n3301), .Y(n1803) );
  OAI21X1 U624 ( .A(n4540), .B(n4579), .C(n3235), .Y(n1804) );
  OAI21X1 U626 ( .A(n4540), .B(n4578), .C(n3168), .Y(n1805) );
  OAI21X1 U628 ( .A(n4540), .B(n4577), .C(n3167), .Y(n1806) );
  OAI21X1 U630 ( .A(n4540), .B(n4576), .C(n3366), .Y(n1807) );
  OAI21X1 U632 ( .A(n4540), .B(n4575), .C(n3300), .Y(n1808) );
  OAI21X1 U634 ( .A(n4540), .B(n4574), .C(n3097), .Y(n1809) );
  OAI21X1 U636 ( .A(n4540), .B(n4573), .C(n3234), .Y(n1810) );
  OAI21X1 U638 ( .A(n4540), .B(n4572), .C(n3030), .Y(n1811) );
  OAI21X1 U640 ( .A(n4540), .B(n4571), .C(n2962), .Y(n1812) );
  OAI21X1 U642 ( .A(n4540), .B(n4570), .C(n2895), .Y(n1813) );
  OAI21X1 U644 ( .A(n4540), .B(n4569), .C(n2831), .Y(n1814) );
  OAI21X1 U646 ( .A(n4540), .B(n4568), .C(n2766), .Y(n1815) );
  OAI21X1 U648 ( .A(n4540), .B(n4567), .C(n2702), .Y(n1816) );
  OAI21X1 U650 ( .A(n4540), .B(n4566), .C(n2638), .Y(n1817) );
  OAI21X1 U652 ( .A(n4540), .B(n4565), .C(n354), .Y(n1818) );
  OAI21X1 U654 ( .A(n4540), .B(n4564), .C(n287), .Y(n1819) );
  OAI21X1 U656 ( .A(n4540), .B(n4563), .C(n223), .Y(n1820) );
  OAI21X1 U658 ( .A(n4540), .B(n4562), .C(n159), .Y(n1821) );
  OAI21X1 U660 ( .A(n4540), .B(n4561), .C(n3096), .Y(n1822) );
  OAI21X1 U662 ( .A(n4540), .B(n4560), .C(n3029), .Y(n1823) );
  OAI21X1 U664 ( .A(n4540), .B(n4559), .C(n2961), .Y(n1824) );
  OAI21X1 U666 ( .A(n4540), .B(n4558), .C(n2894), .Y(n1825) );
  OAI21X1 U668 ( .A(n4540), .B(n4557), .C(n2830), .Y(n1826) );
  OAI21X1 U670 ( .A(n4540), .B(n4556), .C(n2765), .Y(n1827) );
  OAI21X1 U672 ( .A(n4540), .B(n4555), .C(n2701), .Y(n1828) );
  OAI21X1 U674 ( .A(n4540), .B(n4554), .C(n2637), .Y(n1829) );
  OAI21X1 U676 ( .A(n4540), .B(n4553), .C(n352), .Y(n1830) );
  OAI21X1 U678 ( .A(n4540), .B(n4552), .C(n286), .Y(n1831) );
  OAI21X1 U680 ( .A(n4540), .B(n4551), .C(n222), .Y(n1832) );
  OAI21X1 U682 ( .A(n4540), .B(n4550), .C(n158), .Y(n1833) );
  OAI21X1 U684 ( .A(n4540), .B(n4549), .C(n103), .Y(n1834) );
  OAI21X1 U686 ( .A(n3118), .B(n3387), .C(reset), .Y(n695) );
  OAI21X1 U687 ( .A(n4539), .B(n4581), .C(n3299), .Y(n1835) );
  OAI21X1 U689 ( .A(n4539), .B(n4580), .C(n3365), .Y(n1836) );
  OAI21X1 U691 ( .A(n4539), .B(n4579), .C(n3166), .Y(n1837) );
  OAI21X1 U693 ( .A(n4539), .B(n4578), .C(n3233), .Y(n1838) );
  OAI21X1 U695 ( .A(n4539), .B(n4577), .C(n3232), .Y(n1839) );
  OAI21X1 U697 ( .A(n4539), .B(n4576), .C(n3298), .Y(n1840) );
  OAI21X1 U699 ( .A(n4539), .B(n4575), .C(n3364), .Y(n1841) );
  OAI21X1 U701 ( .A(n4539), .B(n4574), .C(n3028), .Y(n1842) );
  OAI21X1 U703 ( .A(n4539), .B(n4573), .C(n3165), .Y(n1843) );
  OAI21X1 U705 ( .A(n4539), .B(n4572), .C(n3095), .Y(n1844) );
  OAI21X1 U707 ( .A(n4539), .B(n4571), .C(n2893), .Y(n1845) );
  OAI21X1 U709 ( .A(n4539), .B(n4570), .C(n2960), .Y(n1846) );
  OAI21X1 U711 ( .A(n4539), .B(n4569), .C(n2764), .Y(n1847) );
  OAI21X1 U713 ( .A(n4539), .B(n4568), .C(n2829), .Y(n1848) );
  OAI21X1 U715 ( .A(n4539), .B(n4567), .C(n2636), .Y(n1849) );
  OAI21X1 U717 ( .A(n4539), .B(n4566), .C(n2700), .Y(n1850) );
  OAI21X1 U719 ( .A(n4539), .B(n4565), .C(n285), .Y(n1851) );
  OAI21X1 U721 ( .A(n4539), .B(n4564), .C(n350), .Y(n1852) );
  OAI21X1 U723 ( .A(n4539), .B(n4563), .C(n157), .Y(n1853) );
  OAI21X1 U725 ( .A(n4539), .B(n4562), .C(n221), .Y(n1854) );
  OAI21X1 U727 ( .A(n4539), .B(n4561), .C(n3027), .Y(n1855) );
  OAI21X1 U729 ( .A(n4539), .B(n4560), .C(n3094), .Y(n1856) );
  OAI21X1 U731 ( .A(n4539), .B(n4559), .C(n2892), .Y(n1857) );
  OAI21X1 U733 ( .A(n4539), .B(n4558), .C(n2959), .Y(n1858) );
  OAI21X1 U735 ( .A(n4539), .B(n4557), .C(n2763), .Y(n1859) );
  OAI21X1 U737 ( .A(n4539), .B(n4556), .C(n2828), .Y(n1860) );
  OAI21X1 U739 ( .A(n4539), .B(n4555), .C(n2635), .Y(n1861) );
  OAI21X1 U741 ( .A(n4539), .B(n4554), .C(n2699), .Y(n1862) );
  OAI21X1 U743 ( .A(n4539), .B(n4553), .C(n284), .Y(n1863) );
  OAI21X1 U745 ( .A(n4539), .B(n4552), .C(n348), .Y(n1864) );
  OAI21X1 U747 ( .A(n4539), .B(n4551), .C(n156), .Y(n1865) );
  OAI21X1 U749 ( .A(n4539), .B(n4550), .C(n220), .Y(n1866) );
  OAI21X1 U751 ( .A(n4539), .B(n4549), .C(n102), .Y(n1867) );
  OAI21X1 U753 ( .A(n3048), .B(n3387), .C(reset), .Y(n730) );
  OAI21X1 U754 ( .A(n4538), .B(n4581), .C(n3231), .Y(n1868) );
  OAI21X1 U756 ( .A(n4538), .B(n4580), .C(n3164), .Y(n1869) );
  OAI21X1 U758 ( .A(n4538), .B(n4579), .C(n3363), .Y(n1870) );
  OAI21X1 U760 ( .A(n4538), .B(n4578), .C(n3297), .Y(n1871) );
  OAI21X1 U762 ( .A(n4538), .B(n4577), .C(n3296), .Y(n1872) );
  OAI21X1 U764 ( .A(n4538), .B(n4576), .C(n3230), .Y(n1873) );
  OAI21X1 U766 ( .A(n4538), .B(n4575), .C(n3163), .Y(n1874) );
  OAI21X1 U768 ( .A(n4538), .B(n4574), .C(n2958), .Y(n1875) );
  OAI21X1 U770 ( .A(n4538), .B(n4573), .C(n3362), .Y(n1876) );
  OAI21X1 U772 ( .A(n4538), .B(n4572), .C(n2891), .Y(n1877) );
  OAI21X1 U774 ( .A(n4538), .B(n4571), .C(n3093), .Y(n1878) );
  OAI21X1 U776 ( .A(n4538), .B(n4570), .C(n3026), .Y(n1879) );
  OAI21X1 U778 ( .A(n4538), .B(n4569), .C(n2698), .Y(n1880) );
  OAI21X1 U780 ( .A(n4538), .B(n4568), .C(n2634), .Y(n1881) );
  OAI21X1 U782 ( .A(n4538), .B(n4567), .C(n2827), .Y(n1882) );
  OAI21X1 U784 ( .A(n4538), .B(n4566), .C(n2762), .Y(n1883) );
  OAI21X1 U786 ( .A(n4538), .B(n4565), .C(n219), .Y(n1884) );
  OAI21X1 U788 ( .A(n4538), .B(n4564), .C(n155), .Y(n1885) );
  OAI21X1 U790 ( .A(n4538), .B(n4563), .C(n347), .Y(n1886) );
  OAI21X1 U792 ( .A(n4538), .B(n4562), .C(n283), .Y(n1887) );
  OAI21X1 U794 ( .A(n4538), .B(n4561), .C(n2957), .Y(n1888) );
  OAI21X1 U796 ( .A(n4538), .B(n4560), .C(n2890), .Y(n1889) );
  OAI21X1 U798 ( .A(n4538), .B(n4559), .C(n3092), .Y(n1890) );
  OAI21X1 U800 ( .A(n4538), .B(n4558), .C(n3025), .Y(n1891) );
  OAI21X1 U802 ( .A(n4538), .B(n4557), .C(n2697), .Y(n1892) );
  OAI21X1 U804 ( .A(n4538), .B(n4556), .C(n2633), .Y(n1893) );
  OAI21X1 U806 ( .A(n4538), .B(n4555), .C(n2826), .Y(n1894) );
  OAI21X1 U808 ( .A(n4538), .B(n4554), .C(n2761), .Y(n1895) );
  OAI21X1 U810 ( .A(n4538), .B(n4553), .C(n218), .Y(n1896) );
  OAI21X1 U812 ( .A(n4538), .B(n4552), .C(n154), .Y(n1897) );
  OAI21X1 U814 ( .A(n4538), .B(n4551), .C(n346), .Y(n1898) );
  OAI21X1 U816 ( .A(n4538), .B(n4550), .C(n282), .Y(n1899) );
  OAI21X1 U818 ( .A(n4538), .B(n4549), .C(n101), .Y(n1900) );
  OAI21X1 U820 ( .A(n2980), .B(n3387), .C(reset), .Y(n764) );
  OAI21X1 U821 ( .A(n4537), .B(n4581), .C(n3162), .Y(n1901) );
  OAI21X1 U823 ( .A(n4537), .B(n4580), .C(n3229), .Y(n1902) );
  OAI21X1 U825 ( .A(n4537), .B(n4579), .C(n3295), .Y(n1903) );
  OAI21X1 U827 ( .A(n4537), .B(n4578), .C(n3361), .Y(n1904) );
  OAI21X1 U829 ( .A(n4537), .B(n4577), .C(n3360), .Y(n1905) );
  OAI21X1 U831 ( .A(n4537), .B(n4576), .C(n3161), .Y(n1906) );
  OAI21X1 U833 ( .A(n4537), .B(n4575), .C(n3228), .Y(n1907) );
  OAI21X1 U835 ( .A(n4537), .B(n4574), .C(n2889), .Y(n1908) );
  OAI21X1 U837 ( .A(n4537), .B(n4573), .C(n3294), .Y(n1909) );
  OAI21X1 U839 ( .A(n4537), .B(n4572), .C(n2956), .Y(n1910) );
  OAI21X1 U841 ( .A(n4537), .B(n4571), .C(n3024), .Y(n1911) );
  OAI21X1 U843 ( .A(n4537), .B(n4570), .C(n3091), .Y(n1912) );
  OAI21X1 U845 ( .A(n4537), .B(n4569), .C(n2632), .Y(n1913) );
  OAI21X1 U847 ( .A(n4537), .B(n4568), .C(n2696), .Y(n1914) );
  OAI21X1 U849 ( .A(n4537), .B(n4567), .C(n2760), .Y(n1915) );
  OAI21X1 U851 ( .A(n4537), .B(n4566), .C(n2825), .Y(n1916) );
  OAI21X1 U853 ( .A(n4537), .B(n4565), .C(n153), .Y(n1917) );
  OAI21X1 U855 ( .A(n4537), .B(n4564), .C(n217), .Y(n1918) );
  OAI21X1 U857 ( .A(n4537), .B(n4563), .C(n281), .Y(n1919) );
  OAI21X1 U859 ( .A(n4537), .B(n4562), .C(n345), .Y(n1920) );
  OAI21X1 U861 ( .A(n4537), .B(n4561), .C(n2888), .Y(n1921) );
  OAI21X1 U863 ( .A(n4537), .B(n4560), .C(n2955), .Y(n1922) );
  OAI21X1 U865 ( .A(n4537), .B(n4559), .C(n3023), .Y(n1923) );
  OAI21X1 U867 ( .A(n4537), .B(n4558), .C(n3090), .Y(n1924) );
  OAI21X1 U869 ( .A(n4537), .B(n4557), .C(n2631), .Y(n1925) );
  OAI21X1 U871 ( .A(n4537), .B(n4556), .C(n2695), .Y(n1926) );
  OAI21X1 U873 ( .A(n4537), .B(n4555), .C(n2759), .Y(n1927) );
  OAI21X1 U875 ( .A(n4537), .B(n4554), .C(n2824), .Y(n1928) );
  OAI21X1 U877 ( .A(n4537), .B(n4553), .C(n152), .Y(n1929) );
  OAI21X1 U879 ( .A(n4537), .B(n4552), .C(n216), .Y(n1930) );
  OAI21X1 U881 ( .A(n4537), .B(n4551), .C(n280), .Y(n1931) );
  OAI21X1 U883 ( .A(n4537), .B(n4550), .C(n344), .Y(n1932) );
  OAI21X1 U885 ( .A(n4537), .B(n4549), .C(n100), .Y(n1933) );
  OAI21X1 U887 ( .A(n2913), .B(n3387), .C(reset), .Y(n798) );
  OAI21X1 U888 ( .A(n4536), .B(n4581), .C(n3089), .Y(n1934) );
  OAI21X1 U890 ( .A(n4536), .B(n4580), .C(n3022), .Y(n1935) );
  OAI21X1 U892 ( .A(n4536), .B(n4579), .C(n2954), .Y(n1936) );
  OAI21X1 U894 ( .A(n4536), .B(n4578), .C(n2887), .Y(n1937) );
  OAI21X1 U896 ( .A(n4536), .B(n4577), .C(n2886), .Y(n1938) );
  OAI21X1 U898 ( .A(n4536), .B(n4576), .C(n3088), .Y(n1939) );
  OAI21X1 U900 ( .A(n4536), .B(n4575), .C(n3021), .Y(n1940) );
  OAI21X1 U902 ( .A(n4536), .B(n4574), .C(n3359), .Y(n1941) );
  OAI21X1 U904 ( .A(n4536), .B(n4573), .C(n2953), .Y(n1942) );
  OAI21X1 U906 ( .A(n4536), .B(n4572), .C(n3293), .Y(n1943) );
  OAI21X1 U908 ( .A(n4536), .B(n4571), .C(n3227), .Y(n1944) );
  OAI21X1 U910 ( .A(n4536), .B(n4570), .C(n3160), .Y(n1945) );
  OAI21X1 U912 ( .A(n4536), .B(n4569), .C(n343), .Y(n1946) );
  OAI21X1 U914 ( .A(n4536), .B(n4568), .C(n279), .Y(n1947) );
  OAI21X1 U916 ( .A(n4536), .B(n4567), .C(n215), .Y(n1948) );
  OAI21X1 U918 ( .A(n4536), .B(n4566), .C(n151), .Y(n1949) );
  OAI21X1 U920 ( .A(n4536), .B(n4565), .C(n2823), .Y(n1950) );
  OAI21X1 U922 ( .A(n4536), .B(n4564), .C(n2758), .Y(n1951) );
  OAI21X1 U924 ( .A(n4536), .B(n4563), .C(n2694), .Y(n1952) );
  OAI21X1 U926 ( .A(n4536), .B(n4562), .C(n2630), .Y(n1953) );
  OAI21X1 U928 ( .A(n4536), .B(n4561), .C(n3358), .Y(n1954) );
  OAI21X1 U930 ( .A(n4536), .B(n4560), .C(n3292), .Y(n1955) );
  OAI21X1 U932 ( .A(n4536), .B(n4559), .C(n3226), .Y(n1956) );
  OAI21X1 U934 ( .A(n4536), .B(n4558), .C(n3159), .Y(n1957) );
  OAI21X1 U936 ( .A(n4536), .B(n4557), .C(n342), .Y(n1958) );
  OAI21X1 U938 ( .A(n4536), .B(n4556), .C(n278), .Y(n1959) );
  OAI21X1 U940 ( .A(n4536), .B(n4555), .C(n214), .Y(n1960) );
  OAI21X1 U942 ( .A(n4536), .B(n4554), .C(n150), .Y(n1961) );
  OAI21X1 U944 ( .A(n4536), .B(n4553), .C(n2822), .Y(n1962) );
  OAI21X1 U946 ( .A(n4536), .B(n4552), .C(n2757), .Y(n1963) );
  OAI21X1 U948 ( .A(n4536), .B(n4551), .C(n2693), .Y(n1964) );
  OAI21X1 U950 ( .A(n4536), .B(n4550), .C(n2629), .Y(n1965) );
  OAI21X1 U952 ( .A(n4536), .B(n4549), .C(n99), .Y(n1966) );
  OAI21X1 U954 ( .A(n2912), .B(n3387), .C(reset), .Y(n832) );
  OAI21X1 U955 ( .A(n4535), .B(n4581), .C(n3020), .Y(n1967) );
  OAI21X1 U957 ( .A(n4535), .B(n4580), .C(n3087), .Y(n1968) );
  OAI21X1 U959 ( .A(n4535), .B(n4579), .C(n2885), .Y(n1969) );
  OAI21X1 U961 ( .A(n4535), .B(n4578), .C(n2952), .Y(n1970) );
  OAI21X1 U963 ( .A(n4535), .B(n4577), .C(n2951), .Y(n1971) );
  OAI21X1 U965 ( .A(n4535), .B(n4576), .C(n3019), .Y(n1972) );
  OAI21X1 U967 ( .A(n4535), .B(n4575), .C(n3086), .Y(n1973) );
  OAI21X1 U969 ( .A(n4535), .B(n4574), .C(n3291), .Y(n1974) );
  OAI21X1 U971 ( .A(n4535), .B(n4573), .C(n2884), .Y(n1975) );
  OAI21X1 U973 ( .A(n4535), .B(n4572), .C(n3357), .Y(n1976) );
  OAI21X1 U975 ( .A(n4535), .B(n4571), .C(n3158), .Y(n1977) );
  OAI21X1 U977 ( .A(n4535), .B(n4570), .C(n3225), .Y(n1978) );
  OAI21X1 U979 ( .A(n4535), .B(n4569), .C(n277), .Y(n1979) );
  OAI21X1 U981 ( .A(n4535), .B(n4568), .C(n341), .Y(n1980) );
  OAI21X1 U983 ( .A(n4535), .B(n4567), .C(n149), .Y(n1981) );
  OAI21X1 U985 ( .A(n4535), .B(n4566), .C(n213), .Y(n1982) );
  OAI21X1 U987 ( .A(n4535), .B(n4565), .C(n2756), .Y(n1983) );
  OAI21X1 U989 ( .A(n4535), .B(n4564), .C(n2821), .Y(n1984) );
  OAI21X1 U991 ( .A(n4535), .B(n4563), .C(n2628), .Y(n1985) );
  OAI21X1 U993 ( .A(n4535), .B(n4562), .C(n2692), .Y(n1986) );
  OAI21X1 U995 ( .A(n4535), .B(n4561), .C(n3290), .Y(n1987) );
  OAI21X1 U997 ( .A(n4535), .B(n4560), .C(n3356), .Y(n1988) );
  OAI21X1 U999 ( .A(n4535), .B(n4559), .C(n3157), .Y(n1989) );
  OAI21X1 U1001 ( .A(n4535), .B(n4558), .C(n3224), .Y(n1990) );
  OAI21X1 U1003 ( .A(n4535), .B(n4557), .C(n276), .Y(n1991) );
  OAI21X1 U1005 ( .A(n4535), .B(n4556), .C(n340), .Y(n1992) );
  OAI21X1 U1007 ( .A(n4535), .B(n4555), .C(n148), .Y(n1993) );
  OAI21X1 U1009 ( .A(n4535), .B(n4554), .C(n212), .Y(n1994) );
  OAI21X1 U1011 ( .A(n4535), .B(n4553), .C(n2755), .Y(n1995) );
  OAI21X1 U1013 ( .A(n4535), .B(n4552), .C(n2820), .Y(n1996) );
  OAI21X1 U1015 ( .A(n4535), .B(n4551), .C(n2627), .Y(n1997) );
  OAI21X1 U1017 ( .A(n4535), .B(n4550), .C(n2691), .Y(n1998) );
  OAI21X1 U1019 ( .A(n4535), .B(n4549), .C(n98), .Y(n1999) );
  OAI21X1 U1021 ( .A(n2979), .B(n3387), .C(reset), .Y(n866) );
  OAI21X1 U1022 ( .A(n4534), .B(n4581), .C(n2950), .Y(n2000) );
  OAI21X1 U1024 ( .A(n4534), .B(n4580), .C(n2883), .Y(n2001) );
  OAI21X1 U1026 ( .A(n4534), .B(n4579), .C(n3085), .Y(n2002) );
  OAI21X1 U1028 ( .A(n4534), .B(n4578), .C(n3018), .Y(n2003) );
  OAI21X1 U1030 ( .A(n4534), .B(n4577), .C(n3017), .Y(n2004) );
  OAI21X1 U1032 ( .A(n4534), .B(n4576), .C(n2949), .Y(n2005) );
  OAI21X1 U1034 ( .A(n4534), .B(n4575), .C(n2882), .Y(n2006) );
  OAI21X1 U1036 ( .A(n4534), .B(n4574), .C(n3223), .Y(n2007) );
  OAI21X1 U1038 ( .A(n4534), .B(n4573), .C(n3084), .Y(n2008) );
  OAI21X1 U1040 ( .A(n4534), .B(n4572), .C(n3156), .Y(n2009) );
  OAI21X1 U1042 ( .A(n4534), .B(n4571), .C(n3355), .Y(n2010) );
  OAI21X1 U1044 ( .A(n4534), .B(n4570), .C(n3289), .Y(n2011) );
  OAI21X1 U1046 ( .A(n4534), .B(n4569), .C(n211), .Y(n2012) );
  OAI21X1 U1048 ( .A(n4534), .B(n4568), .C(n147), .Y(n2013) );
  OAI21X1 U1050 ( .A(n4534), .B(n4567), .C(n339), .Y(n2014) );
  OAI21X1 U1052 ( .A(n4534), .B(n4566), .C(n275), .Y(n2015) );
  OAI21X1 U1054 ( .A(n4534), .B(n4565), .C(n2690), .Y(n2016) );
  OAI21X1 U1056 ( .A(n4534), .B(n4564), .C(n2626), .Y(n2017) );
  OAI21X1 U1058 ( .A(n4534), .B(n4563), .C(n2819), .Y(n2018) );
  OAI21X1 U1060 ( .A(n4534), .B(n4562), .C(n2754), .Y(n2019) );
  OAI21X1 U1062 ( .A(n4534), .B(n4561), .C(n3222), .Y(n2020) );
  OAI21X1 U1064 ( .A(n4534), .B(n4560), .C(n3155), .Y(n2021) );
  OAI21X1 U1066 ( .A(n4534), .B(n4559), .C(n3354), .Y(n2022) );
  OAI21X1 U1068 ( .A(n4534), .B(n4558), .C(n3288), .Y(n2023) );
  OAI21X1 U1070 ( .A(n4534), .B(n4557), .C(n210), .Y(n2024) );
  OAI21X1 U1072 ( .A(n4534), .B(n4556), .C(n146), .Y(n2025) );
  OAI21X1 U1074 ( .A(n4534), .B(n4555), .C(n338), .Y(n2026) );
  OAI21X1 U1076 ( .A(n4534), .B(n4554), .C(n274), .Y(n2027) );
  OAI21X1 U1078 ( .A(n4534), .B(n4553), .C(n2689), .Y(n2028) );
  OAI21X1 U1080 ( .A(n4534), .B(n4552), .C(n2625), .Y(n2029) );
  OAI21X1 U1082 ( .A(n4534), .B(n4551), .C(n2818), .Y(n2030) );
  OAI21X1 U1084 ( .A(n4534), .B(n4550), .C(n2753), .Y(n2031) );
  OAI21X1 U1086 ( .A(n4534), .B(n4549), .C(n97), .Y(n2032) );
  OAI21X1 U1088 ( .A(n3047), .B(n3387), .C(reset), .Y(n900) );
  OAI21X1 U1089 ( .A(n4533), .B(n4581), .C(n2881), .Y(n2033) );
  OAI21X1 U1091 ( .A(n4533), .B(n4580), .C(n2948), .Y(n2034) );
  OAI21X1 U1093 ( .A(n4533), .B(n4579), .C(n3016), .Y(n2035) );
  OAI21X1 U1095 ( .A(n4533), .B(n4578), .C(n3083), .Y(n2036) );
  OAI21X1 U1097 ( .A(n4533), .B(n4577), .C(n3082), .Y(n2037) );
  OAI21X1 U1099 ( .A(n4533), .B(n4576), .C(n2880), .Y(n2038) );
  OAI21X1 U1101 ( .A(n4533), .B(n4575), .C(n2947), .Y(n2039) );
  OAI21X1 U1103 ( .A(n4533), .B(n4574), .C(n3154), .Y(n2040) );
  OAI21X1 U1105 ( .A(n4533), .B(n4573), .C(n3015), .Y(n2041) );
  OAI21X1 U1107 ( .A(n4533), .B(n4572), .C(n3221), .Y(n2042) );
  OAI21X1 U1109 ( .A(n4533), .B(n4571), .C(n3287), .Y(n2043) );
  OAI21X1 U1111 ( .A(n4533), .B(n4570), .C(n3353), .Y(n2044) );
  OAI21X1 U1113 ( .A(n4533), .B(n4569), .C(n145), .Y(n2045) );
  OAI21X1 U1115 ( .A(n4533), .B(n4568), .C(n209), .Y(n2046) );
  OAI21X1 U1117 ( .A(n4533), .B(n4567), .C(n273), .Y(n2047) );
  OAI21X1 U1119 ( .A(n4533), .B(n4566), .C(n337), .Y(n2048) );
  OAI21X1 U1121 ( .A(n4533), .B(n4565), .C(n2624), .Y(n2049) );
  OAI21X1 U1123 ( .A(n4533), .B(n4564), .C(n2688), .Y(n2050) );
  OAI21X1 U1125 ( .A(n4533), .B(n4563), .C(n2752), .Y(n2051) );
  OAI21X1 U1127 ( .A(n4533), .B(n4562), .C(n2817), .Y(n2052) );
  OAI21X1 U1129 ( .A(n4533), .B(n4561), .C(n3153), .Y(n2053) );
  OAI21X1 U1131 ( .A(n4533), .B(n4560), .C(n3220), .Y(n2054) );
  OAI21X1 U1133 ( .A(n4533), .B(n4559), .C(n3286), .Y(n2055) );
  OAI21X1 U1135 ( .A(n4533), .B(n4558), .C(n3352), .Y(n2056) );
  OAI21X1 U1137 ( .A(n4533), .B(n4557), .C(n144), .Y(n2057) );
  OAI21X1 U1139 ( .A(n4533), .B(n4556), .C(n208), .Y(n2058) );
  OAI21X1 U1141 ( .A(n4533), .B(n4555), .C(n272), .Y(n2059) );
  OAI21X1 U1143 ( .A(n4533), .B(n4554), .C(n336), .Y(n2060) );
  OAI21X1 U1145 ( .A(n4533), .B(n4553), .C(n2623), .Y(n2061) );
  OAI21X1 U1147 ( .A(n4533), .B(n4552), .C(n2687), .Y(n2062) );
  OAI21X1 U1149 ( .A(n4533), .B(n4551), .C(n2751), .Y(n2063) );
  OAI21X1 U1151 ( .A(n4533), .B(n4550), .C(n2816), .Y(n2064) );
  OAI21X1 U1153 ( .A(n4533), .B(n4549), .C(n96), .Y(n2065) );
  OAI21X1 U1155 ( .A(n3117), .B(n3387), .C(reset), .Y(n934) );
  NAND3X1 U1156 ( .A(n1481), .B(n4620), .C(wr_ptr[3]), .Y(n696) );
  OAI21X1 U1157 ( .A(n4532), .B(n4581), .C(n2815), .Y(n2066) );
  OAI21X1 U1159 ( .A(n4532), .B(n4580), .C(n2750), .Y(n2067) );
  OAI21X1 U1161 ( .A(n4532), .B(n4579), .C(n2686), .Y(n2068) );
  OAI21X1 U1163 ( .A(n4532), .B(n4578), .C(n2622), .Y(n2069) );
  OAI21X1 U1165 ( .A(n4532), .B(n4577), .C(n2621), .Y(n2070) );
  OAI21X1 U1167 ( .A(n4532), .B(n4576), .C(n2814), .Y(n2071) );
  OAI21X1 U1169 ( .A(n4532), .B(n4575), .C(n2749), .Y(n2072) );
  OAI21X1 U1171 ( .A(n4532), .B(n4574), .C(n335), .Y(n2073) );
  OAI21X1 U1173 ( .A(n4532), .B(n4573), .C(n2685), .Y(n2074) );
  OAI21X1 U1175 ( .A(n4532), .B(n4572), .C(n271), .Y(n2075) );
  OAI21X1 U1177 ( .A(n4532), .B(n4571), .C(n207), .Y(n2076) );
  OAI21X1 U1179 ( .A(n4532), .B(n4570), .C(n143), .Y(n2077) );
  OAI21X1 U1181 ( .A(n4532), .B(n4569), .C(n3351), .Y(n2078) );
  OAI21X1 U1183 ( .A(n4532), .B(n4568), .C(n3285), .Y(n2079) );
  OAI21X1 U1185 ( .A(n4532), .B(n4567), .C(n3219), .Y(n2080) );
  OAI21X1 U1187 ( .A(n4532), .B(n4566), .C(n3152), .Y(n2081) );
  OAI21X1 U1189 ( .A(n4532), .B(n4565), .C(n3081), .Y(n2082) );
  OAI21X1 U1191 ( .A(n4532), .B(n4564), .C(n3014), .Y(n2083) );
  OAI21X1 U1193 ( .A(n4532), .B(n4563), .C(n2946), .Y(n2084) );
  OAI21X1 U1195 ( .A(n4532), .B(n4562), .C(n2879), .Y(n2085) );
  OAI21X1 U1197 ( .A(n4532), .B(n4561), .C(n334), .Y(n2086) );
  OAI21X1 U1199 ( .A(n4532), .B(n4560), .C(n270), .Y(n2087) );
  OAI21X1 U1201 ( .A(n4532), .B(n4559), .C(n206), .Y(n2088) );
  OAI21X1 U1203 ( .A(n4532), .B(n4558), .C(n142), .Y(n2089) );
  OAI21X1 U1205 ( .A(n4532), .B(n4557), .C(n3350), .Y(n2090) );
  OAI21X1 U1207 ( .A(n4532), .B(n4556), .C(n3284), .Y(n2091) );
  OAI21X1 U1209 ( .A(n4532), .B(n4555), .C(n3218), .Y(n2092) );
  OAI21X1 U1211 ( .A(n4532), .B(n4554), .C(n3151), .Y(n2093) );
  OAI21X1 U1213 ( .A(n4532), .B(n4553), .C(n3080), .Y(n2094) );
  OAI21X1 U1215 ( .A(n4532), .B(n4552), .C(n3013), .Y(n2095) );
  OAI21X1 U1217 ( .A(n4532), .B(n4551), .C(n2945), .Y(n2096) );
  OAI21X1 U1219 ( .A(n4532), .B(n4550), .C(n2878), .Y(n2097) );
  OAI21X1 U1221 ( .A(n4532), .B(n4549), .C(n95), .Y(n2098) );
  OAI21X1 U1223 ( .A(n3118), .B(n3319), .C(reset), .Y(n968) );
  OAI21X1 U1224 ( .A(n4531), .B(n4581), .C(n2748), .Y(n2099) );
  OAI21X1 U1226 ( .A(n4531), .B(n4580), .C(n2813), .Y(n2100) );
  OAI21X1 U1228 ( .A(n4531), .B(n4579), .C(n2620), .Y(n2101) );
  OAI21X1 U1230 ( .A(n4531), .B(n4578), .C(n2684), .Y(n2102) );
  OAI21X1 U1232 ( .A(n4531), .B(n4577), .C(n2683), .Y(n2103) );
  OAI21X1 U1234 ( .A(n4531), .B(n4576), .C(n2747), .Y(n2104) );
  OAI21X1 U1236 ( .A(n4531), .B(n4575), .C(n2812), .Y(n2105) );
  OAI21X1 U1238 ( .A(n4531), .B(n4574), .C(n269), .Y(n2106) );
  OAI21X1 U1240 ( .A(n4531), .B(n4573), .C(n2619), .Y(n2107) );
  OAI21X1 U1242 ( .A(n4531), .B(n4572), .C(n333), .Y(n2108) );
  OAI21X1 U1244 ( .A(n4531), .B(n4571), .C(n141), .Y(n2109) );
  OAI21X1 U1246 ( .A(n4531), .B(n4570), .C(n205), .Y(n2110) );
  OAI21X1 U1248 ( .A(n4531), .B(n4569), .C(n3283), .Y(n2111) );
  OAI21X1 U1250 ( .A(n4531), .B(n4568), .C(n3349), .Y(n2112) );
  OAI21X1 U1252 ( .A(n4531), .B(n4567), .C(n3150), .Y(n2113) );
  OAI21X1 U1254 ( .A(n4531), .B(n4566), .C(n3217), .Y(n2114) );
  OAI21X1 U1256 ( .A(n4531), .B(n4565), .C(n3012), .Y(n2115) );
  OAI21X1 U1258 ( .A(n4531), .B(n4564), .C(n3079), .Y(n2116) );
  OAI21X1 U1260 ( .A(n4531), .B(n4563), .C(n2877), .Y(n2117) );
  OAI21X1 U1262 ( .A(n4531), .B(n4562), .C(n2944), .Y(n2118) );
  OAI21X1 U1264 ( .A(n4531), .B(n4561), .C(n268), .Y(n2119) );
  OAI21X1 U1266 ( .A(n4531), .B(n4560), .C(n332), .Y(n2120) );
  OAI21X1 U1268 ( .A(n4531), .B(n4559), .C(n140), .Y(n2121) );
  OAI21X1 U1270 ( .A(n4531), .B(n4558), .C(n204), .Y(n2122) );
  OAI21X1 U1272 ( .A(n4531), .B(n4557), .C(n3282), .Y(n2123) );
  OAI21X1 U1274 ( .A(n4531), .B(n4556), .C(n3348), .Y(n2124) );
  OAI21X1 U1276 ( .A(n4531), .B(n4555), .C(n3149), .Y(n2125) );
  OAI21X1 U1278 ( .A(n4531), .B(n4554), .C(n3216), .Y(n2126) );
  OAI21X1 U1280 ( .A(n4531), .B(n4553), .C(n3011), .Y(n2127) );
  OAI21X1 U1282 ( .A(n4531), .B(n4552), .C(n3078), .Y(n2128) );
  OAI21X1 U1284 ( .A(n4531), .B(n4551), .C(n2876), .Y(n2129) );
  OAI21X1 U1286 ( .A(n4531), .B(n4550), .C(n2943), .Y(n2130) );
  OAI21X1 U1288 ( .A(n4531), .B(n4549), .C(n94), .Y(n2131) );
  OAI21X1 U1290 ( .A(n3048), .B(n3319), .C(reset), .Y(n1003) );
  OAI21X1 U1291 ( .A(n4530), .B(n4581), .C(n2682), .Y(n2132) );
  OAI21X1 U1293 ( .A(n4530), .B(n4580), .C(n2618), .Y(n2133) );
  OAI21X1 U1295 ( .A(n4530), .B(n4579), .C(n2811), .Y(n2134) );
  OAI21X1 U1297 ( .A(n4530), .B(n4578), .C(n2746), .Y(n2135) );
  OAI21X1 U1299 ( .A(n4530), .B(n4577), .C(n2745), .Y(n2136) );
  OAI21X1 U1301 ( .A(n4530), .B(n4576), .C(n2681), .Y(n2137) );
  OAI21X1 U1303 ( .A(n4530), .B(n4575), .C(n2617), .Y(n2138) );
  OAI21X1 U1305 ( .A(n4530), .B(n4574), .C(n203), .Y(n2139) );
  OAI21X1 U1307 ( .A(n4530), .B(n4573), .C(n2810), .Y(n2140) );
  OAI21X1 U1309 ( .A(n4530), .B(n4572), .C(n139), .Y(n2141) );
  OAI21X1 U1311 ( .A(n4530), .B(n4571), .C(n331), .Y(n2142) );
  OAI21X1 U1313 ( .A(n4530), .B(n4570), .C(n267), .Y(n2143) );
  OAI21X1 U1315 ( .A(n4530), .B(n4569), .C(n3215), .Y(n2144) );
  OAI21X1 U1317 ( .A(n4530), .B(n4568), .C(n3148), .Y(n2145) );
  OAI21X1 U1319 ( .A(n4530), .B(n4567), .C(n3347), .Y(n2146) );
  OAI21X1 U1321 ( .A(n4530), .B(n4566), .C(n3281), .Y(n2147) );
  OAI21X1 U1323 ( .A(n4530), .B(n4565), .C(n2942), .Y(n2148) );
  OAI21X1 U1325 ( .A(n4530), .B(n4564), .C(n2875), .Y(n2149) );
  OAI21X1 U1327 ( .A(n4530), .B(n4563), .C(n3077), .Y(n2150) );
  OAI21X1 U1329 ( .A(n4530), .B(n4562), .C(n3010), .Y(n2151) );
  OAI21X1 U1331 ( .A(n4530), .B(n4561), .C(n202), .Y(n2152) );
  OAI21X1 U1333 ( .A(n4530), .B(n4560), .C(n138), .Y(n2153) );
  OAI21X1 U1335 ( .A(n4530), .B(n4559), .C(n330), .Y(n2154) );
  OAI21X1 U1337 ( .A(n4530), .B(n4558), .C(n266), .Y(n2155) );
  OAI21X1 U1339 ( .A(n4530), .B(n4557), .C(n3214), .Y(n2156) );
  OAI21X1 U1341 ( .A(n4530), .B(n4556), .C(n3147), .Y(n2157) );
  OAI21X1 U1343 ( .A(n4530), .B(n4555), .C(n3346), .Y(n2158) );
  OAI21X1 U1345 ( .A(n4530), .B(n4554), .C(n3280), .Y(n2159) );
  OAI21X1 U1347 ( .A(n4530), .B(n4553), .C(n2941), .Y(n2160) );
  OAI21X1 U1349 ( .A(n4530), .B(n4552), .C(n2874), .Y(n2161) );
  OAI21X1 U1351 ( .A(n4530), .B(n4551), .C(n3076), .Y(n2162) );
  OAI21X1 U1353 ( .A(n4530), .B(n4550), .C(n3009), .Y(n2163) );
  OAI21X1 U1355 ( .A(n4530), .B(n4549), .C(n89), .Y(n2164) );
  OAI21X1 U1357 ( .A(n2980), .B(n3319), .C(reset), .Y(n1037) );
  OAI21X1 U1358 ( .A(n4529), .B(n4581), .C(n2616), .Y(n2165) );
  OAI21X1 U1360 ( .A(n4529), .B(n4580), .C(n2680), .Y(n2166) );
  OAI21X1 U1362 ( .A(n4529), .B(n4579), .C(n2744), .Y(n2167) );
  OAI21X1 U1364 ( .A(n4529), .B(n4578), .C(n2809), .Y(n2168) );
  OAI21X1 U1366 ( .A(n4529), .B(n4577), .C(n2808), .Y(n2169) );
  OAI21X1 U1368 ( .A(n4529), .B(n4576), .C(n2615), .Y(n2170) );
  OAI21X1 U1370 ( .A(n4529), .B(n4575), .C(n2679), .Y(n2171) );
  OAI21X1 U1372 ( .A(n4529), .B(n4574), .C(n137), .Y(n2172) );
  OAI21X1 U1374 ( .A(n4529), .B(n4573), .C(n2743), .Y(n2173) );
  OAI21X1 U1376 ( .A(n4529), .B(n4572), .C(n201), .Y(n2174) );
  OAI21X1 U1378 ( .A(n4529), .B(n4571), .C(n265), .Y(n2175) );
  OAI21X1 U1380 ( .A(n4529), .B(n4570), .C(n329), .Y(n2176) );
  OAI21X1 U1382 ( .A(n4529), .B(n4569), .C(n3146), .Y(n2177) );
  OAI21X1 U1384 ( .A(n4529), .B(n4568), .C(n3213), .Y(n2178) );
  OAI21X1 U1386 ( .A(n4529), .B(n4567), .C(n3279), .Y(n2179) );
  OAI21X1 U1388 ( .A(n4529), .B(n4566), .C(n3345), .Y(n2180) );
  OAI21X1 U1390 ( .A(n4529), .B(n4565), .C(n2873), .Y(n2181) );
  OAI21X1 U1392 ( .A(n4529), .B(n4564), .C(n2940), .Y(n2182) );
  OAI21X1 U1394 ( .A(n4529), .B(n4563), .C(n3008), .Y(n2183) );
  OAI21X1 U1396 ( .A(n4529), .B(n4562), .C(n3075), .Y(n2184) );
  OAI21X1 U1398 ( .A(n4529), .B(n4561), .C(n136), .Y(n2185) );
  OAI21X1 U1400 ( .A(n4529), .B(n4560), .C(n200), .Y(n2186) );
  OAI21X1 U1402 ( .A(n4529), .B(n4559), .C(n264), .Y(n2187) );
  OAI21X1 U1404 ( .A(n4529), .B(n4558), .C(n328), .Y(n2188) );
  OAI21X1 U1406 ( .A(n4529), .B(n4557), .C(n3145), .Y(n2189) );
  OAI21X1 U1408 ( .A(n4529), .B(n4556), .C(n3212), .Y(n2190) );
  OAI21X1 U1410 ( .A(n4529), .B(n4555), .C(n3278), .Y(n2191) );
  OAI21X1 U1412 ( .A(n4529), .B(n4554), .C(n3344), .Y(n2192) );
  OAI21X1 U1414 ( .A(n4529), .B(n4553), .C(n2872), .Y(n2193) );
  OAI21X1 U1416 ( .A(n4529), .B(n4552), .C(n2939), .Y(n2194) );
  OAI21X1 U1418 ( .A(n4529), .B(n4551), .C(n3007), .Y(n2195) );
  OAI21X1 U1420 ( .A(n4529), .B(n4550), .C(n3074), .Y(n2196) );
  OAI21X1 U1422 ( .A(n4529), .B(n4549), .C(n55), .Y(n2197) );
  OAI21X1 U1424 ( .A(n2913), .B(n3319), .C(reset), .Y(n1071) );
  OAI21X1 U1425 ( .A(n4528), .B(n4581), .C(n3343), .Y(n2198) );
  OAI21X1 U1427 ( .A(n4528), .B(n4580), .C(n3277), .Y(n2199) );
  OAI21X1 U1429 ( .A(n4528), .B(n4579), .C(n3211), .Y(n2200) );
  OAI21X1 U1431 ( .A(n4528), .B(n4578), .C(n3144), .Y(n2201) );
  OAI21X1 U1433 ( .A(n4528), .B(n4577), .C(n3143), .Y(n2202) );
  OAI21X1 U1435 ( .A(n4528), .B(n4576), .C(n3342), .Y(n2203) );
  OAI21X1 U1437 ( .A(n4528), .B(n4575), .C(n3276), .Y(n2204) );
  OAI21X1 U1439 ( .A(n4528), .B(n4574), .C(n3073), .Y(n2205) );
  OAI21X1 U1441 ( .A(n4528), .B(n4573), .C(n3210), .Y(n2206) );
  OAI21X1 U1443 ( .A(n4528), .B(n4572), .C(n3006), .Y(n2207) );
  OAI21X1 U1445 ( .A(n4528), .B(n4571), .C(n2938), .Y(n2208) );
  OAI21X1 U1447 ( .A(n4528), .B(n4570), .C(n2871), .Y(n2209) );
  OAI21X1 U1449 ( .A(n4528), .B(n4569), .C(n2807), .Y(n2210) );
  OAI21X1 U1451 ( .A(n4528), .B(n4568), .C(n2742), .Y(n2211) );
  OAI21X1 U1453 ( .A(n4528), .B(n4567), .C(n2678), .Y(n2212) );
  OAI21X1 U1455 ( .A(n4528), .B(n4566), .C(n2614), .Y(n2213) );
  OAI21X1 U1457 ( .A(n4528), .B(n4565), .C(n327), .Y(n2214) );
  OAI21X1 U1459 ( .A(n4528), .B(n4564), .C(n263), .Y(n2215) );
  OAI21X1 U1461 ( .A(n4528), .B(n4563), .C(n199), .Y(n2216) );
  OAI21X1 U1463 ( .A(n4528), .B(n4562), .C(n135), .Y(n2217) );
  OAI21X1 U1465 ( .A(n4528), .B(n4561), .C(n3072), .Y(n2218) );
  OAI21X1 U1467 ( .A(n4528), .B(n4560), .C(n3005), .Y(n2219) );
  OAI21X1 U1469 ( .A(n4528), .B(n4559), .C(n2937), .Y(n2220) );
  OAI21X1 U1471 ( .A(n4528), .B(n4558), .C(n2870), .Y(n2221) );
  OAI21X1 U1473 ( .A(n4528), .B(n4557), .C(n2806), .Y(n2222) );
  OAI21X1 U1475 ( .A(n4528), .B(n4556), .C(n2741), .Y(n2223) );
  OAI21X1 U1477 ( .A(n4528), .B(n4555), .C(n2677), .Y(n2224) );
  OAI21X1 U1479 ( .A(n4528), .B(n4554), .C(n2613), .Y(n2225) );
  OAI21X1 U1481 ( .A(n4528), .B(n4553), .C(n326), .Y(n2226) );
  OAI21X1 U1483 ( .A(n4528), .B(n4552), .C(n262), .Y(n2227) );
  OAI21X1 U1485 ( .A(n4528), .B(n4551), .C(n198), .Y(n2228) );
  OAI21X1 U1487 ( .A(n4528), .B(n4550), .C(n134), .Y(n2229) );
  OAI21X1 U1489 ( .A(n4528), .B(n4549), .C(n54), .Y(n2230) );
  OAI21X1 U1491 ( .A(n2912), .B(n3319), .C(reset), .Y(n1105) );
  OAI21X1 U1492 ( .A(n4527), .B(n4581), .C(n3275), .Y(n2231) );
  OAI21X1 U1494 ( .A(n4527), .B(n4580), .C(n3341), .Y(n2232) );
  OAI21X1 U1496 ( .A(n4527), .B(n4579), .C(n3142), .Y(n2233) );
  OAI21X1 U1498 ( .A(n4527), .B(n4578), .C(n3209), .Y(n2234) );
  OAI21X1 U1500 ( .A(n4527), .B(n4577), .C(n3208), .Y(n2235) );
  OAI21X1 U1502 ( .A(n4527), .B(n4576), .C(n3274), .Y(n2236) );
  OAI21X1 U1504 ( .A(n4527), .B(n4575), .C(n3340), .Y(n2237) );
  OAI21X1 U1506 ( .A(n4527), .B(n4574), .C(n3004), .Y(n2238) );
  OAI21X1 U1508 ( .A(n4527), .B(n4573), .C(n3141), .Y(n2239) );
  OAI21X1 U1510 ( .A(n4527), .B(n4572), .C(n3071), .Y(n2240) );
  OAI21X1 U1512 ( .A(n4527), .B(n4571), .C(n2869), .Y(n2241) );
  OAI21X1 U1514 ( .A(n4527), .B(n4570), .C(n2936), .Y(n2242) );
  OAI21X1 U1516 ( .A(n4527), .B(n4569), .C(n2740), .Y(n2243) );
  OAI21X1 U1518 ( .A(n4527), .B(n4568), .C(n2805), .Y(n2244) );
  OAI21X1 U1520 ( .A(n4527), .B(n4567), .C(n2612), .Y(n2245) );
  OAI21X1 U1522 ( .A(n4527), .B(n4566), .C(n2676), .Y(n2246) );
  OAI21X1 U1524 ( .A(n4527), .B(n4565), .C(n261), .Y(n2247) );
  OAI21X1 U1526 ( .A(n4527), .B(n4564), .C(n325), .Y(n2248) );
  OAI21X1 U1528 ( .A(n4527), .B(n4563), .C(n133), .Y(n2249) );
  OAI21X1 U1530 ( .A(n4527), .B(n4562), .C(n197), .Y(n2250) );
  OAI21X1 U1532 ( .A(n4527), .B(n4561), .C(n3003), .Y(n2251) );
  OAI21X1 U1534 ( .A(n4527), .B(n4560), .C(n3070), .Y(n2252) );
  OAI21X1 U1536 ( .A(n4527), .B(n4559), .C(n2868), .Y(n2253) );
  OAI21X1 U1538 ( .A(n4527), .B(n4558), .C(n2935), .Y(n2254) );
  OAI21X1 U1540 ( .A(n4527), .B(n4557), .C(n2739), .Y(n2255) );
  OAI21X1 U1542 ( .A(n4527), .B(n4556), .C(n2804), .Y(n2256) );
  OAI21X1 U1544 ( .A(n4527), .B(n4555), .C(n2611), .Y(n2257) );
  OAI21X1 U1546 ( .A(n4527), .B(n4554), .C(n2675), .Y(n2258) );
  OAI21X1 U1548 ( .A(n4527), .B(n4553), .C(n260), .Y(n2259) );
  OAI21X1 U1550 ( .A(n4527), .B(n4552), .C(n324), .Y(n2260) );
  OAI21X1 U1552 ( .A(n4527), .B(n4551), .C(n132), .Y(n2261) );
  OAI21X1 U1554 ( .A(n4527), .B(n4550), .C(n196), .Y(n2262) );
  OAI21X1 U1556 ( .A(n4527), .B(n4549), .C(n53), .Y(n2263) );
  OAI21X1 U1558 ( .A(n2979), .B(n3319), .C(reset), .Y(n1139) );
  OAI21X1 U1559 ( .A(n4526), .B(n4581), .C(n3207), .Y(n2264) );
  OAI21X1 U1561 ( .A(n4526), .B(n4580), .C(n3140), .Y(n2265) );
  OAI21X1 U1563 ( .A(n4526), .B(n4579), .C(n3339), .Y(n2266) );
  OAI21X1 U1565 ( .A(n4526), .B(n4578), .C(n3273), .Y(n2267) );
  OAI21X1 U1567 ( .A(n4526), .B(n4577), .C(n3272), .Y(n2268) );
  OAI21X1 U1569 ( .A(n4526), .B(n4576), .C(n3206), .Y(n2269) );
  OAI21X1 U1571 ( .A(n4526), .B(n4575), .C(n3139), .Y(n2270) );
  OAI21X1 U1573 ( .A(n4526), .B(n4574), .C(n2934), .Y(n2271) );
  OAI21X1 U1575 ( .A(n4526), .B(n4573), .C(n3338), .Y(n2272) );
  OAI21X1 U1577 ( .A(n4526), .B(n4572), .C(n2867), .Y(n2273) );
  OAI21X1 U1579 ( .A(n4526), .B(n4571), .C(n3069), .Y(n2274) );
  OAI21X1 U1581 ( .A(n4526), .B(n4570), .C(n3002), .Y(n2275) );
  OAI21X1 U1583 ( .A(n4526), .B(n4569), .C(n2674), .Y(n2276) );
  OAI21X1 U1585 ( .A(n4526), .B(n4568), .C(n2610), .Y(n2277) );
  OAI21X1 U1587 ( .A(n4526), .B(n4567), .C(n2803), .Y(n2278) );
  OAI21X1 U1589 ( .A(n4526), .B(n4566), .C(n2738), .Y(n2279) );
  OAI21X1 U1591 ( .A(n4526), .B(n4565), .C(n195), .Y(n2280) );
  OAI21X1 U1593 ( .A(n4526), .B(n4564), .C(n131), .Y(n2281) );
  OAI21X1 U1595 ( .A(n4526), .B(n4563), .C(n323), .Y(n2282) );
  OAI21X1 U1597 ( .A(n4526), .B(n4562), .C(n259), .Y(n2283) );
  OAI21X1 U1599 ( .A(n4526), .B(n4561), .C(n2933), .Y(n2284) );
  OAI21X1 U1601 ( .A(n4526), .B(n4560), .C(n2866), .Y(n2285) );
  OAI21X1 U1603 ( .A(n4526), .B(n4559), .C(n3068), .Y(n2286) );
  OAI21X1 U1605 ( .A(n4526), .B(n4558), .C(n3001), .Y(n2287) );
  OAI21X1 U1607 ( .A(n4526), .B(n4557), .C(n2673), .Y(n2288) );
  OAI21X1 U1609 ( .A(n4526), .B(n4556), .C(n2609), .Y(n2289) );
  OAI21X1 U1611 ( .A(n4526), .B(n4555), .C(n2802), .Y(n2290) );
  OAI21X1 U1613 ( .A(n4526), .B(n4554), .C(n2737), .Y(n2291) );
  OAI21X1 U1615 ( .A(n4526), .B(n4553), .C(n194), .Y(n2292) );
  OAI21X1 U1617 ( .A(n4526), .B(n4552), .C(n130), .Y(n2293) );
  OAI21X1 U1619 ( .A(n4526), .B(n4551), .C(n322), .Y(n2294) );
  OAI21X1 U1621 ( .A(n4526), .B(n4550), .C(n258), .Y(n2295) );
  OAI21X1 U1623 ( .A(n4526), .B(n4549), .C(n52), .Y(n2296) );
  OAI21X1 U1625 ( .A(n3047), .B(n3319), .C(reset), .Y(n1173) );
  OAI21X1 U1626 ( .A(n4525), .B(n4581), .C(n3138), .Y(n2297) );
  OAI21X1 U1628 ( .A(n4525), .B(n4580), .C(n3205), .Y(n2298) );
  OAI21X1 U1630 ( .A(n4525), .B(n4579), .C(n3271), .Y(n2299) );
  OAI21X1 U1632 ( .A(n4525), .B(n4578), .C(n3337), .Y(n2300) );
  OAI21X1 U1634 ( .A(n4525), .B(n4577), .C(n3336), .Y(n2301) );
  OAI21X1 U1636 ( .A(n4525), .B(n4576), .C(n3137), .Y(n2302) );
  OAI21X1 U1638 ( .A(n4525), .B(n4575), .C(n3204), .Y(n2303) );
  OAI21X1 U1640 ( .A(n4525), .B(n4574), .C(n2865), .Y(n2304) );
  OAI21X1 U1642 ( .A(n4525), .B(n4573), .C(n3270), .Y(n2305) );
  OAI21X1 U1644 ( .A(n4525), .B(n4572), .C(n2932), .Y(n2306) );
  OAI21X1 U1646 ( .A(n4525), .B(n4571), .C(n3000), .Y(n2307) );
  OAI21X1 U1648 ( .A(n4525), .B(n4570), .C(n3067), .Y(n2308) );
  OAI21X1 U1650 ( .A(n4525), .B(n4569), .C(n2608), .Y(n2309) );
  OAI21X1 U1652 ( .A(n4525), .B(n4568), .C(n2672), .Y(n2310) );
  OAI21X1 U1654 ( .A(n4525), .B(n4567), .C(n2736), .Y(n2311) );
  OAI21X1 U1656 ( .A(n4525), .B(n4566), .C(n2801), .Y(n2312) );
  OAI21X1 U1658 ( .A(n4525), .B(n4565), .C(n129), .Y(n2313) );
  OAI21X1 U1660 ( .A(n4525), .B(n4564), .C(n193), .Y(n2314) );
  OAI21X1 U1662 ( .A(n4525), .B(n4563), .C(n257), .Y(n2315) );
  OAI21X1 U1664 ( .A(n4525), .B(n4562), .C(n321), .Y(n2316) );
  OAI21X1 U1666 ( .A(n4525), .B(n4561), .C(n2864), .Y(n2317) );
  OAI21X1 U1668 ( .A(n4525), .B(n4560), .C(n2931), .Y(n2318) );
  OAI21X1 U1670 ( .A(n4525), .B(n4559), .C(n2999), .Y(n2319) );
  OAI21X1 U1672 ( .A(n4525), .B(n4558), .C(n3066), .Y(n2320) );
  OAI21X1 U1674 ( .A(n4525), .B(n4557), .C(n2607), .Y(n2321) );
  OAI21X1 U1676 ( .A(n4525), .B(n4556), .C(n2671), .Y(n2322) );
  OAI21X1 U1678 ( .A(n4525), .B(n4555), .C(n2735), .Y(n2323) );
  OAI21X1 U1680 ( .A(n4525), .B(n4554), .C(n2800), .Y(n2324) );
  OAI21X1 U1682 ( .A(n4525), .B(n4553), .C(n128), .Y(n2325) );
  OAI21X1 U1684 ( .A(n4525), .B(n4552), .C(n192), .Y(n2326) );
  OAI21X1 U1686 ( .A(n4525), .B(n4551), .C(n256), .Y(n2327) );
  OAI21X1 U1688 ( .A(n4525), .B(n4550), .C(n320), .Y(n2328) );
  OAI21X1 U1690 ( .A(n4525), .B(n4549), .C(n51), .Y(n2329) );
  OAI21X1 U1692 ( .A(n3117), .B(n3319), .C(reset), .Y(n1207) );
  NAND3X1 U1693 ( .A(n1481), .B(n4623), .C(wr_ptr[4]), .Y(n969) );
  OAI21X1 U1694 ( .A(n4524), .B(n4581), .C(n3065), .Y(n2330) );
  OAI21X1 U1696 ( .A(n4524), .B(n4580), .C(n2998), .Y(n2331) );
  OAI21X1 U1698 ( .A(n4524), .B(n4579), .C(n2930), .Y(n2332) );
  OAI21X1 U1700 ( .A(n4524), .B(n4578), .C(n2863), .Y(n2333) );
  OAI21X1 U1702 ( .A(n4524), .B(n4577), .C(n2862), .Y(n2334) );
  OAI21X1 U1704 ( .A(n4524), .B(n4576), .C(n3064), .Y(n2335) );
  OAI21X1 U1706 ( .A(n4524), .B(n4575), .C(n2997), .Y(n2336) );
  OAI21X1 U1708 ( .A(n4524), .B(n4574), .C(n3335), .Y(n2337) );
  OAI21X1 U1710 ( .A(n4524), .B(n4573), .C(n2929), .Y(n2338) );
  OAI21X1 U1712 ( .A(n4524), .B(n4572), .C(n3269), .Y(n2339) );
  OAI21X1 U1714 ( .A(n4524), .B(n4571), .C(n3203), .Y(n2340) );
  OAI21X1 U1716 ( .A(n4524), .B(n4570), .C(n3136), .Y(n2341) );
  OAI21X1 U1718 ( .A(n4524), .B(n4569), .C(n319), .Y(n2342) );
  OAI21X1 U1720 ( .A(n4524), .B(n4568), .C(n255), .Y(n2343) );
  OAI21X1 U1722 ( .A(n4524), .B(n4567), .C(n191), .Y(n2344) );
  OAI21X1 U1724 ( .A(n4524), .B(n4566), .C(n127), .Y(n2345) );
  OAI21X1 U1726 ( .A(n4524), .B(n4565), .C(n2799), .Y(n2346) );
  OAI21X1 U1728 ( .A(n4524), .B(n4564), .C(n2734), .Y(n2347) );
  OAI21X1 U1730 ( .A(n4524), .B(n4563), .C(n2670), .Y(n2348) );
  OAI21X1 U1732 ( .A(n4524), .B(n4562), .C(n2606), .Y(n2349) );
  OAI21X1 U1734 ( .A(n4524), .B(n4561), .C(n3334), .Y(n2350) );
  OAI21X1 U1736 ( .A(n4524), .B(n4560), .C(n3268), .Y(n2351) );
  OAI21X1 U1738 ( .A(n4524), .B(n4559), .C(n3202), .Y(n2352) );
  OAI21X1 U1740 ( .A(n4524), .B(n4558), .C(n3135), .Y(n2353) );
  OAI21X1 U1742 ( .A(n4524), .B(n4557), .C(n318), .Y(n2354) );
  OAI21X1 U1744 ( .A(n4524), .B(n4556), .C(n254), .Y(n2355) );
  OAI21X1 U1746 ( .A(n4524), .B(n4555), .C(n190), .Y(n2356) );
  OAI21X1 U1748 ( .A(n4524), .B(n4554), .C(n126), .Y(n2357) );
  OAI21X1 U1750 ( .A(n4524), .B(n4553), .C(n2798), .Y(n2358) );
  OAI21X1 U1752 ( .A(n4524), .B(n4552), .C(n2733), .Y(n2359) );
  OAI21X1 U1754 ( .A(n4524), .B(n4551), .C(n2669), .Y(n2360) );
  OAI21X1 U1756 ( .A(n4524), .B(n4550), .C(n2605), .Y(n2361) );
  OAI21X1 U1758 ( .A(n4524), .B(n4549), .C(n50), .Y(n2362) );
  OAI21X1 U1760 ( .A(n3118), .B(n3252), .C(reset), .Y(n1241) );
  NAND3X1 U1761 ( .A(n4621), .B(n4622), .C(n4619), .Y(n416) );
  OAI21X1 U1762 ( .A(n4523), .B(n4581), .C(n2996), .Y(n2363) );
  OAI21X1 U1764 ( .A(n4523), .B(n4580), .C(n3063), .Y(n2364) );
  OAI21X1 U1766 ( .A(n4523), .B(n4579), .C(n2861), .Y(n2365) );
  OAI21X1 U1768 ( .A(n4523), .B(n4578), .C(n2928), .Y(n2366) );
  OAI21X1 U1770 ( .A(n4523), .B(n4577), .C(n2927), .Y(n2367) );
  OAI21X1 U1772 ( .A(n4523), .B(n4576), .C(n2995), .Y(n2368) );
  OAI21X1 U1774 ( .A(n4523), .B(n4575), .C(n3062), .Y(n2369) );
  OAI21X1 U1776 ( .A(n4523), .B(n4574), .C(n3267), .Y(n2370) );
  OAI21X1 U1778 ( .A(n4523), .B(n4573), .C(n2860), .Y(n2371) );
  OAI21X1 U1780 ( .A(n4523), .B(n4572), .C(n3333), .Y(n2372) );
  OAI21X1 U1782 ( .A(n4523), .B(n4571), .C(n3134), .Y(n2373) );
  OAI21X1 U1784 ( .A(n4523), .B(n4570), .C(n3201), .Y(n2374) );
  OAI21X1 U1786 ( .A(n4523), .B(n4569), .C(n253), .Y(n2375) );
  OAI21X1 U1788 ( .A(n4523), .B(n4568), .C(n317), .Y(n2376) );
  OAI21X1 U1790 ( .A(n4523), .B(n4567), .C(n125), .Y(n2377) );
  OAI21X1 U1792 ( .A(n4523), .B(n4566), .C(n189), .Y(n2378) );
  OAI21X1 U1794 ( .A(n4523), .B(n4565), .C(n2732), .Y(n2379) );
  OAI21X1 U1796 ( .A(n4523), .B(n4564), .C(n2797), .Y(n2380) );
  OAI21X1 U1798 ( .A(n4523), .B(n4563), .C(n2604), .Y(n2381) );
  OAI21X1 U1800 ( .A(n4523), .B(n4562), .C(n2668), .Y(n2382) );
  OAI21X1 U1802 ( .A(n4523), .B(n4561), .C(n3266), .Y(n2383) );
  OAI21X1 U1804 ( .A(n4523), .B(n4560), .C(n3332), .Y(n2384) );
  OAI21X1 U1806 ( .A(n4523), .B(n4559), .C(n3133), .Y(n2385) );
  OAI21X1 U1808 ( .A(n4523), .B(n4558), .C(n3200), .Y(n2386) );
  OAI21X1 U1810 ( .A(n4523), .B(n4557), .C(n252), .Y(n2387) );
  OAI21X1 U1812 ( .A(n4523), .B(n4556), .C(n316), .Y(n2388) );
  OAI21X1 U1814 ( .A(n4523), .B(n4555), .C(n124), .Y(n2389) );
  OAI21X1 U1816 ( .A(n4523), .B(n4554), .C(n188), .Y(n2390) );
  OAI21X1 U1818 ( .A(n4523), .B(n4553), .C(n2731), .Y(n2391) );
  OAI21X1 U1820 ( .A(n4523), .B(n4552), .C(n2796), .Y(n2392) );
  OAI21X1 U1822 ( .A(n4523), .B(n4551), .C(n412), .Y(n2393) );
  OAI21X1 U1824 ( .A(n4523), .B(n4550), .C(n2667), .Y(n2394) );
  OAI21X1 U1826 ( .A(n4523), .B(n4549), .C(n49), .Y(n2395) );
  OAI21X1 U1828 ( .A(n3048), .B(n3252), .C(reset), .Y(n1276) );
  NAND3X1 U1829 ( .A(n4621), .B(n4622), .C(wr_ptr[0]), .Y(n451) );
  OAI21X1 U1830 ( .A(n4522), .B(n4581), .C(n2926), .Y(n2396) );
  OAI21X1 U1832 ( .A(n4522), .B(n4580), .C(n2859), .Y(n2397) );
  OAI21X1 U1834 ( .A(n4522), .B(n4579), .C(n3061), .Y(n2398) );
  OAI21X1 U1836 ( .A(n4522), .B(n4578), .C(n2994), .Y(n2399) );
  OAI21X1 U1838 ( .A(n4522), .B(n4577), .C(n2993), .Y(n2400) );
  OAI21X1 U1840 ( .A(n4522), .B(n4576), .C(n2925), .Y(n2401) );
  OAI21X1 U1842 ( .A(n4522), .B(n4575), .C(n2858), .Y(n2402) );
  OAI21X1 U1844 ( .A(n4522), .B(n4574), .C(n3199), .Y(n2403) );
  OAI21X1 U1846 ( .A(n4522), .B(n4573), .C(n3060), .Y(n2404) );
  OAI21X1 U1848 ( .A(n4522), .B(n4572), .C(n3132), .Y(n2405) );
  OAI21X1 U1850 ( .A(n4522), .B(n4571), .C(n3331), .Y(n2406) );
  OAI21X1 U1852 ( .A(n4522), .B(n4570), .C(n3265), .Y(n2407) );
  OAI21X1 U1854 ( .A(n4522), .B(n4569), .C(n187), .Y(n2408) );
  OAI21X1 U1856 ( .A(n4522), .B(n4568), .C(n123), .Y(n2409) );
  OAI21X1 U1858 ( .A(n4522), .B(n4567), .C(n315), .Y(n2410) );
  OAI21X1 U1860 ( .A(n4522), .B(n4566), .C(n251), .Y(n2411) );
  OAI21X1 U1862 ( .A(n4522), .B(n4565), .C(n2666), .Y(n2412) );
  OAI21X1 U1864 ( .A(n4522), .B(n4564), .C(n410), .Y(n2413) );
  OAI21X1 U1866 ( .A(n4522), .B(n4563), .C(n2795), .Y(n2414) );
  OAI21X1 U1868 ( .A(n4522), .B(n4562), .C(n2730), .Y(n2415) );
  OAI21X1 U1870 ( .A(n4522), .B(n4561), .C(n3198), .Y(n2416) );
  OAI21X1 U1872 ( .A(n4522), .B(n4560), .C(n3131), .Y(n2417) );
  OAI21X1 U1874 ( .A(n4522), .B(n4559), .C(n3330), .Y(n2418) );
  OAI21X1 U1876 ( .A(n4522), .B(n4558), .C(n3264), .Y(n2419) );
  OAI21X1 U1878 ( .A(n4522), .B(n4557), .C(n186), .Y(n2420) );
  OAI21X1 U1880 ( .A(n4522), .B(n4556), .C(n122), .Y(n2421) );
  OAI21X1 U1882 ( .A(n4522), .B(n4555), .C(n314), .Y(n2422) );
  OAI21X1 U1884 ( .A(n4522), .B(n4554), .C(n250), .Y(n2423) );
  OAI21X1 U1886 ( .A(n4522), .B(n4553), .C(n2665), .Y(n2424) );
  OAI21X1 U1888 ( .A(n4522), .B(n4552), .C(n408), .Y(n2425) );
  OAI21X1 U1890 ( .A(n4522), .B(n4551), .C(n2794), .Y(n2426) );
  OAI21X1 U1892 ( .A(n4522), .B(n4550), .C(n2729), .Y(n2427) );
  OAI21X1 U1894 ( .A(n4522), .B(n4549), .C(n48), .Y(n2428) );
  OAI21X1 U1896 ( .A(n2980), .B(n3252), .C(reset), .Y(n1310) );
  NAND3X1 U1897 ( .A(n4619), .B(n4622), .C(wr_ptr[1]), .Y(n486) );
  OAI21X1 U1898 ( .A(n4521), .B(n4581), .C(n2857), .Y(n2429) );
  OAI21X1 U1900 ( .A(n4521), .B(n4580), .C(n2924), .Y(n2430) );
  OAI21X1 U1902 ( .A(n4521), .B(n4579), .C(n2992), .Y(n2431) );
  OAI21X1 U1904 ( .A(n4521), .B(n4578), .C(n3059), .Y(n2432) );
  OAI21X1 U1906 ( .A(n4521), .B(n4577), .C(n3058), .Y(n2433) );
  OAI21X1 U1908 ( .A(n4521), .B(n4576), .C(n2856), .Y(n2434) );
  OAI21X1 U1910 ( .A(n4521), .B(n4575), .C(n2923), .Y(n2435) );
  OAI21X1 U1912 ( .A(n4521), .B(n4574), .C(n3130), .Y(n2436) );
  OAI21X1 U1914 ( .A(n4521), .B(n4573), .C(n2991), .Y(n2437) );
  OAI21X1 U1916 ( .A(n4521), .B(n4572), .C(n3197), .Y(n2438) );
  OAI21X1 U1918 ( .A(n4521), .B(n4571), .C(n3263), .Y(n2439) );
  OAI21X1 U1920 ( .A(n4521), .B(n4570), .C(n3329), .Y(n2440) );
  OAI21X1 U1922 ( .A(n4521), .B(n4569), .C(n121), .Y(n2441) );
  OAI21X1 U1924 ( .A(n4521), .B(n4568), .C(n185), .Y(n2442) );
  OAI21X1 U1926 ( .A(n4521), .B(n4567), .C(n249), .Y(n2443) );
  OAI21X1 U1928 ( .A(n4521), .B(n4566), .C(n313), .Y(n2444) );
  OAI21X1 U1930 ( .A(n4521), .B(n4565), .C(n406), .Y(n2445) );
  OAI21X1 U1932 ( .A(n4521), .B(n4564), .C(n2664), .Y(n2446) );
  OAI21X1 U1934 ( .A(n4521), .B(n4563), .C(n2728), .Y(n2447) );
  OAI21X1 U1936 ( .A(n4521), .B(n4562), .C(n2793), .Y(n2448) );
  OAI21X1 U1938 ( .A(n4521), .B(n4561), .C(n3129), .Y(n2449) );
  OAI21X1 U1940 ( .A(n4521), .B(n4560), .C(n3196), .Y(n2450) );
  OAI21X1 U1942 ( .A(n4521), .B(n4559), .C(n3262), .Y(n2451) );
  OAI21X1 U1944 ( .A(n4521), .B(n4558), .C(n3328), .Y(n2452) );
  OAI21X1 U1946 ( .A(n4521), .B(n4557), .C(n120), .Y(n2453) );
  OAI21X1 U1948 ( .A(n4521), .B(n4556), .C(n184), .Y(n2454) );
  OAI21X1 U1950 ( .A(n4521), .B(n4555), .C(n248), .Y(n2455) );
  OAI21X1 U1952 ( .A(n4521), .B(n4554), .C(n312), .Y(n2456) );
  OAI21X1 U1954 ( .A(n4521), .B(n4553), .C(n404), .Y(n2457) );
  OAI21X1 U1956 ( .A(n4521), .B(n4552), .C(n2663), .Y(n2458) );
  OAI21X1 U1958 ( .A(n4521), .B(n4551), .C(n2727), .Y(n2459) );
  OAI21X1 U1960 ( .A(n4521), .B(n4550), .C(n2792), .Y(n2460) );
  OAI21X1 U1962 ( .A(n4521), .B(n4549), .C(n47), .Y(n2461) );
  OAI21X1 U1964 ( .A(n2913), .B(n3252), .C(reset), .Y(n1344) );
  NAND3X1 U1965 ( .A(wr_ptr[0]), .B(n4622), .C(wr_ptr[1]), .Y(n521) );
  OAI21X1 U1966 ( .A(n4520), .B(n4581), .C(n2791), .Y(n2462) );
  OAI21X1 U1968 ( .A(n4520), .B(n4580), .C(n2726), .Y(n2463) );
  OAI21X1 U1970 ( .A(n4520), .B(n4579), .C(n2662), .Y(n2464) );
  OAI21X1 U1972 ( .A(n4520), .B(n4578), .C(n402), .Y(n2465) );
  OAI21X1 U1974 ( .A(n4520), .B(n4577), .C(n400), .Y(n2466) );
  OAI21X1 U1976 ( .A(n4520), .B(n4576), .C(n2790), .Y(n2467) );
  OAI21X1 U1978 ( .A(n4520), .B(n4575), .C(n2725), .Y(n2468) );
  OAI21X1 U1980 ( .A(n4520), .B(n4574), .C(n311), .Y(n2469) );
  OAI21X1 U1982 ( .A(n4520), .B(n4573), .C(n2661), .Y(n2470) );
  OAI21X1 U1984 ( .A(n4520), .B(n4572), .C(n247), .Y(n2471) );
  OAI21X1 U1986 ( .A(n4520), .B(n4571), .C(n183), .Y(n2472) );
  OAI21X1 U1988 ( .A(n4520), .B(n4570), .C(n119), .Y(n2473) );
  OAI21X1 U1990 ( .A(n4520), .B(n4569), .C(n3327), .Y(n2474) );
  OAI21X1 U1992 ( .A(n4520), .B(n4568), .C(n3261), .Y(n2475) );
  OAI21X1 U1994 ( .A(n4520), .B(n4567), .C(n3195), .Y(n2476) );
  OAI21X1 U1996 ( .A(n4520), .B(n4566), .C(n3128), .Y(n2477) );
  OAI21X1 U1998 ( .A(n4520), .B(n4565), .C(n3057), .Y(n2478) );
  OAI21X1 U2000 ( .A(n4520), .B(n4564), .C(n2990), .Y(n2479) );
  OAI21X1 U2002 ( .A(n4520), .B(n4563), .C(n2922), .Y(n2480) );
  OAI21X1 U2004 ( .A(n4520), .B(n4562), .C(n2855), .Y(n2481) );
  OAI21X1 U2006 ( .A(n4520), .B(n4561), .C(n310), .Y(n2482) );
  OAI21X1 U2008 ( .A(n4520), .B(n4560), .C(n246), .Y(n2483) );
  OAI21X1 U2010 ( .A(n4520), .B(n4559), .C(n182), .Y(n2484) );
  OAI21X1 U2012 ( .A(n4520), .B(n4558), .C(n118), .Y(n2485) );
  OAI21X1 U2014 ( .A(n4520), .B(n4557), .C(n3326), .Y(n2486) );
  OAI21X1 U2016 ( .A(n4520), .B(n4556), .C(n3260), .Y(n2487) );
  OAI21X1 U2018 ( .A(n4520), .B(n4555), .C(n3194), .Y(n2488) );
  OAI21X1 U2020 ( .A(n4520), .B(n4554), .C(n3127), .Y(n2489) );
  OAI21X1 U2022 ( .A(n4520), .B(n4553), .C(n3056), .Y(n2490) );
  OAI21X1 U2024 ( .A(n4520), .B(n4552), .C(n2989), .Y(n2491) );
  OAI21X1 U2026 ( .A(n4520), .B(n4551), .C(n2921), .Y(n2492) );
  OAI21X1 U2028 ( .A(n4520), .B(n4550), .C(n2854), .Y(n2493) );
  OAI21X1 U2030 ( .A(n4520), .B(n4549), .C(n46), .Y(n2494) );
  OAI21X1 U2032 ( .A(n2912), .B(n3252), .C(reset), .Y(n1378) );
  NAND3X1 U2033 ( .A(n4619), .B(n4621), .C(wr_ptr[2]), .Y(n556) );
  OAI21X1 U2034 ( .A(n4519), .B(n4581), .C(n2724), .Y(n2495) );
  OAI21X1 U2036 ( .A(n4519), .B(n4580), .C(n2789), .Y(n2496) );
  OAI21X1 U2038 ( .A(n4519), .B(n4579), .C(n398), .Y(n2497) );
  OAI21X1 U2040 ( .A(n4519), .B(n4578), .C(n2660), .Y(n2498) );
  OAI21X1 U2042 ( .A(n4519), .B(n4577), .C(n2659), .Y(n2499) );
  OAI21X1 U2044 ( .A(n4519), .B(n4576), .C(n2723), .Y(n2500) );
  OAI21X1 U2046 ( .A(n4519), .B(n4575), .C(n2788), .Y(n2501) );
  OAI21X1 U2048 ( .A(n4519), .B(n4574), .C(n245), .Y(n2502) );
  OAI21X1 U2050 ( .A(n4519), .B(n4573), .C(n396), .Y(n2503) );
  OAI21X1 U2052 ( .A(n4519), .B(n4572), .C(n309), .Y(n2504) );
  OAI21X1 U2054 ( .A(n4519), .B(n4571), .C(n117), .Y(n2505) );
  OAI21X1 U2056 ( .A(n4519), .B(n4570), .C(n181), .Y(n2506) );
  OAI21X1 U2058 ( .A(n4519), .B(n4569), .C(n3259), .Y(n2507) );
  OAI21X1 U2060 ( .A(n4519), .B(n4568), .C(n3325), .Y(n2508) );
  OAI21X1 U2062 ( .A(n4519), .B(n4567), .C(n3126), .Y(n2509) );
  OAI21X1 U2064 ( .A(n4519), .B(n4566), .C(n3193), .Y(n2510) );
  OAI21X1 U2066 ( .A(n4519), .B(n4565), .C(n2988), .Y(n2511) );
  OAI21X1 U2068 ( .A(n4519), .B(n4564), .C(n3055), .Y(n2512) );
  OAI21X1 U2070 ( .A(n4519), .B(n4563), .C(n2853), .Y(n2513) );
  OAI21X1 U2072 ( .A(n4519), .B(n4562), .C(n2920), .Y(n2514) );
  OAI21X1 U2074 ( .A(n4519), .B(n4561), .C(n244), .Y(n2515) );
  OAI21X1 U2076 ( .A(n4519), .B(n4560), .C(n308), .Y(n2516) );
  OAI21X1 U2078 ( .A(n4519), .B(n4559), .C(n116), .Y(n2517) );
  OAI21X1 U2080 ( .A(n4519), .B(n4558), .C(n180), .Y(n2518) );
  OAI21X1 U2082 ( .A(n4519), .B(n4557), .C(n3258), .Y(n2519) );
  OAI21X1 U2084 ( .A(n4519), .B(n4556), .C(n3324), .Y(n2520) );
  OAI21X1 U2086 ( .A(n4519), .B(n4555), .C(n3125), .Y(n2521) );
  OAI21X1 U2088 ( .A(n4519), .B(n4554), .C(n3192), .Y(n2522) );
  OAI21X1 U2090 ( .A(n4519), .B(n4553), .C(n2987), .Y(n2523) );
  OAI21X1 U2092 ( .A(n4519), .B(n4552), .C(n3054), .Y(n2524) );
  OAI21X1 U2094 ( .A(n4519), .B(n4551), .C(n2852), .Y(n2525) );
  OAI21X1 U2096 ( .A(n4519), .B(n4550), .C(n2919), .Y(n2526) );
  OAI21X1 U2098 ( .A(n4519), .B(n4549), .C(n45), .Y(n2527) );
  OAI21X1 U2100 ( .A(n2979), .B(n3252), .C(reset), .Y(n1412) );
  NAND3X1 U2101 ( .A(wr_ptr[0]), .B(n4621), .C(wr_ptr[2]), .Y(n591) );
  OAI21X1 U2102 ( .A(n4518), .B(n4581), .C(n2658), .Y(n2528) );
  OAI21X1 U2104 ( .A(n4518), .B(n4580), .C(n394), .Y(n2529) );
  OAI21X1 U2106 ( .A(n4518), .B(n4579), .C(n2787), .Y(n2530) );
  OAI21X1 U2108 ( .A(n4518), .B(n4578), .C(n2722), .Y(n2531) );
  OAI21X1 U2110 ( .A(n4518), .B(n4577), .C(n2721), .Y(n2532) );
  OAI21X1 U2112 ( .A(n4518), .B(n4576), .C(n2657), .Y(n2533) );
  OAI21X1 U2114 ( .A(n4518), .B(n4575), .C(n392), .Y(n2534) );
  OAI21X1 U2116 ( .A(n4518), .B(n4574), .C(n179), .Y(n2535) );
  OAI21X1 U2118 ( .A(n4518), .B(n4573), .C(n2786), .Y(n2536) );
  OAI21X1 U2120 ( .A(n4518), .B(n4572), .C(n115), .Y(n2537) );
  OAI21X1 U2122 ( .A(n4518), .B(n4571), .C(n307), .Y(n2538) );
  OAI21X1 U2124 ( .A(n4518), .B(n4570), .C(n243), .Y(n2539) );
  OAI21X1 U2126 ( .A(n4518), .B(n4569), .C(n3191), .Y(n2540) );
  OAI21X1 U2128 ( .A(n4518), .B(n4568), .C(n3124), .Y(n2541) );
  OAI21X1 U2130 ( .A(n4518), .B(n4567), .C(n3323), .Y(n2542) );
  OAI21X1 U2132 ( .A(n4518), .B(n4566), .C(n3257), .Y(n2543) );
  OAI21X1 U2134 ( .A(n4518), .B(n4565), .C(n2918), .Y(n2544) );
  OAI21X1 U2136 ( .A(n4518), .B(n4564), .C(n2851), .Y(n2545) );
  OAI21X1 U2138 ( .A(n4518), .B(n4563), .C(n3053), .Y(n2546) );
  OAI21X1 U2140 ( .A(n4518), .B(n4562), .C(n2986), .Y(n2547) );
  OAI21X1 U2142 ( .A(n4518), .B(n4561), .C(n178), .Y(n2548) );
  OAI21X1 U2144 ( .A(n4518), .B(n4560), .C(n114), .Y(n2549) );
  OAI21X1 U2146 ( .A(n4518), .B(n4559), .C(n306), .Y(n2550) );
  OAI21X1 U2148 ( .A(n4518), .B(n4558), .C(n242), .Y(n2551) );
  OAI21X1 U2150 ( .A(n4518), .B(n4557), .C(n3190), .Y(n2552) );
  OAI21X1 U2152 ( .A(n4518), .B(n4556), .C(n3123), .Y(n2553) );
  OAI21X1 U2154 ( .A(n4518), .B(n4555), .C(n3322), .Y(n2554) );
  OAI21X1 U2156 ( .A(n4518), .B(n4554), .C(n3256), .Y(n2555) );
  OAI21X1 U2158 ( .A(n4518), .B(n4553), .C(n2917), .Y(n2556) );
  OAI21X1 U2160 ( .A(n4518), .B(n4552), .C(n2850), .Y(n2557) );
  OAI21X1 U2162 ( .A(n4518), .B(n4551), .C(n3052), .Y(n2558) );
  OAI21X1 U2164 ( .A(n4518), .B(n4550), .C(n2985), .Y(n2559) );
  OAI21X1 U2166 ( .A(n4518), .B(n4549), .C(n44), .Y(n2560) );
  OAI21X1 U2168 ( .A(n3047), .B(n3252), .C(reset), .Y(n1446) );
  NAND3X1 U2169 ( .A(wr_ptr[1]), .B(n4619), .C(wr_ptr[2]), .Y(n626) );
  OAI21X1 U2170 ( .A(n4517), .B(n4581), .C(n390), .Y(n2561) );
  OAI21X1 U2173 ( .A(n4517), .B(n4580), .C(n2656), .Y(n2562) );
  OAI21X1 U2176 ( .A(n4517), .B(n4579), .C(n2720), .Y(n2563) );
  OAI21X1 U2179 ( .A(n4517), .B(n4578), .C(n2785), .Y(n2564) );
  OAI21X1 U2182 ( .A(n4517), .B(n4577), .C(n2784), .Y(n2565) );
  OAI21X1 U2185 ( .A(n4517), .B(n4576), .C(n388), .Y(n2566) );
  OAI21X1 U2188 ( .A(n4517), .B(n4575), .C(n2655), .Y(n2567) );
  OAI21X1 U2191 ( .A(n4517), .B(n4574), .C(n113), .Y(n2568) );
  OAI21X1 U2194 ( .A(n4517), .B(n4573), .C(n2719), .Y(n2569) );
  OAI21X1 U2197 ( .A(n4517), .B(n4572), .C(n177), .Y(n2570) );
  OAI21X1 U2200 ( .A(n4517), .B(n4571), .C(n241), .Y(n2571) );
  OAI21X1 U2203 ( .A(n4517), .B(n4570), .C(n305), .Y(n2572) );
  OAI21X1 U2206 ( .A(n4517), .B(n4569), .C(n3122), .Y(n2573) );
  OAI21X1 U2209 ( .A(n4517), .B(n4568), .C(n3189), .Y(n2574) );
  OAI21X1 U2212 ( .A(n4517), .B(n4567), .C(n3255), .Y(n2575) );
  OAI21X1 U2215 ( .A(n4517), .B(n4566), .C(n3321), .Y(n2576) );
  OAI21X1 U2218 ( .A(n4517), .B(n4565), .C(n2849), .Y(n2577) );
  OAI21X1 U2221 ( .A(n4517), .B(n4564), .C(n2916), .Y(n2578) );
  OAI21X1 U2224 ( .A(n4517), .B(n4563), .C(n2984), .Y(n2579) );
  OAI21X1 U2227 ( .A(n4517), .B(n4562), .C(n3051), .Y(n2580) );
  OAI21X1 U2230 ( .A(n4517), .B(n4561), .C(n112), .Y(n2581) );
  OAI21X1 U2233 ( .A(n4517), .B(n4560), .C(n176), .Y(n2582) );
  OAI21X1 U2236 ( .A(n4517), .B(n4559), .C(n240), .Y(n2583) );
  OAI21X1 U2239 ( .A(n4517), .B(n4558), .C(n304), .Y(n2584) );
  OAI21X1 U2242 ( .A(n4517), .B(n4557), .C(n3121), .Y(n2585) );
  OAI21X1 U2245 ( .A(n4517), .B(n4556), .C(n3188), .Y(n2586) );
  OAI21X1 U2248 ( .A(n4517), .B(n4555), .C(n3254), .Y(n2587) );
  OAI21X1 U2251 ( .A(n4517), .B(n4554), .C(n3320), .Y(n2588) );
  OAI21X1 U2254 ( .A(n4517), .B(n4553), .C(n2848), .Y(n2589) );
  OAI21X1 U2257 ( .A(n4517), .B(n4552), .C(n2915), .Y(n2590) );
  OAI21X1 U2260 ( .A(n4517), .B(n4551), .C(n2983), .Y(n2591) );
  OAI21X1 U2263 ( .A(n4517), .B(n4550), .C(n3050), .Y(n2592) );
  OAI21X1 U2266 ( .A(n4517), .B(n4549), .C(n43), .Y(n2593) );
  OAI21X1 U2269 ( .A(n3117), .B(n3252), .C(reset), .Y(n1480) );
  NAND3X1 U2270 ( .A(wr_ptr[3]), .B(n1481), .C(wr_ptr[4]), .Y(n1242) );
  NAND3X1 U2271 ( .A(wr_ptr[1]), .B(wr_ptr[0]), .C(wr_ptr[2]), .Y(n661) );
  OAI21X1 U2272 ( .A(n4623), .B(n3318), .C(n2982), .Y(n2594) );
  OAI21X1 U2274 ( .A(n4622), .B(n3318), .C(n3187), .Y(n2595) );
  OAI21X1 U2276 ( .A(n4621), .B(n3318), .C(n3120), .Y(n2596) );
  OAI21X1 U2278 ( .A(n4620), .B(n3318), .C(n2914), .Y(n2597) );
  OAI21X1 U2280 ( .A(n4583), .B(n3384), .C(n3253), .Y(n2598) );
  OAI21X1 U2282 ( .A(n4514), .B(n3384), .C(n3186), .Y(n2599) );
  OAI21X1 U2284 ( .A(n4584), .B(n3384), .C(n3119), .Y(n2600) );
  OAI21X1 U2286 ( .A(n4585), .B(n3384), .C(n3049), .Y(n2601) );
  OAI21X1 U2288 ( .A(n4582), .B(n3384), .C(n2981), .Y(n2602) );
  AOI22X1 U2290 ( .A(n56), .B(n1490), .C(data_out[32]), .D(n1488), .Y(n1495)
         );
  AOI22X1 U2291 ( .A(n57), .B(n1490), .C(data_out[31]), .D(n1488), .Y(n1496)
         );
  AOI22X1 U2292 ( .A(n58), .B(n1490), .C(data_out[30]), .D(n1488), .Y(n1497)
         );
  AOI22X1 U2293 ( .A(n59), .B(n1490), .C(data_out[29]), .D(n1488), .Y(n1498)
         );
  AOI22X1 U2294 ( .A(n60), .B(n1490), .C(data_out[28]), .D(n1488), .Y(n1499)
         );
  AOI22X1 U2295 ( .A(n61), .B(n1490), .C(data_out[27]), .D(n1488), .Y(n1500)
         );
  AOI22X1 U2296 ( .A(n62), .B(n1490), .C(data_out[26]), .D(n1488), .Y(n1501)
         );
  AOI22X1 U2297 ( .A(n63), .B(n1490), .C(data_out[25]), .D(n1488), .Y(n1502)
         );
  AOI22X1 U2298 ( .A(n64), .B(n1490), .C(data_out[24]), .D(n1488), .Y(n1503)
         );
  AOI22X1 U2299 ( .A(n65), .B(n1490), .C(data_out[23]), .D(n1488), .Y(n1504)
         );
  AOI22X1 U2300 ( .A(n66), .B(n1490), .C(data_out[22]), .D(n1488), .Y(n1505)
         );
  AOI22X1 U2301 ( .A(n67), .B(n1490), .C(data_out[21]), .D(n1488), .Y(n1506)
         );
  AOI22X1 U2302 ( .A(n68), .B(n1490), .C(data_out[20]), .D(n1488), .Y(n1507)
         );
  AOI22X1 U2303 ( .A(n69), .B(n1490), .C(data_out[19]), .D(n1488), .Y(n1508)
         );
  AOI22X1 U2304 ( .A(n70), .B(n1490), .C(data_out[18]), .D(n1488), .Y(n1509)
         );
  AOI22X1 U2305 ( .A(n71), .B(n1490), .C(data_out[17]), .D(n1488), .Y(n1510)
         );
  AOI22X1 U2306 ( .A(n72), .B(n1490), .C(data_out[16]), .D(n1488), .Y(n1511)
         );
  AOI22X1 U2307 ( .A(n73), .B(n1490), .C(data_out[15]), .D(n1488), .Y(n1512)
         );
  AOI22X1 U2308 ( .A(n74), .B(n1490), .C(data_out[14]), .D(n1488), .Y(n1513)
         );
  AOI22X1 U2309 ( .A(n75), .B(n1490), .C(data_out[13]), .D(n1488), .Y(n1514)
         );
  AOI22X1 U2310 ( .A(n76), .B(n1490), .C(data_out[12]), .D(n1488), .Y(n1515)
         );
  AOI22X1 U2311 ( .A(n77), .B(n1490), .C(data_out[11]), .D(n1488), .Y(n1516)
         );
  AOI22X1 U2312 ( .A(n78), .B(n1490), .C(data_out[10]), .D(n1488), .Y(n1517)
         );
  AOI22X1 U2313 ( .A(n79), .B(n1490), .C(data_out[9]), .D(n1488), .Y(n1518) );
  AOI22X1 U2314 ( .A(n80), .B(n1490), .C(data_out[8]), .D(n1488), .Y(n1519) );
  AOI22X1 U2315 ( .A(n81), .B(n1490), .C(data_out[7]), .D(n1488), .Y(n1520) );
  AOI22X1 U2316 ( .A(n82), .B(n1490), .C(data_out[6]), .D(n1488), .Y(n1521) );
  AOI22X1 U2317 ( .A(n83), .B(n1490), .C(data_out[5]), .D(n1488), .Y(n1522) );
  AOI22X1 U2318 ( .A(n84), .B(n1490), .C(data_out[4]), .D(n1488), .Y(n1523) );
  AOI22X1 U2319 ( .A(n85), .B(n1490), .C(data_out[3]), .D(n1488), .Y(n1524) );
  AOI22X1 U2320 ( .A(n86), .B(n1490), .C(data_out[2]), .D(n1488), .Y(n1525) );
  AOI22X1 U2321 ( .A(n87), .B(n1490), .C(data_out[1]), .D(n1488), .Y(n1526) );
  AOI22X1 U2322 ( .A(n88), .B(n1490), .C(data_out[0]), .D(n1488), .Y(n1527) );
  OAI21X1 U2325 ( .A(n4619), .B(n3318), .C(n2783), .Y(n2603) );
  NAND3X1 U2329 ( .A(n3116), .B(fillcount[5]), .C(n1531), .Y(n4625) );
  NOR3X1 U2330 ( .A(fillcount[2]), .B(fillcount[4]), .C(fillcount[3]), .Y(
        n1531) );
  NAND3X1 U2332 ( .A(n1532), .B(n1533), .C(n1534), .Y(n4624) );
  NOR3X1 U2333 ( .A(n1535), .B(n1536), .C(n1537), .Y(n1534) );
  XNOR2X1 U2334 ( .A(n4622), .B(n14), .Y(n1537) );
  XNOR2X1 U2335 ( .A(n4623), .B(n15), .Y(n1536) );
  XNOR2X1 U2336 ( .A(n4619), .B(n4452), .Y(n1535) );
  XNOR2X1 U2337 ( .A(n4509), .B(wr_ptr[1]), .Y(n1533) );
  XNOR2X1 U2338 ( .A(n16), .B(wr_ptr[4]), .Y(n1532) );
  HAX1 add_57_U1_1_1 ( .A(n4502), .B(n4460), .YC(add_57_carry[2]), .YS(n90) );
  HAX1 add_57_U1_1_2 ( .A(n14), .B(add_57_carry[2]), .YC(add_57_carry[3]), 
        .YS(n91) );
  HAX1 add_57_U1_1_3 ( .A(n15), .B(add_57_carry[3]), .YC(add_57_carry[4]), 
        .YS(n92) );
  HAX1 add_51_U1_1_1 ( .A(wr_ptr[1]), .B(wr_ptr[0]), .YC(add_51_carry[2]), 
        .YS(n20) );
  HAX1 add_51_U1_1_2 ( .A(wr_ptr[2]), .B(add_51_carry[2]), .YC(add_51_carry[3]), .YS(n21) );
  HAX1 add_51_U1_1_3 ( .A(wr_ptr[3]), .B(add_51_carry[3]), .YC(add_51_carry[4]), .YS(n22) );
  FAX1 sub_93_U2_1 ( .A(wr_ptr[1]), .B(n4584), .C(sub_93_carry[1]), .YC(
        sub_93_carry[2]), .YS(fillcount[1]) );
  FAX1 sub_93_U2_2 ( .A(wr_ptr[2]), .B(n4514), .C(sub_93_carry[2]), .YC(
        sub_93_carry[3]), .YS(fillcount[2]) );
  FAX1 sub_93_U2_3 ( .A(wr_ptr[3]), .B(n4583), .C(sub_93_carry[3]), .YC(
        sub_93_carry[4]), .YS(fillcount[3]) );
  FAX1 sub_93_U2_4 ( .A(wr_ptr[4]), .B(n4582), .C(sub_93_carry[4]), .YC(
        sub_93_carry[5]), .YS(fillcount[4]) );
  AND2X1 U3 ( .A(reset), .B(n3114), .Y(n1482) );
  AND2X1 U4 ( .A(reset), .B(n3385), .Y(n1488) );
  AND2X1 U5 ( .A(reset), .B(n3384), .Y(n1490) );
  AND2X1 U6 ( .A(put), .B(full_bar), .Y(n1481) );
  BUFX2 U7 ( .A(n1527), .Y(n1) );
  BUFX2 U8 ( .A(n1526), .Y(n2) );
  BUFX2 U9 ( .A(n1525), .Y(n3) );
  BUFX2 U10 ( .A(n1524), .Y(n4) );
  BUFX2 U11 ( .A(n1523), .Y(n5) );
  BUFX2 U12 ( .A(n1522), .Y(n6) );
  BUFX2 U13 ( .A(n1521), .Y(n7) );
  BUFX2 U14 ( .A(n1520), .Y(n8) );
  BUFX2 U15 ( .A(n1519), .Y(n9) );
  BUFX2 U16 ( .A(n1518), .Y(n10) );
  BUFX2 U17 ( .A(n1517), .Y(n11) );
  BUFX2 U18 ( .A(n1516), .Y(n17) );
  BUFX2 U19 ( .A(n1515), .Y(n18) );
  BUFX2 U20 ( .A(n1514), .Y(n19) );
  BUFX2 U21 ( .A(n1513), .Y(n24) );
  BUFX2 U22 ( .A(n1512), .Y(n25) );
  BUFX2 U23 ( .A(n1511), .Y(n26) );
  BUFX2 U24 ( .A(n1510), .Y(n27) );
  BUFX2 U25 ( .A(n1509), .Y(n28) );
  BUFX2 U26 ( .A(n1508), .Y(n29) );
  BUFX2 U27 ( .A(n1507), .Y(n30) );
  BUFX2 U28 ( .A(n1506), .Y(n31) );
  BUFX2 U29 ( .A(n1505), .Y(n32) );
  BUFX2 U30 ( .A(n1504), .Y(n33) );
  BUFX2 U31 ( .A(n1503), .Y(n34) );
  BUFX2 U32 ( .A(n1502), .Y(n35) );
  BUFX2 U33 ( .A(n1501), .Y(n36) );
  BUFX2 U34 ( .A(n1500), .Y(n37) );
  BUFX2 U35 ( .A(n1499), .Y(n38) );
  BUFX2 U36 ( .A(n1498), .Y(n39) );
  BUFX2 U37 ( .A(n1497), .Y(n40) );
  BUFX2 U38 ( .A(n1496), .Y(n41) );
  BUFX2 U39 ( .A(n1495), .Y(n42) );
  AND2X1 U40 ( .A(mem[1055]), .B(n4517), .Y(n1479) );
  INVX1 U41 ( .A(n1479), .Y(n43) );
  AND2X1 U42 ( .A(mem[1022]), .B(n4518), .Y(n1445) );
  INVX1 U43 ( .A(n1445), .Y(n44) );
  AND2X1 U44 ( .A(mem[989]), .B(n4519), .Y(n1411) );
  INVX1 U45 ( .A(n1411), .Y(n45) );
  AND2X1 U46 ( .A(mem[956]), .B(n4520), .Y(n1377) );
  INVX1 U47 ( .A(n1377), .Y(n46) );
  AND2X1 U48 ( .A(mem[923]), .B(n4521), .Y(n1343) );
  INVX1 U49 ( .A(n1343), .Y(n47) );
  AND2X1 U50 ( .A(mem[890]), .B(n4522), .Y(n1309) );
  INVX1 U51 ( .A(n1309), .Y(n48) );
  AND2X1 U52 ( .A(mem[857]), .B(n4523), .Y(n1275) );
  INVX1 U53 ( .A(n1275), .Y(n49) );
  AND2X1 U54 ( .A(mem[824]), .B(n4524), .Y(n1240) );
  INVX1 U55 ( .A(n1240), .Y(n50) );
  AND2X1 U56 ( .A(mem[791]), .B(n4525), .Y(n1206) );
  INVX1 U57 ( .A(n1206), .Y(n51) );
  AND2X1 U58 ( .A(mem[758]), .B(n4526), .Y(n1172) );
  INVX1 U59 ( .A(n1172), .Y(n52) );
  AND2X1 U60 ( .A(mem[725]), .B(n4527), .Y(n1138) );
  INVX1 U61 ( .A(n1138), .Y(n53) );
  AND2X1 U62 ( .A(mem[692]), .B(n4528), .Y(n1104) );
  INVX1 U63 ( .A(n1104), .Y(n54) );
  AND2X1 U64 ( .A(mem[659]), .B(n4529), .Y(n1070) );
  INVX1 U65 ( .A(n1070), .Y(n55) );
  AND2X1 U66 ( .A(mem[626]), .B(n4530), .Y(n1036) );
  INVX1 U67 ( .A(n1036), .Y(n89) );
  AND2X1 U68 ( .A(mem[593]), .B(n4531), .Y(n1002) );
  INVX1 U69 ( .A(n1002), .Y(n94) );
  AND2X1 U70 ( .A(mem[560]), .B(n4532), .Y(n967) );
  INVX1 U71 ( .A(n967), .Y(n95) );
  AND2X1 U72 ( .A(mem[527]), .B(n4533), .Y(n933) );
  INVX1 U73 ( .A(n933), .Y(n96) );
  AND2X1 U74 ( .A(mem[494]), .B(n4534), .Y(n899) );
  INVX1 U75 ( .A(n899), .Y(n97) );
  AND2X1 U76 ( .A(mem[461]), .B(n4535), .Y(n865) );
  INVX1 U77 ( .A(n865), .Y(n98) );
  AND2X1 U78 ( .A(mem[428]), .B(n4536), .Y(n831) );
  INVX1 U79 ( .A(n831), .Y(n99) );
  AND2X1 U80 ( .A(mem[395]), .B(n4537), .Y(n797) );
  INVX1 U81 ( .A(n797), .Y(n100) );
  AND2X1 U82 ( .A(mem[362]), .B(n4538), .Y(n763) );
  INVX1 U84 ( .A(n763), .Y(n101) );
  AND2X1 U86 ( .A(mem[329]), .B(n4539), .Y(n729) );
  INVX1 U88 ( .A(n729), .Y(n102) );
  AND2X1 U90 ( .A(mem[296]), .B(n4540), .Y(n694) );
  INVX1 U92 ( .A(n694), .Y(n103) );
  AND2X1 U94 ( .A(mem[263]), .B(n4541), .Y(n659) );
  INVX1 U96 ( .A(n659), .Y(n104) );
  AND2X1 U98 ( .A(mem[230]), .B(n4542), .Y(n624) );
  INVX1 U100 ( .A(n624), .Y(n105) );
  AND2X1 U102 ( .A(mem[197]), .B(n4543), .Y(n589) );
  INVX1 U104 ( .A(n589), .Y(n106) );
  AND2X1 U106 ( .A(mem[164]), .B(n4544), .Y(n554) );
  INVX1 U108 ( .A(n554), .Y(n107) );
  AND2X1 U110 ( .A(mem[131]), .B(n4545), .Y(n519) );
  INVX1 U112 ( .A(n519), .Y(n108) );
  AND2X1 U114 ( .A(mem[98]), .B(n4546), .Y(n484) );
  INVX1 U116 ( .A(n484), .Y(n109) );
  AND2X1 U118 ( .A(mem[65]), .B(n4547), .Y(n449) );
  INVX1 U120 ( .A(n449), .Y(n110) );
  AND2X1 U122 ( .A(mem[32]), .B(n4548), .Y(n413) );
  INVX1 U124 ( .A(n413), .Y(n111) );
  AND2X1 U126 ( .A(mem[1043]), .B(n4517), .Y(n1467) );
  INVX1 U128 ( .A(n1467), .Y(n112) );
  AND2X1 U130 ( .A(mem[1030]), .B(n4517), .Y(n1454) );
  INVX1 U132 ( .A(n1454), .Y(n113) );
  AND2X1 U134 ( .A(mem[1011]), .B(n4518), .Y(n1434) );
  INVX1 U136 ( .A(n1434), .Y(n114) );
  AND2X1 U138 ( .A(mem[999]), .B(n4518), .Y(n1422) );
  INVX1 U140 ( .A(n1422), .Y(n115) );
  AND2X1 U142 ( .A(mem[979]), .B(n4519), .Y(n1401) );
  INVX1 U144 ( .A(n1401), .Y(n116) );
  AND2X1 U146 ( .A(mem[967]), .B(n4519), .Y(n1389) );
  INVX1 U148 ( .A(n1389), .Y(n117) );
  AND2X1 U151 ( .A(mem[947]), .B(n4520), .Y(n1368) );
  INVX1 U153 ( .A(n1368), .Y(n118) );
  AND2X1 U155 ( .A(mem[935]), .B(n4520), .Y(n1356) );
  INVX1 U157 ( .A(n1356), .Y(n119) );
  AND2X1 U159 ( .A(mem[915]), .B(n4521), .Y(n1335) );
  INVX1 U161 ( .A(n1335), .Y(n120) );
  AND2X1 U163 ( .A(mem[903]), .B(n4521), .Y(n1323) );
  INVX1 U165 ( .A(n1323), .Y(n121) );
  AND2X1 U167 ( .A(mem[883]), .B(n4522), .Y(n1302) );
  INVX1 U169 ( .A(n1302), .Y(n122) );
  AND2X1 U171 ( .A(mem[871]), .B(n4522), .Y(n1290) );
  INVX1 U173 ( .A(n1290), .Y(n123) );
  AND2X1 U175 ( .A(mem[851]), .B(n4523), .Y(n1269) );
  INVX1 U177 ( .A(n1269), .Y(n124) );
  AND2X1 U179 ( .A(mem[839]), .B(n4523), .Y(n1257) );
  INVX1 U181 ( .A(n1257), .Y(n125) );
  AND2X1 U183 ( .A(mem[819]), .B(n4524), .Y(n1235) );
  INVX1 U185 ( .A(n1235), .Y(n126) );
  AND2X1 U187 ( .A(mem[807]), .B(n4524), .Y(n1223) );
  INVX1 U189 ( .A(n1223), .Y(n127) );
  AND2X1 U191 ( .A(mem[787]), .B(n4525), .Y(n1202) );
  INVX1 U193 ( .A(n1202), .Y(n128) );
  AND2X1 U195 ( .A(mem[775]), .B(n4525), .Y(n1190) );
  INVX1 U197 ( .A(n1190), .Y(n129) );
  AND2X1 U199 ( .A(mem[755]), .B(n4526), .Y(n1169) );
  INVX1 U201 ( .A(n1169), .Y(n130) );
  AND2X1 U203 ( .A(mem[743]), .B(n4526), .Y(n1157) );
  INVX1 U205 ( .A(n1157), .Y(n131) );
  AND2X1 U207 ( .A(mem[723]), .B(n4527), .Y(n1136) );
  INVX1 U209 ( .A(n1136), .Y(n132) );
  AND2X1 U211 ( .A(mem[711]), .B(n4527), .Y(n1124) );
  INVX1 U213 ( .A(n1124), .Y(n133) );
  AND2X1 U215 ( .A(mem[691]), .B(n4528), .Y(n1103) );
  INVX1 U218 ( .A(n1103), .Y(n134) );
  AND2X1 U220 ( .A(mem[679]), .B(n4528), .Y(n1091) );
  INVX1 U222 ( .A(n1091), .Y(n135) );
  AND2X1 U224 ( .A(mem[647]), .B(n4529), .Y(n1058) );
  INVX1 U226 ( .A(n1058), .Y(n136) );
  AND2X1 U228 ( .A(mem[634]), .B(n4529), .Y(n1045) );
  INVX1 U230 ( .A(n1045), .Y(n137) );
  AND2X1 U232 ( .A(mem[615]), .B(n4530), .Y(n1025) );
  INVX1 U234 ( .A(n1025), .Y(n138) );
  AND2X1 U236 ( .A(mem[603]), .B(n4530), .Y(n1013) );
  INVX1 U238 ( .A(n1013), .Y(n139) );
  AND2X1 U240 ( .A(mem[583]), .B(n4531), .Y(n992) );
  INVX1 U242 ( .A(n992), .Y(n140) );
  AND2X1 U244 ( .A(mem[571]), .B(n4531), .Y(n980) );
  INVX1 U246 ( .A(n980), .Y(n141) );
  AND2X1 U248 ( .A(mem[551]), .B(n4532), .Y(n958) );
  INVX1 U250 ( .A(n958), .Y(n142) );
  AND2X1 U252 ( .A(mem[539]), .B(n4532), .Y(n946) );
  INVX1 U254 ( .A(n946), .Y(n143) );
  AND2X1 U256 ( .A(mem[519]), .B(n4533), .Y(n925) );
  INVX1 U258 ( .A(n925), .Y(n144) );
  AND2X1 U260 ( .A(mem[507]), .B(n4533), .Y(n913) );
  INVX1 U262 ( .A(n913), .Y(n145) );
  AND2X1 U264 ( .A(mem[487]), .B(n4534), .Y(n892) );
  INVX1 U266 ( .A(n892), .Y(n146) );
  AND2X1 U268 ( .A(mem[475]), .B(n4534), .Y(n880) );
  INVX1 U270 ( .A(n880), .Y(n147) );
  AND2X1 U272 ( .A(mem[455]), .B(n4535), .Y(n859) );
  INVX1 U274 ( .A(n859), .Y(n148) );
  AND2X1 U276 ( .A(mem[443]), .B(n4535), .Y(n847) );
  INVX1 U278 ( .A(n847), .Y(n149) );
  AND2X1 U280 ( .A(mem[423]), .B(n4536), .Y(n826) );
  INVX1 U282 ( .A(n826), .Y(n150) );
  AND2X1 U285 ( .A(mem[411]), .B(n4536), .Y(n814) );
  INVX1 U287 ( .A(n814), .Y(n151) );
  AND2X1 U289 ( .A(mem[391]), .B(n4537), .Y(n793) );
  INVX1 U291 ( .A(n793), .Y(n152) );
  AND2X1 U293 ( .A(mem[379]), .B(n4537), .Y(n781) );
  INVX1 U295 ( .A(n781), .Y(n153) );
  AND2X1 U297 ( .A(mem[359]), .B(n4538), .Y(n760) );
  INVX1 U299 ( .A(n760), .Y(n154) );
  AND2X1 U301 ( .A(mem[347]), .B(n4538), .Y(n748) );
  INVX1 U303 ( .A(n748), .Y(n155) );
  AND2X1 U305 ( .A(mem[327]), .B(n4539), .Y(n727) );
  INVX1 U307 ( .A(n727), .Y(n156) );
  AND2X1 U309 ( .A(mem[315]), .B(n4539), .Y(n715) );
  INVX1 U311 ( .A(n715), .Y(n157) );
  AND2X1 U313 ( .A(mem[295]), .B(n4540), .Y(n693) );
  INVX1 U315 ( .A(n693), .Y(n158) );
  AND2X1 U317 ( .A(mem[283]), .B(n4540), .Y(n681) );
  INVX1 U319 ( .A(n681), .Y(n159) );
  AND2X1 U321 ( .A(mem[255]), .B(n4541), .Y(n651) );
  INVX1 U323 ( .A(n651), .Y(n160) );
  AND2X1 U325 ( .A(mem[243]), .B(n4541), .Y(n639) );
  INVX1 U327 ( .A(n639), .Y(n161) );
  AND2X1 U329 ( .A(mem[223]), .B(n4542), .Y(n617) );
  INVX1 U331 ( .A(n617), .Y(n162) );
  AND2X1 U333 ( .A(mem[211]), .B(n4542), .Y(n605) );
  INVX1 U335 ( .A(n605), .Y(n163) );
  AND2X1 U337 ( .A(mem[191]), .B(n4543), .Y(n583) );
  INVX1 U339 ( .A(n583), .Y(n164) );
  AND2X1 U341 ( .A(mem[179]), .B(n4543), .Y(n571) );
  INVX1 U343 ( .A(n571), .Y(n165) );
  AND2X1 U345 ( .A(mem[159]), .B(n4544), .Y(n549) );
  INVX1 U347 ( .A(n549), .Y(n166) );
  AND2X1 U349 ( .A(mem[147]), .B(n4544), .Y(n537) );
  INVX1 U352 ( .A(n537), .Y(n167) );
  AND2X1 U354 ( .A(mem[127]), .B(n4545), .Y(n515) );
  INVX1 U356 ( .A(n515), .Y(n168) );
  AND2X1 U358 ( .A(mem[115]), .B(n4545), .Y(n503) );
  INVX1 U360 ( .A(n503), .Y(n169) );
  AND2X1 U362 ( .A(mem[95]), .B(n4546), .Y(n481) );
  INVX1 U364 ( .A(n481), .Y(n170) );
  AND2X1 U366 ( .A(mem[83]), .B(n4546), .Y(n469) );
  INVX1 U368 ( .A(n469), .Y(n171) );
  AND2X1 U370 ( .A(mem[63]), .B(n4547), .Y(n447) );
  INVX1 U372 ( .A(n447), .Y(n172) );
  AND2X1 U374 ( .A(mem[51]), .B(n4547), .Y(n435) );
  INVX1 U376 ( .A(n435), .Y(n173) );
  AND2X1 U378 ( .A(mem[31]), .B(n4548), .Y(n411) );
  INVX1 U380 ( .A(n411), .Y(n174) );
  AND2X1 U382 ( .A(mem[19]), .B(n4548), .Y(n387) );
  INVX1 U384 ( .A(n387), .Y(n175) );
  AND2X1 U386 ( .A(mem[1044]), .B(n4517), .Y(n1468) );
  INVX1 U388 ( .A(n1468), .Y(n176) );
  AND2X1 U390 ( .A(mem[1032]), .B(n4517), .Y(n1456) );
  INVX1 U392 ( .A(n1456), .Y(n177) );
  AND2X1 U394 ( .A(mem[1010]), .B(n4518), .Y(n1433) );
  INVX1 U396 ( .A(n1433), .Y(n178) );
  AND2X1 U398 ( .A(mem[997]), .B(n4518), .Y(n1420) );
  INVX1 U400 ( .A(n1420), .Y(n179) );
  AND2X1 U402 ( .A(mem[980]), .B(n4519), .Y(n1402) );
  INVX1 U404 ( .A(n1402), .Y(n180) );
  AND2X1 U406 ( .A(mem[968]), .B(n4519), .Y(n1390) );
  INVX1 U408 ( .A(n1390), .Y(n181) );
  AND2X1 U410 ( .A(mem[946]), .B(n4520), .Y(n1367) );
  INVX1 U412 ( .A(n1367), .Y(n182) );
  AND2X1 U414 ( .A(mem[934]), .B(n4520), .Y(n1355) );
  INVX1 U416 ( .A(n1355), .Y(n183) );
  AND2X1 U419 ( .A(mem[916]), .B(n4521), .Y(n1336) );
  INVX1 U421 ( .A(n1336), .Y(n184) );
  AND2X1 U423 ( .A(mem[904]), .B(n4521), .Y(n1324) );
  INVX1 U425 ( .A(n1324), .Y(n185) );
  AND2X1 U427 ( .A(mem[882]), .B(n4522), .Y(n1301) );
  INVX1 U429 ( .A(n1301), .Y(n186) );
  AND2X1 U431 ( .A(mem[870]), .B(n4522), .Y(n1289) );
  INVX1 U433 ( .A(n1289), .Y(n187) );
  AND2X1 U435 ( .A(mem[852]), .B(n4523), .Y(n1270) );
  INVX1 U437 ( .A(n1270), .Y(n188) );
  AND2X1 U439 ( .A(mem[840]), .B(n4523), .Y(n1258) );
  INVX1 U441 ( .A(n1258), .Y(n189) );
  AND2X1 U443 ( .A(mem[818]), .B(n4524), .Y(n1234) );
  INVX1 U445 ( .A(n1234), .Y(n190) );
  AND2X1 U447 ( .A(mem[806]), .B(n4524), .Y(n1222) );
  INVX1 U449 ( .A(n1222), .Y(n191) );
  AND2X1 U451 ( .A(mem[788]), .B(n4525), .Y(n1203) );
  INVX1 U453 ( .A(n1203), .Y(n192) );
  AND2X1 U455 ( .A(mem[776]), .B(n4525), .Y(n1191) );
  INVX1 U457 ( .A(n1191), .Y(n193) );
  AND2X1 U459 ( .A(mem[754]), .B(n4526), .Y(n1168) );
  INVX1 U461 ( .A(n1168), .Y(n194) );
  AND2X1 U463 ( .A(mem[742]), .B(n4526), .Y(n1156) );
  INVX1 U465 ( .A(n1156), .Y(n195) );
  AND2X1 U467 ( .A(mem[724]), .B(n4527), .Y(n1137) );
  INVX1 U469 ( .A(n1137), .Y(n196) );
  AND2X1 U471 ( .A(mem[712]), .B(n4527), .Y(n1125) );
  INVX1 U473 ( .A(n1125), .Y(n197) );
  AND2X1 U475 ( .A(mem[690]), .B(n4528), .Y(n1102) );
  INVX1 U477 ( .A(n1102), .Y(n198) );
  AND2X1 U479 ( .A(mem[678]), .B(n4528), .Y(n1090) );
  INVX1 U481 ( .A(n1090), .Y(n199) );
  AND2X1 U483 ( .A(mem[648]), .B(n4529), .Y(n1059) );
  INVX1 U486 ( .A(n1059), .Y(n200) );
  AND2X1 U488 ( .A(mem[636]), .B(n4529), .Y(n1047) );
  INVX1 U490 ( .A(n1047), .Y(n201) );
  AND2X1 U492 ( .A(mem[614]), .B(n4530), .Y(n1024) );
  INVX1 U494 ( .A(n1024), .Y(n202) );
  AND2X1 U496 ( .A(mem[601]), .B(n4530), .Y(n1011) );
  INVX1 U498 ( .A(n1011), .Y(n203) );
  AND2X1 U500 ( .A(mem[584]), .B(n4531), .Y(n993) );
  INVX1 U502 ( .A(n993), .Y(n204) );
  AND2X1 U504 ( .A(mem[572]), .B(n4531), .Y(n981) );
  INVX1 U506 ( .A(n981), .Y(n205) );
  AND2X1 U508 ( .A(mem[550]), .B(n4532), .Y(n957) );
  INVX1 U510 ( .A(n957), .Y(n206) );
  AND2X1 U512 ( .A(mem[538]), .B(n4532), .Y(n945) );
  INVX1 U514 ( .A(n945), .Y(n207) );
  AND2X1 U516 ( .A(mem[520]), .B(n4533), .Y(n926) );
  INVX1 U518 ( .A(n926), .Y(n208) );
  AND2X1 U520 ( .A(mem[508]), .B(n4533), .Y(n914) );
  INVX1 U522 ( .A(n914), .Y(n209) );
  AND2X1 U524 ( .A(mem[486]), .B(n4534), .Y(n891) );
  INVX1 U526 ( .A(n891), .Y(n210) );
  AND2X1 U528 ( .A(mem[474]), .B(n4534), .Y(n879) );
  INVX1 U530 ( .A(n879), .Y(n211) );
  AND2X1 U532 ( .A(mem[456]), .B(n4535), .Y(n860) );
  INVX1 U534 ( .A(n860), .Y(n212) );
  AND2X1 U536 ( .A(mem[444]), .B(n4535), .Y(n848) );
  INVX1 U538 ( .A(n848), .Y(n213) );
  AND2X1 U540 ( .A(mem[422]), .B(n4536), .Y(n825) );
  INVX1 U542 ( .A(n825), .Y(n214) );
  AND2X1 U544 ( .A(mem[410]), .B(n4536), .Y(n813) );
  INVX1 U546 ( .A(n813), .Y(n215) );
  AND2X1 U548 ( .A(mem[392]), .B(n4537), .Y(n794) );
  INVX1 U550 ( .A(n794), .Y(n216) );
  AND2X1 U553 ( .A(mem[380]), .B(n4537), .Y(n782) );
  INVX1 U555 ( .A(n782), .Y(n217) );
  AND2X1 U557 ( .A(mem[358]), .B(n4538), .Y(n759) );
  INVX1 U559 ( .A(n759), .Y(n218) );
  AND2X1 U561 ( .A(mem[346]), .B(n4538), .Y(n747) );
  INVX1 U563 ( .A(n747), .Y(n219) );
  AND2X1 U565 ( .A(mem[328]), .B(n4539), .Y(n728) );
  INVX1 U567 ( .A(n728), .Y(n220) );
  AND2X1 U569 ( .A(mem[316]), .B(n4539), .Y(n716) );
  INVX1 U571 ( .A(n716), .Y(n221) );
  AND2X1 U573 ( .A(mem[294]), .B(n4540), .Y(n692) );
  INVX1 U575 ( .A(n692), .Y(n222) );
  AND2X1 U577 ( .A(mem[282]), .B(n4540), .Y(n680) );
  INVX1 U579 ( .A(n680), .Y(n223) );
  AND2X1 U581 ( .A(mem[256]), .B(n4541), .Y(n652) );
  INVX1 U583 ( .A(n652), .Y(n224) );
  AND2X1 U585 ( .A(mem[244]), .B(n4541), .Y(n640) );
  INVX1 U587 ( .A(n640), .Y(n225) );
  AND2X1 U589 ( .A(mem[222]), .B(n4542), .Y(n616) );
  INVX1 U591 ( .A(n616), .Y(n226) );
  AND2X1 U593 ( .A(mem[210]), .B(n4542), .Y(n604) );
  INVX1 U595 ( .A(n604), .Y(n227) );
  AND2X1 U597 ( .A(mem[192]), .B(n4543), .Y(n584) );
  INVX1 U599 ( .A(n584), .Y(n228) );
  AND2X1 U601 ( .A(mem[180]), .B(n4543), .Y(n572) );
  INVX1 U603 ( .A(n572), .Y(n229) );
  AND2X1 U605 ( .A(mem[158]), .B(n4544), .Y(n548) );
  INVX1 U607 ( .A(n548), .Y(n230) );
  AND2X1 U609 ( .A(mem[146]), .B(n4544), .Y(n536) );
  INVX1 U611 ( .A(n536), .Y(n231) );
  AND2X1 U613 ( .A(mem[128]), .B(n4545), .Y(n516) );
  INVX1 U615 ( .A(n516), .Y(n232) );
  AND2X1 U617 ( .A(mem[116]), .B(n4545), .Y(n504) );
  INVX1 U621 ( .A(n504), .Y(n233) );
  AND2X1 U623 ( .A(mem[94]), .B(n4546), .Y(n480) );
  INVX1 U625 ( .A(n480), .Y(n234) );
  AND2X1 U627 ( .A(mem[82]), .B(n4546), .Y(n468) );
  INVX1 U629 ( .A(n468), .Y(n235) );
  AND2X1 U631 ( .A(mem[64]), .B(n4547), .Y(n448) );
  INVX1 U633 ( .A(n448), .Y(n236) );
  AND2X1 U635 ( .A(mem[52]), .B(n4547), .Y(n436) );
  INVX1 U637 ( .A(n436), .Y(n237) );
  AND2X1 U639 ( .A(mem[30]), .B(n4548), .Y(n409) );
  INVX1 U641 ( .A(n409), .Y(n238) );
  AND2X1 U643 ( .A(mem[18]), .B(n4548), .Y(n385) );
  INVX1 U645 ( .A(n385), .Y(n239) );
  AND2X1 U647 ( .A(mem[1045]), .B(n4517), .Y(n1469) );
  INVX1 U649 ( .A(n1469), .Y(n240) );
  AND2X1 U651 ( .A(mem[1033]), .B(n4517), .Y(n1457) );
  INVX1 U653 ( .A(n1457), .Y(n241) );
  AND2X1 U655 ( .A(mem[1013]), .B(n4518), .Y(n1436) );
  INVX1 U657 ( .A(n1436), .Y(n242) );
  AND2X1 U659 ( .A(mem[1001]), .B(n4518), .Y(n1424) );
  INVX1 U661 ( .A(n1424), .Y(n243) );
  AND2X1 U663 ( .A(mem[977]), .B(n4519), .Y(n1399) );
  INVX1 U665 ( .A(n1399), .Y(n244) );
  AND2X1 U667 ( .A(mem[964]), .B(n4519), .Y(n1386) );
  INVX1 U669 ( .A(n1386), .Y(n245) );
  AND2X1 U671 ( .A(mem[945]), .B(n4520), .Y(n1366) );
  INVX1 U673 ( .A(n1366), .Y(n246) );
  AND2X1 U675 ( .A(mem[933]), .B(n4520), .Y(n1354) );
  INVX1 U677 ( .A(n1354), .Y(n247) );
  AND2X1 U679 ( .A(mem[917]), .B(n4521), .Y(n1337) );
  INVX1 U681 ( .A(n1337), .Y(n248) );
  AND2X1 U683 ( .A(mem[905]), .B(n4521), .Y(n1325) );
  INVX1 U685 ( .A(n1325), .Y(n249) );
  AND2X1 U688 ( .A(mem[885]), .B(n4522), .Y(n1304) );
  INVX1 U690 ( .A(n1304), .Y(n250) );
  AND2X1 U692 ( .A(mem[873]), .B(n4522), .Y(n1292) );
  INVX1 U694 ( .A(n1292), .Y(n251) );
  AND2X1 U696 ( .A(mem[849]), .B(n4523), .Y(n1267) );
  INVX1 U698 ( .A(n1267), .Y(n252) );
  AND2X1 U700 ( .A(mem[837]), .B(n4523), .Y(n1255) );
  INVX1 U702 ( .A(n1255), .Y(n253) );
  AND2X1 U704 ( .A(mem[817]), .B(n4524), .Y(n1233) );
  INVX1 U706 ( .A(n1233), .Y(n254) );
  AND2X1 U708 ( .A(mem[805]), .B(n4524), .Y(n1221) );
  INVX1 U710 ( .A(n1221), .Y(n255) );
  AND2X1 U712 ( .A(mem[789]), .B(n4525), .Y(n1204) );
  INVX1 U714 ( .A(n1204), .Y(n256) );
  AND2X1 U716 ( .A(mem[777]), .B(n4525), .Y(n1192) );
  INVX1 U718 ( .A(n1192), .Y(n257) );
  AND2X1 U720 ( .A(mem[757]), .B(n4526), .Y(n1171) );
  INVX1 U722 ( .A(n1171), .Y(n258) );
  AND2X1 U724 ( .A(mem[745]), .B(n4526), .Y(n1159) );
  INVX1 U726 ( .A(n1159), .Y(n259) );
  AND2X1 U728 ( .A(mem[721]), .B(n4527), .Y(n1134) );
  INVX1 U730 ( .A(n1134), .Y(n260) );
  AND2X1 U732 ( .A(mem[709]), .B(n4527), .Y(n1122) );
  INVX1 U734 ( .A(n1122), .Y(n261) );
  AND2X1 U736 ( .A(mem[689]), .B(n4528), .Y(n1101) );
  INVX1 U738 ( .A(n1101), .Y(n262) );
  AND2X1 U740 ( .A(mem[677]), .B(n4528), .Y(n1089) );
  INVX1 U742 ( .A(n1089), .Y(n263) );
  AND2X1 U744 ( .A(mem[649]), .B(n4529), .Y(n1060) );
  INVX1 U746 ( .A(n1060), .Y(n264) );
  AND2X1 U748 ( .A(mem[637]), .B(n4529), .Y(n1048) );
  INVX1 U750 ( .A(n1048), .Y(n265) );
  AND2X1 U752 ( .A(mem[617]), .B(n4530), .Y(n1027) );
  INVX1 U755 ( .A(n1027), .Y(n266) );
  AND2X1 U757 ( .A(mem[605]), .B(n4530), .Y(n1015) );
  INVX1 U759 ( .A(n1015), .Y(n267) );
  AND2X1 U761 ( .A(mem[581]), .B(n4531), .Y(n990) );
  INVX1 U763 ( .A(n990), .Y(n268) );
  AND2X1 U765 ( .A(mem[568]), .B(n4531), .Y(n977) );
  INVX1 U767 ( .A(n977), .Y(n269) );
  AND2X1 U769 ( .A(mem[549]), .B(n4532), .Y(n956) );
  INVX1 U771 ( .A(n956), .Y(n270) );
  AND2X1 U773 ( .A(mem[537]), .B(n4532), .Y(n944) );
  INVX1 U775 ( .A(n944), .Y(n271) );
  AND2X1 U777 ( .A(mem[521]), .B(n4533), .Y(n927) );
  INVX1 U779 ( .A(n927), .Y(n272) );
  AND2X1 U781 ( .A(mem[509]), .B(n4533), .Y(n915) );
  INVX1 U783 ( .A(n915), .Y(n273) );
  AND2X1 U785 ( .A(mem[489]), .B(n4534), .Y(n894) );
  INVX1 U787 ( .A(n894), .Y(n274) );
  AND2X1 U789 ( .A(mem[477]), .B(n4534), .Y(n882) );
  INVX1 U791 ( .A(n882), .Y(n275) );
  AND2X1 U793 ( .A(mem[453]), .B(n4535), .Y(n857) );
  INVX1 U795 ( .A(n857), .Y(n276) );
  AND2X1 U797 ( .A(mem[441]), .B(n4535), .Y(n845) );
  INVX1 U799 ( .A(n845), .Y(n277) );
  AND2X1 U801 ( .A(mem[421]), .B(n4536), .Y(n824) );
  INVX1 U803 ( .A(n824), .Y(n278) );
  AND2X1 U805 ( .A(mem[409]), .B(n4536), .Y(n812) );
  INVX1 U807 ( .A(n812), .Y(n279) );
  AND2X1 U809 ( .A(mem[393]), .B(n4537), .Y(n795) );
  INVX1 U811 ( .A(n795), .Y(n280) );
  AND2X1 U813 ( .A(mem[381]), .B(n4537), .Y(n783) );
  INVX1 U815 ( .A(n783), .Y(n281) );
  AND2X1 U817 ( .A(mem[361]), .B(n4538), .Y(n762) );
  INVX1 U819 ( .A(n762), .Y(n282) );
  AND2X1 U822 ( .A(mem[349]), .B(n4538), .Y(n750) );
  INVX1 U824 ( .A(n750), .Y(n283) );
  AND2X1 U826 ( .A(mem[325]), .B(n4539), .Y(n725) );
  INVX1 U828 ( .A(n725), .Y(n284) );
  AND2X1 U830 ( .A(mem[313]), .B(n4539), .Y(n713) );
  INVX1 U832 ( .A(n713), .Y(n285) );
  AND2X1 U834 ( .A(mem[293]), .B(n4540), .Y(n691) );
  INVX1 U836 ( .A(n691), .Y(n286) );
  AND2X1 U838 ( .A(mem[281]), .B(n4540), .Y(n679) );
  INVX1 U840 ( .A(n679), .Y(n287) );
  AND2X1 U842 ( .A(mem[257]), .B(n4541), .Y(n653) );
  INVX1 U844 ( .A(n653), .Y(n288) );
  AND2X1 U846 ( .A(mem[245]), .B(n4541), .Y(n641) );
  INVX1 U848 ( .A(n641), .Y(n289) );
  AND2X1 U850 ( .A(mem[225]), .B(n4542), .Y(n619) );
  INVX1 U852 ( .A(n619), .Y(n290) );
  AND2X1 U854 ( .A(mem[213]), .B(n4542), .Y(n607) );
  INVX1 U856 ( .A(n607), .Y(n291) );
  AND2X1 U858 ( .A(mem[189]), .B(n4543), .Y(n581) );
  INVX1 U860 ( .A(n581), .Y(n292) );
  AND2X1 U862 ( .A(mem[177]), .B(n4543), .Y(n569) );
  INVX1 U864 ( .A(n569), .Y(n293) );
  AND2X1 U866 ( .A(mem[157]), .B(n4544), .Y(n547) );
  INVX1 U868 ( .A(n547), .Y(n294) );
  AND2X1 U870 ( .A(mem[145]), .B(n4544), .Y(n535) );
  INVX1 U872 ( .A(n535), .Y(n295) );
  AND2X1 U874 ( .A(mem[129]), .B(n4545), .Y(n517) );
  INVX1 U876 ( .A(n517), .Y(n296) );
  AND2X1 U878 ( .A(mem[117]), .B(n4545), .Y(n505) );
  INVX1 U880 ( .A(n505), .Y(n297) );
  AND2X1 U882 ( .A(mem[97]), .B(n4546), .Y(n483) );
  INVX1 U884 ( .A(n483), .Y(n298) );
  AND2X1 U886 ( .A(mem[85]), .B(n4546), .Y(n471) );
  INVX1 U889 ( .A(n471), .Y(n299) );
  AND2X1 U891 ( .A(mem[61]), .B(n4547), .Y(n445) );
  INVX1 U893 ( .A(n445), .Y(n300) );
  AND2X1 U895 ( .A(mem[49]), .B(n4547), .Y(n433) );
  INVX1 U897 ( .A(n433), .Y(n301) );
  AND2X1 U899 ( .A(mem[29]), .B(n4548), .Y(n407) );
  INVX1 U901 ( .A(n407), .Y(n302) );
  AND2X1 U903 ( .A(mem[17]), .B(n4548), .Y(n383) );
  INVX1 U905 ( .A(n383), .Y(n303) );
  AND2X1 U907 ( .A(mem[1046]), .B(n4517), .Y(n1470) );
  INVX1 U909 ( .A(n1470), .Y(n304) );
  AND2X1 U911 ( .A(mem[1034]), .B(n4517), .Y(n1458) );
  INVX1 U913 ( .A(n1458), .Y(n305) );
  AND2X1 U915 ( .A(mem[1012]), .B(n4518), .Y(n1435) );
  INVX1 U917 ( .A(n1435), .Y(n306) );
  AND2X1 U919 ( .A(mem[1000]), .B(n4518), .Y(n1423) );
  INVX1 U921 ( .A(n1423), .Y(n307) );
  AND2X1 U923 ( .A(mem[978]), .B(n4519), .Y(n1400) );
  INVX1 U925 ( .A(n1400), .Y(n308) );
  AND2X1 U927 ( .A(mem[966]), .B(n4519), .Y(n1388) );
  INVX1 U929 ( .A(n1388), .Y(n309) );
  AND2X1 U931 ( .A(mem[944]), .B(n4520), .Y(n1365) );
  INVX1 U933 ( .A(n1365), .Y(n310) );
  AND2X1 U935 ( .A(mem[931]), .B(n4520), .Y(n1352) );
  INVX1 U937 ( .A(n1352), .Y(n311) );
  AND2X1 U939 ( .A(mem[918]), .B(n4521), .Y(n1338) );
  INVX1 U941 ( .A(n1338), .Y(n312) );
  AND2X1 U943 ( .A(mem[906]), .B(n4521), .Y(n1326) );
  INVX1 U945 ( .A(n1326), .Y(n313) );
  AND2X1 U947 ( .A(mem[884]), .B(n4522), .Y(n1303) );
  INVX1 U949 ( .A(n1303), .Y(n314) );
  AND2X1 U951 ( .A(mem[872]), .B(n4522), .Y(n1291) );
  INVX1 U953 ( .A(n1291), .Y(n315) );
  AND2X1 U956 ( .A(mem[850]), .B(n4523), .Y(n1268) );
  INVX1 U958 ( .A(n1268), .Y(n316) );
  AND2X1 U960 ( .A(mem[838]), .B(n4523), .Y(n1256) );
  INVX1 U962 ( .A(n1256), .Y(n317) );
  AND2X1 U964 ( .A(mem[816]), .B(n4524), .Y(n1232) );
  INVX1 U966 ( .A(n1232), .Y(n318) );
  AND2X1 U968 ( .A(mem[804]), .B(n4524), .Y(n1220) );
  INVX1 U970 ( .A(n1220), .Y(n319) );
  AND2X1 U972 ( .A(mem[790]), .B(n4525), .Y(n1205) );
  INVX1 U974 ( .A(n1205), .Y(n320) );
  AND2X1 U976 ( .A(mem[778]), .B(n4525), .Y(n1193) );
  INVX1 U978 ( .A(n1193), .Y(n321) );
  AND2X1 U980 ( .A(mem[756]), .B(n4526), .Y(n1170) );
  INVX1 U982 ( .A(n1170), .Y(n322) );
  AND2X1 U984 ( .A(mem[744]), .B(n4526), .Y(n1158) );
  INVX1 U986 ( .A(n1158), .Y(n323) );
  AND2X1 U988 ( .A(mem[722]), .B(n4527), .Y(n1135) );
  INVX1 U990 ( .A(n1135), .Y(n324) );
  AND2X1 U992 ( .A(mem[710]), .B(n4527), .Y(n1123) );
  INVX1 U994 ( .A(n1123), .Y(n325) );
  AND2X1 U996 ( .A(mem[688]), .B(n4528), .Y(n1100) );
  INVX1 U998 ( .A(n1100), .Y(n326) );
  AND2X1 U1000 ( .A(mem[676]), .B(n4528), .Y(n1088) );
  INVX1 U1002 ( .A(n1088), .Y(n327) );
  AND2X1 U1004 ( .A(mem[650]), .B(n4529), .Y(n1061) );
  INVX1 U1006 ( .A(n1061), .Y(n328) );
  AND2X1 U1008 ( .A(mem[638]), .B(n4529), .Y(n1049) );
  INVX1 U1010 ( .A(n1049), .Y(n329) );
  AND2X1 U1012 ( .A(mem[616]), .B(n4530), .Y(n1026) );
  INVX1 U1014 ( .A(n1026), .Y(n330) );
  AND2X1 U1016 ( .A(mem[604]), .B(n4530), .Y(n1014) );
  INVX1 U1018 ( .A(n1014), .Y(n331) );
  AND2X1 U1020 ( .A(mem[582]), .B(n4531), .Y(n991) );
  INVX1 U1023 ( .A(n991), .Y(n332) );
  AND2X1 U1025 ( .A(mem[570]), .B(n4531), .Y(n979) );
  INVX1 U1027 ( .A(n979), .Y(n333) );
  AND2X1 U1029 ( .A(mem[548]), .B(n4532), .Y(n955) );
  INVX1 U1031 ( .A(n955), .Y(n334) );
  AND2X1 U1033 ( .A(mem[535]), .B(n4532), .Y(n942) );
  INVX1 U1035 ( .A(n942), .Y(n335) );
  AND2X1 U1037 ( .A(mem[522]), .B(n4533), .Y(n928) );
  INVX1 U1039 ( .A(n928), .Y(n336) );
  AND2X1 U1041 ( .A(mem[510]), .B(n4533), .Y(n916) );
  INVX1 U1043 ( .A(n916), .Y(n337) );
  AND2X1 U1045 ( .A(mem[488]), .B(n4534), .Y(n893) );
  INVX1 U1047 ( .A(n893), .Y(n338) );
  AND2X1 U1049 ( .A(mem[476]), .B(n4534), .Y(n881) );
  INVX1 U1051 ( .A(n881), .Y(n339) );
  AND2X1 U1053 ( .A(mem[454]), .B(n4535), .Y(n858) );
  INVX1 U1055 ( .A(n858), .Y(n340) );
  AND2X1 U1057 ( .A(mem[442]), .B(n4535), .Y(n846) );
  INVX1 U1059 ( .A(n846), .Y(n341) );
  AND2X1 U1061 ( .A(mem[420]), .B(n4536), .Y(n823) );
  INVX1 U1063 ( .A(n823), .Y(n342) );
  AND2X1 U1065 ( .A(mem[408]), .B(n4536), .Y(n811) );
  INVX1 U1067 ( .A(n811), .Y(n343) );
  AND2X1 U1069 ( .A(mem[394]), .B(n4537), .Y(n796) );
  INVX1 U1071 ( .A(n796), .Y(n344) );
  AND2X1 U1073 ( .A(mem[382]), .B(n4537), .Y(n784) );
  INVX1 U1075 ( .A(n784), .Y(n345) );
  AND2X1 U1077 ( .A(mem[360]), .B(n4538), .Y(n761) );
  INVX1 U1079 ( .A(n761), .Y(n346) );
  AND2X1 U1081 ( .A(mem[348]), .B(n4538), .Y(n749) );
  INVX1 U1083 ( .A(n749), .Y(n347) );
  AND2X1 U1085 ( .A(mem[326]), .B(n4539), .Y(n726) );
  INVX1 U1087 ( .A(n726), .Y(n348) );
  AND2X1 U1090 ( .A(mem[314]), .B(n4539), .Y(n714) );
  INVX1 U1092 ( .A(n714), .Y(n350) );
  AND2X1 U1094 ( .A(mem[292]), .B(n4540), .Y(n690) );
  INVX1 U1096 ( .A(n690), .Y(n352) );
  AND2X1 U1098 ( .A(mem[280]), .B(n4540), .Y(n678) );
  INVX1 U1100 ( .A(n678), .Y(n354) );
  AND2X1 U1102 ( .A(mem[258]), .B(n4541), .Y(n654) );
  INVX1 U1104 ( .A(n654), .Y(n356) );
  AND2X1 U1106 ( .A(mem[246]), .B(n4541), .Y(n642) );
  INVX1 U1108 ( .A(n642), .Y(n358) );
  AND2X1 U1110 ( .A(mem[224]), .B(n4542), .Y(n618) );
  INVX1 U1112 ( .A(n618), .Y(n360) );
  AND2X1 U1114 ( .A(mem[212]), .B(n4542), .Y(n606) );
  INVX1 U1116 ( .A(n606), .Y(n362) );
  AND2X1 U1118 ( .A(mem[190]), .B(n4543), .Y(n582) );
  INVX1 U1120 ( .A(n582), .Y(n364) );
  AND2X1 U1122 ( .A(mem[178]), .B(n4543), .Y(n570) );
  INVX1 U1124 ( .A(n570), .Y(n366) );
  AND2X1 U1126 ( .A(mem[156]), .B(n4544), .Y(n546) );
  INVX1 U1128 ( .A(n546), .Y(n368) );
  AND2X1 U1130 ( .A(mem[144]), .B(n4544), .Y(n534) );
  INVX1 U1132 ( .A(n534), .Y(n370) );
  AND2X1 U1134 ( .A(mem[130]), .B(n4545), .Y(n518) );
  INVX1 U1136 ( .A(n518), .Y(n372) );
  AND2X1 U1138 ( .A(mem[118]), .B(n4545), .Y(n506) );
  INVX1 U1140 ( .A(n506), .Y(n374) );
  AND2X1 U1142 ( .A(mem[96]), .B(n4546), .Y(n482) );
  INVX1 U1144 ( .A(n482), .Y(n376) );
  AND2X1 U1146 ( .A(mem[84]), .B(n4546), .Y(n470) );
  INVX1 U1148 ( .A(n470), .Y(n378) );
  AND2X1 U1150 ( .A(mem[62]), .B(n4547), .Y(n446) );
  INVX1 U1152 ( .A(n446), .Y(n380) );
  AND2X1 U1154 ( .A(mem[50]), .B(n4547), .Y(n434) );
  INVX1 U1158 ( .A(n434), .Y(n382) );
  AND2X1 U1160 ( .A(mem[28]), .B(n4548), .Y(n405) );
  INVX1 U1162 ( .A(n405), .Y(n384) );
  AND2X1 U1164 ( .A(mem[16]), .B(n4548), .Y(n381) );
  INVX1 U1166 ( .A(n381), .Y(n386) );
  AND2X1 U1168 ( .A(mem[1028]), .B(n4517), .Y(n1452) );
  INVX1 U1170 ( .A(n1452), .Y(n388) );
  AND2X1 U1172 ( .A(mem[1023]), .B(n4517), .Y(n1447) );
  INVX1 U1174 ( .A(n1447), .Y(n390) );
  AND2X1 U1176 ( .A(mem[996]), .B(n4518), .Y(n1419) );
  INVX1 U1178 ( .A(n1419), .Y(n392) );
  AND2X1 U1180 ( .A(mem[991]), .B(n4518), .Y(n1414) );
  INVX1 U1182 ( .A(n1414), .Y(n394) );
  AND2X1 U1184 ( .A(mem[965]), .B(n4519), .Y(n1387) );
  INVX1 U1186 ( .A(n1387), .Y(n396) );
  AND2X1 U1188 ( .A(mem[959]), .B(n4519), .Y(n1381) );
  INVX1 U1190 ( .A(n1381), .Y(n398) );
  AND2X1 U1192 ( .A(mem[928]), .B(n4520), .Y(n1349) );
  INVX1 U1194 ( .A(n1349), .Y(n400) );
  AND2X1 U1196 ( .A(mem[927]), .B(n4520), .Y(n1348) );
  INVX1 U1198 ( .A(n1348), .Y(n402) );
  AND2X1 U1200 ( .A(mem[919]), .B(n4521), .Y(n1339) );
  INVX1 U1202 ( .A(n1339), .Y(n404) );
  AND2X1 U1204 ( .A(mem[907]), .B(n4521), .Y(n1327) );
  INVX1 U1206 ( .A(n1327), .Y(n406) );
  AND2X1 U1208 ( .A(mem[887]), .B(n4522), .Y(n1306) );
  INVX1 U1210 ( .A(n1306), .Y(n408) );
  AND2X1 U1212 ( .A(mem[875]), .B(n4522), .Y(n1294) );
  INVX1 U1214 ( .A(n1294), .Y(n410) );
  AND2X1 U1216 ( .A(mem[855]), .B(n4523), .Y(n1273) );
  INVX1 U1218 ( .A(n1273), .Y(n412) );
  AND2X1 U1220 ( .A(mem[843]), .B(n4523), .Y(n1261) );
  INVX1 U1222 ( .A(n1261), .Y(n2604) );
  AND2X1 U1225 ( .A(mem[823]), .B(n4524), .Y(n1239) );
  INVX1 U1227 ( .A(n1239), .Y(n2605) );
  AND2X1 U1229 ( .A(mem[811]), .B(n4524), .Y(n1227) );
  INVX1 U1231 ( .A(n1227), .Y(n2606) );
  AND2X1 U1233 ( .A(mem[783]), .B(n4525), .Y(n1198) );
  INVX1 U1235 ( .A(n1198), .Y(n2607) );
  AND2X1 U1237 ( .A(mem[771]), .B(n4525), .Y(n1186) );
  INVX1 U1239 ( .A(n1186), .Y(n2608) );
  AND2X1 U1241 ( .A(mem[751]), .B(n4526), .Y(n1165) );
  INVX1 U1243 ( .A(n1165), .Y(n2609) );
  AND2X1 U1245 ( .A(mem[739]), .B(n4526), .Y(n1153) );
  INVX1 U1247 ( .A(n1153), .Y(n2610) );
  AND2X1 U1249 ( .A(mem[719]), .B(n4527), .Y(n1132) );
  INVX1 U1251 ( .A(n1132), .Y(n2611) );
  AND2X1 U1253 ( .A(mem[707]), .B(n4527), .Y(n1120) );
  INVX1 U1255 ( .A(n1120), .Y(n2612) );
  AND2X1 U1257 ( .A(mem[687]), .B(n4528), .Y(n1099) );
  INVX1 U1259 ( .A(n1099), .Y(n2613) );
  AND2X1 U1261 ( .A(mem[675]), .B(n4528), .Y(n1087) );
  INVX1 U1263 ( .A(n1087), .Y(n2614) );
  AND2X1 U1265 ( .A(mem[632]), .B(n4529), .Y(n1043) );
  INVX1 U1267 ( .A(n1043), .Y(n2615) );
  AND2X1 U1269 ( .A(mem[627]), .B(n4529), .Y(n1038) );
  INVX1 U1271 ( .A(n1038), .Y(n2616) );
  AND2X1 U1273 ( .A(mem[600]), .B(n4530), .Y(n1010) );
  INVX1 U1275 ( .A(n1010), .Y(n2617) );
  AND2X1 U1277 ( .A(mem[595]), .B(n4530), .Y(n1005) );
  INVX1 U1279 ( .A(n1005), .Y(n2618) );
  AND2X1 U1281 ( .A(mem[569]), .B(n4531), .Y(n978) );
  INVX1 U1283 ( .A(n978), .Y(n2619) );
  AND2X1 U1285 ( .A(mem[563]), .B(n4531), .Y(n972) );
  INVX1 U1287 ( .A(n972), .Y(n2620) );
  AND2X1 U1289 ( .A(mem[532]), .B(n4532), .Y(n939) );
  INVX1 U1292 ( .A(n939), .Y(n2621) );
  AND2X1 U1294 ( .A(mem[531]), .B(n4532), .Y(n938) );
  INVX1 U1296 ( .A(n938), .Y(n2622) );
  AND2X1 U1298 ( .A(mem[523]), .B(n4533), .Y(n929) );
  INVX1 U1300 ( .A(n929), .Y(n2623) );
  AND2X1 U1302 ( .A(mem[511]), .B(n4533), .Y(n917) );
  INVX1 U1304 ( .A(n917), .Y(n2624) );
  AND2X1 U1306 ( .A(mem[491]), .B(n4534), .Y(n896) );
  INVX1 U1308 ( .A(n896), .Y(n2625) );
  AND2X1 U1310 ( .A(mem[479]), .B(n4534), .Y(n884) );
  INVX1 U1312 ( .A(n884), .Y(n2626) );
  AND2X1 U1314 ( .A(mem[459]), .B(n4535), .Y(n863) );
  INVX1 U1316 ( .A(n863), .Y(n2627) );
  AND2X1 U1318 ( .A(mem[447]), .B(n4535), .Y(n851) );
  INVX1 U1320 ( .A(n851), .Y(n2628) );
  AND2X1 U1322 ( .A(mem[427]), .B(n4536), .Y(n830) );
  INVX1 U1324 ( .A(n830), .Y(n2629) );
  AND2X1 U1326 ( .A(mem[415]), .B(n4536), .Y(n818) );
  INVX1 U1328 ( .A(n818), .Y(n2630) );
  AND2X1 U1330 ( .A(mem[387]), .B(n4537), .Y(n789) );
  INVX1 U1332 ( .A(n789), .Y(n2631) );
  AND2X1 U1334 ( .A(mem[375]), .B(n4537), .Y(n777) );
  INVX1 U1336 ( .A(n777), .Y(n2632) );
  AND2X1 U1338 ( .A(mem[355]), .B(n4538), .Y(n756) );
  INVX1 U1340 ( .A(n756), .Y(n2633) );
  AND2X1 U1342 ( .A(mem[343]), .B(n4538), .Y(n744) );
  INVX1 U1344 ( .A(n744), .Y(n2634) );
  AND2X1 U1346 ( .A(mem[323]), .B(n4539), .Y(n723) );
  INVX1 U1348 ( .A(n723), .Y(n2635) );
  AND2X1 U1350 ( .A(mem[311]), .B(n4539), .Y(n711) );
  INVX1 U1352 ( .A(n711), .Y(n2636) );
  AND2X1 U1354 ( .A(mem[291]), .B(n4540), .Y(n689) );
  INVX1 U1356 ( .A(n689), .Y(n2637) );
  AND2X1 U1359 ( .A(mem[279]), .B(n4540), .Y(n677) );
  INVX1 U1361 ( .A(n677), .Y(n2638) );
  AND2X1 U1363 ( .A(mem[259]), .B(n4541), .Y(n655) );
  INVX1 U1365 ( .A(n655), .Y(n2639) );
  AND2X1 U1367 ( .A(mem[247]), .B(n4541), .Y(n643) );
  INVX1 U1369 ( .A(n643), .Y(n2640) );
  AND2X1 U1371 ( .A(mem[227]), .B(n4542), .Y(n621) );
  INVX1 U1373 ( .A(n621), .Y(n2641) );
  AND2X1 U1375 ( .A(mem[215]), .B(n4542), .Y(n609) );
  INVX1 U1377 ( .A(n609), .Y(n2642) );
  AND2X1 U1379 ( .A(mem[195]), .B(n4543), .Y(n587) );
  INVX1 U1381 ( .A(n587), .Y(n2643) );
  AND2X1 U1383 ( .A(mem[183]), .B(n4543), .Y(n575) );
  INVX1 U1385 ( .A(n575), .Y(n2644) );
  AND2X1 U1387 ( .A(mem[163]), .B(n4544), .Y(n553) );
  INVX1 U1389 ( .A(n553), .Y(n2645) );
  AND2X1 U1391 ( .A(mem[151]), .B(n4544), .Y(n541) );
  INVX1 U1393 ( .A(n541), .Y(n2646) );
  AND2X1 U1395 ( .A(mem[123]), .B(n4545), .Y(n511) );
  INVX1 U1397 ( .A(n511), .Y(n2647) );
  AND2X1 U1399 ( .A(mem[111]), .B(n4545), .Y(n499) );
  INVX1 U1401 ( .A(n499), .Y(n2648) );
  AND2X1 U1403 ( .A(mem[91]), .B(n4546), .Y(n477) );
  INVX1 U1405 ( .A(n477), .Y(n2649) );
  AND2X1 U1407 ( .A(mem[79]), .B(n4546), .Y(n465) );
  INVX1 U1409 ( .A(n465), .Y(n2650) );
  AND2X1 U1411 ( .A(mem[59]), .B(n4547), .Y(n443) );
  INVX1 U1413 ( .A(n443), .Y(n2651) );
  AND2X1 U1415 ( .A(mem[47]), .B(n4547), .Y(n431) );
  INVX1 U1417 ( .A(n431), .Y(n2652) );
  AND2X1 U1419 ( .A(mem[27]), .B(n4548), .Y(n403) );
  INVX1 U1421 ( .A(n403), .Y(n2653) );
  AND2X1 U1423 ( .A(mem[15]), .B(n4548), .Y(n379) );
  INVX1 U1426 ( .A(n379), .Y(n2654) );
  AND2X1 U1428 ( .A(mem[1029]), .B(n4517), .Y(n1453) );
  INVX1 U1430 ( .A(n1453), .Y(n2655) );
  AND2X1 U1432 ( .A(mem[1024]), .B(n4517), .Y(n1448) );
  INVX1 U1434 ( .A(n1448), .Y(n2656) );
  AND2X1 U1436 ( .A(mem[995]), .B(n4518), .Y(n1418) );
  INVX1 U1438 ( .A(n1418), .Y(n2657) );
  AND2X1 U1440 ( .A(mem[990]), .B(n4518), .Y(n1413) );
  INVX1 U1442 ( .A(n1413), .Y(n2658) );
  AND2X1 U1444 ( .A(mem[961]), .B(n4519), .Y(n1383) );
  INVX1 U1446 ( .A(n1383), .Y(n2659) );
  AND2X1 U1448 ( .A(mem[960]), .B(n4519), .Y(n1382) );
  INVX1 U1450 ( .A(n1382), .Y(n2660) );
  AND2X1 U1452 ( .A(mem[932]), .B(n4520), .Y(n1353) );
  INVX1 U1454 ( .A(n1353), .Y(n2661) );
  AND2X1 U1456 ( .A(mem[926]), .B(n4520), .Y(n1347) );
  INVX1 U1458 ( .A(n1347), .Y(n2662) );
  AND2X1 U1460 ( .A(mem[920]), .B(n4521), .Y(n1340) );
  INVX1 U1462 ( .A(n1340), .Y(n2663) );
  AND2X1 U1464 ( .A(mem[908]), .B(n4521), .Y(n1328) );
  INVX1 U1466 ( .A(n1328), .Y(n2664) );
  AND2X1 U1468 ( .A(mem[886]), .B(n4522), .Y(n1305) );
  INVX1 U1470 ( .A(n1305), .Y(n2665) );
  AND2X1 U1472 ( .A(mem[874]), .B(n4522), .Y(n1293) );
  INVX1 U1474 ( .A(n1293), .Y(n2666) );
  AND2X1 U1476 ( .A(mem[856]), .B(n4523), .Y(n1274) );
  INVX1 U1478 ( .A(n1274), .Y(n2667) );
  AND2X1 U1480 ( .A(mem[844]), .B(n4523), .Y(n1262) );
  INVX1 U1482 ( .A(n1262), .Y(n2668) );
  AND2X1 U1484 ( .A(mem[822]), .B(n4524), .Y(n1238) );
  INVX1 U1486 ( .A(n1238), .Y(n2669) );
  AND2X1 U1488 ( .A(mem[810]), .B(n4524), .Y(n1226) );
  INVX1 U1490 ( .A(n1226), .Y(n2670) );
  AND2X1 U1493 ( .A(mem[784]), .B(n4525), .Y(n1199) );
  INVX1 U1495 ( .A(n1199), .Y(n2671) );
  AND2X1 U1497 ( .A(mem[772]), .B(n4525), .Y(n1187) );
  INVX1 U1499 ( .A(n1187), .Y(n2672) );
  AND2X1 U1501 ( .A(mem[750]), .B(n4526), .Y(n1164) );
  INVX1 U1503 ( .A(n1164), .Y(n2673) );
  AND2X1 U1505 ( .A(mem[738]), .B(n4526), .Y(n1152) );
  INVX1 U1507 ( .A(n1152), .Y(n2674) );
  AND2X1 U1509 ( .A(mem[720]), .B(n4527), .Y(n1133) );
  INVX1 U1511 ( .A(n1133), .Y(n2675) );
  AND2X1 U1513 ( .A(mem[708]), .B(n4527), .Y(n1121) );
  INVX1 U1515 ( .A(n1121), .Y(n2676) );
  AND2X1 U1517 ( .A(mem[686]), .B(n4528), .Y(n1098) );
  INVX1 U1519 ( .A(n1098), .Y(n2677) );
  AND2X1 U1521 ( .A(mem[674]), .B(n4528), .Y(n1086) );
  INVX1 U1523 ( .A(n1086), .Y(n2678) );
  AND2X1 U1525 ( .A(mem[633]), .B(n4529), .Y(n1044) );
  INVX1 U1527 ( .A(n1044), .Y(n2679) );
  AND2X1 U1529 ( .A(mem[628]), .B(n4529), .Y(n1039) );
  INVX1 U1531 ( .A(n1039), .Y(n2680) );
  AND2X1 U1533 ( .A(mem[599]), .B(n4530), .Y(n1009) );
  INVX1 U1535 ( .A(n1009), .Y(n2681) );
  AND2X1 U1537 ( .A(mem[594]), .B(n4530), .Y(n1004) );
  INVX1 U1539 ( .A(n1004), .Y(n2682) );
  AND2X1 U1541 ( .A(mem[565]), .B(n4531), .Y(n974) );
  INVX1 U1543 ( .A(n974), .Y(n2683) );
  AND2X1 U1545 ( .A(mem[564]), .B(n4531), .Y(n973) );
  INVX1 U1547 ( .A(n973), .Y(n2684) );
  AND2X1 U1549 ( .A(mem[536]), .B(n4532), .Y(n943) );
  INVX1 U1551 ( .A(n943), .Y(n2685) );
  AND2X1 U1553 ( .A(mem[530]), .B(n4532), .Y(n937) );
  INVX1 U1555 ( .A(n937), .Y(n2686) );
  AND2X1 U1557 ( .A(mem[524]), .B(n4533), .Y(n930) );
  INVX1 U1560 ( .A(n930), .Y(n2687) );
  AND2X1 U1562 ( .A(mem[512]), .B(n4533), .Y(n918) );
  INVX1 U1564 ( .A(n918), .Y(n2688) );
  AND2X1 U1566 ( .A(mem[490]), .B(n4534), .Y(n895) );
  INVX1 U1568 ( .A(n895), .Y(n2689) );
  AND2X1 U1570 ( .A(mem[478]), .B(n4534), .Y(n883) );
  INVX1 U1572 ( .A(n883), .Y(n2690) );
  AND2X1 U1574 ( .A(mem[460]), .B(n4535), .Y(n864) );
  INVX1 U1576 ( .A(n864), .Y(n2691) );
  AND2X1 U1578 ( .A(mem[448]), .B(n4535), .Y(n852) );
  INVX1 U1580 ( .A(n852), .Y(n2692) );
  AND2X1 U1582 ( .A(mem[426]), .B(n4536), .Y(n829) );
  INVX1 U1584 ( .A(n829), .Y(n2693) );
  AND2X1 U1586 ( .A(mem[414]), .B(n4536), .Y(n817) );
  INVX1 U1588 ( .A(n817), .Y(n2694) );
  AND2X1 U1590 ( .A(mem[388]), .B(n4537), .Y(n790) );
  INVX1 U1592 ( .A(n790), .Y(n2695) );
  AND2X1 U1594 ( .A(mem[376]), .B(n4537), .Y(n778) );
  INVX1 U1596 ( .A(n778), .Y(n2696) );
  AND2X1 U1598 ( .A(mem[354]), .B(n4538), .Y(n755) );
  INVX1 U1600 ( .A(n755), .Y(n2697) );
  AND2X1 U1602 ( .A(mem[342]), .B(n4538), .Y(n743) );
  INVX1 U1604 ( .A(n743), .Y(n2698) );
  AND2X1 U1606 ( .A(mem[324]), .B(n4539), .Y(n724) );
  INVX1 U1608 ( .A(n724), .Y(n2699) );
  AND2X1 U1610 ( .A(mem[312]), .B(n4539), .Y(n712) );
  INVX1 U1612 ( .A(n712), .Y(n2700) );
  AND2X1 U1614 ( .A(mem[290]), .B(n4540), .Y(n688) );
  INVX1 U1616 ( .A(n688), .Y(n2701) );
  AND2X1 U1618 ( .A(mem[278]), .B(n4540), .Y(n676) );
  INVX1 U1620 ( .A(n676), .Y(n2702) );
  AND2X1 U1622 ( .A(mem[260]), .B(n4541), .Y(n656) );
  INVX1 U1624 ( .A(n656), .Y(n2703) );
  AND2X1 U1627 ( .A(mem[248]), .B(n4541), .Y(n644) );
  INVX1 U1629 ( .A(n644), .Y(n2704) );
  AND2X1 U1631 ( .A(mem[226]), .B(n4542), .Y(n620) );
  INVX1 U1633 ( .A(n620), .Y(n2705) );
  AND2X1 U1635 ( .A(mem[214]), .B(n4542), .Y(n608) );
  INVX1 U1637 ( .A(n608), .Y(n2706) );
  AND2X1 U1639 ( .A(mem[196]), .B(n4543), .Y(n588) );
  INVX1 U1641 ( .A(n588), .Y(n2707) );
  AND2X1 U1643 ( .A(mem[184]), .B(n4543), .Y(n576) );
  INVX1 U1645 ( .A(n576), .Y(n2708) );
  AND2X1 U1647 ( .A(mem[162]), .B(n4544), .Y(n552) );
  INVX1 U1649 ( .A(n552), .Y(n2709) );
  AND2X1 U1651 ( .A(mem[150]), .B(n4544), .Y(n540) );
  INVX1 U1653 ( .A(n540), .Y(n2710) );
  AND2X1 U1655 ( .A(mem[124]), .B(n4545), .Y(n512) );
  INVX1 U1657 ( .A(n512), .Y(n2711) );
  AND2X1 U1659 ( .A(mem[112]), .B(n4545), .Y(n500) );
  INVX1 U1661 ( .A(n500), .Y(n2712) );
  AND2X1 U1663 ( .A(mem[90]), .B(n4546), .Y(n476) );
  INVX1 U1665 ( .A(n476), .Y(n2713) );
  AND2X1 U1667 ( .A(mem[78]), .B(n4546), .Y(n464) );
  INVX1 U1669 ( .A(n464), .Y(n2714) );
  AND2X1 U1671 ( .A(mem[60]), .B(n4547), .Y(n444) );
  INVX1 U1673 ( .A(n444), .Y(n2715) );
  AND2X1 U1675 ( .A(mem[48]), .B(n4547), .Y(n432) );
  INVX1 U1677 ( .A(n432), .Y(n2716) );
  AND2X1 U1679 ( .A(mem[26]), .B(n4548), .Y(n401) );
  INVX1 U1681 ( .A(n401), .Y(n2717) );
  AND2X1 U1683 ( .A(mem[14]), .B(n4548), .Y(n377) );
  INVX1 U1685 ( .A(n377), .Y(n2718) );
  AND2X1 U1687 ( .A(mem[1031]), .B(n4517), .Y(n1455) );
  INVX1 U1689 ( .A(n1455), .Y(n2719) );
  AND2X1 U1691 ( .A(mem[1025]), .B(n4517), .Y(n1449) );
  INVX1 U1695 ( .A(n1449), .Y(n2720) );
  AND2X1 U1697 ( .A(mem[994]), .B(n4518), .Y(n1417) );
  INVX1 U1699 ( .A(n1417), .Y(n2721) );
  AND2X1 U1701 ( .A(mem[993]), .B(n4518), .Y(n1416) );
  INVX1 U1703 ( .A(n1416), .Y(n2722) );
  AND2X1 U1705 ( .A(mem[962]), .B(n4519), .Y(n1384) );
  INVX1 U1707 ( .A(n1384), .Y(n2723) );
  AND2X1 U1709 ( .A(mem[957]), .B(n4519), .Y(n1379) );
  INVX1 U1711 ( .A(n1379), .Y(n2724) );
  AND2X1 U1713 ( .A(mem[930]), .B(n4520), .Y(n1351) );
  INVX1 U1715 ( .A(n1351), .Y(n2725) );
  AND2X1 U1717 ( .A(mem[925]), .B(n4520), .Y(n1346) );
  INVX1 U1719 ( .A(n1346), .Y(n2726) );
  AND2X1 U1721 ( .A(mem[921]), .B(n4521), .Y(n1341) );
  INVX1 U1723 ( .A(n1341), .Y(n2727) );
  AND2X1 U1725 ( .A(mem[909]), .B(n4521), .Y(n1329) );
  INVX1 U1727 ( .A(n1329), .Y(n2728) );
  AND2X1 U1729 ( .A(mem[889]), .B(n4522), .Y(n1308) );
  INVX1 U1731 ( .A(n1308), .Y(n2729) );
  AND2X1 U1733 ( .A(mem[877]), .B(n4522), .Y(n1296) );
  INVX1 U1735 ( .A(n1296), .Y(n2730) );
  AND2X1 U1737 ( .A(mem[853]), .B(n4523), .Y(n1271) );
  INVX1 U1739 ( .A(n1271), .Y(n2731) );
  AND2X1 U1741 ( .A(mem[841]), .B(n4523), .Y(n1259) );
  INVX1 U1743 ( .A(n1259), .Y(n2732) );
  AND2X1 U1745 ( .A(mem[821]), .B(n4524), .Y(n1237) );
  INVX1 U1747 ( .A(n1237), .Y(n2733) );
  AND2X1 U1749 ( .A(mem[809]), .B(n4524), .Y(n1225) );
  INVX1 U1751 ( .A(n1225), .Y(n2734) );
  AND2X1 U1753 ( .A(mem[785]), .B(n4525), .Y(n1200) );
  INVX1 U1755 ( .A(n1200), .Y(n2735) );
  AND2X1 U1757 ( .A(mem[773]), .B(n4525), .Y(n1188) );
  INVX1 U1759 ( .A(n1188), .Y(n2736) );
  AND2X1 U1763 ( .A(mem[753]), .B(n4526), .Y(n1167) );
  INVX1 U1765 ( .A(n1167), .Y(n2737) );
  AND2X1 U1767 ( .A(mem[741]), .B(n4526), .Y(n1155) );
  INVX1 U1769 ( .A(n1155), .Y(n2738) );
  AND2X1 U1771 ( .A(mem[717]), .B(n4527), .Y(n1130) );
  INVX1 U1773 ( .A(n1130), .Y(n2739) );
  AND2X1 U1775 ( .A(mem[705]), .B(n4527), .Y(n1118) );
  INVX1 U1777 ( .A(n1118), .Y(n2740) );
  AND2X1 U1779 ( .A(mem[685]), .B(n4528), .Y(n1097) );
  INVX1 U1781 ( .A(n1097), .Y(n2741) );
  AND2X1 U1783 ( .A(mem[673]), .B(n4528), .Y(n1085) );
  INVX1 U1785 ( .A(n1085), .Y(n2742) );
  AND2X1 U1787 ( .A(mem[635]), .B(n4529), .Y(n1046) );
  INVX1 U1789 ( .A(n1046), .Y(n2743) );
  AND2X1 U1791 ( .A(mem[629]), .B(n4529), .Y(n1040) );
  INVX1 U1793 ( .A(n1040), .Y(n2744) );
  AND2X1 U1795 ( .A(mem[598]), .B(n4530), .Y(n1008) );
  INVX1 U1797 ( .A(n1008), .Y(n2745) );
  AND2X1 U1799 ( .A(mem[597]), .B(n4530), .Y(n1007) );
  INVX1 U1801 ( .A(n1007), .Y(n2746) );
  AND2X1 U1803 ( .A(mem[566]), .B(n4531), .Y(n975) );
  INVX1 U1805 ( .A(n975), .Y(n2747) );
  AND2X1 U1807 ( .A(mem[561]), .B(n4531), .Y(n970) );
  INVX1 U1809 ( .A(n970), .Y(n2748) );
  AND2X1 U1811 ( .A(mem[534]), .B(n4532), .Y(n941) );
  INVX1 U1813 ( .A(n941), .Y(n2749) );
  AND2X1 U1815 ( .A(mem[529]), .B(n4532), .Y(n936) );
  INVX1 U1817 ( .A(n936), .Y(n2750) );
  AND2X1 U1819 ( .A(mem[525]), .B(n4533), .Y(n931) );
  INVX1 U1821 ( .A(n931), .Y(n2751) );
  AND2X1 U1823 ( .A(mem[513]), .B(n4533), .Y(n919) );
  INVX1 U1825 ( .A(n919), .Y(n2752) );
  AND2X1 U1827 ( .A(mem[493]), .B(n4534), .Y(n898) );
  INVX1 U1831 ( .A(n898), .Y(n2753) );
  AND2X1 U1833 ( .A(mem[481]), .B(n4534), .Y(n886) );
  INVX1 U1835 ( .A(n886), .Y(n2754) );
  AND2X1 U1837 ( .A(mem[457]), .B(n4535), .Y(n861) );
  INVX1 U1839 ( .A(n861), .Y(n2755) );
  AND2X1 U1841 ( .A(mem[445]), .B(n4535), .Y(n849) );
  INVX1 U1843 ( .A(n849), .Y(n2756) );
  AND2X1 U1845 ( .A(mem[425]), .B(n4536), .Y(n828) );
  INVX1 U1847 ( .A(n828), .Y(n2757) );
  AND2X1 U1849 ( .A(mem[413]), .B(n4536), .Y(n816) );
  INVX1 U1851 ( .A(n816), .Y(n2758) );
  AND2X1 U1853 ( .A(mem[389]), .B(n4537), .Y(n791) );
  INVX1 U1855 ( .A(n791), .Y(n2759) );
  AND2X1 U1857 ( .A(mem[377]), .B(n4537), .Y(n779) );
  INVX1 U1859 ( .A(n779), .Y(n2760) );
  AND2X1 U1861 ( .A(mem[357]), .B(n4538), .Y(n758) );
  INVX1 U1863 ( .A(n758), .Y(n2761) );
  AND2X1 U1865 ( .A(mem[345]), .B(n4538), .Y(n746) );
  INVX1 U1867 ( .A(n746), .Y(n2762) );
  AND2X1 U1869 ( .A(mem[321]), .B(n4539), .Y(n721) );
  INVX1 U1871 ( .A(n721), .Y(n2763) );
  AND2X1 U1873 ( .A(mem[309]), .B(n4539), .Y(n709) );
  INVX1 U1875 ( .A(n709), .Y(n2764) );
  AND2X1 U1877 ( .A(mem[289]), .B(n4540), .Y(n687) );
  INVX1 U1879 ( .A(n687), .Y(n2765) );
  AND2X1 U1881 ( .A(mem[277]), .B(n4540), .Y(n675) );
  INVX1 U1883 ( .A(n675), .Y(n2766) );
  AND2X1 U1885 ( .A(mem[261]), .B(n4541), .Y(n657) );
  INVX1 U1887 ( .A(n657), .Y(n2767) );
  AND2X1 U1889 ( .A(mem[249]), .B(n4541), .Y(n645) );
  INVX1 U1891 ( .A(n645), .Y(n2768) );
  AND2X1 U1893 ( .A(mem[229]), .B(n4542), .Y(n623) );
  INVX1 U1895 ( .A(n623), .Y(n2769) );
  AND2X1 U1899 ( .A(mem[217]), .B(n4542), .Y(n611) );
  INVX1 U1901 ( .A(n611), .Y(n2770) );
  AND2X1 U1903 ( .A(mem[193]), .B(n4543), .Y(n585) );
  INVX1 U1905 ( .A(n585), .Y(n2771) );
  AND2X1 U1907 ( .A(mem[181]), .B(n4543), .Y(n573) );
  INVX1 U1909 ( .A(n573), .Y(n2772) );
  AND2X1 U1911 ( .A(mem[161]), .B(n4544), .Y(n551) );
  INVX1 U1913 ( .A(n551), .Y(n2773) );
  AND2X1 U1915 ( .A(mem[149]), .B(n4544), .Y(n539) );
  INVX1 U1917 ( .A(n539), .Y(n2774) );
  AND2X1 U1919 ( .A(mem[125]), .B(n4545), .Y(n513) );
  INVX1 U1921 ( .A(n513), .Y(n2775) );
  AND2X1 U1923 ( .A(mem[113]), .B(n4545), .Y(n501) );
  INVX1 U1925 ( .A(n501), .Y(n2776) );
  AND2X1 U1927 ( .A(mem[93]), .B(n4546), .Y(n479) );
  INVX1 U1929 ( .A(n479), .Y(n2777) );
  AND2X1 U1931 ( .A(mem[81]), .B(n4546), .Y(n467) );
  INVX1 U1933 ( .A(n467), .Y(n2778) );
  AND2X1 U1935 ( .A(mem[57]), .B(n4547), .Y(n441) );
  INVX1 U1937 ( .A(n441), .Y(n2779) );
  AND2X1 U1939 ( .A(mem[45]), .B(n4547), .Y(n429) );
  INVX1 U1941 ( .A(n429), .Y(n2780) );
  AND2X1 U1943 ( .A(mem[25]), .B(n4548), .Y(n399) );
  INVX1 U1945 ( .A(n399), .Y(n2781) );
  AND2X1 U1947 ( .A(mem[13]), .B(n4548), .Y(n375) );
  INVX1 U1949 ( .A(n375), .Y(n2782) );
  AND2X1 U1951 ( .A(n4619), .B(n1484), .Y(n1529) );
  INVX1 U1953 ( .A(n1529), .Y(n2783) );
  AND2X1 U1955 ( .A(mem[1027]), .B(n4517), .Y(n1451) );
  INVX1 U1957 ( .A(n1451), .Y(n2784) );
  AND2X1 U1959 ( .A(mem[1026]), .B(n4517), .Y(n1450) );
  INVX1 U1961 ( .A(n1450), .Y(n2785) );
  AND2X1 U1963 ( .A(mem[998]), .B(n4518), .Y(n1421) );
  INVX1 U1967 ( .A(n1421), .Y(n2786) );
  AND2X1 U1969 ( .A(mem[992]), .B(n4518), .Y(n1415) );
  INVX1 U1971 ( .A(n1415), .Y(n2787) );
  AND2X1 U1973 ( .A(mem[963]), .B(n4519), .Y(n1385) );
  INVX1 U1975 ( .A(n1385), .Y(n2788) );
  AND2X1 U1977 ( .A(mem[958]), .B(n4519), .Y(n1380) );
  INVX1 U1979 ( .A(n1380), .Y(n2789) );
  AND2X1 U1981 ( .A(mem[929]), .B(n4520), .Y(n1350) );
  INVX1 U1983 ( .A(n1350), .Y(n2790) );
  AND2X1 U1985 ( .A(mem[924]), .B(n4520), .Y(n1345) );
  INVX1 U1987 ( .A(n1345), .Y(n2791) );
  AND2X1 U1989 ( .A(mem[922]), .B(n4521), .Y(n1342) );
  INVX1 U1991 ( .A(n1342), .Y(n2792) );
  AND2X1 U1993 ( .A(mem[910]), .B(n4521), .Y(n1330) );
  INVX1 U1995 ( .A(n1330), .Y(n2793) );
  AND2X1 U1997 ( .A(mem[888]), .B(n4522), .Y(n1307) );
  INVX1 U1999 ( .A(n1307), .Y(n2794) );
  AND2X1 U2001 ( .A(mem[876]), .B(n4522), .Y(n1295) );
  INVX1 U2003 ( .A(n1295), .Y(n2795) );
  AND2X1 U2005 ( .A(mem[854]), .B(n4523), .Y(n1272) );
  INVX1 U2007 ( .A(n1272), .Y(n2796) );
  AND2X1 U2009 ( .A(mem[842]), .B(n4523), .Y(n1260) );
  INVX1 U2011 ( .A(n1260), .Y(n2797) );
  AND2X1 U2013 ( .A(mem[820]), .B(n4524), .Y(n1236) );
  INVX1 U2015 ( .A(n1236), .Y(n2798) );
  AND2X1 U2017 ( .A(mem[808]), .B(n4524), .Y(n1224) );
  INVX1 U2019 ( .A(n1224), .Y(n2799) );
  AND2X1 U2021 ( .A(mem[786]), .B(n4525), .Y(n1201) );
  INVX1 U2023 ( .A(n1201), .Y(n2800) );
  AND2X1 U2025 ( .A(mem[774]), .B(n4525), .Y(n1189) );
  INVX1 U2027 ( .A(n1189), .Y(n2801) );
  AND2X1 U2029 ( .A(mem[752]), .B(n4526), .Y(n1166) );
  INVX1 U2031 ( .A(n1166), .Y(n2802) );
  AND2X1 U2035 ( .A(mem[740]), .B(n4526), .Y(n1154) );
  INVX1 U2037 ( .A(n1154), .Y(n2803) );
  AND2X1 U2039 ( .A(mem[718]), .B(n4527), .Y(n1131) );
  INVX1 U2041 ( .A(n1131), .Y(n2804) );
  AND2X1 U2043 ( .A(mem[706]), .B(n4527), .Y(n1119) );
  INVX1 U2045 ( .A(n1119), .Y(n2805) );
  AND2X1 U2047 ( .A(mem[684]), .B(n4528), .Y(n1096) );
  INVX1 U2049 ( .A(n1096), .Y(n2806) );
  AND2X1 U2051 ( .A(mem[672]), .B(n4528), .Y(n1084) );
  INVX1 U2053 ( .A(n1084), .Y(n2807) );
  AND2X1 U2055 ( .A(mem[631]), .B(n4529), .Y(n1042) );
  INVX1 U2057 ( .A(n1042), .Y(n2808) );
  AND2X1 U2059 ( .A(mem[630]), .B(n4529), .Y(n1041) );
  INVX1 U2061 ( .A(n1041), .Y(n2809) );
  AND2X1 U2063 ( .A(mem[602]), .B(n4530), .Y(n1012) );
  INVX1 U2065 ( .A(n1012), .Y(n2810) );
  AND2X1 U2067 ( .A(mem[596]), .B(n4530), .Y(n1006) );
  INVX1 U2069 ( .A(n1006), .Y(n2811) );
  AND2X1 U2071 ( .A(mem[567]), .B(n4531), .Y(n976) );
  INVX1 U2073 ( .A(n976), .Y(n2812) );
  AND2X1 U2075 ( .A(mem[562]), .B(n4531), .Y(n971) );
  INVX1 U2077 ( .A(n971), .Y(n2813) );
  AND2X1 U2079 ( .A(mem[533]), .B(n4532), .Y(n940) );
  INVX1 U2081 ( .A(n940), .Y(n2814) );
  AND2X1 U2083 ( .A(mem[528]), .B(n4532), .Y(n935) );
  INVX1 U2085 ( .A(n935), .Y(n2815) );
  AND2X1 U2087 ( .A(mem[526]), .B(n4533), .Y(n932) );
  INVX1 U2089 ( .A(n932), .Y(n2816) );
  AND2X1 U2091 ( .A(mem[514]), .B(n4533), .Y(n920) );
  INVX1 U2093 ( .A(n920), .Y(n2817) );
  AND2X1 U2095 ( .A(mem[492]), .B(n4534), .Y(n897) );
  INVX1 U2097 ( .A(n897), .Y(n2818) );
  AND2X1 U2099 ( .A(mem[480]), .B(n4534), .Y(n885) );
  INVX1 U2103 ( .A(n885), .Y(n2819) );
  AND2X1 U2105 ( .A(mem[458]), .B(n4535), .Y(n862) );
  INVX1 U2107 ( .A(n862), .Y(n2820) );
  AND2X1 U2109 ( .A(mem[446]), .B(n4535), .Y(n850) );
  INVX1 U2111 ( .A(n850), .Y(n2821) );
  AND2X1 U2113 ( .A(mem[424]), .B(n4536), .Y(n827) );
  INVX1 U2115 ( .A(n827), .Y(n2822) );
  AND2X1 U2117 ( .A(mem[412]), .B(n4536), .Y(n815) );
  INVX1 U2119 ( .A(n815), .Y(n2823) );
  AND2X1 U2121 ( .A(mem[390]), .B(n4537), .Y(n792) );
  INVX1 U2123 ( .A(n792), .Y(n2824) );
  AND2X1 U2125 ( .A(mem[378]), .B(n4537), .Y(n780) );
  INVX1 U2127 ( .A(n780), .Y(n2825) );
  AND2X1 U2129 ( .A(mem[356]), .B(n4538), .Y(n757) );
  INVX1 U2131 ( .A(n757), .Y(n2826) );
  AND2X1 U2133 ( .A(mem[344]), .B(n4538), .Y(n745) );
  INVX1 U2135 ( .A(n745), .Y(n2827) );
  AND2X1 U2137 ( .A(mem[322]), .B(n4539), .Y(n722) );
  INVX1 U2139 ( .A(n722), .Y(n2828) );
  AND2X1 U2141 ( .A(mem[310]), .B(n4539), .Y(n710) );
  INVX1 U2143 ( .A(n710), .Y(n2829) );
  AND2X1 U2145 ( .A(mem[288]), .B(n4540), .Y(n686) );
  INVX1 U2147 ( .A(n686), .Y(n2830) );
  AND2X1 U2149 ( .A(mem[276]), .B(n4540), .Y(n674) );
  INVX1 U2151 ( .A(n674), .Y(n2831) );
  AND2X1 U2153 ( .A(mem[262]), .B(n4541), .Y(n658) );
  INVX1 U2155 ( .A(n658), .Y(n2832) );
  AND2X1 U2157 ( .A(mem[250]), .B(n4541), .Y(n646) );
  INVX1 U2159 ( .A(n646), .Y(n2833) );
  AND2X1 U2161 ( .A(mem[228]), .B(n4542), .Y(n622) );
  INVX1 U2163 ( .A(n622), .Y(n2834) );
  AND2X1 U2165 ( .A(mem[216]), .B(n4542), .Y(n610) );
  INVX1 U2167 ( .A(n610), .Y(n2835) );
  AND2X1 U2171 ( .A(mem[194]), .B(n4543), .Y(n586) );
  INVX1 U2172 ( .A(n586), .Y(n2836) );
  AND2X1 U2174 ( .A(mem[182]), .B(n4543), .Y(n574) );
  INVX1 U2175 ( .A(n574), .Y(n2837) );
  AND2X1 U2177 ( .A(mem[160]), .B(n4544), .Y(n550) );
  INVX1 U2178 ( .A(n550), .Y(n2838) );
  AND2X1 U2180 ( .A(mem[148]), .B(n4544), .Y(n538) );
  INVX1 U2181 ( .A(n538), .Y(n2839) );
  AND2X1 U2183 ( .A(mem[126]), .B(n4545), .Y(n514) );
  INVX1 U2184 ( .A(n514), .Y(n2840) );
  AND2X1 U2186 ( .A(mem[114]), .B(n4545), .Y(n502) );
  INVX1 U2187 ( .A(n502), .Y(n2841) );
  AND2X1 U2189 ( .A(mem[92]), .B(n4546), .Y(n478) );
  INVX1 U2190 ( .A(n478), .Y(n2842) );
  AND2X1 U2192 ( .A(mem[80]), .B(n4546), .Y(n466) );
  INVX1 U2193 ( .A(n466), .Y(n2843) );
  AND2X1 U2195 ( .A(mem[58]), .B(n4547), .Y(n442) );
  INVX1 U2196 ( .A(n442), .Y(n2844) );
  AND2X1 U2198 ( .A(mem[46]), .B(n4547), .Y(n430) );
  INVX1 U2199 ( .A(n430), .Y(n2845) );
  AND2X1 U2201 ( .A(mem[24]), .B(n4548), .Y(n397) );
  INVX1 U2202 ( .A(n397), .Y(n2846) );
  AND2X1 U2204 ( .A(mem[12]), .B(n4548), .Y(n373) );
  INVX1 U2205 ( .A(n373), .Y(n2847) );
  AND2X1 U2207 ( .A(mem[1051]), .B(n4517), .Y(n1475) );
  INVX1 U2208 ( .A(n1475), .Y(n2848) );
  AND2X1 U2210 ( .A(mem[1039]), .B(n4517), .Y(n1463) );
  INVX1 U2211 ( .A(n1463), .Y(n2849) );
  AND2X1 U2213 ( .A(mem[1019]), .B(n4518), .Y(n1442) );
  INVX1 U2214 ( .A(n1442), .Y(n2850) );
  AND2X1 U2216 ( .A(mem[1007]), .B(n4518), .Y(n1430) );
  INVX1 U2217 ( .A(n1430), .Y(n2851) );
  AND2X1 U2219 ( .A(mem[987]), .B(n4519), .Y(n1409) );
  INVX1 U2220 ( .A(n1409), .Y(n2852) );
  AND2X1 U2222 ( .A(mem[975]), .B(n4519), .Y(n1397) );
  INVX1 U2223 ( .A(n1397), .Y(n2853) );
  AND2X1 U2225 ( .A(mem[955]), .B(n4520), .Y(n1376) );
  INVX1 U2226 ( .A(n1376), .Y(n2854) );
  AND2X1 U2228 ( .A(mem[943]), .B(n4520), .Y(n1364) );
  INVX1 U2229 ( .A(n1364), .Y(n2855) );
  AND2X1 U2231 ( .A(mem[896]), .B(n4521), .Y(n1316) );
  INVX1 U2232 ( .A(n1316), .Y(n2856) );
  AND2X1 U2234 ( .A(mem[891]), .B(n4521), .Y(n1311) );
  INVX1 U2235 ( .A(n1311), .Y(n2857) );
  AND2X1 U2237 ( .A(mem[864]), .B(n4522), .Y(n1283) );
  INVX1 U2238 ( .A(n1283), .Y(n2858) );
  AND2X1 U2240 ( .A(mem[859]), .B(n4522), .Y(n1278) );
  INVX1 U2241 ( .A(n1278), .Y(n2859) );
  AND2X1 U2243 ( .A(mem[833]), .B(n4523), .Y(n1251) );
  INVX1 U2244 ( .A(n1251), .Y(n2860) );
  AND2X1 U2246 ( .A(mem[827]), .B(n4523), .Y(n1245) );
  INVX1 U2247 ( .A(n1245), .Y(n2861) );
  AND2X1 U2249 ( .A(mem[796]), .B(n4524), .Y(n1212) );
  INVX1 U2250 ( .A(n1212), .Y(n2862) );
  AND2X1 U2252 ( .A(mem[795]), .B(n4524), .Y(n1211) );
  INVX1 U2253 ( .A(n1211), .Y(n2863) );
  AND2X1 U2255 ( .A(mem[779]), .B(n4525), .Y(n1194) );
  INVX1 U2256 ( .A(n1194), .Y(n2864) );
  AND2X1 U2258 ( .A(mem[766]), .B(n4525), .Y(n1181) );
  INVX1 U2259 ( .A(n1181), .Y(n2865) );
  AND2X1 U2261 ( .A(mem[747]), .B(n4526), .Y(n1161) );
  INVX1 U2262 ( .A(n1161), .Y(n2866) );
  AND2X1 U2264 ( .A(mem[735]), .B(n4526), .Y(n1149) );
  INVX1 U2265 ( .A(n1149), .Y(n2867) );
  AND2X1 U2267 ( .A(mem[715]), .B(n4527), .Y(n1128) );
  INVX1 U2268 ( .A(n1128), .Y(n2868) );
  AND2X1 U2273 ( .A(mem[703]), .B(n4527), .Y(n1116) );
  INVX1 U2275 ( .A(n1116), .Y(n2869) );
  AND2X1 U2277 ( .A(mem[683]), .B(n4528), .Y(n1095) );
  INVX1 U2279 ( .A(n1095), .Y(n2870) );
  AND2X1 U2281 ( .A(mem[671]), .B(n4528), .Y(n1083) );
  INVX1 U2283 ( .A(n1083), .Y(n2871) );
  AND2X1 U2285 ( .A(mem[655]), .B(n4529), .Y(n1066) );
  INVX1 U2287 ( .A(n1066), .Y(n2872) );
  AND2X1 U2289 ( .A(mem[643]), .B(n4529), .Y(n1054) );
  INVX1 U2323 ( .A(n1054), .Y(n2873) );
  AND2X1 U2324 ( .A(mem[623]), .B(n4530), .Y(n1033) );
  INVX1 U2326 ( .A(n1033), .Y(n2874) );
  AND2X1 U2327 ( .A(mem[611]), .B(n4530), .Y(n1021) );
  INVX1 U2328 ( .A(n1021), .Y(n2875) );
  AND2X1 U2331 ( .A(mem[591]), .B(n4531), .Y(n1000) );
  INVX1 U2339 ( .A(n1000), .Y(n2876) );
  AND2X1 U2340 ( .A(mem[579]), .B(n4531), .Y(n988) );
  INVX1 U2341 ( .A(n988), .Y(n2877) );
  AND2X1 U2342 ( .A(mem[559]), .B(n4532), .Y(n966) );
  INVX1 U2343 ( .A(n966), .Y(n2878) );
  AND2X1 U2344 ( .A(mem[547]), .B(n4532), .Y(n954) );
  INVX1 U2345 ( .A(n954), .Y(n2879) );
  AND2X1 U2346 ( .A(mem[500]), .B(n4533), .Y(n906) );
  INVX1 U2347 ( .A(n906), .Y(n2880) );
  AND2X1 U2348 ( .A(mem[495]), .B(n4533), .Y(n901) );
  INVX1 U2349 ( .A(n901), .Y(n2881) );
  AND2X1 U2350 ( .A(mem[468]), .B(n4534), .Y(n873) );
  INVX1 U2351 ( .A(n873), .Y(n2882) );
  AND2X1 U2352 ( .A(mem[463]), .B(n4534), .Y(n868) );
  INVX1 U2353 ( .A(n868), .Y(n2883) );
  AND2X1 U2354 ( .A(mem[437]), .B(n4535), .Y(n841) );
  INVX1 U2355 ( .A(n841), .Y(n2884) );
  AND2X1 U2356 ( .A(mem[431]), .B(n4535), .Y(n835) );
  INVX1 U2357 ( .A(n835), .Y(n2885) );
  AND2X1 U2358 ( .A(mem[400]), .B(n4536), .Y(n803) );
  INVX1 U2359 ( .A(n803), .Y(n2886) );
  AND2X1 U2360 ( .A(mem[399]), .B(n4536), .Y(n802) );
  INVX1 U2361 ( .A(n802), .Y(n2887) );
  AND2X1 U2362 ( .A(mem[383]), .B(n4537), .Y(n785) );
  INVX1 U2363 ( .A(n785), .Y(n2888) );
  AND2X1 U2364 ( .A(mem[370]), .B(n4537), .Y(n772) );
  INVX1 U2365 ( .A(n772), .Y(n2889) );
  AND2X1 U2366 ( .A(mem[351]), .B(n4538), .Y(n752) );
  INVX1 U2367 ( .A(n752), .Y(n2890) );
  AND2X1 U2368 ( .A(mem[339]), .B(n4538), .Y(n740) );
  INVX1 U2369 ( .A(n740), .Y(n2891) );
  AND2X1 U2370 ( .A(mem[319]), .B(n4539), .Y(n719) );
  INVX1 U2371 ( .A(n719), .Y(n2892) );
  AND2X1 U2372 ( .A(mem[307]), .B(n4539), .Y(n707) );
  INVX1 U2373 ( .A(n707), .Y(n2893) );
  AND2X1 U2374 ( .A(mem[287]), .B(n4540), .Y(n685) );
  INVX1 U2375 ( .A(n685), .Y(n2894) );
  AND2X1 U2376 ( .A(mem[275]), .B(n4540), .Y(n673) );
  INVX1 U2377 ( .A(n673), .Y(n2895) );
  AND2X1 U2378 ( .A(mem[236]), .B(n4541), .Y(n632) );
  INVX1 U2379 ( .A(n632), .Y(n2896) );
  AND2X1 U2380 ( .A(mem[231]), .B(n4541), .Y(n627) );
  INVX1 U2381 ( .A(n627), .Y(n2897) );
  AND2X1 U2382 ( .A(mem[204]), .B(n4542), .Y(n598) );
  INVX1 U2383 ( .A(n598), .Y(n2898) );
  AND2X1 U2384 ( .A(mem[199]), .B(n4542), .Y(n593) );
  INVX1 U2385 ( .A(n593), .Y(n2899) );
  AND2X1 U2386 ( .A(mem[173]), .B(n4543), .Y(n565) );
  INVX1 U2387 ( .A(n565), .Y(n2900) );
  AND2X1 U2388 ( .A(mem[167]), .B(n4543), .Y(n559) );
  INVX1 U2389 ( .A(n559), .Y(n2901) );
  AND2X1 U2390 ( .A(mem[136]), .B(n4544), .Y(n526) );
  INVX1 U2391 ( .A(n526), .Y(n2902) );
  AND2X1 U2392 ( .A(mem[135]), .B(n4544), .Y(n525) );
  INVX1 U2393 ( .A(n525), .Y(n2903) );
  AND2X1 U2394 ( .A(mem[119]), .B(n4545), .Y(n507) );
  INVX1 U2395 ( .A(n507), .Y(n2904) );
  AND2X1 U2396 ( .A(mem[106]), .B(n4545), .Y(n494) );
  INVX1 U2397 ( .A(n494), .Y(n2905) );
  AND2X1 U2398 ( .A(mem[87]), .B(n4546), .Y(n473) );
  INVX1 U2399 ( .A(n473), .Y(n2906) );
  AND2X1 U2400 ( .A(mem[75]), .B(n4546), .Y(n461) );
  INVX1 U2401 ( .A(n461), .Y(n2907) );
  AND2X1 U2402 ( .A(mem[55]), .B(n4547), .Y(n439) );
  INVX1 U2403 ( .A(n439), .Y(n2908) );
  AND2X1 U2404 ( .A(mem[43]), .B(n4547), .Y(n427) );
  INVX1 U2405 ( .A(n427), .Y(n2909) );
  AND2X1 U2406 ( .A(mem[23]), .B(n4548), .Y(n395) );
  INVX1 U2407 ( .A(n395), .Y(n2910) );
  AND2X1 U2408 ( .A(mem[11]), .B(n4548), .Y(n371) );
  INVX1 U2409 ( .A(n371), .Y(n2911) );
  BUFX2 U2410 ( .A(n556), .Y(n2912) );
  BUFX2 U2411 ( .A(n521), .Y(n2913) );
  AND2X1 U2412 ( .A(n23), .B(n1484), .Y(n1487) );
  INVX1 U2413 ( .A(n1487), .Y(n2914) );
  AND2X1 U2414 ( .A(mem[1052]), .B(n4517), .Y(n1476) );
  INVX1 U2415 ( .A(n1476), .Y(n2915) );
  AND2X1 U2416 ( .A(mem[1040]), .B(n4517), .Y(n1464) );
  INVX1 U2417 ( .A(n1464), .Y(n2916) );
  AND2X1 U2418 ( .A(mem[1018]), .B(n4518), .Y(n1441) );
  INVX1 U2419 ( .A(n1441), .Y(n2917) );
  AND2X1 U2420 ( .A(mem[1006]), .B(n4518), .Y(n1429) );
  INVX1 U2421 ( .A(n1429), .Y(n2918) );
  AND2X1 U2422 ( .A(mem[988]), .B(n4519), .Y(n1410) );
  INVX1 U2423 ( .A(n1410), .Y(n2919) );
  AND2X1 U2424 ( .A(mem[976]), .B(n4519), .Y(n1398) );
  INVX1 U2425 ( .A(n1398), .Y(n2920) );
  AND2X1 U2426 ( .A(mem[954]), .B(n4520), .Y(n1375) );
  INVX1 U2427 ( .A(n1375), .Y(n2921) );
  AND2X1 U2428 ( .A(mem[942]), .B(n4520), .Y(n1363) );
  INVX1 U2429 ( .A(n1363), .Y(n2922) );
  AND2X1 U2430 ( .A(mem[897]), .B(n4521), .Y(n1317) );
  INVX1 U2431 ( .A(n1317), .Y(n2923) );
  AND2X1 U2432 ( .A(mem[892]), .B(n4521), .Y(n1312) );
  INVX1 U2433 ( .A(n1312), .Y(n2924) );
  AND2X1 U2434 ( .A(mem[863]), .B(n4522), .Y(n1282) );
  INVX1 U2435 ( .A(n1282), .Y(n2925) );
  AND2X1 U2436 ( .A(mem[858]), .B(n4522), .Y(n1277) );
  INVX1 U2437 ( .A(n1277), .Y(n2926) );
  AND2X1 U2438 ( .A(mem[829]), .B(n4523), .Y(n1247) );
  INVX1 U2439 ( .A(n1247), .Y(n2927) );
  AND2X1 U2440 ( .A(mem[828]), .B(n4523), .Y(n1246) );
  INVX1 U2441 ( .A(n1246), .Y(n2928) );
  AND2X1 U2442 ( .A(mem[800]), .B(n4524), .Y(n1216) );
  INVX1 U2443 ( .A(n1216), .Y(n2929) );
  AND2X1 U2444 ( .A(mem[794]), .B(n4524), .Y(n1210) );
  INVX1 U2445 ( .A(n1210), .Y(n2930) );
  AND2X1 U2446 ( .A(mem[780]), .B(n4525), .Y(n1195) );
  INVX1 U2447 ( .A(n1195), .Y(n2931) );
  AND2X1 U2448 ( .A(mem[768]), .B(n4525), .Y(n1183) );
  INVX1 U2449 ( .A(n1183), .Y(n2932) );
  AND2X1 U2450 ( .A(mem[746]), .B(n4526), .Y(n1160) );
  INVX1 U2451 ( .A(n1160), .Y(n2933) );
  AND2X1 U2452 ( .A(mem[733]), .B(n4526), .Y(n1147) );
  INVX1 U2453 ( .A(n1147), .Y(n2934) );
  AND2X1 U2454 ( .A(mem[716]), .B(n4527), .Y(n1129) );
  INVX1 U2455 ( .A(n1129), .Y(n2935) );
  AND2X1 U2456 ( .A(mem[704]), .B(n4527), .Y(n1117) );
  INVX1 U2457 ( .A(n1117), .Y(n2936) );
  AND2X1 U2458 ( .A(mem[682]), .B(n4528), .Y(n1094) );
  INVX1 U2459 ( .A(n1094), .Y(n2937) );
  AND2X1 U2460 ( .A(mem[670]), .B(n4528), .Y(n1082) );
  INVX1 U2461 ( .A(n1082), .Y(n2938) );
  AND2X1 U2462 ( .A(mem[656]), .B(n4529), .Y(n1067) );
  INVX1 U2463 ( .A(n1067), .Y(n2939) );
  AND2X1 U2464 ( .A(mem[644]), .B(n4529), .Y(n1055) );
  INVX1 U2465 ( .A(n1055), .Y(n2940) );
  AND2X1 U2466 ( .A(mem[622]), .B(n4530), .Y(n1032) );
  INVX1 U2467 ( .A(n1032), .Y(n2941) );
  AND2X1 U2468 ( .A(mem[610]), .B(n4530), .Y(n1020) );
  INVX1 U2469 ( .A(n1020), .Y(n2942) );
  AND2X1 U2470 ( .A(mem[592]), .B(n4531), .Y(n1001) );
  INVX1 U2471 ( .A(n1001), .Y(n2943) );
  AND2X1 U2472 ( .A(mem[580]), .B(n4531), .Y(n989) );
  INVX1 U2473 ( .A(n989), .Y(n2944) );
  AND2X1 U2474 ( .A(mem[558]), .B(n4532), .Y(n965) );
  INVX1 U2475 ( .A(n965), .Y(n2945) );
  AND2X1 U2476 ( .A(mem[546]), .B(n4532), .Y(n953) );
  INVX1 U2477 ( .A(n953), .Y(n2946) );
  AND2X1 U2478 ( .A(mem[501]), .B(n4533), .Y(n907) );
  INVX1 U2479 ( .A(n907), .Y(n2947) );
  AND2X1 U2480 ( .A(mem[496]), .B(n4533), .Y(n902) );
  INVX1 U2481 ( .A(n902), .Y(n2948) );
  AND2X1 U2482 ( .A(mem[467]), .B(n4534), .Y(n872) );
  INVX1 U2483 ( .A(n872), .Y(n2949) );
  AND2X1 U2484 ( .A(mem[462]), .B(n4534), .Y(n867) );
  INVX1 U2485 ( .A(n867), .Y(n2950) );
  AND2X1 U2486 ( .A(mem[433]), .B(n4535), .Y(n837) );
  INVX1 U2487 ( .A(n837), .Y(n2951) );
  AND2X1 U2488 ( .A(mem[432]), .B(n4535), .Y(n836) );
  INVX1 U2489 ( .A(n836), .Y(n2952) );
  AND2X1 U2490 ( .A(mem[404]), .B(n4536), .Y(n807) );
  INVX1 U2491 ( .A(n807), .Y(n2953) );
  AND2X1 U2492 ( .A(mem[398]), .B(n4536), .Y(n801) );
  INVX1 U2493 ( .A(n801), .Y(n2954) );
  AND2X1 U2494 ( .A(mem[384]), .B(n4537), .Y(n786) );
  INVX1 U2495 ( .A(n786), .Y(n2955) );
  AND2X1 U2496 ( .A(mem[372]), .B(n4537), .Y(n774) );
  INVX1 U2497 ( .A(n774), .Y(n2956) );
  AND2X1 U2498 ( .A(mem[350]), .B(n4538), .Y(n751) );
  INVX1 U2499 ( .A(n751), .Y(n2957) );
  AND2X1 U2500 ( .A(mem[337]), .B(n4538), .Y(n738) );
  INVX1 U2501 ( .A(n738), .Y(n2958) );
  AND2X1 U2502 ( .A(mem[320]), .B(n4539), .Y(n720) );
  INVX1 U2503 ( .A(n720), .Y(n2959) );
  AND2X1 U2504 ( .A(mem[308]), .B(n4539), .Y(n708) );
  INVX1 U2505 ( .A(n708), .Y(n2960) );
  AND2X1 U2506 ( .A(mem[286]), .B(n4540), .Y(n684) );
  INVX1 U2507 ( .A(n684), .Y(n2961) );
  AND2X1 U2508 ( .A(mem[274]), .B(n4540), .Y(n672) );
  INVX1 U2509 ( .A(n672), .Y(n2962) );
  AND2X1 U2510 ( .A(mem[237]), .B(n4541), .Y(n633) );
  INVX1 U2511 ( .A(n633), .Y(n2963) );
  AND2X1 U2512 ( .A(mem[232]), .B(n4541), .Y(n628) );
  INVX1 U2513 ( .A(n628), .Y(n2964) );
  AND2X1 U2514 ( .A(mem[203]), .B(n4542), .Y(n597) );
  INVX1 U2515 ( .A(n597), .Y(n2965) );
  AND2X1 U2516 ( .A(mem[198]), .B(n4542), .Y(n592) );
  INVX1 U2517 ( .A(n592), .Y(n2966) );
  AND2X1 U2518 ( .A(mem[169]), .B(n4543), .Y(n561) );
  INVX1 U2519 ( .A(n561), .Y(n2967) );
  AND2X1 U2520 ( .A(mem[168]), .B(n4543), .Y(n560) );
  INVX1 U2521 ( .A(n560), .Y(n2968) );
  AND2X1 U2522 ( .A(mem[140]), .B(n4544), .Y(n530) );
  INVX1 U2523 ( .A(n530), .Y(n2969) );
  AND2X1 U2524 ( .A(mem[134]), .B(n4544), .Y(n524) );
  INVX1 U2525 ( .A(n524), .Y(n2970) );
  AND2X1 U2526 ( .A(mem[120]), .B(n4545), .Y(n508) );
  INVX1 U2527 ( .A(n508), .Y(n2971) );
  AND2X1 U2528 ( .A(mem[108]), .B(n4545), .Y(n496) );
  INVX1 U2529 ( .A(n496), .Y(n2972) );
  AND2X1 U2530 ( .A(mem[86]), .B(n4546), .Y(n472) );
  INVX1 U2531 ( .A(n472), .Y(n2973) );
  AND2X1 U2532 ( .A(mem[73]), .B(n4546), .Y(n459) );
  INVX1 U2533 ( .A(n459), .Y(n2974) );
  AND2X1 U2534 ( .A(mem[56]), .B(n4547), .Y(n440) );
  INVX1 U2535 ( .A(n440), .Y(n2975) );
  AND2X1 U2536 ( .A(mem[44]), .B(n4547), .Y(n428) );
  INVX1 U2537 ( .A(n428), .Y(n2976) );
  AND2X1 U2538 ( .A(mem[22]), .B(n4548), .Y(n393) );
  INVX1 U2539 ( .A(n393), .Y(n2977) );
  AND2X1 U2540 ( .A(mem[10]), .B(n4548), .Y(n369) );
  INVX1 U2541 ( .A(n369), .Y(n2978) );
  BUFX2 U2542 ( .A(n591), .Y(n2979) );
  BUFX2 U2543 ( .A(n486), .Y(n2980) );
  AND2X1 U2544 ( .A(n93), .B(n1490), .Y(n1494) );
  INVX1 U2545 ( .A(n1494), .Y(n2981) );
  AND2X1 U2546 ( .A(n22), .B(n1484), .Y(n1483) );
  INVX1 U2547 ( .A(n1483), .Y(n2982) );
  AND2X1 U2548 ( .A(mem[1053]), .B(n4517), .Y(n1477) );
  INVX1 U2549 ( .A(n1477), .Y(n2983) );
  AND2X1 U2550 ( .A(mem[1041]), .B(n4517), .Y(n1465) );
  INVX1 U2551 ( .A(n1465), .Y(n2984) );
  AND2X1 U2552 ( .A(mem[1021]), .B(n4518), .Y(n1444) );
  INVX1 U2553 ( .A(n1444), .Y(n2985) );
  AND2X1 U2554 ( .A(mem[1009]), .B(n4518), .Y(n1432) );
  INVX1 U2555 ( .A(n1432), .Y(n2986) );
  AND2X1 U2556 ( .A(mem[985]), .B(n4519), .Y(n1407) );
  INVX1 U2557 ( .A(n1407), .Y(n2987) );
  AND2X1 U2558 ( .A(mem[973]), .B(n4519), .Y(n1395) );
  INVX1 U2559 ( .A(n1395), .Y(n2988) );
  AND2X1 U2560 ( .A(mem[953]), .B(n4520), .Y(n1374) );
  INVX1 U2561 ( .A(n1374), .Y(n2989) );
  AND2X1 U2562 ( .A(mem[941]), .B(n4520), .Y(n1362) );
  INVX1 U2563 ( .A(n1362), .Y(n2990) );
  AND2X1 U2564 ( .A(mem[899]), .B(n4521), .Y(n1319) );
  INVX1 U2565 ( .A(n1319), .Y(n2991) );
  AND2X1 U2566 ( .A(mem[893]), .B(n4521), .Y(n1313) );
  INVX1 U2567 ( .A(n1313), .Y(n2992) );
  AND2X1 U2568 ( .A(mem[862]), .B(n4522), .Y(n1281) );
  INVX1 U2569 ( .A(n1281), .Y(n2993) );
  AND2X1 U2570 ( .A(mem[861]), .B(n4522), .Y(n1280) );
  INVX1 U2571 ( .A(n1280), .Y(n2994) );
  AND2X1 U2572 ( .A(mem[830]), .B(n4523), .Y(n1248) );
  INVX1 U2573 ( .A(n1248), .Y(n2995) );
  AND2X1 U2574 ( .A(mem[825]), .B(n4523), .Y(n1243) );
  INVX1 U2575 ( .A(n1243), .Y(n2996) );
  AND2X1 U2576 ( .A(mem[798]), .B(n4524), .Y(n1214) );
  INVX1 U2577 ( .A(n1214), .Y(n2997) );
  AND2X1 U2578 ( .A(mem[793]), .B(n4524), .Y(n1209) );
  INVX1 U2579 ( .A(n1209), .Y(n2998) );
  AND2X1 U2580 ( .A(mem[781]), .B(n4525), .Y(n1196) );
  INVX1 U2581 ( .A(n1196), .Y(n2999) );
  AND2X1 U2582 ( .A(mem[769]), .B(n4525), .Y(n1184) );
  INVX1 U2583 ( .A(n1184), .Y(n3000) );
  AND2X1 U2584 ( .A(mem[749]), .B(n4526), .Y(n1163) );
  INVX1 U2585 ( .A(n1163), .Y(n3001) );
  AND2X1 U2586 ( .A(mem[737]), .B(n4526), .Y(n1151) );
  INVX1 U2587 ( .A(n1151), .Y(n3002) );
  AND2X1 U2588 ( .A(mem[713]), .B(n4527), .Y(n1126) );
  INVX1 U2589 ( .A(n1126), .Y(n3003) );
  AND2X1 U2590 ( .A(mem[700]), .B(n4527), .Y(n1113) );
  INVX1 U2591 ( .A(n1113), .Y(n3004) );
  AND2X1 U2592 ( .A(mem[681]), .B(n4528), .Y(n1093) );
  INVX1 U2593 ( .A(n1093), .Y(n3005) );
  AND2X1 U2594 ( .A(mem[669]), .B(n4528), .Y(n1081) );
  INVX1 U2595 ( .A(n1081), .Y(n3006) );
  AND2X1 U2596 ( .A(mem[657]), .B(n4529), .Y(n1068) );
  INVX1 U2597 ( .A(n1068), .Y(n3007) );
  AND2X1 U2598 ( .A(mem[645]), .B(n4529), .Y(n1056) );
  INVX1 U2599 ( .A(n1056), .Y(n3008) );
  AND2X1 U2600 ( .A(mem[625]), .B(n4530), .Y(n1035) );
  INVX1 U2601 ( .A(n1035), .Y(n3009) );
  AND2X1 U2602 ( .A(mem[613]), .B(n4530), .Y(n1023) );
  INVX1 U2603 ( .A(n1023), .Y(n3010) );
  AND2X1 U2604 ( .A(mem[589]), .B(n4531), .Y(n998) );
  INVX1 U2605 ( .A(n998), .Y(n3011) );
  AND2X1 U2606 ( .A(mem[577]), .B(n4531), .Y(n986) );
  INVX1 U2607 ( .A(n986), .Y(n3012) );
  AND2X1 U2608 ( .A(mem[557]), .B(n4532), .Y(n964) );
  INVX1 U2609 ( .A(n964), .Y(n3013) );
  AND2X1 U2610 ( .A(mem[545]), .B(n4532), .Y(n952) );
  INVX1 U2611 ( .A(n952), .Y(n3014) );
  AND2X1 U2612 ( .A(mem[503]), .B(n4533), .Y(n909) );
  INVX1 U2613 ( .A(n909), .Y(n3015) );
  AND2X1 U2614 ( .A(mem[497]), .B(n4533), .Y(n903) );
  INVX1 U2615 ( .A(n903), .Y(n3016) );
  AND2X1 U2616 ( .A(mem[466]), .B(n4534), .Y(n871) );
  INVX1 U2617 ( .A(n871), .Y(n3017) );
  AND2X1 U2618 ( .A(mem[465]), .B(n4534), .Y(n870) );
  INVX1 U2619 ( .A(n870), .Y(n3018) );
  AND2X1 U2620 ( .A(mem[434]), .B(n4535), .Y(n838) );
  INVX1 U2621 ( .A(n838), .Y(n3019) );
  AND2X1 U2622 ( .A(mem[429]), .B(n4535), .Y(n833) );
  INVX1 U2623 ( .A(n833), .Y(n3020) );
  AND2X1 U2624 ( .A(mem[402]), .B(n4536), .Y(n805) );
  INVX1 U2625 ( .A(n805), .Y(n3021) );
  AND2X1 U2626 ( .A(mem[397]), .B(n4536), .Y(n800) );
  INVX1 U2627 ( .A(n800), .Y(n3022) );
  AND2X1 U2628 ( .A(mem[385]), .B(n4537), .Y(n787) );
  INVX1 U2629 ( .A(n787), .Y(n3023) );
  AND2X1 U2630 ( .A(mem[373]), .B(n4537), .Y(n775) );
  INVX1 U2631 ( .A(n775), .Y(n3024) );
  AND2X1 U2632 ( .A(mem[353]), .B(n4538), .Y(n754) );
  INVX1 U2633 ( .A(n754), .Y(n3025) );
  AND2X1 U2634 ( .A(mem[341]), .B(n4538), .Y(n742) );
  INVX1 U2635 ( .A(n742), .Y(n3026) );
  AND2X1 U2636 ( .A(mem[317]), .B(n4539), .Y(n717) );
  INVX1 U2637 ( .A(n717), .Y(n3027) );
  AND2X1 U2638 ( .A(mem[304]), .B(n4539), .Y(n704) );
  INVX1 U2639 ( .A(n704), .Y(n3028) );
  AND2X1 U2640 ( .A(mem[285]), .B(n4540), .Y(n683) );
  INVX1 U2641 ( .A(n683), .Y(n3029) );
  AND2X1 U2642 ( .A(mem[273]), .B(n4540), .Y(n671) );
  INVX1 U2643 ( .A(n671), .Y(n3030) );
  AND2X1 U2644 ( .A(mem[239]), .B(n4541), .Y(n635) );
  INVX1 U2645 ( .A(n635), .Y(n3031) );
  AND2X1 U2646 ( .A(mem[233]), .B(n4541), .Y(n629) );
  INVX1 U2647 ( .A(n629), .Y(n3032) );
  AND2X1 U2648 ( .A(mem[202]), .B(n4542), .Y(n596) );
  INVX1 U2649 ( .A(n596), .Y(n3033) );
  AND2X1 U2650 ( .A(mem[201]), .B(n4542), .Y(n595) );
  INVX1 U2651 ( .A(n595), .Y(n3034) );
  AND2X1 U2652 ( .A(mem[170]), .B(n4543), .Y(n562) );
  INVX1 U2653 ( .A(n562), .Y(n3035) );
  AND2X1 U2654 ( .A(mem[165]), .B(n4543), .Y(n557) );
  INVX1 U2655 ( .A(n557), .Y(n3036) );
  AND2X1 U2656 ( .A(mem[138]), .B(n4544), .Y(n528) );
  INVX1 U2657 ( .A(n528), .Y(n3037) );
  AND2X1 U2658 ( .A(mem[133]), .B(n4544), .Y(n523) );
  INVX1 U2659 ( .A(n523), .Y(n3038) );
  AND2X1 U2660 ( .A(mem[121]), .B(n4545), .Y(n509) );
  INVX1 U2661 ( .A(n509), .Y(n3039) );
  AND2X1 U2662 ( .A(mem[109]), .B(n4545), .Y(n497) );
  INVX1 U2663 ( .A(n497), .Y(n3040) );
  AND2X1 U2664 ( .A(mem[89]), .B(n4546), .Y(n475) );
  INVX1 U2665 ( .A(n475), .Y(n3041) );
  AND2X1 U2666 ( .A(mem[77]), .B(n4546), .Y(n463) );
  INVX1 U2667 ( .A(n463), .Y(n3042) );
  AND2X1 U2668 ( .A(mem[53]), .B(n4547), .Y(n437) );
  INVX1 U2669 ( .A(n437), .Y(n3043) );
  AND2X1 U2670 ( .A(mem[40]), .B(n4547), .Y(n424) );
  INVX1 U2671 ( .A(n424), .Y(n3044) );
  AND2X1 U2672 ( .A(mem[21]), .B(n4548), .Y(n391) );
  INVX1 U2673 ( .A(n391), .Y(n3045) );
  AND2X1 U2674 ( .A(mem[9]), .B(n4548), .Y(n367) );
  INVX1 U2675 ( .A(n367), .Y(n3046) );
  BUFX2 U2676 ( .A(n626), .Y(n3047) );
  BUFX2 U2677 ( .A(n451), .Y(n3048) );
  AND2X1 U2678 ( .A(n4585), .B(n1490), .Y(n1493) );
  INVX1 U2679 ( .A(n1493), .Y(n3049) );
  AND2X1 U2680 ( .A(mem[1054]), .B(n4517), .Y(n1478) );
  INVX1 U2681 ( .A(n1478), .Y(n3050) );
  AND2X1 U2682 ( .A(mem[1042]), .B(n4517), .Y(n1466) );
  INVX1 U2683 ( .A(n1466), .Y(n3051) );
  AND2X1 U2684 ( .A(mem[1020]), .B(n4518), .Y(n1443) );
  INVX1 U2685 ( .A(n1443), .Y(n3052) );
  AND2X1 U2686 ( .A(mem[1008]), .B(n4518), .Y(n1431) );
  INVX1 U2687 ( .A(n1431), .Y(n3053) );
  AND2X1 U2688 ( .A(mem[986]), .B(n4519), .Y(n1408) );
  INVX1 U2689 ( .A(n1408), .Y(n3054) );
  AND2X1 U2690 ( .A(mem[974]), .B(n4519), .Y(n1396) );
  INVX1 U2691 ( .A(n1396), .Y(n3055) );
  AND2X1 U2692 ( .A(mem[952]), .B(n4520), .Y(n1373) );
  INVX1 U2693 ( .A(n1373), .Y(n3056) );
  AND2X1 U2694 ( .A(mem[940]), .B(n4520), .Y(n1361) );
  INVX1 U2695 ( .A(n1361), .Y(n3057) );
  AND2X1 U2696 ( .A(mem[895]), .B(n4521), .Y(n1315) );
  INVX1 U2697 ( .A(n1315), .Y(n3058) );
  AND2X1 U2698 ( .A(mem[894]), .B(n4521), .Y(n1314) );
  INVX1 U2699 ( .A(n1314), .Y(n3059) );
  AND2X1 U2700 ( .A(mem[866]), .B(n4522), .Y(n1285) );
  INVX1 U2701 ( .A(n1285), .Y(n3060) );
  AND2X1 U2702 ( .A(mem[860]), .B(n4522), .Y(n1279) );
  INVX1 U2703 ( .A(n1279), .Y(n3061) );
  AND2X1 U2704 ( .A(mem[831]), .B(n4523), .Y(n1249) );
  INVX1 U2705 ( .A(n1249), .Y(n3062) );
  AND2X1 U2706 ( .A(mem[826]), .B(n4523), .Y(n1244) );
  INVX1 U2707 ( .A(n1244), .Y(n3063) );
  AND2X1 U2708 ( .A(mem[797]), .B(n4524), .Y(n1213) );
  INVX1 U2709 ( .A(n1213), .Y(n3064) );
  AND2X1 U2710 ( .A(mem[792]), .B(n4524), .Y(n1208) );
  INVX1 U2711 ( .A(n1208), .Y(n3065) );
  AND2X1 U2712 ( .A(mem[782]), .B(n4525), .Y(n1197) );
  INVX1 U2713 ( .A(n1197), .Y(n3066) );
  AND2X1 U2714 ( .A(mem[770]), .B(n4525), .Y(n1185) );
  INVX1 U2715 ( .A(n1185), .Y(n3067) );
  AND2X1 U2716 ( .A(mem[748]), .B(n4526), .Y(n1162) );
  INVX1 U2717 ( .A(n1162), .Y(n3068) );
  AND2X1 U2718 ( .A(mem[736]), .B(n4526), .Y(n1150) );
  INVX1 U2719 ( .A(n1150), .Y(n3069) );
  AND2X1 U2720 ( .A(mem[714]), .B(n4527), .Y(n1127) );
  INVX1 U2721 ( .A(n1127), .Y(n3070) );
  AND2X1 U2722 ( .A(mem[702]), .B(n4527), .Y(n1115) );
  INVX1 U2723 ( .A(n1115), .Y(n3071) );
  AND2X1 U2724 ( .A(mem[680]), .B(n4528), .Y(n1092) );
  INVX1 U2725 ( .A(n1092), .Y(n3072) );
  AND2X1 U2726 ( .A(mem[667]), .B(n4528), .Y(n1079) );
  INVX1 U2727 ( .A(n1079), .Y(n3073) );
  AND2X1 U2728 ( .A(mem[658]), .B(n4529), .Y(n1069) );
  INVX1 U2729 ( .A(n1069), .Y(n3074) );
  AND2X1 U2730 ( .A(mem[646]), .B(n4529), .Y(n1057) );
  INVX1 U2731 ( .A(n1057), .Y(n3075) );
  AND2X1 U2732 ( .A(mem[624]), .B(n4530), .Y(n1034) );
  INVX1 U2733 ( .A(n1034), .Y(n3076) );
  AND2X1 U2734 ( .A(mem[612]), .B(n4530), .Y(n1022) );
  INVX1 U2735 ( .A(n1022), .Y(n3077) );
  AND2X1 U2736 ( .A(mem[590]), .B(n4531), .Y(n999) );
  INVX1 U2737 ( .A(n999), .Y(n3078) );
  AND2X1 U2738 ( .A(mem[578]), .B(n4531), .Y(n987) );
  INVX1 U2739 ( .A(n987), .Y(n3079) );
  AND2X1 U2740 ( .A(mem[556]), .B(n4532), .Y(n963) );
  INVX1 U2741 ( .A(n963), .Y(n3080) );
  AND2X1 U2742 ( .A(mem[544]), .B(n4532), .Y(n951) );
  INVX1 U2743 ( .A(n951), .Y(n3081) );
  AND2X1 U2744 ( .A(mem[499]), .B(n4533), .Y(n905) );
  INVX1 U2745 ( .A(n905), .Y(n3082) );
  AND2X1 U2746 ( .A(mem[498]), .B(n4533), .Y(n904) );
  INVX1 U2747 ( .A(n904), .Y(n3083) );
  AND2X1 U2748 ( .A(mem[470]), .B(n4534), .Y(n875) );
  INVX1 U2749 ( .A(n875), .Y(n3084) );
  AND2X1 U2750 ( .A(mem[464]), .B(n4534), .Y(n869) );
  INVX1 U2751 ( .A(n869), .Y(n3085) );
  AND2X1 U2752 ( .A(mem[435]), .B(n4535), .Y(n839) );
  INVX1 U2753 ( .A(n839), .Y(n3086) );
  AND2X1 U2754 ( .A(mem[430]), .B(n4535), .Y(n834) );
  INVX1 U2755 ( .A(n834), .Y(n3087) );
  AND2X1 U2756 ( .A(mem[401]), .B(n4536), .Y(n804) );
  INVX1 U2757 ( .A(n804), .Y(n3088) );
  AND2X1 U2758 ( .A(mem[396]), .B(n4536), .Y(n799) );
  INVX1 U2759 ( .A(n799), .Y(n3089) );
  AND2X1 U2760 ( .A(mem[386]), .B(n4537), .Y(n788) );
  INVX1 U2761 ( .A(n788), .Y(n3090) );
  AND2X1 U2762 ( .A(mem[374]), .B(n4537), .Y(n776) );
  INVX1 U2763 ( .A(n776), .Y(n3091) );
  AND2X1 U2764 ( .A(mem[352]), .B(n4538), .Y(n753) );
  INVX1 U2765 ( .A(n753), .Y(n3092) );
  AND2X1 U2766 ( .A(mem[340]), .B(n4538), .Y(n741) );
  INVX1 U2767 ( .A(n741), .Y(n3093) );
  AND2X1 U2768 ( .A(mem[318]), .B(n4539), .Y(n718) );
  INVX1 U2769 ( .A(n718), .Y(n3094) );
  AND2X1 U2770 ( .A(mem[306]), .B(n4539), .Y(n706) );
  INVX1 U2771 ( .A(n706), .Y(n3095) );
  AND2X1 U2772 ( .A(mem[284]), .B(n4540), .Y(n682) );
  INVX1 U2773 ( .A(n682), .Y(n3096) );
  AND2X1 U2774 ( .A(mem[271]), .B(n4540), .Y(n669) );
  INVX1 U2775 ( .A(n669), .Y(n3097) );
  AND2X1 U2776 ( .A(mem[235]), .B(n4541), .Y(n631) );
  INVX1 U2777 ( .A(n631), .Y(n3098) );
  AND2X1 U2778 ( .A(mem[234]), .B(n4541), .Y(n630) );
  INVX1 U2779 ( .A(n630), .Y(n3099) );
  AND2X1 U2780 ( .A(mem[206]), .B(n4542), .Y(n600) );
  INVX1 U2781 ( .A(n600), .Y(n3100) );
  AND2X1 U2782 ( .A(mem[200]), .B(n4542), .Y(n594) );
  INVX1 U2783 ( .A(n594), .Y(n3101) );
  AND2X1 U2784 ( .A(mem[171]), .B(n4543), .Y(n563) );
  INVX1 U2785 ( .A(n563), .Y(n3102) );
  AND2X1 U2786 ( .A(mem[166]), .B(n4543), .Y(n558) );
  INVX1 U2787 ( .A(n558), .Y(n3103) );
  AND2X1 U2788 ( .A(mem[137]), .B(n4544), .Y(n527) );
  INVX1 U2789 ( .A(n527), .Y(n3104) );
  AND2X1 U2790 ( .A(mem[132]), .B(n4544), .Y(n522) );
  INVX1 U2791 ( .A(n522), .Y(n3105) );
  AND2X1 U2792 ( .A(mem[122]), .B(n4545), .Y(n510) );
  INVX1 U2793 ( .A(n510), .Y(n3106) );
  AND2X1 U2794 ( .A(mem[110]), .B(n4545), .Y(n498) );
  INVX1 U2795 ( .A(n498), .Y(n3107) );
  AND2X1 U2796 ( .A(mem[88]), .B(n4546), .Y(n474) );
  INVX1 U2797 ( .A(n474), .Y(n3108) );
  AND2X1 U2798 ( .A(mem[76]), .B(n4546), .Y(n462) );
  INVX1 U2799 ( .A(n462), .Y(n3109) );
  AND2X1 U2800 ( .A(mem[54]), .B(n4547), .Y(n438) );
  INVX1 U2801 ( .A(n438), .Y(n3110) );
  AND2X1 U2802 ( .A(mem[42]), .B(n4547), .Y(n426) );
  INVX1 U2803 ( .A(n426), .Y(n3111) );
  AND2X1 U2804 ( .A(mem[20]), .B(n4548), .Y(n389) );
  INVX1 U2805 ( .A(n389), .Y(n3112) );
  AND2X1 U2806 ( .A(mem[7]), .B(n4548), .Y(n363) );
  INVX1 U2807 ( .A(n363), .Y(n3113) );
  INVX1 U2808 ( .A(n1481), .Y(n3114) );
  BUFX2 U2809 ( .A(n4625), .Y(full_bar) );
  OR2X1 U2810 ( .A(fillcount[1]), .B(fillcount[0]), .Y(n1530) );
  INVX1 U2811 ( .A(n1530), .Y(n3116) );
  BUFX2 U2812 ( .A(n661), .Y(n3117) );
  BUFX2 U2813 ( .A(n416), .Y(n3118) );
  AND2X1 U2814 ( .A(n90), .B(n1490), .Y(n1492) );
  INVX1 U2815 ( .A(n1492), .Y(n3119) );
  AND2X1 U2816 ( .A(n20), .B(n1484), .Y(n1486) );
  INVX1 U2817 ( .A(n1486), .Y(n3120) );
  AND2X1 U2818 ( .A(mem[1047]), .B(n4517), .Y(n1471) );
  INVX1 U2819 ( .A(n1471), .Y(n3121) );
  AND2X1 U2820 ( .A(mem[1035]), .B(n4517), .Y(n1459) );
  INVX1 U2821 ( .A(n1459), .Y(n3122) );
  AND2X1 U2822 ( .A(mem[1015]), .B(n4518), .Y(n1438) );
  INVX1 U2823 ( .A(n1438), .Y(n3123) );
  AND2X1 U2824 ( .A(mem[1003]), .B(n4518), .Y(n1426) );
  INVX1 U2825 ( .A(n1426), .Y(n3124) );
  AND2X1 U2826 ( .A(mem[983]), .B(n4519), .Y(n1405) );
  INVX1 U2827 ( .A(n1405), .Y(n3125) );
  AND2X1 U2828 ( .A(mem[971]), .B(n4519), .Y(n1393) );
  INVX1 U2829 ( .A(n1393), .Y(n3126) );
  AND2X1 U2830 ( .A(mem[951]), .B(n4520), .Y(n1372) );
  INVX1 U2831 ( .A(n1372), .Y(n3127) );
  AND2X1 U2832 ( .A(mem[939]), .B(n4520), .Y(n1360) );
  INVX1 U2833 ( .A(n1360), .Y(n3128) );
  AND2X1 U2834 ( .A(mem[911]), .B(n4521), .Y(n1331) );
  INVX1 U2835 ( .A(n1331), .Y(n3129) );
  AND2X1 U2836 ( .A(mem[898]), .B(n4521), .Y(n1318) );
  INVX1 U2837 ( .A(n1318), .Y(n3130) );
  AND2X1 U2838 ( .A(mem[879]), .B(n4522), .Y(n1298) );
  INVX1 U2839 ( .A(n1298), .Y(n3131) );
  AND2X1 U2840 ( .A(mem[867]), .B(n4522), .Y(n1286) );
  INVX1 U2841 ( .A(n1286), .Y(n3132) );
  AND2X1 U2842 ( .A(mem[847]), .B(n4523), .Y(n1265) );
  INVX1 U2843 ( .A(n1265), .Y(n3133) );
  AND2X1 U2844 ( .A(mem[835]), .B(n4523), .Y(n1253) );
  INVX1 U2845 ( .A(n1253), .Y(n3134) );
  AND2X1 U2846 ( .A(mem[815]), .B(n4524), .Y(n1231) );
  INVX1 U2847 ( .A(n1231), .Y(n3135) );
  AND2X1 U2848 ( .A(mem[803]), .B(n4524), .Y(n1219) );
  INVX1 U2849 ( .A(n1219), .Y(n3136) );
  AND2X1 U2850 ( .A(mem[764]), .B(n4525), .Y(n1179) );
  INVX1 U2851 ( .A(n1179), .Y(n3137) );
  AND2X1 U2852 ( .A(mem[759]), .B(n4525), .Y(n1174) );
  INVX1 U2853 ( .A(n1174), .Y(n3138) );
  AND2X1 U2854 ( .A(mem[732]), .B(n4526), .Y(n1146) );
  INVX1 U2855 ( .A(n1146), .Y(n3139) );
  AND2X1 U2856 ( .A(mem[727]), .B(n4526), .Y(n1141) );
  INVX1 U2857 ( .A(n1141), .Y(n3140) );
  AND2X1 U2858 ( .A(mem[701]), .B(n4527), .Y(n1114) );
  INVX1 U2859 ( .A(n1114), .Y(n3141) );
  AND2X1 U2860 ( .A(mem[695]), .B(n4527), .Y(n1108) );
  INVX1 U2861 ( .A(n1108), .Y(n3142) );
  AND2X1 U2862 ( .A(mem[664]), .B(n4528), .Y(n1076) );
  INVX1 U2863 ( .A(n1076), .Y(n3143) );
  AND2X1 U2864 ( .A(mem[663]), .B(n4528), .Y(n1075) );
  INVX1 U2865 ( .A(n1075), .Y(n3144) );
  AND2X1 U2866 ( .A(mem[651]), .B(n4529), .Y(n1062) );
  INVX1 U2867 ( .A(n1062), .Y(n3145) );
  AND2X1 U2868 ( .A(mem[639]), .B(n4529), .Y(n1050) );
  INVX1 U2869 ( .A(n1050), .Y(n3146) );
  AND2X1 U2870 ( .A(mem[619]), .B(n4530), .Y(n1029) );
  INVX1 U2871 ( .A(n1029), .Y(n3147) );
  AND2X1 U2872 ( .A(mem[607]), .B(n4530), .Y(n1017) );
  INVX1 U2873 ( .A(n1017), .Y(n3148) );
  AND2X1 U2874 ( .A(mem[587]), .B(n4531), .Y(n996) );
  INVX1 U2875 ( .A(n996), .Y(n3149) );
  AND2X1 U2876 ( .A(mem[575]), .B(n4531), .Y(n984) );
  INVX1 U2877 ( .A(n984), .Y(n3150) );
  AND2X1 U2878 ( .A(mem[555]), .B(n4532), .Y(n962) );
  INVX1 U2879 ( .A(n962), .Y(n3151) );
  AND2X1 U2880 ( .A(mem[543]), .B(n4532), .Y(n950) );
  INVX1 U2881 ( .A(n950), .Y(n3152) );
  AND2X1 U2882 ( .A(mem[515]), .B(n4533), .Y(n921) );
  INVX1 U2883 ( .A(n921), .Y(n3153) );
  AND2X1 U2884 ( .A(mem[502]), .B(n4533), .Y(n908) );
  INVX1 U2885 ( .A(n908), .Y(n3154) );
  AND2X1 U2886 ( .A(mem[483]), .B(n4534), .Y(n888) );
  INVX1 U2887 ( .A(n888), .Y(n3155) );
  AND2X1 U2888 ( .A(mem[471]), .B(n4534), .Y(n876) );
  INVX1 U2889 ( .A(n876), .Y(n3156) );
  AND2X1 U2890 ( .A(mem[451]), .B(n4535), .Y(n855) );
  INVX1 U2891 ( .A(n855), .Y(n3157) );
  AND2X1 U2892 ( .A(mem[439]), .B(n4535), .Y(n843) );
  INVX1 U2893 ( .A(n843), .Y(n3158) );
  AND2X1 U2894 ( .A(mem[419]), .B(n4536), .Y(n822) );
  INVX1 U2895 ( .A(n822), .Y(n3159) );
  AND2X1 U2896 ( .A(mem[407]), .B(n4536), .Y(n810) );
  INVX1 U2897 ( .A(n810), .Y(n3160) );
  AND2X1 U2898 ( .A(mem[368]), .B(n4537), .Y(n770) );
  INVX1 U2899 ( .A(n770), .Y(n3161) );
  AND2X1 U2900 ( .A(mem[363]), .B(n4537), .Y(n765) );
  INVX1 U2901 ( .A(n765), .Y(n3162) );
  AND2X1 U2902 ( .A(mem[336]), .B(n4538), .Y(n737) );
  INVX1 U2903 ( .A(n737), .Y(n3163) );
  AND2X1 U2904 ( .A(mem[331]), .B(n4538), .Y(n732) );
  INVX1 U2905 ( .A(n732), .Y(n3164) );
  AND2X1 U2906 ( .A(mem[305]), .B(n4539), .Y(n705) );
  INVX1 U2907 ( .A(n705), .Y(n3165) );
  AND2X1 U2908 ( .A(mem[299]), .B(n4539), .Y(n699) );
  INVX1 U2909 ( .A(n699), .Y(n3166) );
  AND2X1 U2910 ( .A(mem[268]), .B(n4540), .Y(n666) );
  INVX1 U2911 ( .A(n666), .Y(n3167) );
  AND2X1 U2912 ( .A(mem[267]), .B(n4540), .Y(n665) );
  INVX1 U2913 ( .A(n665), .Y(n3168) );
  AND2X1 U2914 ( .A(mem[251]), .B(n4541), .Y(n647) );
  INVX1 U2915 ( .A(n647), .Y(n3169) );
  AND2X1 U2916 ( .A(mem[238]), .B(n4541), .Y(n634) );
  INVX1 U2917 ( .A(n634), .Y(n3170) );
  AND2X1 U2918 ( .A(mem[219]), .B(n4542), .Y(n613) );
  INVX1 U2919 ( .A(n613), .Y(n3171) );
  AND2X1 U2920 ( .A(mem[207]), .B(n4542), .Y(n601) );
  INVX1 U2921 ( .A(n601), .Y(n3172) );
  AND2X1 U2922 ( .A(mem[187]), .B(n4543), .Y(n579) );
  INVX1 U2923 ( .A(n579), .Y(n3173) );
  AND2X1 U2924 ( .A(mem[175]), .B(n4543), .Y(n567) );
  INVX1 U2925 ( .A(n567), .Y(n3174) );
  AND2X1 U2926 ( .A(mem[155]), .B(n4544), .Y(n545) );
  INVX1 U2927 ( .A(n545), .Y(n3175) );
  AND2X1 U2928 ( .A(mem[143]), .B(n4544), .Y(n533) );
  INVX1 U2929 ( .A(n533), .Y(n3176) );
  AND2X1 U2930 ( .A(mem[104]), .B(n4545), .Y(n492) );
  INVX1 U2931 ( .A(n492), .Y(n3177) );
  AND2X1 U2932 ( .A(mem[99]), .B(n4545), .Y(n487) );
  INVX1 U2933 ( .A(n487), .Y(n3178) );
  AND2X1 U2934 ( .A(mem[72]), .B(n4546), .Y(n458) );
  INVX1 U2935 ( .A(n458), .Y(n3179) );
  AND2X1 U2936 ( .A(mem[67]), .B(n4546), .Y(n453) );
  INVX1 U2937 ( .A(n453), .Y(n3180) );
  AND2X1 U2938 ( .A(mem[41]), .B(n4547), .Y(n425) );
  INVX1 U2939 ( .A(n425), .Y(n3181) );
  AND2X1 U2940 ( .A(mem[35]), .B(n4547), .Y(n419) );
  INVX1 U2941 ( .A(n419), .Y(n3182) );
  AND2X1 U2942 ( .A(mem[4]), .B(n4548), .Y(n357) );
  INVX1 U2943 ( .A(n357), .Y(n3183) );
  AND2X1 U2944 ( .A(mem[3]), .B(n4548), .Y(n355) );
  INVX1 U2945 ( .A(n355), .Y(n3184) );
  BUFX2 U2946 ( .A(n415), .Y(n3185) );
  AND2X1 U2947 ( .A(n91), .B(n1490), .Y(n1491) );
  INVX1 U2948 ( .A(n1491), .Y(n3186) );
  AND2X1 U2949 ( .A(n21), .B(n1484), .Y(n1485) );
  INVX1 U2950 ( .A(n1485), .Y(n3187) );
  AND2X1 U2951 ( .A(reset), .B(n3318), .Y(n1484) );
  AND2X1 U2952 ( .A(mem[1048]), .B(n4517), .Y(n1472) );
  INVX1 U2953 ( .A(n1472), .Y(n3188) );
  AND2X1 U2954 ( .A(mem[1036]), .B(n4517), .Y(n1460) );
  INVX1 U2955 ( .A(n1460), .Y(n3189) );
  AND2X1 U2956 ( .A(mem[1014]), .B(n4518), .Y(n1437) );
  INVX1 U2957 ( .A(n1437), .Y(n3190) );
  AND2X1 U2958 ( .A(mem[1002]), .B(n4518), .Y(n1425) );
  INVX1 U2959 ( .A(n1425), .Y(n3191) );
  AND2X1 U2960 ( .A(mem[984]), .B(n4519), .Y(n1406) );
  INVX1 U2961 ( .A(n1406), .Y(n3192) );
  AND2X1 U2962 ( .A(mem[972]), .B(n4519), .Y(n1394) );
  INVX1 U2963 ( .A(n1394), .Y(n3193) );
  AND2X1 U2964 ( .A(mem[950]), .B(n4520), .Y(n1371) );
  INVX1 U2965 ( .A(n1371), .Y(n3194) );
  AND2X1 U2966 ( .A(mem[938]), .B(n4520), .Y(n1359) );
  INVX1 U2967 ( .A(n1359), .Y(n3195) );
  AND2X1 U2968 ( .A(mem[912]), .B(n4521), .Y(n1332) );
  INVX1 U2969 ( .A(n1332), .Y(n3196) );
  AND2X1 U2970 ( .A(mem[900]), .B(n4521), .Y(n1320) );
  INVX1 U2971 ( .A(n1320), .Y(n3197) );
  AND2X1 U2972 ( .A(mem[878]), .B(n4522), .Y(n1297) );
  INVX1 U2973 ( .A(n1297), .Y(n3198) );
  AND2X1 U2974 ( .A(mem[865]), .B(n4522), .Y(n1284) );
  INVX1 U2975 ( .A(n1284), .Y(n3199) );
  AND2X1 U2976 ( .A(mem[848]), .B(n4523), .Y(n1266) );
  INVX1 U2977 ( .A(n1266), .Y(n3200) );
  AND2X1 U2978 ( .A(mem[836]), .B(n4523), .Y(n1254) );
  INVX1 U2979 ( .A(n1254), .Y(n3201) );
  AND2X1 U2980 ( .A(mem[814]), .B(n4524), .Y(n1230) );
  INVX1 U2981 ( .A(n1230), .Y(n3202) );
  AND2X1 U2982 ( .A(mem[802]), .B(n4524), .Y(n1218) );
  INVX1 U2983 ( .A(n1218), .Y(n3203) );
  AND2X1 U2984 ( .A(mem[765]), .B(n4525), .Y(n1180) );
  INVX1 U2985 ( .A(n1180), .Y(n3204) );
  AND2X1 U2986 ( .A(mem[760]), .B(n4525), .Y(n1175) );
  INVX1 U2987 ( .A(n1175), .Y(n3205) );
  AND2X1 U2988 ( .A(mem[731]), .B(n4526), .Y(n1145) );
  INVX1 U2989 ( .A(n1145), .Y(n3206) );
  AND2X1 U2990 ( .A(mem[726]), .B(n4526), .Y(n1140) );
  INVX1 U2991 ( .A(n1140), .Y(n3207) );
  AND2X1 U2992 ( .A(mem[697]), .B(n4527), .Y(n1110) );
  INVX1 U2993 ( .A(n1110), .Y(n3208) );
  AND2X1 U2994 ( .A(mem[696]), .B(n4527), .Y(n1109) );
  INVX1 U2995 ( .A(n1109), .Y(n3209) );
  AND2X1 U2996 ( .A(mem[668]), .B(n4528), .Y(n1080) );
  INVX1 U2997 ( .A(n1080), .Y(n3210) );
  AND2X1 U2998 ( .A(mem[662]), .B(n4528), .Y(n1074) );
  INVX1 U2999 ( .A(n1074), .Y(n3211) );
  AND2X1 U3000 ( .A(mem[652]), .B(n4529), .Y(n1063) );
  INVX1 U3001 ( .A(n1063), .Y(n3212) );
  AND2X1 U3002 ( .A(mem[640]), .B(n4529), .Y(n1051) );
  INVX1 U3003 ( .A(n1051), .Y(n3213) );
  AND2X1 U3004 ( .A(mem[618]), .B(n4530), .Y(n1028) );
  INVX1 U3005 ( .A(n1028), .Y(n3214) );
  AND2X1 U3006 ( .A(mem[606]), .B(n4530), .Y(n1016) );
  INVX1 U3007 ( .A(n1016), .Y(n3215) );
  AND2X1 U3008 ( .A(mem[588]), .B(n4531), .Y(n997) );
  INVX1 U3009 ( .A(n997), .Y(n3216) );
  AND2X1 U3010 ( .A(mem[576]), .B(n4531), .Y(n985) );
  INVX1 U3011 ( .A(n985), .Y(n3217) );
  AND2X1 U3012 ( .A(mem[554]), .B(n4532), .Y(n961) );
  INVX1 U3013 ( .A(n961), .Y(n3218) );
  AND2X1 U3014 ( .A(mem[542]), .B(n4532), .Y(n949) );
  INVX1 U3015 ( .A(n949), .Y(n3219) );
  AND2X1 U3016 ( .A(mem[516]), .B(n4533), .Y(n922) );
  INVX1 U3017 ( .A(n922), .Y(n3220) );
  AND2X1 U3018 ( .A(mem[504]), .B(n4533), .Y(n910) );
  INVX1 U3019 ( .A(n910), .Y(n3221) );
  AND2X1 U3020 ( .A(mem[482]), .B(n4534), .Y(n887) );
  INVX1 U3021 ( .A(n887), .Y(n3222) );
  AND2X1 U3022 ( .A(mem[469]), .B(n4534), .Y(n874) );
  INVX1 U3023 ( .A(n874), .Y(n3223) );
  AND2X1 U3024 ( .A(mem[452]), .B(n4535), .Y(n856) );
  INVX1 U3025 ( .A(n856), .Y(n3224) );
  AND2X1 U3026 ( .A(mem[440]), .B(n4535), .Y(n844) );
  INVX1 U3027 ( .A(n844), .Y(n3225) );
  AND2X1 U3028 ( .A(mem[418]), .B(n4536), .Y(n821) );
  INVX1 U3029 ( .A(n821), .Y(n3226) );
  AND2X1 U3030 ( .A(mem[406]), .B(n4536), .Y(n809) );
  INVX1 U3031 ( .A(n809), .Y(n3227) );
  AND2X1 U3032 ( .A(mem[369]), .B(n4537), .Y(n771) );
  INVX1 U3033 ( .A(n771), .Y(n3228) );
  AND2X1 U3034 ( .A(mem[364]), .B(n4537), .Y(n766) );
  INVX1 U3035 ( .A(n766), .Y(n3229) );
  AND2X1 U3036 ( .A(mem[335]), .B(n4538), .Y(n736) );
  INVX1 U3037 ( .A(n736), .Y(n3230) );
  AND2X1 U3038 ( .A(mem[330]), .B(n4538), .Y(n731) );
  INVX1 U3039 ( .A(n731), .Y(n3231) );
  AND2X1 U3040 ( .A(mem[301]), .B(n4539), .Y(n701) );
  INVX1 U3041 ( .A(n701), .Y(n3232) );
  AND2X1 U3042 ( .A(mem[300]), .B(n4539), .Y(n700) );
  INVX1 U3043 ( .A(n700), .Y(n3233) );
  AND2X1 U3044 ( .A(mem[272]), .B(n4540), .Y(n670) );
  INVX1 U3045 ( .A(n670), .Y(n3234) );
  AND2X1 U3046 ( .A(mem[266]), .B(n4540), .Y(n664) );
  INVX1 U3047 ( .A(n664), .Y(n3235) );
  AND2X1 U3048 ( .A(mem[252]), .B(n4541), .Y(n648) );
  INVX1 U3049 ( .A(n648), .Y(n3236) );
  AND2X1 U3050 ( .A(mem[240]), .B(n4541), .Y(n636) );
  INVX1 U3051 ( .A(n636), .Y(n3237) );
  AND2X1 U3052 ( .A(mem[218]), .B(n4542), .Y(n612) );
  INVX1 U3053 ( .A(n612), .Y(n3238) );
  AND2X1 U3054 ( .A(mem[205]), .B(n4542), .Y(n599) );
  INVX1 U3055 ( .A(n599), .Y(n3239) );
  AND2X1 U3056 ( .A(mem[188]), .B(n4543), .Y(n580) );
  INVX1 U3057 ( .A(n580), .Y(n3240) );
  AND2X1 U3058 ( .A(mem[176]), .B(n4543), .Y(n568) );
  INVX1 U3059 ( .A(n568), .Y(n3241) );
  AND2X1 U3060 ( .A(mem[154]), .B(n4544), .Y(n544) );
  INVX1 U3061 ( .A(n544), .Y(n3242) );
  AND2X1 U3062 ( .A(mem[142]), .B(n4544), .Y(n532) );
  INVX1 U3063 ( .A(n532), .Y(n3243) );
  AND2X1 U3064 ( .A(mem[105]), .B(n4545), .Y(n493) );
  INVX1 U3065 ( .A(n493), .Y(n3244) );
  AND2X1 U3066 ( .A(mem[100]), .B(n4545), .Y(n488) );
  INVX1 U3067 ( .A(n488), .Y(n3245) );
  AND2X1 U3068 ( .A(mem[71]), .B(n4546), .Y(n457) );
  INVX1 U3069 ( .A(n457), .Y(n3246) );
  AND2X1 U3070 ( .A(mem[66]), .B(n4546), .Y(n452) );
  INVX1 U3071 ( .A(n452), .Y(n3247) );
  AND2X1 U3072 ( .A(mem[37]), .B(n4547), .Y(n421) );
  INVX1 U3073 ( .A(n421), .Y(n3248) );
  AND2X1 U3074 ( .A(mem[36]), .B(n4547), .Y(n420) );
  INVX1 U3075 ( .A(n420), .Y(n3249) );
  AND2X1 U3076 ( .A(mem[8]), .B(n4548), .Y(n365) );
  INVX1 U3077 ( .A(n365), .Y(n3250) );
  AND2X1 U3078 ( .A(mem[2]), .B(n4548), .Y(n353) );
  INVX1 U3079 ( .A(n353), .Y(n3251) );
  BUFX2 U3080 ( .A(n1242), .Y(n3252) );
  AND2X1 U3081 ( .A(n92), .B(n1490), .Y(n1489) );
  INVX1 U3082 ( .A(n1489), .Y(n3253) );
  AND2X1 U3083 ( .A(mem[1049]), .B(n4517), .Y(n1473) );
  INVX1 U3084 ( .A(n1473), .Y(n3254) );
  AND2X1 U3085 ( .A(mem[1037]), .B(n4517), .Y(n1461) );
  INVX1 U3086 ( .A(n1461), .Y(n3255) );
  AND2X1 U3087 ( .A(mem[1017]), .B(n4518), .Y(n1440) );
  INVX1 U3088 ( .A(n1440), .Y(n3256) );
  AND2X1 U3089 ( .A(mem[1005]), .B(n4518), .Y(n1428) );
  INVX1 U3090 ( .A(n1428), .Y(n3257) );
  AND2X1 U3091 ( .A(mem[981]), .B(n4519), .Y(n1403) );
  INVX1 U3092 ( .A(n1403), .Y(n3258) );
  AND2X1 U3093 ( .A(mem[969]), .B(n4519), .Y(n1391) );
  INVX1 U3094 ( .A(n1391), .Y(n3259) );
  AND2X1 U3095 ( .A(mem[949]), .B(n4520), .Y(n1370) );
  INVX1 U3096 ( .A(n1370), .Y(n3260) );
  AND2X1 U3097 ( .A(mem[937]), .B(n4520), .Y(n1358) );
  INVX1 U3098 ( .A(n1358), .Y(n3261) );
  AND2X1 U3099 ( .A(mem[913]), .B(n4521), .Y(n1333) );
  INVX1 U3100 ( .A(n1333), .Y(n3262) );
  AND2X1 U3101 ( .A(mem[901]), .B(n4521), .Y(n1321) );
  INVX1 U3102 ( .A(n1321), .Y(n3263) );
  AND2X1 U3103 ( .A(mem[881]), .B(n4522), .Y(n1300) );
  INVX1 U3104 ( .A(n1300), .Y(n3264) );
  AND2X1 U3105 ( .A(mem[869]), .B(n4522), .Y(n1288) );
  INVX1 U3106 ( .A(n1288), .Y(n3265) );
  AND2X1 U3107 ( .A(mem[845]), .B(n4523), .Y(n1263) );
  INVX1 U3108 ( .A(n1263), .Y(n3266) );
  AND2X1 U3109 ( .A(mem[832]), .B(n4523), .Y(n1250) );
  INVX1 U3110 ( .A(n1250), .Y(n3267) );
  AND2X1 U3111 ( .A(mem[813]), .B(n4524), .Y(n1229) );
  INVX1 U3112 ( .A(n1229), .Y(n3268) );
  AND2X1 U3113 ( .A(mem[801]), .B(n4524), .Y(n1217) );
  INVX1 U3114 ( .A(n1217), .Y(n3269) );
  AND2X1 U3115 ( .A(mem[767]), .B(n4525), .Y(n1182) );
  INVX1 U3116 ( .A(n1182), .Y(n3270) );
  AND2X1 U3117 ( .A(mem[761]), .B(n4525), .Y(n1176) );
  INVX1 U3118 ( .A(n1176), .Y(n3271) );
  AND2X1 U3119 ( .A(mem[730]), .B(n4526), .Y(n1144) );
  INVX1 U3120 ( .A(n1144), .Y(n3272) );
  AND2X1 U3121 ( .A(mem[729]), .B(n4526), .Y(n1143) );
  INVX1 U3122 ( .A(n1143), .Y(n3273) );
  AND2X1 U3123 ( .A(mem[698]), .B(n4527), .Y(n1111) );
  INVX1 U3124 ( .A(n1111), .Y(n3274) );
  AND2X1 U3125 ( .A(mem[693]), .B(n4527), .Y(n1106) );
  INVX1 U3126 ( .A(n1106), .Y(n3275) );
  AND2X1 U3127 ( .A(mem[666]), .B(n4528), .Y(n1078) );
  INVX1 U3128 ( .A(n1078), .Y(n3276) );
  AND2X1 U3129 ( .A(mem[661]), .B(n4528), .Y(n1073) );
  INVX1 U3130 ( .A(n1073), .Y(n3277) );
  AND2X1 U3131 ( .A(mem[653]), .B(n4529), .Y(n1064) );
  INVX1 U3132 ( .A(n1064), .Y(n3278) );
  AND2X1 U3133 ( .A(mem[641]), .B(n4529), .Y(n1052) );
  INVX1 U3134 ( .A(n1052), .Y(n3279) );
  AND2X1 U3135 ( .A(mem[621]), .B(n4530), .Y(n1031) );
  INVX1 U3136 ( .A(n1031), .Y(n3280) );
  AND2X1 U3137 ( .A(mem[609]), .B(n4530), .Y(n1019) );
  INVX1 U3138 ( .A(n1019), .Y(n3281) );
  AND2X1 U3139 ( .A(mem[585]), .B(n4531), .Y(n994) );
  INVX1 U3140 ( .A(n994), .Y(n3282) );
  AND2X1 U3141 ( .A(mem[573]), .B(n4531), .Y(n982) );
  INVX1 U3142 ( .A(n982), .Y(n3283) );
  AND2X1 U3143 ( .A(mem[553]), .B(n4532), .Y(n960) );
  INVX1 U3144 ( .A(n960), .Y(n3284) );
  AND2X1 U3145 ( .A(mem[541]), .B(n4532), .Y(n948) );
  INVX1 U3146 ( .A(n948), .Y(n3285) );
  AND2X1 U3147 ( .A(mem[517]), .B(n4533), .Y(n923) );
  INVX1 U3148 ( .A(n923), .Y(n3286) );
  AND2X1 U3149 ( .A(mem[505]), .B(n4533), .Y(n911) );
  INVX1 U3150 ( .A(n911), .Y(n3287) );
  AND2X1 U3151 ( .A(mem[485]), .B(n4534), .Y(n890) );
  INVX1 U3152 ( .A(n890), .Y(n3288) );
  AND2X1 U3153 ( .A(mem[473]), .B(n4534), .Y(n878) );
  INVX1 U3154 ( .A(n878), .Y(n3289) );
  AND2X1 U3155 ( .A(mem[449]), .B(n4535), .Y(n853) );
  INVX1 U3156 ( .A(n853), .Y(n3290) );
  AND2X1 U3157 ( .A(mem[436]), .B(n4535), .Y(n840) );
  INVX1 U3158 ( .A(n840), .Y(n3291) );
  AND2X1 U3159 ( .A(mem[417]), .B(n4536), .Y(n820) );
  INVX1 U3160 ( .A(n820), .Y(n3292) );
  AND2X1 U3161 ( .A(mem[405]), .B(n4536), .Y(n808) );
  INVX1 U3162 ( .A(n808), .Y(n3293) );
  AND2X1 U3163 ( .A(mem[371]), .B(n4537), .Y(n773) );
  INVX1 U3164 ( .A(n773), .Y(n3294) );
  AND2X1 U3165 ( .A(mem[365]), .B(n4537), .Y(n767) );
  INVX1 U3166 ( .A(n767), .Y(n3295) );
  AND2X1 U3167 ( .A(mem[334]), .B(n4538), .Y(n735) );
  INVX1 U3168 ( .A(n735), .Y(n3296) );
  AND2X1 U3169 ( .A(mem[333]), .B(n4538), .Y(n734) );
  INVX1 U3170 ( .A(n734), .Y(n3297) );
  AND2X1 U3171 ( .A(mem[302]), .B(n4539), .Y(n702) );
  INVX1 U3172 ( .A(n702), .Y(n3298) );
  AND2X1 U3173 ( .A(mem[297]), .B(n4539), .Y(n697) );
  INVX1 U3174 ( .A(n697), .Y(n3299) );
  AND2X1 U3175 ( .A(mem[270]), .B(n4540), .Y(n668) );
  INVX1 U3176 ( .A(n668), .Y(n3300) );
  AND2X1 U3177 ( .A(mem[265]), .B(n4540), .Y(n663) );
  INVX1 U3178 ( .A(n663), .Y(n3301) );
  AND2X1 U3179 ( .A(mem[253]), .B(n4541), .Y(n649) );
  INVX1 U3180 ( .A(n649), .Y(n3302) );
  AND2X1 U3181 ( .A(mem[241]), .B(n4541), .Y(n637) );
  INVX1 U3182 ( .A(n637), .Y(n3303) );
  AND2X1 U3183 ( .A(mem[221]), .B(n4542), .Y(n615) );
  INVX1 U3184 ( .A(n615), .Y(n3304) );
  AND2X1 U3185 ( .A(mem[209]), .B(n4542), .Y(n603) );
  INVX1 U3186 ( .A(n603), .Y(n3305) );
  AND2X1 U3187 ( .A(mem[185]), .B(n4543), .Y(n577) );
  INVX1 U3188 ( .A(n577), .Y(n3306) );
  AND2X1 U3189 ( .A(mem[172]), .B(n4543), .Y(n564) );
  INVX1 U3190 ( .A(n564), .Y(n3307) );
  AND2X1 U3191 ( .A(mem[153]), .B(n4544), .Y(n543) );
  INVX1 U3192 ( .A(n543), .Y(n3308) );
  AND2X1 U3193 ( .A(mem[141]), .B(n4544), .Y(n531) );
  INVX1 U3194 ( .A(n531), .Y(n3309) );
  AND2X1 U3195 ( .A(mem[107]), .B(n4545), .Y(n495) );
  INVX1 U3196 ( .A(n495), .Y(n3310) );
  AND2X1 U3197 ( .A(mem[101]), .B(n4545), .Y(n489) );
  INVX1 U3198 ( .A(n489), .Y(n3311) );
  AND2X1 U3199 ( .A(mem[70]), .B(n4546), .Y(n456) );
  INVX1 U3200 ( .A(n456), .Y(n3312) );
  AND2X1 U3201 ( .A(mem[69]), .B(n4546), .Y(n455) );
  INVX1 U3202 ( .A(n455), .Y(n3313) );
  AND2X1 U3203 ( .A(mem[38]), .B(n4547), .Y(n422) );
  INVX1 U3204 ( .A(n422), .Y(n3314) );
  AND2X1 U3205 ( .A(mem[33]), .B(n4547), .Y(n417) );
  INVX1 U3206 ( .A(n417), .Y(n3315) );
  AND2X1 U3207 ( .A(mem[6]), .B(n4548), .Y(n361) );
  INVX1 U3208 ( .A(n361), .Y(n3316) );
  AND2X1 U3209 ( .A(mem[1]), .B(n4548), .Y(n351) );
  INVX1 U3210 ( .A(n351), .Y(n3317) );
  INVX1 U3211 ( .A(n1482), .Y(n3318) );
  BUFX2 U3212 ( .A(n969), .Y(n3319) );
  AND2X1 U3213 ( .A(mem[1050]), .B(n4517), .Y(n1474) );
  INVX1 U3214 ( .A(n1474), .Y(n3320) );
  AND2X1 U3215 ( .A(mem[1038]), .B(n4517), .Y(n1462) );
  INVX1 U3216 ( .A(n1462), .Y(n3321) );
  AND2X1 U3217 ( .A(mem[1016]), .B(n4518), .Y(n1439) );
  INVX1 U3218 ( .A(n1439), .Y(n3322) );
  AND2X1 U3219 ( .A(mem[1004]), .B(n4518), .Y(n1427) );
  INVX1 U3220 ( .A(n1427), .Y(n3323) );
  AND2X1 U3221 ( .A(mem[982]), .B(n4519), .Y(n1404) );
  INVX1 U3222 ( .A(n1404), .Y(n3324) );
  AND2X1 U3223 ( .A(mem[970]), .B(n4519), .Y(n1392) );
  INVX1 U3224 ( .A(n1392), .Y(n3325) );
  AND2X1 U3225 ( .A(mem[948]), .B(n4520), .Y(n1369) );
  INVX1 U3226 ( .A(n1369), .Y(n3326) );
  AND2X1 U3227 ( .A(mem[936]), .B(n4520), .Y(n1357) );
  INVX1 U3228 ( .A(n1357), .Y(n3327) );
  AND2X1 U3229 ( .A(mem[914]), .B(n4521), .Y(n1334) );
  INVX1 U3230 ( .A(n1334), .Y(n3328) );
  AND2X1 U3231 ( .A(mem[902]), .B(n4521), .Y(n1322) );
  INVX1 U3232 ( .A(n1322), .Y(n3329) );
  AND2X1 U3233 ( .A(mem[880]), .B(n4522), .Y(n1299) );
  INVX1 U3234 ( .A(n1299), .Y(n3330) );
  AND2X1 U3235 ( .A(mem[868]), .B(n4522), .Y(n1287) );
  INVX1 U3236 ( .A(n1287), .Y(n3331) );
  AND2X1 U3237 ( .A(mem[846]), .B(n4523), .Y(n1264) );
  INVX1 U3238 ( .A(n1264), .Y(n3332) );
  AND2X1 U3239 ( .A(mem[834]), .B(n4523), .Y(n1252) );
  INVX1 U3240 ( .A(n1252), .Y(n3333) );
  AND2X1 U3241 ( .A(mem[812]), .B(n4524), .Y(n1228) );
  INVX1 U3242 ( .A(n1228), .Y(n3334) );
  AND2X1 U3243 ( .A(mem[799]), .B(n4524), .Y(n1215) );
  INVX1 U3244 ( .A(n1215), .Y(n3335) );
  AND2X1 U3245 ( .A(mem[763]), .B(n4525), .Y(n1178) );
  INVX1 U3246 ( .A(n1178), .Y(n3336) );
  AND2X1 U3247 ( .A(mem[762]), .B(n4525), .Y(n1177) );
  INVX1 U3248 ( .A(n1177), .Y(n3337) );
  AND2X1 U3249 ( .A(mem[734]), .B(n4526), .Y(n1148) );
  INVX1 U3250 ( .A(n1148), .Y(n3338) );
  AND2X1 U3251 ( .A(mem[728]), .B(n4526), .Y(n1142) );
  INVX1 U3252 ( .A(n1142), .Y(n3339) );
  AND2X1 U3253 ( .A(mem[699]), .B(n4527), .Y(n1112) );
  INVX1 U3254 ( .A(n1112), .Y(n3340) );
  AND2X1 U3255 ( .A(mem[694]), .B(n4527), .Y(n1107) );
  INVX1 U3256 ( .A(n1107), .Y(n3341) );
  AND2X1 U3257 ( .A(mem[665]), .B(n4528), .Y(n1077) );
  INVX1 U3258 ( .A(n1077), .Y(n3342) );
  AND2X1 U3259 ( .A(mem[660]), .B(n4528), .Y(n1072) );
  INVX1 U3260 ( .A(n1072), .Y(n3343) );
  AND2X1 U3261 ( .A(mem[654]), .B(n4529), .Y(n1065) );
  INVX1 U3262 ( .A(n1065), .Y(n3344) );
  AND2X1 U3263 ( .A(mem[642]), .B(n4529), .Y(n1053) );
  INVX1 U3264 ( .A(n1053), .Y(n3345) );
  AND2X1 U3265 ( .A(mem[620]), .B(n4530), .Y(n1030) );
  INVX1 U3266 ( .A(n1030), .Y(n3346) );
  AND2X1 U3267 ( .A(mem[608]), .B(n4530), .Y(n1018) );
  INVX1 U3268 ( .A(n1018), .Y(n3347) );
  AND2X1 U3269 ( .A(mem[586]), .B(n4531), .Y(n995) );
  INVX1 U3270 ( .A(n995), .Y(n3348) );
  AND2X1 U3271 ( .A(mem[574]), .B(n4531), .Y(n983) );
  INVX1 U3272 ( .A(n983), .Y(n3349) );
  AND2X1 U3273 ( .A(mem[552]), .B(n4532), .Y(n959) );
  INVX1 U3274 ( .A(n959), .Y(n3350) );
  AND2X1 U3275 ( .A(mem[540]), .B(n4532), .Y(n947) );
  INVX1 U3276 ( .A(n947), .Y(n3351) );
  AND2X1 U3277 ( .A(mem[518]), .B(n4533), .Y(n924) );
  INVX1 U3278 ( .A(n924), .Y(n3352) );
  AND2X1 U3279 ( .A(mem[506]), .B(n4533), .Y(n912) );
  INVX1 U3280 ( .A(n912), .Y(n3353) );
  AND2X1 U3281 ( .A(mem[484]), .B(n4534), .Y(n889) );
  INVX1 U3282 ( .A(n889), .Y(n3354) );
  AND2X1 U3283 ( .A(mem[472]), .B(n4534), .Y(n877) );
  INVX1 U3284 ( .A(n877), .Y(n3355) );
  AND2X1 U3285 ( .A(mem[450]), .B(n4535), .Y(n854) );
  INVX1 U3286 ( .A(n854), .Y(n3356) );
  AND2X1 U3287 ( .A(mem[438]), .B(n4535), .Y(n842) );
  INVX1 U3288 ( .A(n842), .Y(n3357) );
  AND2X1 U3289 ( .A(mem[416]), .B(n4536), .Y(n819) );
  INVX1 U3290 ( .A(n819), .Y(n3358) );
  AND2X1 U3291 ( .A(mem[403]), .B(n4536), .Y(n806) );
  INVX1 U3292 ( .A(n806), .Y(n3359) );
  AND2X1 U3293 ( .A(mem[367]), .B(n4537), .Y(n769) );
  INVX1 U3294 ( .A(n769), .Y(n3360) );
  AND2X1 U3295 ( .A(mem[366]), .B(n4537), .Y(n768) );
  INVX1 U3296 ( .A(n768), .Y(n3361) );
  AND2X1 U3297 ( .A(mem[338]), .B(n4538), .Y(n739) );
  INVX1 U3298 ( .A(n739), .Y(n3362) );
  AND2X1 U3299 ( .A(mem[332]), .B(n4538), .Y(n733) );
  INVX1 U3300 ( .A(n733), .Y(n3363) );
  AND2X1 U3301 ( .A(mem[303]), .B(n4539), .Y(n703) );
  INVX1 U3302 ( .A(n703), .Y(n3364) );
  AND2X1 U3303 ( .A(mem[298]), .B(n4539), .Y(n698) );
  INVX1 U3304 ( .A(n698), .Y(n3365) );
  AND2X1 U3305 ( .A(mem[269]), .B(n4540), .Y(n667) );
  INVX1 U3306 ( .A(n667), .Y(n3366) );
  AND2X1 U3307 ( .A(mem[264]), .B(n4540), .Y(n662) );
  INVX1 U3308 ( .A(n662), .Y(n3367) );
  AND2X1 U3309 ( .A(mem[254]), .B(n4541), .Y(n650) );
  INVX1 U3310 ( .A(n650), .Y(n3368) );
  AND2X1 U3311 ( .A(mem[242]), .B(n4541), .Y(n638) );
  INVX1 U3312 ( .A(n638), .Y(n3369) );
  AND2X1 U3313 ( .A(mem[220]), .B(n4542), .Y(n614) );
  INVX1 U3314 ( .A(n614), .Y(n3370) );
  AND2X1 U3315 ( .A(mem[208]), .B(n4542), .Y(n602) );
  INVX1 U3316 ( .A(n602), .Y(n3371) );
  AND2X1 U3317 ( .A(mem[186]), .B(n4543), .Y(n578) );
  INVX1 U3318 ( .A(n578), .Y(n3372) );
  AND2X1 U3319 ( .A(mem[174]), .B(n4543), .Y(n566) );
  INVX1 U3320 ( .A(n566), .Y(n3373) );
  AND2X1 U3321 ( .A(mem[152]), .B(n4544), .Y(n542) );
  INVX1 U3322 ( .A(n542), .Y(n3374) );
  AND2X1 U3323 ( .A(mem[139]), .B(n4544), .Y(n529) );
  INVX1 U3324 ( .A(n529), .Y(n3375) );
  AND2X1 U3325 ( .A(mem[103]), .B(n4545), .Y(n491) );
  INVX1 U3326 ( .A(n491), .Y(n3376) );
  AND2X1 U3327 ( .A(mem[102]), .B(n4545), .Y(n490) );
  INVX1 U3328 ( .A(n490), .Y(n3377) );
  AND2X1 U3329 ( .A(mem[74]), .B(n4546), .Y(n460) );
  INVX1 U3330 ( .A(n460), .Y(n3378) );
  AND2X1 U3331 ( .A(mem[68]), .B(n4546), .Y(n454) );
  INVX1 U3332 ( .A(n454), .Y(n3379) );
  AND2X1 U3333 ( .A(mem[39]), .B(n4547), .Y(n423) );
  INVX1 U3334 ( .A(n423), .Y(n3380) );
  AND2X1 U3335 ( .A(mem[34]), .B(n4547), .Y(n418) );
  INVX1 U3336 ( .A(n418), .Y(n3381) );
  AND2X1 U3337 ( .A(mem[5]), .B(n4548), .Y(n359) );
  INVX1 U3338 ( .A(n359), .Y(n3382) );
  AND2X1 U3339 ( .A(mem[0]), .B(n4548), .Y(n349) );
  INVX1 U3340 ( .A(n349), .Y(n3383) );
  INVX1 U3341 ( .A(n1488), .Y(n3384) );
  AND2X2 U3342 ( .A(get), .B(empty_bar), .Y(n1528) );
  INVX1 U3343 ( .A(n1528), .Y(n3385) );
  BUFX2 U3344 ( .A(n4624), .Y(empty_bar) );
  BUFX2 U3345 ( .A(n696), .Y(n3387) );
  INVX1 U3346 ( .A(n4444), .Y(n4469) );
  INVX1 U3347 ( .A(n4444), .Y(n4470) );
  INVX1 U3348 ( .A(n4444), .Y(n4471) );
  INVX1 U3349 ( .A(n4447), .Y(n4472) );
  INVX1 U3350 ( .A(n4444), .Y(n4473) );
  INVX1 U3351 ( .A(n4450), .Y(n4474) );
  INVX1 U3352 ( .A(n4449), .Y(n4475) );
  INVX1 U3353 ( .A(n4449), .Y(n4476) );
  INVX1 U3354 ( .A(n4448), .Y(n4477) );
  INVX1 U3355 ( .A(n4449), .Y(n4478) );
  INVX1 U3356 ( .A(n4448), .Y(n4479) );
  INVX1 U3357 ( .A(n4450), .Y(n4480) );
  INVX1 U3358 ( .A(n4446), .Y(n4481) );
  INVX1 U3359 ( .A(n4445), .Y(n4482) );
  INVX1 U3360 ( .A(n4448), .Y(n4483) );
  INVX1 U3361 ( .A(n4450), .Y(n4484) );
  INVX1 U3362 ( .A(n4444), .Y(n4485) );
  INVX1 U3363 ( .A(n4444), .Y(n4486) );
  INVX1 U3364 ( .A(n4446), .Y(n4487) );
  INVX1 U3365 ( .A(n4446), .Y(n4488) );
  INVX1 U3366 ( .A(n4445), .Y(n4489) );
  INVX1 U3367 ( .A(n4447), .Y(n4490) );
  INVX1 U3368 ( .A(n4445), .Y(n4491) );
  INVX1 U3369 ( .A(n4445), .Y(n4492) );
  INVX1 U3370 ( .A(n4584), .Y(n4495) );
  INVX1 U3371 ( .A(n4584), .Y(n4496) );
  INVX1 U3372 ( .A(n4584), .Y(n4497) );
  INVX1 U3373 ( .A(n4584), .Y(n4498) );
  INVX1 U3374 ( .A(n4584), .Y(n4499) );
  INVX1 U3375 ( .A(n4584), .Y(n4500) );
  INVX1 U3376 ( .A(n4584), .Y(n4501) );
  INVX1 U3377 ( .A(n4584), .Y(n4502) );
  INVX1 U3378 ( .A(n4584), .Y(n4503) );
  INVX1 U3379 ( .A(n4584), .Y(n4504) );
  INVX1 U3380 ( .A(n4584), .Y(n4505) );
  INVX1 U3381 ( .A(n4584), .Y(n4506) );
  INVX1 U3382 ( .A(n4584), .Y(n4507) );
  INVX1 U3383 ( .A(n4584), .Y(n4508) );
  INVX1 U3384 ( .A(n4584), .Y(n4509) );
  INVX1 U3385 ( .A(n4584), .Y(n4510) );
  INVX1 U3386 ( .A(n4584), .Y(n4511) );
  INVX1 U3387 ( .A(n4584), .Y(n4512) );
  INVX1 U3388 ( .A(n4450), .Y(n4451) );
  INVX1 U3389 ( .A(n4450), .Y(n4452) );
  INVX1 U3390 ( .A(n4450), .Y(n4453) );
  INVX1 U3391 ( .A(n4449), .Y(n4454) );
  INVX1 U3392 ( .A(n4449), .Y(n4455) );
  INVX1 U3393 ( .A(n4449), .Y(n4456) );
  INVX1 U3394 ( .A(n4448), .Y(n4457) );
  INVX1 U3395 ( .A(n4448), .Y(n4458) );
  INVX1 U3396 ( .A(n4448), .Y(n4459) );
  INVX1 U3397 ( .A(n4447), .Y(n4460) );
  INVX1 U3398 ( .A(n4447), .Y(n4461) );
  INVX1 U3399 ( .A(n4447), .Y(n4462) );
  INVX1 U3400 ( .A(n4446), .Y(n4463) );
  INVX1 U3401 ( .A(n4446), .Y(n4464) );
  INVX1 U3402 ( .A(n4446), .Y(n4465) );
  INVX1 U3403 ( .A(n4445), .Y(n4466) );
  INVX1 U3404 ( .A(n4445), .Y(n4467) );
  INVX1 U3405 ( .A(n4445), .Y(n4468) );
  INVX1 U3406 ( .A(n4514), .Y(n4515) );
  INVX1 U3407 ( .A(n4514), .Y(n4516) );
  INVX1 U3408 ( .A(n4447), .Y(n4493) );
  INVX1 U3409 ( .A(n4446), .Y(n4494) );
  INVX1 U3410 ( .A(n4584), .Y(n4513) );
  INVX1 U3411 ( .A(n414), .Y(n4548) );
  INVX1 U3412 ( .A(n12), .Y(n4444) );
  INVX1 U3413 ( .A(n12), .Y(n4450) );
  INVX1 U3414 ( .A(n12), .Y(n4449) );
  INVX1 U3415 ( .A(n12), .Y(n4448) );
  INVX1 U3416 ( .A(n12), .Y(n4447) );
  INVX1 U3417 ( .A(n12), .Y(n4446) );
  INVX1 U3418 ( .A(n12), .Y(n4445) );
  INVX1 U3419 ( .A(n14), .Y(n4514) );
  INVX1 U3420 ( .A(n450), .Y(n4547) );
  INVX1 U3421 ( .A(n485), .Y(n4546) );
  INVX1 U3422 ( .A(n520), .Y(n4545) );
  INVX1 U3423 ( .A(n555), .Y(n4544) );
  INVX1 U3424 ( .A(n590), .Y(n4543) );
  INVX1 U3425 ( .A(n625), .Y(n4542) );
  INVX1 U3426 ( .A(n660), .Y(n4541) );
  INVX1 U3427 ( .A(n695), .Y(n4540) );
  INVX1 U3428 ( .A(n730), .Y(n4539) );
  INVX1 U3429 ( .A(n764), .Y(n4538) );
  INVX1 U3430 ( .A(n798), .Y(n4537) );
  INVX1 U3431 ( .A(n832), .Y(n4536) );
  INVX1 U3432 ( .A(n866), .Y(n4535) );
  INVX1 U3433 ( .A(n900), .Y(n4534) );
  INVX1 U3434 ( .A(n934), .Y(n4533) );
  INVX1 U3435 ( .A(n968), .Y(n4532) );
  INVX1 U3436 ( .A(n1003), .Y(n4531) );
  INVX1 U3437 ( .A(n1037), .Y(n4530) );
  INVX1 U3438 ( .A(n1071), .Y(n4529) );
  INVX1 U3439 ( .A(n1105), .Y(n4528) );
  INVX1 U3440 ( .A(n1139), .Y(n4527) );
  INVX1 U3441 ( .A(n1173), .Y(n4526) );
  INVX1 U3442 ( .A(n1207), .Y(n4525) );
  INVX1 U3443 ( .A(n1241), .Y(n4524) );
  INVX1 U3444 ( .A(n1276), .Y(n4523) );
  INVX1 U3445 ( .A(n1310), .Y(n4522) );
  INVX1 U3446 ( .A(n1344), .Y(n4521) );
  INVX1 U3447 ( .A(n1378), .Y(n4520) );
  INVX1 U3448 ( .A(n1412), .Y(n4519) );
  INVX1 U3449 ( .A(n1446), .Y(n4518) );
  INVX1 U3450 ( .A(n1480), .Y(n4517) );
  INVX1 U3451 ( .A(n3388), .Y(n4570) );
  INVX1 U3452 ( .A(n3389), .Y(n4569) );
  INVX1 U3453 ( .A(n3390), .Y(n4568) );
  INVX1 U3454 ( .A(n3391), .Y(n4567) );
  INVX1 U3455 ( .A(n3392), .Y(n4566) );
  INVX1 U3456 ( .A(n3393), .Y(n4565) );
  INVX1 U3457 ( .A(n3394), .Y(n4564) );
  INVX1 U3458 ( .A(n3395), .Y(n4563) );
  INVX1 U3459 ( .A(n3396), .Y(n4562) );
  INVX1 U3460 ( .A(n3397), .Y(n4561) );
  INVX1 U3461 ( .A(n3398), .Y(n4560) );
  INVX1 U3462 ( .A(n3399), .Y(n4559) );
  INVX1 U3463 ( .A(n3400), .Y(n4558) );
  INVX1 U3464 ( .A(n3401), .Y(n4557) );
  INVX1 U3465 ( .A(n3402), .Y(n4556) );
  INVX1 U3466 ( .A(n3403), .Y(n4555) );
  INVX1 U3467 ( .A(n3404), .Y(n4554) );
  INVX1 U3468 ( .A(n3405), .Y(n4553) );
  INVX1 U3469 ( .A(n3406), .Y(n4552) );
  INVX1 U3470 ( .A(n3407), .Y(n4551) );
  INVX1 U3471 ( .A(n3408), .Y(n4550) );
  INVX1 U3472 ( .A(n3409), .Y(n4549) );
  INVX1 U3473 ( .A(n3410), .Y(n4581) );
  INVX1 U3474 ( .A(n3411), .Y(n4580) );
  INVX1 U3475 ( .A(n3412), .Y(n4579) );
  INVX1 U3476 ( .A(n3413), .Y(n4578) );
  INVX1 U3477 ( .A(n3414), .Y(n4577) );
  INVX1 U3478 ( .A(n3415), .Y(n4576) );
  INVX1 U3479 ( .A(n3416), .Y(n4575) );
  INVX1 U3480 ( .A(n3417), .Y(n4574) );
  INVX1 U3481 ( .A(n3418), .Y(n4573) );
  INVX1 U3482 ( .A(n3419), .Y(n4572) );
  INVX1 U3483 ( .A(n3420), .Y(n4571) );
  INVX1 U3484 ( .A(wr_ptr[2]), .Y(n4622) );
  INVX1 U3485 ( .A(wr_ptr[0]), .Y(n4619) );
  INVX1 U3486 ( .A(n1), .Y(n4586) );
  INVX1 U3487 ( .A(n4411), .Y(n88) );
  INVX1 U3488 ( .A(n2), .Y(n4587) );
  INVX1 U3489 ( .A(n4412), .Y(n87) );
  INVX1 U3490 ( .A(n3), .Y(n4588) );
  INVX1 U3491 ( .A(n4413), .Y(n86) );
  INVX1 U3492 ( .A(n4), .Y(n4589) );
  INVX1 U3493 ( .A(n4414), .Y(n85) );
  INVX1 U3494 ( .A(n5), .Y(n4590) );
  INVX1 U3495 ( .A(n4415), .Y(n84) );
  INVX1 U3496 ( .A(n6), .Y(n4591) );
  INVX1 U3497 ( .A(n4416), .Y(n83) );
  INVX1 U3498 ( .A(n7), .Y(n4592) );
  INVX1 U3499 ( .A(n4417), .Y(n82) );
  INVX1 U3500 ( .A(n8), .Y(n4593) );
  INVX1 U3501 ( .A(n4418), .Y(n81) );
  INVX1 U3502 ( .A(n9), .Y(n4594) );
  INVX1 U3503 ( .A(n4419), .Y(n80) );
  INVX1 U3504 ( .A(n10), .Y(n4595) );
  INVX1 U3505 ( .A(n4420), .Y(n79) );
  INVX1 U3506 ( .A(n11), .Y(n4596) );
  INVX1 U3507 ( .A(n4421), .Y(n78) );
  INVX1 U3508 ( .A(n17), .Y(n4597) );
  INVX1 U3509 ( .A(n4422), .Y(n77) );
  INVX1 U3510 ( .A(n18), .Y(n4598) );
  INVX1 U3511 ( .A(n4423), .Y(n76) );
  INVX1 U3512 ( .A(n19), .Y(n4599) );
  INVX1 U3513 ( .A(n4424), .Y(n75) );
  INVX1 U3514 ( .A(n24), .Y(n4600) );
  INVX1 U3515 ( .A(n4425), .Y(n74) );
  INVX1 U3516 ( .A(n25), .Y(n4601) );
  INVX1 U3517 ( .A(n4426), .Y(n73) );
  INVX1 U3518 ( .A(n26), .Y(n4602) );
  INVX1 U3519 ( .A(n4427), .Y(n72) );
  INVX1 U3520 ( .A(n27), .Y(n4603) );
  INVX1 U3521 ( .A(n4428), .Y(n71) );
  INVX1 U3522 ( .A(n28), .Y(n4604) );
  INVX1 U3523 ( .A(n4429), .Y(n70) );
  INVX1 U3524 ( .A(n29), .Y(n4605) );
  INVX1 U3525 ( .A(n4430), .Y(n69) );
  INVX1 U3526 ( .A(n30), .Y(n4606) );
  INVX1 U3527 ( .A(n4431), .Y(n68) );
  INVX1 U3528 ( .A(n31), .Y(n4607) );
  INVX1 U3529 ( .A(n4432), .Y(n67) );
  INVX1 U3530 ( .A(n32), .Y(n4608) );
  INVX1 U3531 ( .A(n4433), .Y(n66) );
  INVX1 U3532 ( .A(n33), .Y(n4609) );
  INVX1 U3533 ( .A(n4434), .Y(n65) );
  INVX1 U3534 ( .A(n34), .Y(n4610) );
  INVX1 U3535 ( .A(n4435), .Y(n64) );
  INVX1 U3536 ( .A(n35), .Y(n4611) );
  INVX1 U3537 ( .A(n4436), .Y(n63) );
  INVX1 U3538 ( .A(n36), .Y(n4612) );
  INVX1 U3539 ( .A(n4437), .Y(n62) );
  INVX1 U3540 ( .A(n37), .Y(n4613) );
  INVX1 U3541 ( .A(n4438), .Y(n61) );
  INVX1 U3542 ( .A(n38), .Y(n4614) );
  INVX1 U3543 ( .A(n4439), .Y(n60) );
  INVX1 U3544 ( .A(n39), .Y(n4615) );
  INVX1 U3545 ( .A(n4440), .Y(n59) );
  INVX1 U3546 ( .A(n40), .Y(n4616) );
  INVX1 U3547 ( .A(n4441), .Y(n58) );
  INVX1 U3548 ( .A(n41), .Y(n4617) );
  INVX1 U3549 ( .A(n4442), .Y(n57) );
  INVX1 U3550 ( .A(n42), .Y(n4618) );
  INVX1 U3551 ( .A(n4443), .Y(n56) );
  INVX1 U3552 ( .A(wr_ptr[1]), .Y(n4621) );
  INVX1 U3553 ( .A(wr_ptr[3]), .Y(n4623) );
  INVX1 U3554 ( .A(wr_ptr[4]), .Y(n4620) );
  INVX1 U3555 ( .A(n13), .Y(n4584) );
  INVX1 U3556 ( .A(n16), .Y(n4582) );
  INVX1 U3557 ( .A(n15), .Y(n4583) );
  INVX1 U3558 ( .A(n12), .Y(n4585) );
  INVX1 U3559 ( .A(sub_93_carry[5]), .Y(fillcount[5]) );
  AND2X1 U3560 ( .A(data_in[11]), .B(reset), .Y(n3388) );
  AND2X1 U3561 ( .A(data_in[12]), .B(reset), .Y(n3389) );
  AND2X1 U3562 ( .A(data_in[13]), .B(reset), .Y(n3390) );
  AND2X1 U3563 ( .A(data_in[14]), .B(reset), .Y(n3391) );
  AND2X1 U3564 ( .A(data_in[15]), .B(reset), .Y(n3392) );
  AND2X1 U3565 ( .A(data_in[16]), .B(reset), .Y(n3393) );
  AND2X1 U3566 ( .A(data_in[17]), .B(reset), .Y(n3394) );
  AND2X1 U3567 ( .A(data_in[18]), .B(reset), .Y(n3395) );
  AND2X1 U3568 ( .A(data_in[19]), .B(reset), .Y(n3396) );
  AND2X1 U3569 ( .A(data_in[20]), .B(reset), .Y(n3397) );
  AND2X1 U3570 ( .A(data_in[21]), .B(reset), .Y(n3398) );
  AND2X1 U3571 ( .A(data_in[22]), .B(reset), .Y(n3399) );
  AND2X1 U3572 ( .A(data_in[23]), .B(reset), .Y(n3400) );
  AND2X1 U3573 ( .A(data_in[24]), .B(reset), .Y(n3401) );
  AND2X1 U3574 ( .A(data_in[25]), .B(reset), .Y(n3402) );
  AND2X1 U3575 ( .A(data_in[26]), .B(reset), .Y(n3403) );
  AND2X1 U3576 ( .A(data_in[27]), .B(reset), .Y(n3404) );
  AND2X1 U3577 ( .A(data_in[28]), .B(reset), .Y(n3405) );
  AND2X1 U3578 ( .A(data_in[29]), .B(reset), .Y(n3406) );
  AND2X1 U3579 ( .A(data_in[30]), .B(reset), .Y(n3407) );
  AND2X1 U3580 ( .A(data_in[31]), .B(reset), .Y(n3408) );
  AND2X1 U3581 ( .A(data_in[32]), .B(reset), .Y(n3409) );
  AND2X1 U3582 ( .A(data_in[0]), .B(reset), .Y(n3410) );
  AND2X1 U3583 ( .A(data_in[1]), .B(reset), .Y(n3411) );
  AND2X1 U3584 ( .A(data_in[2]), .B(reset), .Y(n3412) );
  AND2X1 U3585 ( .A(data_in[3]), .B(reset), .Y(n3413) );
  AND2X1 U3586 ( .A(data_in[4]), .B(reset), .Y(n3414) );
  AND2X1 U3587 ( .A(data_in[5]), .B(reset), .Y(n3415) );
  AND2X1 U3588 ( .A(data_in[6]), .B(reset), .Y(n3416) );
  AND2X1 U3589 ( .A(data_in[7]), .B(reset), .Y(n3417) );
  AND2X1 U3590 ( .A(data_in[8]), .B(reset), .Y(n3418) );
  AND2X1 U3591 ( .A(data_in[9]), .B(reset), .Y(n3419) );
  AND2X1 U3592 ( .A(data_in[10]), .B(reset), .Y(n3420) );
  MUX2X1 U3593 ( .B(n3422), .A(n3423), .S(n4495), .Y(n3421) );
  MUX2X1 U3594 ( .B(n3425), .A(n3426), .S(n4495), .Y(n3424) );
  MUX2X1 U3595 ( .B(n3428), .A(n3429), .S(n4495), .Y(n3427) );
  MUX2X1 U3596 ( .B(n3431), .A(n3432), .S(n4495), .Y(n3430) );
  MUX2X1 U3597 ( .B(n3434), .A(n3435), .S(n15), .Y(n3433) );
  MUX2X1 U3598 ( .B(n3437), .A(n3438), .S(n4495), .Y(n3436) );
  MUX2X1 U3599 ( .B(n3440), .A(n3441), .S(n4495), .Y(n3439) );
  MUX2X1 U3600 ( .B(n3443), .A(n3444), .S(n4495), .Y(n3442) );
  MUX2X1 U3601 ( .B(n3446), .A(n3447), .S(n4495), .Y(n3445) );
  MUX2X1 U3602 ( .B(n3449), .A(n3450), .S(n15), .Y(n3448) );
  MUX2X1 U3603 ( .B(n3452), .A(n3453), .S(n4495), .Y(n3451) );
  MUX2X1 U3604 ( .B(n3455), .A(n3456), .S(n4495), .Y(n3454) );
  MUX2X1 U3605 ( .B(n3458), .A(n3459), .S(n4495), .Y(n3457) );
  MUX2X1 U3606 ( .B(n3461), .A(n3462), .S(n4495), .Y(n3460) );
  MUX2X1 U3607 ( .B(n3464), .A(n3465), .S(n15), .Y(n3463) );
  MUX2X1 U3608 ( .B(n3467), .A(n3468), .S(n4496), .Y(n3466) );
  MUX2X1 U3609 ( .B(n3470), .A(n3471), .S(n4496), .Y(n3469) );
  MUX2X1 U3610 ( .B(n3473), .A(n3474), .S(n4496), .Y(n3472) );
  MUX2X1 U3611 ( .B(n3476), .A(n3477), .S(n4496), .Y(n3475) );
  MUX2X1 U3612 ( .B(n3479), .A(n3480), .S(n15), .Y(n3478) );
  MUX2X1 U3613 ( .B(n3482), .A(n3483), .S(n4496), .Y(n3481) );
  MUX2X1 U3614 ( .B(n3485), .A(n3486), .S(n4496), .Y(n3484) );
  MUX2X1 U3615 ( .B(n3488), .A(n3489), .S(n4496), .Y(n3487) );
  MUX2X1 U3616 ( .B(n3491), .A(n3492), .S(n4496), .Y(n3490) );
  MUX2X1 U3617 ( .B(n3494), .A(n3495), .S(n15), .Y(n3493) );
  MUX2X1 U3618 ( .B(n3497), .A(n3498), .S(n4496), .Y(n3496) );
  MUX2X1 U3619 ( .B(n3500), .A(n3501), .S(n4496), .Y(n3499) );
  MUX2X1 U3620 ( .B(n3503), .A(n3504), .S(n4496), .Y(n3502) );
  MUX2X1 U3621 ( .B(n3506), .A(n3507), .S(n4496), .Y(n3505) );
  MUX2X1 U3622 ( .B(n3509), .A(n3510), .S(n15), .Y(n3508) );
  MUX2X1 U3623 ( .B(n3512), .A(n3513), .S(n4497), .Y(n3511) );
  MUX2X1 U3624 ( .B(n3515), .A(n3516), .S(n4497), .Y(n3514) );
  MUX2X1 U3625 ( .B(n3518), .A(n3519), .S(n4497), .Y(n3517) );
  MUX2X1 U3626 ( .B(n3521), .A(n3522), .S(n4497), .Y(n3520) );
  MUX2X1 U3627 ( .B(n3524), .A(n3525), .S(n15), .Y(n3523) );
  MUX2X1 U3628 ( .B(n3527), .A(n3528), .S(n4497), .Y(n3526) );
  MUX2X1 U3629 ( .B(n3530), .A(n3531), .S(n4497), .Y(n3529) );
  MUX2X1 U3630 ( .B(n3533), .A(n3534), .S(n4497), .Y(n3532) );
  MUX2X1 U3631 ( .B(n3536), .A(n3537), .S(n4497), .Y(n3535) );
  MUX2X1 U3632 ( .B(n3539), .A(n3540), .S(n15), .Y(n3538) );
  MUX2X1 U3633 ( .B(n3542), .A(n3543), .S(n4497), .Y(n3541) );
  MUX2X1 U3634 ( .B(n3545), .A(n3546), .S(n4497), .Y(n3544) );
  MUX2X1 U3635 ( .B(n3548), .A(n3549), .S(n4497), .Y(n3547) );
  MUX2X1 U3636 ( .B(n3551), .A(n3552), .S(n4497), .Y(n3550) );
  MUX2X1 U3637 ( .B(n3554), .A(n3555), .S(n15), .Y(n3553) );
  MUX2X1 U3638 ( .B(n3557), .A(n3558), .S(n4498), .Y(n3556) );
  MUX2X1 U3639 ( .B(n3560), .A(n3561), .S(n4498), .Y(n3559) );
  MUX2X1 U3640 ( .B(n3563), .A(n3564), .S(n4498), .Y(n3562) );
  MUX2X1 U3641 ( .B(n3566), .A(n3567), .S(n4498), .Y(n3565) );
  MUX2X1 U3642 ( .B(n3569), .A(n3570), .S(n15), .Y(n3568) );
  MUX2X1 U3643 ( .B(n3572), .A(n3573), .S(n4498), .Y(n3571) );
  MUX2X1 U3644 ( .B(n3575), .A(n3576), .S(n4498), .Y(n3574) );
  MUX2X1 U3645 ( .B(n3578), .A(n3579), .S(n4498), .Y(n3577) );
  MUX2X1 U3646 ( .B(n3581), .A(n3582), .S(n4498), .Y(n3580) );
  MUX2X1 U3647 ( .B(n3584), .A(n3585), .S(n15), .Y(n3583) );
  MUX2X1 U3648 ( .B(n3587), .A(n3588), .S(n4498), .Y(n3586) );
  MUX2X1 U3649 ( .B(n3590), .A(n3591), .S(n4498), .Y(n3589) );
  MUX2X1 U3650 ( .B(n3593), .A(n3594), .S(n4498), .Y(n3592) );
  MUX2X1 U3651 ( .B(n3596), .A(n3597), .S(n4498), .Y(n3595) );
  MUX2X1 U3652 ( .B(n3599), .A(n3600), .S(n15), .Y(n3598) );
  MUX2X1 U3653 ( .B(n3602), .A(n3603), .S(n4499), .Y(n3601) );
  MUX2X1 U3654 ( .B(n3605), .A(n3606), .S(n4499), .Y(n3604) );
  MUX2X1 U3655 ( .B(n3608), .A(n3609), .S(n4499), .Y(n3607) );
  MUX2X1 U3656 ( .B(n3611), .A(n3612), .S(n4499), .Y(n3610) );
  MUX2X1 U3657 ( .B(n3614), .A(n3615), .S(n15), .Y(n3613) );
  MUX2X1 U3658 ( .B(n3617), .A(n3618), .S(n4499), .Y(n3616) );
  MUX2X1 U3659 ( .B(n3620), .A(n3621), .S(n4499), .Y(n3619) );
  MUX2X1 U3660 ( .B(n3623), .A(n3624), .S(n4499), .Y(n3622) );
  MUX2X1 U3661 ( .B(n3626), .A(n3627), .S(n4499), .Y(n3625) );
  MUX2X1 U3662 ( .B(n3629), .A(n3630), .S(n15), .Y(n3628) );
  MUX2X1 U3663 ( .B(n3632), .A(n3633), .S(n4499), .Y(n3631) );
  MUX2X1 U3664 ( .B(n3635), .A(n3636), .S(n4499), .Y(n3634) );
  MUX2X1 U3665 ( .B(n3638), .A(n3639), .S(n4499), .Y(n3637) );
  MUX2X1 U3666 ( .B(n3641), .A(n3642), .S(n4499), .Y(n3640) );
  MUX2X1 U3667 ( .B(n3644), .A(n3645), .S(n15), .Y(n3643) );
  MUX2X1 U3668 ( .B(n3647), .A(n3648), .S(n4500), .Y(n3646) );
  MUX2X1 U3669 ( .B(n3650), .A(n3651), .S(n4500), .Y(n3649) );
  MUX2X1 U3670 ( .B(n3653), .A(n3654), .S(n4500), .Y(n3652) );
  MUX2X1 U3671 ( .B(n3656), .A(n3657), .S(n4500), .Y(n3655) );
  MUX2X1 U3672 ( .B(n3659), .A(n3660), .S(n15), .Y(n3658) );
  MUX2X1 U3673 ( .B(n3662), .A(n3663), .S(n4500), .Y(n3661) );
  MUX2X1 U3674 ( .B(n3665), .A(n3666), .S(n4500), .Y(n3664) );
  MUX2X1 U3675 ( .B(n3668), .A(n3669), .S(n4500), .Y(n3667) );
  MUX2X1 U3676 ( .B(n3671), .A(n3672), .S(n4500), .Y(n3670) );
  MUX2X1 U3677 ( .B(n3674), .A(n3675), .S(n15), .Y(n3673) );
  MUX2X1 U3678 ( .B(n3677), .A(n3678), .S(n4500), .Y(n3676) );
  MUX2X1 U3679 ( .B(n3680), .A(n3681), .S(n4500), .Y(n3679) );
  MUX2X1 U3680 ( .B(n3683), .A(n3684), .S(n4500), .Y(n3682) );
  MUX2X1 U3681 ( .B(n3686), .A(n3687), .S(n4500), .Y(n3685) );
  MUX2X1 U3682 ( .B(n3689), .A(n3690), .S(n15), .Y(n3688) );
  MUX2X1 U3683 ( .B(n3692), .A(n3693), .S(n4501), .Y(n3691) );
  MUX2X1 U3684 ( .B(n3695), .A(n3696), .S(n4501), .Y(n3694) );
  MUX2X1 U3685 ( .B(n3698), .A(n3699), .S(n4501), .Y(n3697) );
  MUX2X1 U3686 ( .B(n3701), .A(n3702), .S(n4501), .Y(n3700) );
  MUX2X1 U3687 ( .B(n3704), .A(n3705), .S(n15), .Y(n3703) );
  MUX2X1 U3688 ( .B(n3707), .A(n3708), .S(n4501), .Y(n3706) );
  MUX2X1 U3689 ( .B(n3710), .A(n3711), .S(n4501), .Y(n3709) );
  MUX2X1 U3690 ( .B(n3713), .A(n3714), .S(n4501), .Y(n3712) );
  MUX2X1 U3691 ( .B(n3716), .A(n3717), .S(n4501), .Y(n3715) );
  MUX2X1 U3692 ( .B(n3719), .A(n3720), .S(n15), .Y(n3718) );
  MUX2X1 U3693 ( .B(n3722), .A(n3723), .S(n4501), .Y(n3721) );
  MUX2X1 U3694 ( .B(n3725), .A(n3726), .S(n4501), .Y(n3724) );
  MUX2X1 U3695 ( .B(n3728), .A(n3729), .S(n4501), .Y(n3727) );
  MUX2X1 U3696 ( .B(n3731), .A(n3732), .S(n4501), .Y(n3730) );
  MUX2X1 U3697 ( .B(n3734), .A(n3735), .S(n15), .Y(n3733) );
  MUX2X1 U3698 ( .B(n3737), .A(n3738), .S(n4502), .Y(n3736) );
  MUX2X1 U3699 ( .B(n3740), .A(n3741), .S(n4502), .Y(n3739) );
  MUX2X1 U3700 ( .B(n3743), .A(n3744), .S(n4502), .Y(n3742) );
  MUX2X1 U3701 ( .B(n3746), .A(n3747), .S(n4502), .Y(n3745) );
  MUX2X1 U3702 ( .B(n3749), .A(n3750), .S(n15), .Y(n3748) );
  MUX2X1 U3703 ( .B(n3752), .A(n3753), .S(n4502), .Y(n3751) );
  MUX2X1 U3704 ( .B(n3755), .A(n3756), .S(n4502), .Y(n3754) );
  MUX2X1 U3705 ( .B(n3758), .A(n3759), .S(n4502), .Y(n3757) );
  MUX2X1 U3706 ( .B(n3761), .A(n3762), .S(n4502), .Y(n3760) );
  MUX2X1 U3707 ( .B(n3764), .A(n3765), .S(n15), .Y(n3763) );
  MUX2X1 U3708 ( .B(n3767), .A(n3768), .S(n4502), .Y(n3766) );
  MUX2X1 U3709 ( .B(n3770), .A(n3771), .S(n4502), .Y(n3769) );
  MUX2X1 U3710 ( .B(n3773), .A(n3774), .S(n4502), .Y(n3772) );
  MUX2X1 U3711 ( .B(n3776), .A(n3777), .S(n4502), .Y(n3775) );
  MUX2X1 U3712 ( .B(n3779), .A(n3780), .S(n15), .Y(n3778) );
  MUX2X1 U3713 ( .B(n3782), .A(n3783), .S(n4503), .Y(n3781) );
  MUX2X1 U3714 ( .B(n3785), .A(n3786), .S(n4503), .Y(n3784) );
  MUX2X1 U3715 ( .B(n3788), .A(n3789), .S(n4503), .Y(n3787) );
  MUX2X1 U3716 ( .B(n3791), .A(n3792), .S(n4503), .Y(n3790) );
  MUX2X1 U3717 ( .B(n3794), .A(n3795), .S(n15), .Y(n3793) );
  MUX2X1 U3718 ( .B(n3797), .A(n3798), .S(n4503), .Y(n3796) );
  MUX2X1 U3719 ( .B(n3800), .A(n3801), .S(n4503), .Y(n3799) );
  MUX2X1 U3720 ( .B(n3803), .A(n3804), .S(n4503), .Y(n3802) );
  MUX2X1 U3721 ( .B(n3806), .A(n3807), .S(n4503), .Y(n3805) );
  MUX2X1 U3722 ( .B(n3809), .A(n3810), .S(n15), .Y(n3808) );
  MUX2X1 U3723 ( .B(n3812), .A(n3813), .S(n4503), .Y(n3811) );
  MUX2X1 U3724 ( .B(n3815), .A(n3816), .S(n4503), .Y(n3814) );
  MUX2X1 U3725 ( .B(n3818), .A(n3819), .S(n4503), .Y(n3817) );
  MUX2X1 U3726 ( .B(n3821), .A(n3822), .S(n4503), .Y(n3820) );
  MUX2X1 U3727 ( .B(n3824), .A(n3825), .S(n15), .Y(n3823) );
  MUX2X1 U3728 ( .B(n3827), .A(n3828), .S(n4504), .Y(n3826) );
  MUX2X1 U3729 ( .B(n3830), .A(n3831), .S(n4504), .Y(n3829) );
  MUX2X1 U3730 ( .B(n3833), .A(n3834), .S(n4504), .Y(n3832) );
  MUX2X1 U3731 ( .B(n3836), .A(n3837), .S(n4504), .Y(n3835) );
  MUX2X1 U3732 ( .B(n3839), .A(n3840), .S(n15), .Y(n3838) );
  MUX2X1 U3733 ( .B(n3842), .A(n3843), .S(n4504), .Y(n3841) );
  MUX2X1 U3734 ( .B(n3845), .A(n3846), .S(n4504), .Y(n3844) );
  MUX2X1 U3735 ( .B(n3848), .A(n3849), .S(n4504), .Y(n3847) );
  MUX2X1 U3736 ( .B(n3851), .A(n3852), .S(n4504), .Y(n3850) );
  MUX2X1 U3737 ( .B(n3854), .A(n3855), .S(n15), .Y(n3853) );
  MUX2X1 U3738 ( .B(n3857), .A(n3858), .S(n4504), .Y(n3856) );
  MUX2X1 U3739 ( .B(n3860), .A(n3861), .S(n4504), .Y(n3859) );
  MUX2X1 U3740 ( .B(n3863), .A(n3864), .S(n4504), .Y(n3862) );
  MUX2X1 U3741 ( .B(n3866), .A(n3867), .S(n4504), .Y(n3865) );
  MUX2X1 U3742 ( .B(n3869), .A(n3870), .S(n15), .Y(n3868) );
  MUX2X1 U3743 ( .B(n3872), .A(n3873), .S(n4505), .Y(n3871) );
  MUX2X1 U3744 ( .B(n3875), .A(n3876), .S(n4505), .Y(n3874) );
  MUX2X1 U3745 ( .B(n3878), .A(n3879), .S(n4505), .Y(n3877) );
  MUX2X1 U3746 ( .B(n3881), .A(n3882), .S(n4505), .Y(n3880) );
  MUX2X1 U3747 ( .B(n3884), .A(n3885), .S(n15), .Y(n3883) );
  MUX2X1 U3748 ( .B(n3887), .A(n3888), .S(n4505), .Y(n3886) );
  MUX2X1 U3749 ( .B(n3890), .A(n3891), .S(n4505), .Y(n3889) );
  MUX2X1 U3750 ( .B(n3893), .A(n3894), .S(n4505), .Y(n3892) );
  MUX2X1 U3751 ( .B(n3896), .A(n3897), .S(n4505), .Y(n3895) );
  MUX2X1 U3752 ( .B(n3899), .A(n3900), .S(n15), .Y(n3898) );
  MUX2X1 U3753 ( .B(n3902), .A(n3903), .S(n4505), .Y(n3901) );
  MUX2X1 U3754 ( .B(n3905), .A(n3906), .S(n4505), .Y(n3904) );
  MUX2X1 U3755 ( .B(n3908), .A(n3909), .S(n4505), .Y(n3907) );
  MUX2X1 U3756 ( .B(n3911), .A(n3912), .S(n4505), .Y(n3910) );
  MUX2X1 U3757 ( .B(n3914), .A(n3915), .S(n15), .Y(n3913) );
  MUX2X1 U3758 ( .B(n3917), .A(n3918), .S(n4506), .Y(n3916) );
  MUX2X1 U3759 ( .B(n3920), .A(n3921), .S(n4506), .Y(n3919) );
  MUX2X1 U3760 ( .B(n3923), .A(n3924), .S(n4506), .Y(n3922) );
  MUX2X1 U3761 ( .B(n3926), .A(n3927), .S(n4506), .Y(n3925) );
  MUX2X1 U3762 ( .B(n3929), .A(n3930), .S(n15), .Y(n3928) );
  MUX2X1 U3763 ( .B(n3932), .A(n3933), .S(n4506), .Y(n3931) );
  MUX2X1 U3764 ( .B(n3935), .A(n3936), .S(n4506), .Y(n3934) );
  MUX2X1 U3765 ( .B(n3938), .A(n3939), .S(n4506), .Y(n3937) );
  MUX2X1 U3766 ( .B(n3941), .A(n3942), .S(n4506), .Y(n3940) );
  MUX2X1 U3767 ( .B(n3944), .A(n3945), .S(n15), .Y(n3943) );
  MUX2X1 U3768 ( .B(n3947), .A(n3948), .S(n4506), .Y(n3946) );
  MUX2X1 U3769 ( .B(n3950), .A(n3951), .S(n4506), .Y(n3949) );
  MUX2X1 U3770 ( .B(n3953), .A(n3954), .S(n4506), .Y(n3952) );
  MUX2X1 U3771 ( .B(n3956), .A(n3957), .S(n4506), .Y(n3955) );
  MUX2X1 U3772 ( .B(n3959), .A(n3960), .S(n15), .Y(n3958) );
  MUX2X1 U3773 ( .B(n3962), .A(n3963), .S(n4507), .Y(n3961) );
  MUX2X1 U3774 ( .B(n3965), .A(n3966), .S(n4507), .Y(n3964) );
  MUX2X1 U3775 ( .B(n3968), .A(n3969), .S(n4507), .Y(n3967) );
  MUX2X1 U3776 ( .B(n3971), .A(n3972), .S(n4507), .Y(n3970) );
  MUX2X1 U3777 ( .B(n3974), .A(n3975), .S(n15), .Y(n3973) );
  MUX2X1 U3778 ( .B(n3977), .A(n3978), .S(n4507), .Y(n3976) );
  MUX2X1 U3779 ( .B(n3980), .A(n3981), .S(n4507), .Y(n3979) );
  MUX2X1 U3780 ( .B(n3983), .A(n3984), .S(n4507), .Y(n3982) );
  MUX2X1 U3781 ( .B(n3986), .A(n3987), .S(n4507), .Y(n3985) );
  MUX2X1 U3782 ( .B(n3989), .A(n3990), .S(n15), .Y(n3988) );
  MUX2X1 U3783 ( .B(n3992), .A(n3993), .S(n4507), .Y(n3991) );
  MUX2X1 U3784 ( .B(n3995), .A(n3996), .S(n4507), .Y(n3994) );
  MUX2X1 U3785 ( .B(n3998), .A(n3999), .S(n4507), .Y(n3997) );
  MUX2X1 U3786 ( .B(n4001), .A(n4002), .S(n4507), .Y(n4000) );
  MUX2X1 U3787 ( .B(n4004), .A(n4005), .S(n15), .Y(n4003) );
  MUX2X1 U3788 ( .B(n4007), .A(n4008), .S(n4508), .Y(n4006) );
  MUX2X1 U3789 ( .B(n4010), .A(n4011), .S(n4508), .Y(n4009) );
  MUX2X1 U3790 ( .B(n4013), .A(n4014), .S(n4508), .Y(n4012) );
  MUX2X1 U3791 ( .B(n4016), .A(n4017), .S(n4508), .Y(n4015) );
  MUX2X1 U3792 ( .B(n4019), .A(n4020), .S(n15), .Y(n4018) );
  MUX2X1 U3793 ( .B(n4022), .A(n4023), .S(n4508), .Y(n4021) );
  MUX2X1 U3794 ( .B(n4025), .A(n4026), .S(n4508), .Y(n4024) );
  MUX2X1 U3795 ( .B(n4028), .A(n4029), .S(n4508), .Y(n4027) );
  MUX2X1 U3796 ( .B(n4031), .A(n4032), .S(n4508), .Y(n4030) );
  MUX2X1 U3797 ( .B(n4034), .A(n4035), .S(n15), .Y(n4033) );
  MUX2X1 U3798 ( .B(n4037), .A(n4038), .S(n4508), .Y(n4036) );
  MUX2X1 U3799 ( .B(n4040), .A(n4041), .S(n4508), .Y(n4039) );
  MUX2X1 U3800 ( .B(n4043), .A(n4044), .S(n4508), .Y(n4042) );
  MUX2X1 U3801 ( .B(n4046), .A(n4047), .S(n4508), .Y(n4045) );
  MUX2X1 U3802 ( .B(n4049), .A(n4050), .S(n15), .Y(n4048) );
  MUX2X1 U3803 ( .B(n4052), .A(n4053), .S(n4509), .Y(n4051) );
  MUX2X1 U3804 ( .B(n4055), .A(n4056), .S(n4509), .Y(n4054) );
  MUX2X1 U3805 ( .B(n4058), .A(n4059), .S(n4509), .Y(n4057) );
  MUX2X1 U3806 ( .B(n4061), .A(n4062), .S(n4509), .Y(n4060) );
  MUX2X1 U3807 ( .B(n4064), .A(n4065), .S(n15), .Y(n4063) );
  MUX2X1 U3808 ( .B(n4067), .A(n4068), .S(n4509), .Y(n4066) );
  MUX2X1 U3809 ( .B(n4070), .A(n4071), .S(n4509), .Y(n4069) );
  MUX2X1 U3810 ( .B(n4073), .A(n4074), .S(n4509), .Y(n4072) );
  MUX2X1 U3811 ( .B(n4076), .A(n4077), .S(n4509), .Y(n4075) );
  MUX2X1 U3812 ( .B(n4079), .A(n4080), .S(n15), .Y(n4078) );
  MUX2X1 U3813 ( .B(n4082), .A(n4083), .S(n4509), .Y(n4081) );
  MUX2X1 U3814 ( .B(n4085), .A(n4086), .S(n4509), .Y(n4084) );
  MUX2X1 U3815 ( .B(n4088), .A(n4089), .S(n4509), .Y(n4087) );
  MUX2X1 U3816 ( .B(n4091), .A(n4092), .S(n4509), .Y(n4090) );
  MUX2X1 U3817 ( .B(n4094), .A(n4095), .S(n15), .Y(n4093) );
  MUX2X1 U3818 ( .B(n4097), .A(n4098), .S(n4510), .Y(n4096) );
  MUX2X1 U3819 ( .B(n4100), .A(n4101), .S(n4510), .Y(n4099) );
  MUX2X1 U3820 ( .B(n4103), .A(n4104), .S(n4510), .Y(n4102) );
  MUX2X1 U3821 ( .B(n4106), .A(n4107), .S(n4510), .Y(n4105) );
  MUX2X1 U3822 ( .B(n4109), .A(n4110), .S(n15), .Y(n4108) );
  MUX2X1 U3823 ( .B(n4112), .A(n4113), .S(n4510), .Y(n4111) );
  MUX2X1 U3824 ( .B(n4115), .A(n4116), .S(n4510), .Y(n4114) );
  MUX2X1 U3825 ( .B(n4118), .A(n4119), .S(n4510), .Y(n4117) );
  MUX2X1 U3826 ( .B(n4121), .A(n4122), .S(n4510), .Y(n4120) );
  MUX2X1 U3827 ( .B(n4124), .A(n4125), .S(n15), .Y(n4123) );
  MUX2X1 U3828 ( .B(n4127), .A(n4128), .S(n4510), .Y(n4126) );
  MUX2X1 U3829 ( .B(n4130), .A(n4131), .S(n4510), .Y(n4129) );
  MUX2X1 U3830 ( .B(n4133), .A(n4134), .S(n4510), .Y(n4132) );
  MUX2X1 U3831 ( .B(n4136), .A(n4137), .S(n4510), .Y(n4135) );
  MUX2X1 U3832 ( .B(n4139), .A(n4140), .S(n15), .Y(n4138) );
  MUX2X1 U3833 ( .B(n4142), .A(n4143), .S(n4511), .Y(n4141) );
  MUX2X1 U3834 ( .B(n4145), .A(n4146), .S(n4511), .Y(n4144) );
  MUX2X1 U3835 ( .B(n4148), .A(n4149), .S(n4511), .Y(n4147) );
  MUX2X1 U3836 ( .B(n4151), .A(n4152), .S(n4511), .Y(n4150) );
  MUX2X1 U3837 ( .B(n4154), .A(n4155), .S(n15), .Y(n4153) );
  MUX2X1 U3838 ( .B(n4157), .A(n4158), .S(n4511), .Y(n4156) );
  MUX2X1 U3839 ( .B(n4160), .A(n4161), .S(n4511), .Y(n4159) );
  MUX2X1 U3840 ( .B(n4163), .A(n4164), .S(n4511), .Y(n4162) );
  MUX2X1 U3841 ( .B(n4166), .A(n4167), .S(n4511), .Y(n4165) );
  MUX2X1 U3842 ( .B(n4169), .A(n4170), .S(n15), .Y(n4168) );
  MUX2X1 U3843 ( .B(n4172), .A(n4173), .S(n4511), .Y(n4171) );
  MUX2X1 U3844 ( .B(n4175), .A(n4176), .S(n4511), .Y(n4174) );
  MUX2X1 U3845 ( .B(n4178), .A(n4179), .S(n4511), .Y(n4177) );
  MUX2X1 U3846 ( .B(n4181), .A(n4182), .S(n4511), .Y(n4180) );
  MUX2X1 U3847 ( .B(n4184), .A(n4185), .S(n15), .Y(n4183) );
  MUX2X1 U3848 ( .B(n4187), .A(n4188), .S(n4512), .Y(n4186) );
  MUX2X1 U3849 ( .B(n4190), .A(n4191), .S(n4512), .Y(n4189) );
  MUX2X1 U3850 ( .B(n4193), .A(n4194), .S(n4512), .Y(n4192) );
  MUX2X1 U3851 ( .B(n4196), .A(n4197), .S(n4512), .Y(n4195) );
  MUX2X1 U3852 ( .B(n4199), .A(n4200), .S(n15), .Y(n4198) );
  MUX2X1 U3853 ( .B(n4202), .A(n4203), .S(n4512), .Y(n4201) );
  MUX2X1 U3854 ( .B(n4205), .A(n4206), .S(n4512), .Y(n4204) );
  MUX2X1 U3855 ( .B(n4208), .A(n4209), .S(n4512), .Y(n4207) );
  MUX2X1 U3856 ( .B(n4211), .A(n4212), .S(n4512), .Y(n4210) );
  MUX2X1 U3857 ( .B(n4214), .A(n4215), .S(n15), .Y(n4213) );
  MUX2X1 U3858 ( .B(n4217), .A(n4218), .S(n4512), .Y(n4216) );
  MUX2X1 U3859 ( .B(n4220), .A(n4221), .S(n4512), .Y(n4219) );
  MUX2X1 U3860 ( .B(n4223), .A(n4224), .S(n4512), .Y(n4222) );
  MUX2X1 U3861 ( .B(n4226), .A(n4227), .S(n4512), .Y(n4225) );
  MUX2X1 U3862 ( .B(n4229), .A(n4230), .S(n15), .Y(n4228) );
  MUX2X1 U3863 ( .B(n4232), .A(n4233), .S(n4513), .Y(n4231) );
  MUX2X1 U3864 ( .B(n4235), .A(n4236), .S(n4513), .Y(n4234) );
  MUX2X1 U3865 ( .B(n4238), .A(n4239), .S(n4513), .Y(n4237) );
  MUX2X1 U3866 ( .B(n4241), .A(n4242), .S(n4513), .Y(n4240) );
  MUX2X1 U3867 ( .B(n4244), .A(n4245), .S(n15), .Y(n4243) );
  MUX2X1 U3868 ( .B(n4247), .A(n4248), .S(n4513), .Y(n4246) );
  MUX2X1 U3869 ( .B(n4250), .A(n4251), .S(n4513), .Y(n4249) );
  MUX2X1 U3870 ( .B(n4253), .A(n4254), .S(n4513), .Y(n4252) );
  MUX2X1 U3871 ( .B(n4256), .A(n4257), .S(n4513), .Y(n4255) );
  MUX2X1 U3872 ( .B(n4259), .A(n4260), .S(n15), .Y(n4258) );
  MUX2X1 U3873 ( .B(n4262), .A(n4263), .S(n4513), .Y(n4261) );
  MUX2X1 U3874 ( .B(n4265), .A(n4266), .S(n4513), .Y(n4264) );
  MUX2X1 U3875 ( .B(n4268), .A(n4269), .S(n4513), .Y(n4267) );
  MUX2X1 U3876 ( .B(n4271), .A(n4272), .S(n4513), .Y(n4270) );
  MUX2X1 U3877 ( .B(n4274), .A(n4275), .S(n15), .Y(n4273) );
  MUX2X1 U3878 ( .B(n4277), .A(n4278), .S(n4512), .Y(n4276) );
  MUX2X1 U3879 ( .B(n4280), .A(n4281), .S(n4503), .Y(n4279) );
  MUX2X1 U3880 ( .B(n4283), .A(n4284), .S(n4497), .Y(n4282) );
  MUX2X1 U3881 ( .B(n4286), .A(n4287), .S(n4496), .Y(n4285) );
  MUX2X1 U3882 ( .B(n4289), .A(n4290), .S(n15), .Y(n4288) );
  MUX2X1 U3883 ( .B(n4292), .A(n4293), .S(n4510), .Y(n4291) );
  MUX2X1 U3884 ( .B(n4295), .A(n4296), .S(n4504), .Y(n4294) );
  MUX2X1 U3885 ( .B(n4298), .A(n4299), .S(n4513), .Y(n4297) );
  MUX2X1 U3886 ( .B(n4301), .A(n4302), .S(n4505), .Y(n4300) );
  MUX2X1 U3887 ( .B(n4304), .A(n4305), .S(n15), .Y(n4303) );
  MUX2X1 U3888 ( .B(n4307), .A(n4308), .S(n4501), .Y(n4306) );
  MUX2X1 U3889 ( .B(n4310), .A(n4311), .S(n4507), .Y(n4309) );
  MUX2X1 U3890 ( .B(n4313), .A(n4314), .S(n4511), .Y(n4312) );
  MUX2X1 U3891 ( .B(n4316), .A(n4317), .S(n4508), .Y(n4315) );
  MUX2X1 U3892 ( .B(n4319), .A(n4320), .S(n15), .Y(n4318) );
  MUX2X1 U3893 ( .B(n4322), .A(n4323), .S(n4500), .Y(n4321) );
  MUX2X1 U3894 ( .B(n4325), .A(n4326), .S(n4512), .Y(n4324) );
  MUX2X1 U3895 ( .B(n4328), .A(n4329), .S(n4498), .Y(n4327) );
  MUX2X1 U3896 ( .B(n4331), .A(n4332), .S(n4510), .Y(n4330) );
  MUX2X1 U3897 ( .B(n4334), .A(n4335), .S(n15), .Y(n4333) );
  MUX2X1 U3898 ( .B(n4337), .A(n4338), .S(n4506), .Y(n4336) );
  MUX2X1 U3899 ( .B(n4340), .A(n4341), .S(n4505), .Y(n4339) );
  MUX2X1 U3900 ( .B(n4343), .A(n4344), .S(n4502), .Y(n4342) );
  MUX2X1 U3901 ( .B(n4346), .A(n4347), .S(n4506), .Y(n4345) );
  MUX2X1 U3902 ( .B(n4349), .A(n4350), .S(n15), .Y(n4348) );
  MUX2X1 U3903 ( .B(n4352), .A(n4353), .S(n4495), .Y(n4351) );
  MUX2X1 U3904 ( .B(n4355), .A(n4356), .S(n4511), .Y(n4354) );
  MUX2X1 U3905 ( .B(n4358), .A(n4359), .S(n4499), .Y(n4357) );
  MUX2X1 U3906 ( .B(n4361), .A(n4362), .S(n4513), .Y(n4360) );
  MUX2X1 U3907 ( .B(n4364), .A(n4365), .S(n15), .Y(n4363) );
  MUX2X1 U3908 ( .B(n4367), .A(n4368), .S(n4498), .Y(n4366) );
  MUX2X1 U3909 ( .B(n4370), .A(n4371), .S(n4507), .Y(n4369) );
  MUX2X1 U3910 ( .B(n4373), .A(n4374), .S(n4500), .Y(n4372) );
  MUX2X1 U3911 ( .B(n4376), .A(n4377), .S(n4496), .Y(n4375) );
  MUX2X1 U3912 ( .B(n4379), .A(n4380), .S(n15), .Y(n4378) );
  MUX2X1 U3913 ( .B(n4382), .A(n4383), .S(n4497), .Y(n4381) );
  MUX2X1 U3914 ( .B(n4385), .A(n4386), .S(n4504), .Y(n4384) );
  MUX2X1 U3915 ( .B(n4388), .A(n4389), .S(n4497), .Y(n4387) );
  MUX2X1 U3916 ( .B(n4391), .A(n4392), .S(n4501), .Y(n4390) );
  MUX2X1 U3917 ( .B(n4394), .A(n4395), .S(n15), .Y(n4393) );
  MUX2X1 U3918 ( .B(n4397), .A(n4398), .S(n4499), .Y(n4396) );
  MUX2X1 U3919 ( .B(n4400), .A(n4401), .S(n4508), .Y(n4399) );
  MUX2X1 U3920 ( .B(n4403), .A(n4404), .S(n4495), .Y(n4402) );
  MUX2X1 U3921 ( .B(n4406), .A(n4407), .S(n4503), .Y(n4405) );
  MUX2X1 U3922 ( .B(n4409), .A(n4410), .S(n15), .Y(n4408) );
  MUX2X1 U3923 ( .B(mem[990]), .A(mem[1023]), .S(n4451), .Y(n3423) );
  MUX2X1 U3924 ( .B(mem[924]), .A(mem[957]), .S(n4451), .Y(n3422) );
  MUX2X1 U3925 ( .B(mem[858]), .A(mem[891]), .S(n4451), .Y(n3426) );
  MUX2X1 U3926 ( .B(mem[792]), .A(mem[825]), .S(n4451), .Y(n3425) );
  MUX2X1 U3927 ( .B(n3424), .A(n3421), .S(n4515), .Y(n3435) );
  MUX2X1 U3928 ( .B(mem[726]), .A(mem[759]), .S(n4451), .Y(n3429) );
  MUX2X1 U3929 ( .B(mem[660]), .A(mem[693]), .S(n4451), .Y(n3428) );
  MUX2X1 U3930 ( .B(mem[594]), .A(mem[627]), .S(n4451), .Y(n3432) );
  MUX2X1 U3931 ( .B(mem[528]), .A(mem[561]), .S(n4451), .Y(n3431) );
  MUX2X1 U3932 ( .B(n3430), .A(n3427), .S(n4515), .Y(n3434) );
  MUX2X1 U3933 ( .B(mem[462]), .A(mem[495]), .S(n4451), .Y(n3438) );
  MUX2X1 U3934 ( .B(mem[396]), .A(mem[429]), .S(n4451), .Y(n3437) );
  MUX2X1 U3935 ( .B(mem[330]), .A(mem[363]), .S(n4451), .Y(n3441) );
  MUX2X1 U3936 ( .B(mem[264]), .A(mem[297]), .S(n4451), .Y(n3440) );
  MUX2X1 U3937 ( .B(n3439), .A(n3436), .S(n4515), .Y(n3450) );
  MUX2X1 U3938 ( .B(mem[198]), .A(mem[231]), .S(n4452), .Y(n3444) );
  MUX2X1 U3939 ( .B(mem[132]), .A(mem[165]), .S(n4452), .Y(n3443) );
  MUX2X1 U3940 ( .B(mem[66]), .A(mem[99]), .S(n4452), .Y(n3447) );
  MUX2X1 U3941 ( .B(mem[0]), .A(mem[33]), .S(n4452), .Y(n3446) );
  MUX2X1 U3942 ( .B(n3445), .A(n3442), .S(n4515), .Y(n3449) );
  MUX2X1 U3943 ( .B(n3448), .A(n3433), .S(n16), .Y(n4411) );
  MUX2X1 U3944 ( .B(mem[991]), .A(mem[1024]), .S(n4452), .Y(n3453) );
  MUX2X1 U3945 ( .B(mem[925]), .A(mem[958]), .S(n4452), .Y(n3452) );
  MUX2X1 U3946 ( .B(mem[859]), .A(mem[892]), .S(n4452), .Y(n3456) );
  MUX2X1 U3947 ( .B(mem[793]), .A(mem[826]), .S(n4452), .Y(n3455) );
  MUX2X1 U3948 ( .B(n3454), .A(n3451), .S(n4515), .Y(n3465) );
  MUX2X1 U3949 ( .B(mem[727]), .A(mem[760]), .S(n4452), .Y(n3459) );
  MUX2X1 U3950 ( .B(mem[661]), .A(mem[694]), .S(n4452), .Y(n3458) );
  MUX2X1 U3951 ( .B(mem[595]), .A(mem[628]), .S(n4452), .Y(n3462) );
  MUX2X1 U3952 ( .B(mem[529]), .A(mem[562]), .S(n4452), .Y(n3461) );
  MUX2X1 U3953 ( .B(n3460), .A(n3457), .S(n4515), .Y(n3464) );
  MUX2X1 U3954 ( .B(mem[463]), .A(mem[496]), .S(n4453), .Y(n3468) );
  MUX2X1 U3955 ( .B(mem[397]), .A(mem[430]), .S(n4453), .Y(n3467) );
  MUX2X1 U3956 ( .B(mem[331]), .A(mem[364]), .S(n4453), .Y(n3471) );
  MUX2X1 U3957 ( .B(mem[265]), .A(mem[298]), .S(n4453), .Y(n3470) );
  MUX2X1 U3958 ( .B(n3469), .A(n3466), .S(n4515), .Y(n3480) );
  MUX2X1 U3959 ( .B(mem[199]), .A(mem[232]), .S(n4453), .Y(n3474) );
  MUX2X1 U3960 ( .B(mem[133]), .A(mem[166]), .S(n4453), .Y(n3473) );
  MUX2X1 U3961 ( .B(mem[67]), .A(mem[100]), .S(n4453), .Y(n3477) );
  MUX2X1 U3962 ( .B(mem[1]), .A(mem[34]), .S(n4453), .Y(n3476) );
  MUX2X1 U3963 ( .B(n3475), .A(n3472), .S(n4515), .Y(n3479) );
  MUX2X1 U3964 ( .B(n3478), .A(n3463), .S(n16), .Y(n4412) );
  MUX2X1 U3965 ( .B(mem[992]), .A(mem[1025]), .S(n4453), .Y(n3483) );
  MUX2X1 U3966 ( .B(mem[926]), .A(mem[959]), .S(n4453), .Y(n3482) );
  MUX2X1 U3967 ( .B(mem[860]), .A(mem[893]), .S(n4453), .Y(n3486) );
  MUX2X1 U3968 ( .B(mem[794]), .A(mem[827]), .S(n4453), .Y(n3485) );
  MUX2X1 U3969 ( .B(n3484), .A(n3481), .S(n4515), .Y(n3495) );
  MUX2X1 U3970 ( .B(mem[728]), .A(mem[761]), .S(n4454), .Y(n3489) );
  MUX2X1 U3971 ( .B(mem[662]), .A(mem[695]), .S(n4454), .Y(n3488) );
  MUX2X1 U3972 ( .B(mem[596]), .A(mem[629]), .S(n4454), .Y(n3492) );
  MUX2X1 U3973 ( .B(mem[530]), .A(mem[563]), .S(n4454), .Y(n3491) );
  MUX2X1 U3974 ( .B(n3490), .A(n3487), .S(n4515), .Y(n3494) );
  MUX2X1 U3975 ( .B(mem[464]), .A(mem[497]), .S(n4454), .Y(n3498) );
  MUX2X1 U3976 ( .B(mem[398]), .A(mem[431]), .S(n4454), .Y(n3497) );
  MUX2X1 U3977 ( .B(mem[332]), .A(mem[365]), .S(n4454), .Y(n3501) );
  MUX2X1 U3978 ( .B(mem[266]), .A(mem[299]), .S(n4454), .Y(n3500) );
  MUX2X1 U3979 ( .B(n3499), .A(n3496), .S(n4515), .Y(n3510) );
  MUX2X1 U3980 ( .B(mem[200]), .A(mem[233]), .S(n4454), .Y(n3504) );
  MUX2X1 U3981 ( .B(mem[134]), .A(mem[167]), .S(n4454), .Y(n3503) );
  MUX2X1 U3982 ( .B(mem[68]), .A(mem[101]), .S(n4454), .Y(n3507) );
  MUX2X1 U3983 ( .B(mem[2]), .A(mem[35]), .S(n4454), .Y(n3506) );
  MUX2X1 U3984 ( .B(n3505), .A(n3502), .S(n4515), .Y(n3509) );
  MUX2X1 U3985 ( .B(n3508), .A(n3493), .S(n16), .Y(n4413) );
  MUX2X1 U3986 ( .B(mem[993]), .A(mem[1026]), .S(n4455), .Y(n3513) );
  MUX2X1 U3987 ( .B(mem[927]), .A(mem[960]), .S(n4455), .Y(n3512) );
  MUX2X1 U3988 ( .B(mem[861]), .A(mem[894]), .S(n4455), .Y(n3516) );
  MUX2X1 U3989 ( .B(mem[795]), .A(mem[828]), .S(n4455), .Y(n3515) );
  MUX2X1 U3990 ( .B(n3514), .A(n3511), .S(n4516), .Y(n3525) );
  MUX2X1 U3991 ( .B(mem[729]), .A(mem[762]), .S(n4455), .Y(n3519) );
  MUX2X1 U3992 ( .B(mem[663]), .A(mem[696]), .S(n4455), .Y(n3518) );
  MUX2X1 U3993 ( .B(mem[597]), .A(mem[630]), .S(n4455), .Y(n3522) );
  MUX2X1 U3994 ( .B(mem[531]), .A(mem[564]), .S(n4455), .Y(n3521) );
  MUX2X1 U3995 ( .B(n3520), .A(n3517), .S(n4516), .Y(n3524) );
  MUX2X1 U3996 ( .B(mem[465]), .A(mem[498]), .S(n4455), .Y(n3528) );
  MUX2X1 U3997 ( .B(mem[399]), .A(mem[432]), .S(n4455), .Y(n3527) );
  MUX2X1 U3998 ( .B(mem[333]), .A(mem[366]), .S(n4455), .Y(n3531) );
  MUX2X1 U3999 ( .B(mem[267]), .A(mem[300]), .S(n4455), .Y(n3530) );
  MUX2X1 U4000 ( .B(n3529), .A(n3526), .S(n4516), .Y(n3540) );
  MUX2X1 U4001 ( .B(mem[201]), .A(mem[234]), .S(n4456), .Y(n3534) );
  MUX2X1 U4002 ( .B(mem[135]), .A(mem[168]), .S(n4456), .Y(n3533) );
  MUX2X1 U4003 ( .B(mem[69]), .A(mem[102]), .S(n4456), .Y(n3537) );
  MUX2X1 U4004 ( .B(mem[3]), .A(mem[36]), .S(n4456), .Y(n3536) );
  MUX2X1 U4005 ( .B(n3535), .A(n3532), .S(n4516), .Y(n3539) );
  MUX2X1 U4006 ( .B(n3538), .A(n3523), .S(n16), .Y(n4414) );
  MUX2X1 U4007 ( .B(mem[994]), .A(mem[1027]), .S(n4456), .Y(n3543) );
  MUX2X1 U4008 ( .B(mem[928]), .A(mem[961]), .S(n4456), .Y(n3542) );
  MUX2X1 U4009 ( .B(mem[862]), .A(mem[895]), .S(n4456), .Y(n3546) );
  MUX2X1 U4010 ( .B(mem[796]), .A(mem[829]), .S(n4456), .Y(n3545) );
  MUX2X1 U4011 ( .B(n3544), .A(n3541), .S(n4516), .Y(n3555) );
  MUX2X1 U4012 ( .B(mem[730]), .A(mem[763]), .S(n4456), .Y(n3549) );
  MUX2X1 U4013 ( .B(mem[664]), .A(mem[697]), .S(n4456), .Y(n3548) );
  MUX2X1 U4014 ( .B(mem[598]), .A(mem[631]), .S(n4456), .Y(n3552) );
  MUX2X1 U4015 ( .B(mem[532]), .A(mem[565]), .S(n4456), .Y(n3551) );
  MUX2X1 U4016 ( .B(n3550), .A(n3547), .S(n4516), .Y(n3554) );
  MUX2X1 U4017 ( .B(mem[466]), .A(mem[499]), .S(n4457), .Y(n3558) );
  MUX2X1 U4018 ( .B(mem[400]), .A(mem[433]), .S(n4457), .Y(n3557) );
  MUX2X1 U4019 ( .B(mem[334]), .A(mem[367]), .S(n4457), .Y(n3561) );
  MUX2X1 U4020 ( .B(mem[268]), .A(mem[301]), .S(n4457), .Y(n3560) );
  MUX2X1 U4021 ( .B(n3559), .A(n3556), .S(n4516), .Y(n3570) );
  MUX2X1 U4022 ( .B(mem[202]), .A(mem[235]), .S(n4457), .Y(n3564) );
  MUX2X1 U4023 ( .B(mem[136]), .A(mem[169]), .S(n4457), .Y(n3563) );
  MUX2X1 U4024 ( .B(mem[70]), .A(mem[103]), .S(n4457), .Y(n3567) );
  MUX2X1 U4025 ( .B(mem[4]), .A(mem[37]), .S(n4457), .Y(n3566) );
  MUX2X1 U4026 ( .B(n3565), .A(n3562), .S(n4516), .Y(n3569) );
  MUX2X1 U4027 ( .B(n3568), .A(n3553), .S(n16), .Y(n4415) );
  MUX2X1 U4028 ( .B(mem[995]), .A(mem[1028]), .S(n4457), .Y(n3573) );
  MUX2X1 U4029 ( .B(mem[929]), .A(mem[962]), .S(n4457), .Y(n3572) );
  MUX2X1 U4030 ( .B(mem[863]), .A(mem[896]), .S(n4457), .Y(n3576) );
  MUX2X1 U4031 ( .B(mem[797]), .A(mem[830]), .S(n4457), .Y(n3575) );
  MUX2X1 U4032 ( .B(n3574), .A(n3571), .S(n4516), .Y(n3585) );
  MUX2X1 U4033 ( .B(mem[731]), .A(mem[764]), .S(n4458), .Y(n3579) );
  MUX2X1 U4034 ( .B(mem[665]), .A(mem[698]), .S(n4458), .Y(n3578) );
  MUX2X1 U4035 ( .B(mem[599]), .A(mem[632]), .S(n4458), .Y(n3582) );
  MUX2X1 U4036 ( .B(mem[533]), .A(mem[566]), .S(n4458), .Y(n3581) );
  MUX2X1 U4037 ( .B(n3580), .A(n3577), .S(n4516), .Y(n3584) );
  MUX2X1 U4038 ( .B(mem[467]), .A(mem[500]), .S(n4458), .Y(n3588) );
  MUX2X1 U4039 ( .B(mem[401]), .A(mem[434]), .S(n4458), .Y(n3587) );
  MUX2X1 U4040 ( .B(mem[335]), .A(mem[368]), .S(n4458), .Y(n3591) );
  MUX2X1 U4041 ( .B(mem[269]), .A(mem[302]), .S(n4458), .Y(n3590) );
  MUX2X1 U4042 ( .B(n3589), .A(n3586), .S(n4516), .Y(n3600) );
  MUX2X1 U4043 ( .B(mem[203]), .A(mem[236]), .S(n4458), .Y(n3594) );
  MUX2X1 U4044 ( .B(mem[137]), .A(mem[170]), .S(n4458), .Y(n3593) );
  MUX2X1 U4045 ( .B(mem[71]), .A(mem[104]), .S(n4458), .Y(n3597) );
  MUX2X1 U4046 ( .B(mem[5]), .A(mem[38]), .S(n4458), .Y(n3596) );
  MUX2X1 U4047 ( .B(n3595), .A(n3592), .S(n4516), .Y(n3599) );
  MUX2X1 U4048 ( .B(n3598), .A(n3583), .S(n16), .Y(n4416) );
  MUX2X1 U4049 ( .B(mem[996]), .A(mem[1029]), .S(n4459), .Y(n3603) );
  MUX2X1 U4050 ( .B(mem[930]), .A(mem[963]), .S(n4459), .Y(n3602) );
  MUX2X1 U4051 ( .B(mem[864]), .A(mem[897]), .S(n4459), .Y(n3606) );
  MUX2X1 U4052 ( .B(mem[798]), .A(mem[831]), .S(n4459), .Y(n3605) );
  MUX2X1 U4053 ( .B(n3604), .A(n3601), .S(n14), .Y(n3615) );
  MUX2X1 U4054 ( .B(mem[732]), .A(mem[765]), .S(n4459), .Y(n3609) );
  MUX2X1 U4055 ( .B(mem[666]), .A(mem[699]), .S(n4459), .Y(n3608) );
  MUX2X1 U4056 ( .B(mem[600]), .A(mem[633]), .S(n4459), .Y(n3612) );
  MUX2X1 U4057 ( .B(mem[534]), .A(mem[567]), .S(n4459), .Y(n3611) );
  MUX2X1 U4058 ( .B(n3610), .A(n3607), .S(n14), .Y(n3614) );
  MUX2X1 U4059 ( .B(mem[468]), .A(mem[501]), .S(n4459), .Y(n3618) );
  MUX2X1 U4060 ( .B(mem[402]), .A(mem[435]), .S(n4459), .Y(n3617) );
  MUX2X1 U4061 ( .B(mem[336]), .A(mem[369]), .S(n4459), .Y(n3621) );
  MUX2X1 U4062 ( .B(mem[270]), .A(mem[303]), .S(n4459), .Y(n3620) );
  MUX2X1 U4063 ( .B(n3619), .A(n3616), .S(n14), .Y(n3630) );
  MUX2X1 U4064 ( .B(mem[204]), .A(mem[237]), .S(n4460), .Y(n3624) );
  MUX2X1 U4065 ( .B(mem[138]), .A(mem[171]), .S(n4460), .Y(n3623) );
  MUX2X1 U4066 ( .B(mem[72]), .A(mem[105]), .S(n4460), .Y(n3627) );
  MUX2X1 U4067 ( .B(mem[6]), .A(mem[39]), .S(n4460), .Y(n3626) );
  MUX2X1 U4068 ( .B(n3625), .A(n3622), .S(n14), .Y(n3629) );
  MUX2X1 U4069 ( .B(n3628), .A(n3613), .S(n16), .Y(n4417) );
  MUX2X1 U4070 ( .B(mem[997]), .A(mem[1030]), .S(n4460), .Y(n3633) );
  MUX2X1 U4071 ( .B(mem[931]), .A(mem[964]), .S(n4460), .Y(n3632) );
  MUX2X1 U4072 ( .B(mem[865]), .A(mem[898]), .S(n4460), .Y(n3636) );
  MUX2X1 U4073 ( .B(mem[799]), .A(mem[832]), .S(n4460), .Y(n3635) );
  MUX2X1 U4074 ( .B(n3634), .A(n3631), .S(n14), .Y(n3645) );
  MUX2X1 U4075 ( .B(mem[733]), .A(mem[766]), .S(n4460), .Y(n3639) );
  MUX2X1 U4076 ( .B(mem[667]), .A(mem[700]), .S(n4460), .Y(n3638) );
  MUX2X1 U4077 ( .B(mem[601]), .A(mem[634]), .S(n4460), .Y(n3642) );
  MUX2X1 U4078 ( .B(mem[535]), .A(mem[568]), .S(n4460), .Y(n3641) );
  MUX2X1 U4079 ( .B(n3640), .A(n3637), .S(n14), .Y(n3644) );
  MUX2X1 U4080 ( .B(mem[469]), .A(mem[502]), .S(n4461), .Y(n3648) );
  MUX2X1 U4081 ( .B(mem[403]), .A(mem[436]), .S(n4461), .Y(n3647) );
  MUX2X1 U4082 ( .B(mem[337]), .A(mem[370]), .S(n4461), .Y(n3651) );
  MUX2X1 U4083 ( .B(mem[271]), .A(mem[304]), .S(n4461), .Y(n3650) );
  MUX2X1 U4084 ( .B(n3649), .A(n3646), .S(n14), .Y(n3660) );
  MUX2X1 U4085 ( .B(mem[205]), .A(mem[238]), .S(n4461), .Y(n3654) );
  MUX2X1 U4086 ( .B(mem[139]), .A(mem[172]), .S(n4461), .Y(n3653) );
  MUX2X1 U4087 ( .B(mem[73]), .A(mem[106]), .S(n4461), .Y(n3657) );
  MUX2X1 U4088 ( .B(mem[7]), .A(mem[40]), .S(n4461), .Y(n3656) );
  MUX2X1 U4089 ( .B(n3655), .A(n3652), .S(n14), .Y(n3659) );
  MUX2X1 U4090 ( .B(n3658), .A(n3643), .S(n16), .Y(n4418) );
  MUX2X1 U4091 ( .B(mem[998]), .A(mem[1031]), .S(n4461), .Y(n3663) );
  MUX2X1 U4092 ( .B(mem[932]), .A(mem[965]), .S(n4461), .Y(n3662) );
  MUX2X1 U4093 ( .B(mem[866]), .A(mem[899]), .S(n4461), .Y(n3666) );
  MUX2X1 U4094 ( .B(mem[800]), .A(mem[833]), .S(n4461), .Y(n3665) );
  MUX2X1 U4095 ( .B(n3664), .A(n3661), .S(n14), .Y(n3675) );
  MUX2X1 U4096 ( .B(mem[734]), .A(mem[767]), .S(n4462), .Y(n3669) );
  MUX2X1 U4097 ( .B(mem[668]), .A(mem[701]), .S(n4462), .Y(n3668) );
  MUX2X1 U4098 ( .B(mem[602]), .A(mem[635]), .S(n4462), .Y(n3672) );
  MUX2X1 U4099 ( .B(mem[536]), .A(mem[569]), .S(n4462), .Y(n3671) );
  MUX2X1 U4100 ( .B(n3670), .A(n3667), .S(n14), .Y(n3674) );
  MUX2X1 U4101 ( .B(mem[470]), .A(mem[503]), .S(n4462), .Y(n3678) );
  MUX2X1 U4102 ( .B(mem[404]), .A(mem[437]), .S(n4462), .Y(n3677) );
  MUX2X1 U4103 ( .B(mem[338]), .A(mem[371]), .S(n4462), .Y(n3681) );
  MUX2X1 U4104 ( .B(mem[272]), .A(mem[305]), .S(n4462), .Y(n3680) );
  MUX2X1 U4105 ( .B(n3679), .A(n3676), .S(n14), .Y(n3690) );
  MUX2X1 U4106 ( .B(mem[206]), .A(mem[239]), .S(n4462), .Y(n3684) );
  MUX2X1 U4107 ( .B(mem[140]), .A(mem[173]), .S(n4462), .Y(n3683) );
  MUX2X1 U4108 ( .B(mem[74]), .A(mem[107]), .S(n4462), .Y(n3687) );
  MUX2X1 U4109 ( .B(mem[8]), .A(mem[41]), .S(n4462), .Y(n3686) );
  MUX2X1 U4110 ( .B(n3685), .A(n3682), .S(n14), .Y(n3689) );
  MUX2X1 U4111 ( .B(n3688), .A(n3673), .S(n16), .Y(n4419) );
  MUX2X1 U4112 ( .B(mem[999]), .A(mem[1032]), .S(n4463), .Y(n3693) );
  MUX2X1 U4113 ( .B(mem[933]), .A(mem[966]), .S(n4463), .Y(n3692) );
  MUX2X1 U4114 ( .B(mem[867]), .A(mem[900]), .S(n4463), .Y(n3696) );
  MUX2X1 U4115 ( .B(mem[801]), .A(mem[834]), .S(n4463), .Y(n3695) );
  MUX2X1 U4116 ( .B(n3694), .A(n3691), .S(n14), .Y(n3705) );
  MUX2X1 U4117 ( .B(mem[735]), .A(mem[768]), .S(n4463), .Y(n3699) );
  MUX2X1 U4118 ( .B(mem[669]), .A(mem[702]), .S(n4463), .Y(n3698) );
  MUX2X1 U4119 ( .B(mem[603]), .A(mem[636]), .S(n4463), .Y(n3702) );
  MUX2X1 U4120 ( .B(mem[537]), .A(mem[570]), .S(n4463), .Y(n3701) );
  MUX2X1 U4121 ( .B(n3700), .A(n3697), .S(n14), .Y(n3704) );
  MUX2X1 U4122 ( .B(mem[471]), .A(mem[504]), .S(n4463), .Y(n3708) );
  MUX2X1 U4123 ( .B(mem[405]), .A(mem[438]), .S(n4463), .Y(n3707) );
  MUX2X1 U4124 ( .B(mem[339]), .A(mem[372]), .S(n4463), .Y(n3711) );
  MUX2X1 U4125 ( .B(mem[273]), .A(mem[306]), .S(n4463), .Y(n3710) );
  MUX2X1 U4126 ( .B(n3709), .A(n3706), .S(n14), .Y(n3720) );
  MUX2X1 U4127 ( .B(mem[207]), .A(mem[240]), .S(n4464), .Y(n3714) );
  MUX2X1 U4128 ( .B(mem[141]), .A(mem[174]), .S(n4464), .Y(n3713) );
  MUX2X1 U4129 ( .B(mem[75]), .A(mem[108]), .S(n4464), .Y(n3717) );
  MUX2X1 U4130 ( .B(mem[9]), .A(mem[42]), .S(n4464), .Y(n3716) );
  MUX2X1 U4131 ( .B(n3715), .A(n3712), .S(n14), .Y(n3719) );
  MUX2X1 U4132 ( .B(n3718), .A(n3703), .S(n16), .Y(n4420) );
  MUX2X1 U4133 ( .B(mem[1000]), .A(mem[1033]), .S(n4464), .Y(n3723) );
  MUX2X1 U4134 ( .B(mem[934]), .A(mem[967]), .S(n4464), .Y(n3722) );
  MUX2X1 U4135 ( .B(mem[868]), .A(mem[901]), .S(n4464), .Y(n3726) );
  MUX2X1 U4136 ( .B(mem[802]), .A(mem[835]), .S(n4464), .Y(n3725) );
  MUX2X1 U4137 ( .B(n3724), .A(n3721), .S(n14), .Y(n3735) );
  MUX2X1 U4138 ( .B(mem[736]), .A(mem[769]), .S(n4464), .Y(n3729) );
  MUX2X1 U4139 ( .B(mem[670]), .A(mem[703]), .S(n4464), .Y(n3728) );
  MUX2X1 U4140 ( .B(mem[604]), .A(mem[637]), .S(n4464), .Y(n3732) );
  MUX2X1 U4141 ( .B(mem[538]), .A(mem[571]), .S(n4464), .Y(n3731) );
  MUX2X1 U4142 ( .B(n3730), .A(n3727), .S(n14), .Y(n3734) );
  MUX2X1 U4143 ( .B(mem[472]), .A(mem[505]), .S(n4465), .Y(n3738) );
  MUX2X1 U4144 ( .B(mem[406]), .A(mem[439]), .S(n4465), .Y(n3737) );
  MUX2X1 U4145 ( .B(mem[340]), .A(mem[373]), .S(n4465), .Y(n3741) );
  MUX2X1 U4146 ( .B(mem[274]), .A(mem[307]), .S(n4465), .Y(n3740) );
  MUX2X1 U4147 ( .B(n3739), .A(n3736), .S(n14), .Y(n3750) );
  MUX2X1 U4148 ( .B(mem[208]), .A(mem[241]), .S(n4465), .Y(n3744) );
  MUX2X1 U4149 ( .B(mem[142]), .A(mem[175]), .S(n4465), .Y(n3743) );
  MUX2X1 U4150 ( .B(mem[76]), .A(mem[109]), .S(n4465), .Y(n3747) );
  MUX2X1 U4151 ( .B(mem[10]), .A(mem[43]), .S(n4465), .Y(n3746) );
  MUX2X1 U4152 ( .B(n3745), .A(n3742), .S(n14), .Y(n3749) );
  MUX2X1 U4153 ( .B(n3748), .A(n3733), .S(n16), .Y(n4421) );
  MUX2X1 U4154 ( .B(mem[1001]), .A(mem[1034]), .S(n4465), .Y(n3753) );
  MUX2X1 U4155 ( .B(mem[935]), .A(mem[968]), .S(n4465), .Y(n3752) );
  MUX2X1 U4156 ( .B(mem[869]), .A(mem[902]), .S(n4465), .Y(n3756) );
  MUX2X1 U4157 ( .B(mem[803]), .A(mem[836]), .S(n4465), .Y(n3755) );
  MUX2X1 U4158 ( .B(n3754), .A(n3751), .S(n14), .Y(n3765) );
  MUX2X1 U4159 ( .B(mem[737]), .A(mem[770]), .S(n4466), .Y(n3759) );
  MUX2X1 U4160 ( .B(mem[671]), .A(mem[704]), .S(n4466), .Y(n3758) );
  MUX2X1 U4161 ( .B(mem[605]), .A(mem[638]), .S(n4466), .Y(n3762) );
  MUX2X1 U4162 ( .B(mem[539]), .A(mem[572]), .S(n4466), .Y(n3761) );
  MUX2X1 U4163 ( .B(n3760), .A(n3757), .S(n14), .Y(n3764) );
  MUX2X1 U4164 ( .B(mem[473]), .A(mem[506]), .S(n4466), .Y(n3768) );
  MUX2X1 U4165 ( .B(mem[407]), .A(mem[440]), .S(n4466), .Y(n3767) );
  MUX2X1 U4166 ( .B(mem[341]), .A(mem[374]), .S(n4466), .Y(n3771) );
  MUX2X1 U4167 ( .B(mem[275]), .A(mem[308]), .S(n4466), .Y(n3770) );
  MUX2X1 U4168 ( .B(n3769), .A(n3766), .S(n14), .Y(n3780) );
  MUX2X1 U4169 ( .B(mem[209]), .A(mem[242]), .S(n4466), .Y(n3774) );
  MUX2X1 U4170 ( .B(mem[143]), .A(mem[176]), .S(n4466), .Y(n3773) );
  MUX2X1 U4171 ( .B(mem[77]), .A(mem[110]), .S(n4466), .Y(n3777) );
  MUX2X1 U4172 ( .B(mem[11]), .A(mem[44]), .S(n4466), .Y(n3776) );
  MUX2X1 U4173 ( .B(n3775), .A(n3772), .S(n14), .Y(n3779) );
  MUX2X1 U4174 ( .B(n3778), .A(n3763), .S(n16), .Y(n4422) );
  MUX2X1 U4175 ( .B(mem[1002]), .A(mem[1035]), .S(n4467), .Y(n3783) );
  MUX2X1 U4176 ( .B(mem[936]), .A(mem[969]), .S(n4467), .Y(n3782) );
  MUX2X1 U4177 ( .B(mem[870]), .A(mem[903]), .S(n4467), .Y(n3786) );
  MUX2X1 U4178 ( .B(mem[804]), .A(mem[837]), .S(n4467), .Y(n3785) );
  MUX2X1 U4179 ( .B(n3784), .A(n3781), .S(n14), .Y(n3795) );
  MUX2X1 U4180 ( .B(mem[738]), .A(mem[771]), .S(n4467), .Y(n3789) );
  MUX2X1 U4181 ( .B(mem[672]), .A(mem[705]), .S(n4467), .Y(n3788) );
  MUX2X1 U4182 ( .B(mem[606]), .A(mem[639]), .S(n4467), .Y(n3792) );
  MUX2X1 U4183 ( .B(mem[540]), .A(mem[573]), .S(n4467), .Y(n3791) );
  MUX2X1 U4184 ( .B(n3790), .A(n3787), .S(n14), .Y(n3794) );
  MUX2X1 U4185 ( .B(mem[474]), .A(mem[507]), .S(n4467), .Y(n3798) );
  MUX2X1 U4186 ( .B(mem[408]), .A(mem[441]), .S(n4467), .Y(n3797) );
  MUX2X1 U4187 ( .B(mem[342]), .A(mem[375]), .S(n4467), .Y(n3801) );
  MUX2X1 U4188 ( .B(mem[276]), .A(mem[309]), .S(n4467), .Y(n3800) );
  MUX2X1 U4189 ( .B(n3799), .A(n3796), .S(n14), .Y(n3810) );
  MUX2X1 U4190 ( .B(mem[210]), .A(mem[243]), .S(n4468), .Y(n3804) );
  MUX2X1 U4191 ( .B(mem[144]), .A(mem[177]), .S(n4468), .Y(n3803) );
  MUX2X1 U4192 ( .B(mem[78]), .A(mem[111]), .S(n4468), .Y(n3807) );
  MUX2X1 U4193 ( .B(mem[12]), .A(mem[45]), .S(n4468), .Y(n3806) );
  MUX2X1 U4194 ( .B(n3805), .A(n3802), .S(n14), .Y(n3809) );
  MUX2X1 U4195 ( .B(n3808), .A(n3793), .S(n16), .Y(n4423) );
  MUX2X1 U4196 ( .B(mem[1003]), .A(mem[1036]), .S(n4468), .Y(n3813) );
  MUX2X1 U4197 ( .B(mem[937]), .A(mem[970]), .S(n4468), .Y(n3812) );
  MUX2X1 U4198 ( .B(mem[871]), .A(mem[904]), .S(n4468), .Y(n3816) );
  MUX2X1 U4199 ( .B(mem[805]), .A(mem[838]), .S(n4468), .Y(n3815) );
  MUX2X1 U4200 ( .B(n3814), .A(n3811), .S(n14), .Y(n3825) );
  MUX2X1 U4201 ( .B(mem[739]), .A(mem[772]), .S(n4468), .Y(n3819) );
  MUX2X1 U4202 ( .B(mem[673]), .A(mem[706]), .S(n4468), .Y(n3818) );
  MUX2X1 U4203 ( .B(mem[607]), .A(mem[640]), .S(n4468), .Y(n3822) );
  MUX2X1 U4204 ( .B(mem[541]), .A(mem[574]), .S(n4468), .Y(n3821) );
  MUX2X1 U4205 ( .B(n3820), .A(n3817), .S(n14), .Y(n3824) );
  MUX2X1 U4206 ( .B(mem[475]), .A(mem[508]), .S(n4469), .Y(n3828) );
  MUX2X1 U4207 ( .B(mem[409]), .A(mem[442]), .S(n4469), .Y(n3827) );
  MUX2X1 U4208 ( .B(mem[343]), .A(mem[376]), .S(n4469), .Y(n3831) );
  MUX2X1 U4209 ( .B(mem[277]), .A(mem[310]), .S(n4469), .Y(n3830) );
  MUX2X1 U4210 ( .B(n3829), .A(n3826), .S(n14), .Y(n3840) );
  MUX2X1 U4211 ( .B(mem[211]), .A(mem[244]), .S(n4469), .Y(n3834) );
  MUX2X1 U4212 ( .B(mem[145]), .A(mem[178]), .S(n4469), .Y(n3833) );
  MUX2X1 U4213 ( .B(mem[79]), .A(mem[112]), .S(n4469), .Y(n3837) );
  MUX2X1 U4214 ( .B(mem[13]), .A(mem[46]), .S(n4469), .Y(n3836) );
  MUX2X1 U4215 ( .B(n3835), .A(n3832), .S(n14), .Y(n3839) );
  MUX2X1 U4216 ( .B(n3838), .A(n3823), .S(n16), .Y(n4424) );
  MUX2X1 U4217 ( .B(mem[1004]), .A(mem[1037]), .S(n4469), .Y(n3843) );
  MUX2X1 U4218 ( .B(mem[938]), .A(mem[971]), .S(n4469), .Y(n3842) );
  MUX2X1 U4219 ( .B(mem[872]), .A(mem[905]), .S(n4469), .Y(n3846) );
  MUX2X1 U4220 ( .B(mem[806]), .A(mem[839]), .S(n4469), .Y(n3845) );
  MUX2X1 U4221 ( .B(n3844), .A(n3841), .S(n14), .Y(n3855) );
  MUX2X1 U4222 ( .B(mem[740]), .A(mem[773]), .S(n4470), .Y(n3849) );
  MUX2X1 U4223 ( .B(mem[674]), .A(mem[707]), .S(n4470), .Y(n3848) );
  MUX2X1 U4224 ( .B(mem[608]), .A(mem[641]), .S(n4470), .Y(n3852) );
  MUX2X1 U4225 ( .B(mem[542]), .A(mem[575]), .S(n4470), .Y(n3851) );
  MUX2X1 U4226 ( .B(n3850), .A(n3847), .S(n14), .Y(n3854) );
  MUX2X1 U4227 ( .B(mem[476]), .A(mem[509]), .S(n4470), .Y(n3858) );
  MUX2X1 U4228 ( .B(mem[410]), .A(mem[443]), .S(n4470), .Y(n3857) );
  MUX2X1 U4229 ( .B(mem[344]), .A(mem[377]), .S(n4470), .Y(n3861) );
  MUX2X1 U4230 ( .B(mem[278]), .A(mem[311]), .S(n4470), .Y(n3860) );
  MUX2X1 U4231 ( .B(n3859), .A(n3856), .S(n14), .Y(n3870) );
  MUX2X1 U4232 ( .B(mem[212]), .A(mem[245]), .S(n4470), .Y(n3864) );
  MUX2X1 U4233 ( .B(mem[146]), .A(mem[179]), .S(n4470), .Y(n3863) );
  MUX2X1 U4234 ( .B(mem[80]), .A(mem[113]), .S(n4470), .Y(n3867) );
  MUX2X1 U4235 ( .B(mem[14]), .A(mem[47]), .S(n4470), .Y(n3866) );
  MUX2X1 U4236 ( .B(n3865), .A(n3862), .S(n14), .Y(n3869) );
  MUX2X1 U4237 ( .B(n3868), .A(n3853), .S(n16), .Y(n4425) );
  MUX2X1 U4238 ( .B(mem[1005]), .A(mem[1038]), .S(n4471), .Y(n3873) );
  MUX2X1 U4239 ( .B(mem[939]), .A(mem[972]), .S(n4471), .Y(n3872) );
  MUX2X1 U4240 ( .B(mem[873]), .A(mem[906]), .S(n4471), .Y(n3876) );
  MUX2X1 U4241 ( .B(mem[807]), .A(mem[840]), .S(n4471), .Y(n3875) );
  MUX2X1 U4242 ( .B(n3874), .A(n3871), .S(n14), .Y(n3885) );
  MUX2X1 U4243 ( .B(mem[741]), .A(mem[774]), .S(n4471), .Y(n3879) );
  MUX2X1 U4244 ( .B(mem[675]), .A(mem[708]), .S(n4471), .Y(n3878) );
  MUX2X1 U4245 ( .B(mem[609]), .A(mem[642]), .S(n4471), .Y(n3882) );
  MUX2X1 U4246 ( .B(mem[543]), .A(mem[576]), .S(n4471), .Y(n3881) );
  MUX2X1 U4247 ( .B(n3880), .A(n3877), .S(n14), .Y(n3884) );
  MUX2X1 U4248 ( .B(mem[477]), .A(mem[510]), .S(n4471), .Y(n3888) );
  MUX2X1 U4249 ( .B(mem[411]), .A(mem[444]), .S(n4471), .Y(n3887) );
  MUX2X1 U4250 ( .B(mem[345]), .A(mem[378]), .S(n4471), .Y(n3891) );
  MUX2X1 U4251 ( .B(mem[279]), .A(mem[312]), .S(n4471), .Y(n3890) );
  MUX2X1 U4252 ( .B(n3889), .A(n3886), .S(n14), .Y(n3900) );
  MUX2X1 U4253 ( .B(mem[213]), .A(mem[246]), .S(n4472), .Y(n3894) );
  MUX2X1 U4254 ( .B(mem[147]), .A(mem[180]), .S(n4472), .Y(n3893) );
  MUX2X1 U4255 ( .B(mem[81]), .A(mem[114]), .S(n4472), .Y(n3897) );
  MUX2X1 U4256 ( .B(mem[15]), .A(mem[48]), .S(n4472), .Y(n3896) );
  MUX2X1 U4257 ( .B(n3895), .A(n3892), .S(n14), .Y(n3899) );
  MUX2X1 U4258 ( .B(n3898), .A(n3883), .S(n16), .Y(n4426) );
  MUX2X1 U4259 ( .B(mem[1006]), .A(mem[1039]), .S(n4472), .Y(n3903) );
  MUX2X1 U4260 ( .B(mem[940]), .A(mem[973]), .S(n4472), .Y(n3902) );
  MUX2X1 U4261 ( .B(mem[874]), .A(mem[907]), .S(n4472), .Y(n3906) );
  MUX2X1 U4262 ( .B(mem[808]), .A(mem[841]), .S(n4472), .Y(n3905) );
  MUX2X1 U4263 ( .B(n3904), .A(n3901), .S(n14), .Y(n3915) );
  MUX2X1 U4264 ( .B(mem[742]), .A(mem[775]), .S(n4472), .Y(n3909) );
  MUX2X1 U4265 ( .B(mem[676]), .A(mem[709]), .S(n4472), .Y(n3908) );
  MUX2X1 U4266 ( .B(mem[610]), .A(mem[643]), .S(n4472), .Y(n3912) );
  MUX2X1 U4267 ( .B(mem[544]), .A(mem[577]), .S(n4472), .Y(n3911) );
  MUX2X1 U4268 ( .B(n3910), .A(n3907), .S(n14), .Y(n3914) );
  MUX2X1 U4269 ( .B(mem[478]), .A(mem[511]), .S(n4473), .Y(n3918) );
  MUX2X1 U4270 ( .B(mem[412]), .A(mem[445]), .S(n4473), .Y(n3917) );
  MUX2X1 U4271 ( .B(mem[346]), .A(mem[379]), .S(n4473), .Y(n3921) );
  MUX2X1 U4272 ( .B(mem[280]), .A(mem[313]), .S(n4473), .Y(n3920) );
  MUX2X1 U4273 ( .B(n3919), .A(n3916), .S(n14), .Y(n3930) );
  MUX2X1 U4274 ( .B(mem[214]), .A(mem[247]), .S(n4473), .Y(n3924) );
  MUX2X1 U4275 ( .B(mem[148]), .A(mem[181]), .S(n4473), .Y(n3923) );
  MUX2X1 U4276 ( .B(mem[82]), .A(mem[115]), .S(n4473), .Y(n3927) );
  MUX2X1 U4277 ( .B(mem[16]), .A(mem[49]), .S(n4473), .Y(n3926) );
  MUX2X1 U4278 ( .B(n3925), .A(n3922), .S(n14), .Y(n3929) );
  MUX2X1 U4279 ( .B(n3928), .A(n3913), .S(n16), .Y(n4427) );
  MUX2X1 U4280 ( .B(mem[1007]), .A(mem[1040]), .S(n4473), .Y(n3933) );
  MUX2X1 U4281 ( .B(mem[941]), .A(mem[974]), .S(n4473), .Y(n3932) );
  MUX2X1 U4282 ( .B(mem[875]), .A(mem[908]), .S(n4473), .Y(n3936) );
  MUX2X1 U4283 ( .B(mem[809]), .A(mem[842]), .S(n4473), .Y(n3935) );
  MUX2X1 U4284 ( .B(n3934), .A(n3931), .S(n14), .Y(n3945) );
  MUX2X1 U4285 ( .B(mem[743]), .A(mem[776]), .S(n4474), .Y(n3939) );
  MUX2X1 U4286 ( .B(mem[677]), .A(mem[710]), .S(n4474), .Y(n3938) );
  MUX2X1 U4287 ( .B(mem[611]), .A(mem[644]), .S(n4474), .Y(n3942) );
  MUX2X1 U4288 ( .B(mem[545]), .A(mem[578]), .S(n4474), .Y(n3941) );
  MUX2X1 U4289 ( .B(n3940), .A(n3937), .S(n14), .Y(n3944) );
  MUX2X1 U4290 ( .B(mem[479]), .A(mem[512]), .S(n4474), .Y(n3948) );
  MUX2X1 U4291 ( .B(mem[413]), .A(mem[446]), .S(n4474), .Y(n3947) );
  MUX2X1 U4292 ( .B(mem[347]), .A(mem[380]), .S(n4474), .Y(n3951) );
  MUX2X1 U4293 ( .B(mem[281]), .A(mem[314]), .S(n4474), .Y(n3950) );
  MUX2X1 U4294 ( .B(n3949), .A(n3946), .S(n14), .Y(n3960) );
  MUX2X1 U4295 ( .B(mem[215]), .A(mem[248]), .S(n4474), .Y(n3954) );
  MUX2X1 U4296 ( .B(mem[149]), .A(mem[182]), .S(n4474), .Y(n3953) );
  MUX2X1 U4297 ( .B(mem[83]), .A(mem[116]), .S(n4474), .Y(n3957) );
  MUX2X1 U4298 ( .B(mem[17]), .A(mem[50]), .S(n4474), .Y(n3956) );
  MUX2X1 U4299 ( .B(n3955), .A(n3952), .S(n14), .Y(n3959) );
  MUX2X1 U4300 ( .B(n3958), .A(n3943), .S(n16), .Y(n4428) );
  MUX2X1 U4301 ( .B(mem[1008]), .A(mem[1041]), .S(n4475), .Y(n3963) );
  MUX2X1 U4302 ( .B(mem[942]), .A(mem[975]), .S(n4475), .Y(n3962) );
  MUX2X1 U4303 ( .B(mem[876]), .A(mem[909]), .S(n4475), .Y(n3966) );
  MUX2X1 U4304 ( .B(mem[810]), .A(mem[843]), .S(n4475), .Y(n3965) );
  MUX2X1 U4305 ( .B(n3964), .A(n3961), .S(n14), .Y(n3975) );
  MUX2X1 U4306 ( .B(mem[744]), .A(mem[777]), .S(n4475), .Y(n3969) );
  MUX2X1 U4307 ( .B(mem[678]), .A(mem[711]), .S(n4475), .Y(n3968) );
  MUX2X1 U4308 ( .B(mem[612]), .A(mem[645]), .S(n4475), .Y(n3972) );
  MUX2X1 U4309 ( .B(mem[546]), .A(mem[579]), .S(n4475), .Y(n3971) );
  MUX2X1 U4310 ( .B(n3970), .A(n3967), .S(n14), .Y(n3974) );
  MUX2X1 U4311 ( .B(mem[480]), .A(mem[513]), .S(n4475), .Y(n3978) );
  MUX2X1 U4312 ( .B(mem[414]), .A(mem[447]), .S(n4475), .Y(n3977) );
  MUX2X1 U4313 ( .B(mem[348]), .A(mem[381]), .S(n4475), .Y(n3981) );
  MUX2X1 U4314 ( .B(mem[282]), .A(mem[315]), .S(n4475), .Y(n3980) );
  MUX2X1 U4315 ( .B(n3979), .A(n3976), .S(n14), .Y(n3990) );
  MUX2X1 U4316 ( .B(mem[216]), .A(mem[249]), .S(n4476), .Y(n3984) );
  MUX2X1 U4317 ( .B(mem[150]), .A(mem[183]), .S(n4476), .Y(n3983) );
  MUX2X1 U4318 ( .B(mem[84]), .A(mem[117]), .S(n4476), .Y(n3987) );
  MUX2X1 U4319 ( .B(mem[18]), .A(mem[51]), .S(n4476), .Y(n3986) );
  MUX2X1 U4320 ( .B(n3985), .A(n3982), .S(n14), .Y(n3989) );
  MUX2X1 U4321 ( .B(n3988), .A(n3973), .S(n16), .Y(n4429) );
  MUX2X1 U4322 ( .B(mem[1009]), .A(mem[1042]), .S(n4476), .Y(n3993) );
  MUX2X1 U4323 ( .B(mem[943]), .A(mem[976]), .S(n4476), .Y(n3992) );
  MUX2X1 U4324 ( .B(mem[877]), .A(mem[910]), .S(n4476), .Y(n3996) );
  MUX2X1 U4325 ( .B(mem[811]), .A(mem[844]), .S(n4476), .Y(n3995) );
  MUX2X1 U4326 ( .B(n3994), .A(n3991), .S(n14), .Y(n4005) );
  MUX2X1 U4327 ( .B(mem[745]), .A(mem[778]), .S(n4476), .Y(n3999) );
  MUX2X1 U4328 ( .B(mem[679]), .A(mem[712]), .S(n4476), .Y(n3998) );
  MUX2X1 U4329 ( .B(mem[613]), .A(mem[646]), .S(n4476), .Y(n4002) );
  MUX2X1 U4330 ( .B(mem[547]), .A(mem[580]), .S(n4476), .Y(n4001) );
  MUX2X1 U4331 ( .B(n4000), .A(n3997), .S(n14), .Y(n4004) );
  MUX2X1 U4332 ( .B(mem[481]), .A(mem[514]), .S(n4477), .Y(n4008) );
  MUX2X1 U4333 ( .B(mem[415]), .A(mem[448]), .S(n4477), .Y(n4007) );
  MUX2X1 U4334 ( .B(mem[349]), .A(mem[382]), .S(n4477), .Y(n4011) );
  MUX2X1 U4335 ( .B(mem[283]), .A(mem[316]), .S(n4477), .Y(n4010) );
  MUX2X1 U4336 ( .B(n4009), .A(n4006), .S(n14), .Y(n4020) );
  MUX2X1 U4337 ( .B(mem[217]), .A(mem[250]), .S(n4477), .Y(n4014) );
  MUX2X1 U4338 ( .B(mem[151]), .A(mem[184]), .S(n4477), .Y(n4013) );
  MUX2X1 U4339 ( .B(mem[85]), .A(mem[118]), .S(n4477), .Y(n4017) );
  MUX2X1 U4340 ( .B(mem[19]), .A(mem[52]), .S(n4477), .Y(n4016) );
  MUX2X1 U4341 ( .B(n4015), .A(n4012), .S(n14), .Y(n4019) );
  MUX2X1 U4342 ( .B(n4018), .A(n4003), .S(n16), .Y(n4430) );
  MUX2X1 U4343 ( .B(mem[1010]), .A(mem[1043]), .S(n4477), .Y(n4023) );
  MUX2X1 U4344 ( .B(mem[944]), .A(mem[977]), .S(n4477), .Y(n4022) );
  MUX2X1 U4345 ( .B(mem[878]), .A(mem[911]), .S(n4477), .Y(n4026) );
  MUX2X1 U4346 ( .B(mem[812]), .A(mem[845]), .S(n4477), .Y(n4025) );
  MUX2X1 U4347 ( .B(n4024), .A(n4021), .S(n14), .Y(n4035) );
  MUX2X1 U4348 ( .B(mem[746]), .A(mem[779]), .S(n4478), .Y(n4029) );
  MUX2X1 U4349 ( .B(mem[680]), .A(mem[713]), .S(n4478), .Y(n4028) );
  MUX2X1 U4350 ( .B(mem[614]), .A(mem[647]), .S(n4478), .Y(n4032) );
  MUX2X1 U4351 ( .B(mem[548]), .A(mem[581]), .S(n4478), .Y(n4031) );
  MUX2X1 U4352 ( .B(n4030), .A(n4027), .S(n14), .Y(n4034) );
  MUX2X1 U4353 ( .B(mem[482]), .A(mem[515]), .S(n4478), .Y(n4038) );
  MUX2X1 U4354 ( .B(mem[416]), .A(mem[449]), .S(n4478), .Y(n4037) );
  MUX2X1 U4355 ( .B(mem[350]), .A(mem[383]), .S(n4478), .Y(n4041) );
  MUX2X1 U4356 ( .B(mem[284]), .A(mem[317]), .S(n4478), .Y(n4040) );
  MUX2X1 U4357 ( .B(n4039), .A(n4036), .S(n14), .Y(n4050) );
  MUX2X1 U4358 ( .B(mem[218]), .A(mem[251]), .S(n4478), .Y(n4044) );
  MUX2X1 U4359 ( .B(mem[152]), .A(mem[185]), .S(n4478), .Y(n4043) );
  MUX2X1 U4360 ( .B(mem[86]), .A(mem[119]), .S(n4478), .Y(n4047) );
  MUX2X1 U4361 ( .B(mem[20]), .A(mem[53]), .S(n4478), .Y(n4046) );
  MUX2X1 U4362 ( .B(n4045), .A(n4042), .S(n14), .Y(n4049) );
  MUX2X1 U4363 ( .B(n4048), .A(n4033), .S(n16), .Y(n4431) );
  MUX2X1 U4364 ( .B(mem[1011]), .A(mem[1044]), .S(n4479), .Y(n4053) );
  MUX2X1 U4365 ( .B(mem[945]), .A(mem[978]), .S(n4479), .Y(n4052) );
  MUX2X1 U4366 ( .B(mem[879]), .A(mem[912]), .S(n4479), .Y(n4056) );
  MUX2X1 U4367 ( .B(mem[813]), .A(mem[846]), .S(n4479), .Y(n4055) );
  MUX2X1 U4368 ( .B(n4054), .A(n4051), .S(n14), .Y(n4065) );
  MUX2X1 U4369 ( .B(mem[747]), .A(mem[780]), .S(n4479), .Y(n4059) );
  MUX2X1 U4370 ( .B(mem[681]), .A(mem[714]), .S(n4479), .Y(n4058) );
  MUX2X1 U4371 ( .B(mem[615]), .A(mem[648]), .S(n4479), .Y(n4062) );
  MUX2X1 U4372 ( .B(mem[549]), .A(mem[582]), .S(n4479), .Y(n4061) );
  MUX2X1 U4373 ( .B(n4060), .A(n4057), .S(n14), .Y(n4064) );
  MUX2X1 U4374 ( .B(mem[483]), .A(mem[516]), .S(n4479), .Y(n4068) );
  MUX2X1 U4375 ( .B(mem[417]), .A(mem[450]), .S(n4479), .Y(n4067) );
  MUX2X1 U4376 ( .B(mem[351]), .A(mem[384]), .S(n4479), .Y(n4071) );
  MUX2X1 U4377 ( .B(mem[285]), .A(mem[318]), .S(n4479), .Y(n4070) );
  MUX2X1 U4378 ( .B(n4069), .A(n4066), .S(n14), .Y(n4080) );
  MUX2X1 U4379 ( .B(mem[219]), .A(mem[252]), .S(n4480), .Y(n4074) );
  MUX2X1 U4380 ( .B(mem[153]), .A(mem[186]), .S(n4480), .Y(n4073) );
  MUX2X1 U4381 ( .B(mem[87]), .A(mem[120]), .S(n4480), .Y(n4077) );
  MUX2X1 U4382 ( .B(mem[21]), .A(mem[54]), .S(n4480), .Y(n4076) );
  MUX2X1 U4383 ( .B(n4075), .A(n4072), .S(n14), .Y(n4079) );
  MUX2X1 U4384 ( .B(n4078), .A(n4063), .S(n16), .Y(n4432) );
  MUX2X1 U4385 ( .B(mem[1012]), .A(mem[1045]), .S(n4480), .Y(n4083) );
  MUX2X1 U4386 ( .B(mem[946]), .A(mem[979]), .S(n4480), .Y(n4082) );
  MUX2X1 U4387 ( .B(mem[880]), .A(mem[913]), .S(n4480), .Y(n4086) );
  MUX2X1 U4388 ( .B(mem[814]), .A(mem[847]), .S(n4480), .Y(n4085) );
  MUX2X1 U4389 ( .B(n4084), .A(n4081), .S(n14), .Y(n4095) );
  MUX2X1 U4390 ( .B(mem[748]), .A(mem[781]), .S(n4480), .Y(n4089) );
  MUX2X1 U4391 ( .B(mem[682]), .A(mem[715]), .S(n4480), .Y(n4088) );
  MUX2X1 U4392 ( .B(mem[616]), .A(mem[649]), .S(n4480), .Y(n4092) );
  MUX2X1 U4393 ( .B(mem[550]), .A(mem[583]), .S(n4480), .Y(n4091) );
  MUX2X1 U4394 ( .B(n4090), .A(n4087), .S(n14), .Y(n4094) );
  MUX2X1 U4395 ( .B(mem[484]), .A(mem[517]), .S(n4481), .Y(n4098) );
  MUX2X1 U4396 ( .B(mem[418]), .A(mem[451]), .S(n4481), .Y(n4097) );
  MUX2X1 U4397 ( .B(mem[352]), .A(mem[385]), .S(n4481), .Y(n4101) );
  MUX2X1 U4398 ( .B(mem[286]), .A(mem[319]), .S(n4481), .Y(n4100) );
  MUX2X1 U4399 ( .B(n4099), .A(n4096), .S(n14), .Y(n4110) );
  MUX2X1 U4400 ( .B(mem[220]), .A(mem[253]), .S(n4481), .Y(n4104) );
  MUX2X1 U4401 ( .B(mem[154]), .A(mem[187]), .S(n4481), .Y(n4103) );
  MUX2X1 U4402 ( .B(mem[88]), .A(mem[121]), .S(n4481), .Y(n4107) );
  MUX2X1 U4403 ( .B(mem[22]), .A(mem[55]), .S(n4481), .Y(n4106) );
  MUX2X1 U4404 ( .B(n4105), .A(n4102), .S(n14), .Y(n4109) );
  MUX2X1 U4405 ( .B(n4108), .A(n4093), .S(n16), .Y(n4433) );
  MUX2X1 U4406 ( .B(mem[1013]), .A(mem[1046]), .S(n4481), .Y(n4113) );
  MUX2X1 U4407 ( .B(mem[947]), .A(mem[980]), .S(n4481), .Y(n4112) );
  MUX2X1 U4408 ( .B(mem[881]), .A(mem[914]), .S(n4481), .Y(n4116) );
  MUX2X1 U4409 ( .B(mem[815]), .A(mem[848]), .S(n4481), .Y(n4115) );
  MUX2X1 U4410 ( .B(n4114), .A(n4111), .S(n14), .Y(n4125) );
  MUX2X1 U4411 ( .B(mem[749]), .A(mem[782]), .S(n4482), .Y(n4119) );
  MUX2X1 U4412 ( .B(mem[683]), .A(mem[716]), .S(n4482), .Y(n4118) );
  MUX2X1 U4413 ( .B(mem[617]), .A(mem[650]), .S(n4482), .Y(n4122) );
  MUX2X1 U4414 ( .B(mem[551]), .A(mem[584]), .S(n4482), .Y(n4121) );
  MUX2X1 U4415 ( .B(n4120), .A(n4117), .S(n14), .Y(n4124) );
  MUX2X1 U4416 ( .B(mem[485]), .A(mem[518]), .S(n4482), .Y(n4128) );
  MUX2X1 U4417 ( .B(mem[419]), .A(mem[452]), .S(n4482), .Y(n4127) );
  MUX2X1 U4418 ( .B(mem[353]), .A(mem[386]), .S(n4482), .Y(n4131) );
  MUX2X1 U4419 ( .B(mem[287]), .A(mem[320]), .S(n4482), .Y(n4130) );
  MUX2X1 U4420 ( .B(n4129), .A(n4126), .S(n14), .Y(n4140) );
  MUX2X1 U4421 ( .B(mem[221]), .A(mem[254]), .S(n4482), .Y(n4134) );
  MUX2X1 U4422 ( .B(mem[155]), .A(mem[188]), .S(n4482), .Y(n4133) );
  MUX2X1 U4423 ( .B(mem[89]), .A(mem[122]), .S(n4482), .Y(n4137) );
  MUX2X1 U4424 ( .B(mem[23]), .A(mem[56]), .S(n4482), .Y(n4136) );
  MUX2X1 U4425 ( .B(n4135), .A(n4132), .S(n14), .Y(n4139) );
  MUX2X1 U4426 ( .B(n4138), .A(n4123), .S(n16), .Y(n4434) );
  MUX2X1 U4427 ( .B(mem[1014]), .A(mem[1047]), .S(n4483), .Y(n4143) );
  MUX2X1 U4428 ( .B(mem[948]), .A(mem[981]), .S(n4483), .Y(n4142) );
  MUX2X1 U4429 ( .B(mem[882]), .A(mem[915]), .S(n4483), .Y(n4146) );
  MUX2X1 U4430 ( .B(mem[816]), .A(mem[849]), .S(n4483), .Y(n4145) );
  MUX2X1 U4431 ( .B(n4144), .A(n4141), .S(n14), .Y(n4155) );
  MUX2X1 U4432 ( .B(mem[750]), .A(mem[783]), .S(n4483), .Y(n4149) );
  MUX2X1 U4433 ( .B(mem[684]), .A(mem[717]), .S(n4483), .Y(n4148) );
  MUX2X1 U4434 ( .B(mem[618]), .A(mem[651]), .S(n4483), .Y(n4152) );
  MUX2X1 U4435 ( .B(mem[552]), .A(mem[585]), .S(n4483), .Y(n4151) );
  MUX2X1 U4436 ( .B(n4150), .A(n4147), .S(n14), .Y(n4154) );
  MUX2X1 U4437 ( .B(mem[486]), .A(mem[519]), .S(n4483), .Y(n4158) );
  MUX2X1 U4438 ( .B(mem[420]), .A(mem[453]), .S(n4483), .Y(n4157) );
  MUX2X1 U4439 ( .B(mem[354]), .A(mem[387]), .S(n4483), .Y(n4161) );
  MUX2X1 U4440 ( .B(mem[288]), .A(mem[321]), .S(n4483), .Y(n4160) );
  MUX2X1 U4441 ( .B(n4159), .A(n4156), .S(n14), .Y(n4170) );
  MUX2X1 U4442 ( .B(mem[222]), .A(mem[255]), .S(n4484), .Y(n4164) );
  MUX2X1 U4443 ( .B(mem[156]), .A(mem[189]), .S(n4484), .Y(n4163) );
  MUX2X1 U4444 ( .B(mem[90]), .A(mem[123]), .S(n4484), .Y(n4167) );
  MUX2X1 U4445 ( .B(mem[24]), .A(mem[57]), .S(n4484), .Y(n4166) );
  MUX2X1 U4446 ( .B(n4165), .A(n4162), .S(n14), .Y(n4169) );
  MUX2X1 U4447 ( .B(n4168), .A(n4153), .S(n16), .Y(n4435) );
  MUX2X1 U4448 ( .B(mem[1015]), .A(mem[1048]), .S(n4484), .Y(n4173) );
  MUX2X1 U4449 ( .B(mem[949]), .A(mem[982]), .S(n4484), .Y(n4172) );
  MUX2X1 U4450 ( .B(mem[883]), .A(mem[916]), .S(n4484), .Y(n4176) );
  MUX2X1 U4451 ( .B(mem[817]), .A(mem[850]), .S(n4484), .Y(n4175) );
  MUX2X1 U4452 ( .B(n4174), .A(n4171), .S(n14), .Y(n4185) );
  MUX2X1 U4453 ( .B(mem[751]), .A(mem[784]), .S(n4484), .Y(n4179) );
  MUX2X1 U4454 ( .B(mem[685]), .A(mem[718]), .S(n4484), .Y(n4178) );
  MUX2X1 U4455 ( .B(mem[619]), .A(mem[652]), .S(n4484), .Y(n4182) );
  MUX2X1 U4456 ( .B(mem[553]), .A(mem[586]), .S(n4484), .Y(n4181) );
  MUX2X1 U4457 ( .B(n4180), .A(n4177), .S(n14), .Y(n4184) );
  MUX2X1 U4458 ( .B(mem[487]), .A(mem[520]), .S(n4485), .Y(n4188) );
  MUX2X1 U4459 ( .B(mem[421]), .A(mem[454]), .S(n4485), .Y(n4187) );
  MUX2X1 U4460 ( .B(mem[355]), .A(mem[388]), .S(n4485), .Y(n4191) );
  MUX2X1 U4461 ( .B(mem[289]), .A(mem[322]), .S(n4485), .Y(n4190) );
  MUX2X1 U4462 ( .B(n4189), .A(n4186), .S(n14), .Y(n4200) );
  MUX2X1 U4463 ( .B(mem[223]), .A(mem[256]), .S(n4485), .Y(n4194) );
  MUX2X1 U4464 ( .B(mem[157]), .A(mem[190]), .S(n4485), .Y(n4193) );
  MUX2X1 U4465 ( .B(mem[91]), .A(mem[124]), .S(n4485), .Y(n4197) );
  MUX2X1 U4466 ( .B(mem[25]), .A(mem[58]), .S(n4485), .Y(n4196) );
  MUX2X1 U4467 ( .B(n4195), .A(n4192), .S(n14), .Y(n4199) );
  MUX2X1 U4468 ( .B(n4198), .A(n4183), .S(n16), .Y(n4436) );
  MUX2X1 U4469 ( .B(mem[1016]), .A(mem[1049]), .S(n4485), .Y(n4203) );
  MUX2X1 U4470 ( .B(mem[950]), .A(mem[983]), .S(n4485), .Y(n4202) );
  MUX2X1 U4471 ( .B(mem[884]), .A(mem[917]), .S(n4485), .Y(n4206) );
  MUX2X1 U4472 ( .B(mem[818]), .A(mem[851]), .S(n4485), .Y(n4205) );
  MUX2X1 U4473 ( .B(n4204), .A(n4201), .S(n14), .Y(n4215) );
  MUX2X1 U4474 ( .B(mem[752]), .A(mem[785]), .S(n4486), .Y(n4209) );
  MUX2X1 U4475 ( .B(mem[686]), .A(mem[719]), .S(n4486), .Y(n4208) );
  MUX2X1 U4476 ( .B(mem[620]), .A(mem[653]), .S(n4486), .Y(n4212) );
  MUX2X1 U4477 ( .B(mem[554]), .A(mem[587]), .S(n4486), .Y(n4211) );
  MUX2X1 U4478 ( .B(n4210), .A(n4207), .S(n14), .Y(n4214) );
  MUX2X1 U4479 ( .B(mem[488]), .A(mem[521]), .S(n4486), .Y(n4218) );
  MUX2X1 U4480 ( .B(mem[422]), .A(mem[455]), .S(n4486), .Y(n4217) );
  MUX2X1 U4481 ( .B(mem[356]), .A(mem[389]), .S(n4486), .Y(n4221) );
  MUX2X1 U4482 ( .B(mem[290]), .A(mem[323]), .S(n4486), .Y(n4220) );
  MUX2X1 U4483 ( .B(n4219), .A(n4216), .S(n14), .Y(n4230) );
  MUX2X1 U4484 ( .B(mem[224]), .A(mem[257]), .S(n4486), .Y(n4224) );
  MUX2X1 U4485 ( .B(mem[158]), .A(mem[191]), .S(n4486), .Y(n4223) );
  MUX2X1 U4486 ( .B(mem[92]), .A(mem[125]), .S(n4486), .Y(n4227) );
  MUX2X1 U4487 ( .B(mem[26]), .A(mem[59]), .S(n4486), .Y(n4226) );
  MUX2X1 U4488 ( .B(n4225), .A(n4222), .S(n14), .Y(n4229) );
  MUX2X1 U4489 ( .B(n4228), .A(n4213), .S(n16), .Y(n4437) );
  MUX2X1 U4490 ( .B(mem[1017]), .A(mem[1050]), .S(n4487), .Y(n4233) );
  MUX2X1 U4491 ( .B(mem[951]), .A(mem[984]), .S(n4487), .Y(n4232) );
  MUX2X1 U4492 ( .B(mem[885]), .A(mem[918]), .S(n4487), .Y(n4236) );
  MUX2X1 U4493 ( .B(mem[819]), .A(mem[852]), .S(n4487), .Y(n4235) );
  MUX2X1 U4494 ( .B(n4234), .A(n4231), .S(n14), .Y(n4245) );
  MUX2X1 U4495 ( .B(mem[753]), .A(mem[786]), .S(n4487), .Y(n4239) );
  MUX2X1 U4496 ( .B(mem[687]), .A(mem[720]), .S(n4487), .Y(n4238) );
  MUX2X1 U4497 ( .B(mem[621]), .A(mem[654]), .S(n4487), .Y(n4242) );
  MUX2X1 U4498 ( .B(mem[555]), .A(mem[588]), .S(n4487), .Y(n4241) );
  MUX2X1 U4499 ( .B(n4240), .A(n4237), .S(n14), .Y(n4244) );
  MUX2X1 U4500 ( .B(mem[489]), .A(mem[522]), .S(n4487), .Y(n4248) );
  MUX2X1 U4501 ( .B(mem[423]), .A(mem[456]), .S(n4487), .Y(n4247) );
  MUX2X1 U4502 ( .B(mem[357]), .A(mem[390]), .S(n4487), .Y(n4251) );
  MUX2X1 U4503 ( .B(mem[291]), .A(mem[324]), .S(n4487), .Y(n4250) );
  MUX2X1 U4504 ( .B(n4249), .A(n4246), .S(n14), .Y(n4260) );
  MUX2X1 U4505 ( .B(mem[225]), .A(mem[258]), .S(n4488), .Y(n4254) );
  MUX2X1 U4506 ( .B(mem[159]), .A(mem[192]), .S(n4488), .Y(n4253) );
  MUX2X1 U4507 ( .B(mem[93]), .A(mem[126]), .S(n4488), .Y(n4257) );
  MUX2X1 U4508 ( .B(mem[27]), .A(mem[60]), .S(n4488), .Y(n4256) );
  MUX2X1 U4509 ( .B(n4255), .A(n4252), .S(n14), .Y(n4259) );
  MUX2X1 U4510 ( .B(n4258), .A(n4243), .S(n16), .Y(n4438) );
  MUX2X1 U4511 ( .B(mem[1018]), .A(mem[1051]), .S(n4488), .Y(n4263) );
  MUX2X1 U4512 ( .B(mem[952]), .A(mem[985]), .S(n4488), .Y(n4262) );
  MUX2X1 U4513 ( .B(mem[886]), .A(mem[919]), .S(n4488), .Y(n4266) );
  MUX2X1 U4514 ( .B(mem[820]), .A(mem[853]), .S(n4488), .Y(n4265) );
  MUX2X1 U4515 ( .B(n4264), .A(n4261), .S(n14), .Y(n4275) );
  MUX2X1 U4516 ( .B(mem[754]), .A(mem[787]), .S(n4488), .Y(n4269) );
  MUX2X1 U4517 ( .B(mem[688]), .A(mem[721]), .S(n4488), .Y(n4268) );
  MUX2X1 U4518 ( .B(mem[622]), .A(mem[655]), .S(n4488), .Y(n4272) );
  MUX2X1 U4519 ( .B(mem[556]), .A(mem[589]), .S(n4488), .Y(n4271) );
  MUX2X1 U4520 ( .B(n4270), .A(n4267), .S(n14), .Y(n4274) );
  MUX2X1 U4521 ( .B(mem[490]), .A(mem[523]), .S(n4489), .Y(n4278) );
  MUX2X1 U4522 ( .B(mem[424]), .A(mem[457]), .S(n4489), .Y(n4277) );
  MUX2X1 U4523 ( .B(mem[358]), .A(mem[391]), .S(n4489), .Y(n4281) );
  MUX2X1 U4524 ( .B(mem[292]), .A(mem[325]), .S(n4489), .Y(n4280) );
  MUX2X1 U4525 ( .B(n4279), .A(n4276), .S(n14), .Y(n4290) );
  MUX2X1 U4526 ( .B(mem[226]), .A(mem[259]), .S(n4489), .Y(n4284) );
  MUX2X1 U4527 ( .B(mem[160]), .A(mem[193]), .S(n4489), .Y(n4283) );
  MUX2X1 U4528 ( .B(mem[94]), .A(mem[127]), .S(n4489), .Y(n4287) );
  MUX2X1 U4529 ( .B(mem[28]), .A(mem[61]), .S(n4489), .Y(n4286) );
  MUX2X1 U4530 ( .B(n4285), .A(n4282), .S(n14), .Y(n4289) );
  MUX2X1 U4531 ( .B(n4288), .A(n4273), .S(n16), .Y(n4439) );
  MUX2X1 U4532 ( .B(mem[1019]), .A(mem[1052]), .S(n4489), .Y(n4293) );
  MUX2X1 U4533 ( .B(mem[953]), .A(mem[986]), .S(n4489), .Y(n4292) );
  MUX2X1 U4534 ( .B(mem[887]), .A(mem[920]), .S(n4489), .Y(n4296) );
  MUX2X1 U4535 ( .B(mem[821]), .A(mem[854]), .S(n4489), .Y(n4295) );
  MUX2X1 U4536 ( .B(n4294), .A(n4291), .S(n14), .Y(n4305) );
  MUX2X1 U4537 ( .B(mem[755]), .A(mem[788]), .S(n4490), .Y(n4299) );
  MUX2X1 U4538 ( .B(mem[689]), .A(mem[722]), .S(n4490), .Y(n4298) );
  MUX2X1 U4539 ( .B(mem[623]), .A(mem[656]), .S(n4490), .Y(n4302) );
  MUX2X1 U4540 ( .B(mem[557]), .A(mem[590]), .S(n4490), .Y(n4301) );
  MUX2X1 U4541 ( .B(n4300), .A(n4297), .S(n14), .Y(n4304) );
  MUX2X1 U4542 ( .B(mem[491]), .A(mem[524]), .S(n4490), .Y(n4308) );
  MUX2X1 U4543 ( .B(mem[425]), .A(mem[458]), .S(n4490), .Y(n4307) );
  MUX2X1 U4544 ( .B(mem[359]), .A(mem[392]), .S(n4490), .Y(n4311) );
  MUX2X1 U4545 ( .B(mem[293]), .A(mem[326]), .S(n4490), .Y(n4310) );
  MUX2X1 U4546 ( .B(n4309), .A(n4306), .S(n14), .Y(n4320) );
  MUX2X1 U4547 ( .B(mem[227]), .A(mem[260]), .S(n4490), .Y(n4314) );
  MUX2X1 U4548 ( .B(mem[161]), .A(mem[194]), .S(n4490), .Y(n4313) );
  MUX2X1 U4549 ( .B(mem[95]), .A(mem[128]), .S(n4490), .Y(n4317) );
  MUX2X1 U4550 ( .B(mem[29]), .A(mem[62]), .S(n4490), .Y(n4316) );
  MUX2X1 U4551 ( .B(n4315), .A(n4312), .S(n14), .Y(n4319) );
  MUX2X1 U4552 ( .B(n4318), .A(n4303), .S(n16), .Y(n4440) );
  MUX2X1 U4553 ( .B(mem[1020]), .A(mem[1053]), .S(n4491), .Y(n4323) );
  MUX2X1 U4554 ( .B(mem[954]), .A(mem[987]), .S(n4491), .Y(n4322) );
  MUX2X1 U4555 ( .B(mem[888]), .A(mem[921]), .S(n4491), .Y(n4326) );
  MUX2X1 U4556 ( .B(mem[822]), .A(mem[855]), .S(n4491), .Y(n4325) );
  MUX2X1 U4557 ( .B(n4324), .A(n4321), .S(n14), .Y(n4335) );
  MUX2X1 U4558 ( .B(mem[756]), .A(mem[789]), .S(n4491), .Y(n4329) );
  MUX2X1 U4559 ( .B(mem[690]), .A(mem[723]), .S(n4491), .Y(n4328) );
  MUX2X1 U4560 ( .B(mem[624]), .A(mem[657]), .S(n4491), .Y(n4332) );
  MUX2X1 U4561 ( .B(mem[558]), .A(mem[591]), .S(n4491), .Y(n4331) );
  MUX2X1 U4562 ( .B(n4330), .A(n4327), .S(n14), .Y(n4334) );
  MUX2X1 U4563 ( .B(mem[492]), .A(mem[525]), .S(n4491), .Y(n4338) );
  MUX2X1 U4564 ( .B(mem[426]), .A(mem[459]), .S(n4491), .Y(n4337) );
  MUX2X1 U4565 ( .B(mem[360]), .A(mem[393]), .S(n4491), .Y(n4341) );
  MUX2X1 U4566 ( .B(mem[294]), .A(mem[327]), .S(n4491), .Y(n4340) );
  MUX2X1 U4567 ( .B(n4339), .A(n4336), .S(n14), .Y(n4350) );
  MUX2X1 U4568 ( .B(mem[228]), .A(mem[261]), .S(n4492), .Y(n4344) );
  MUX2X1 U4569 ( .B(mem[162]), .A(mem[195]), .S(n4492), .Y(n4343) );
  MUX2X1 U4570 ( .B(mem[96]), .A(mem[129]), .S(n4492), .Y(n4347) );
  MUX2X1 U4571 ( .B(mem[30]), .A(mem[63]), .S(n4492), .Y(n4346) );
  MUX2X1 U4572 ( .B(n4345), .A(n4342), .S(n14), .Y(n4349) );
  MUX2X1 U4573 ( .B(n4348), .A(n4333), .S(n16), .Y(n4441) );
  MUX2X1 U4574 ( .B(mem[1021]), .A(mem[1054]), .S(n4492), .Y(n4353) );
  MUX2X1 U4575 ( .B(mem[955]), .A(mem[988]), .S(n4492), .Y(n4352) );
  MUX2X1 U4576 ( .B(mem[889]), .A(mem[922]), .S(n4492), .Y(n4356) );
  MUX2X1 U4577 ( .B(mem[823]), .A(mem[856]), .S(n4492), .Y(n4355) );
  MUX2X1 U4578 ( .B(n4354), .A(n4351), .S(n14), .Y(n4365) );
  MUX2X1 U4579 ( .B(mem[757]), .A(mem[790]), .S(n4492), .Y(n4359) );
  MUX2X1 U4580 ( .B(mem[691]), .A(mem[724]), .S(n4492), .Y(n4358) );
  MUX2X1 U4581 ( .B(mem[625]), .A(mem[658]), .S(n4492), .Y(n4362) );
  MUX2X1 U4582 ( .B(mem[559]), .A(mem[592]), .S(n4492), .Y(n4361) );
  MUX2X1 U4583 ( .B(n4360), .A(n4357), .S(n14), .Y(n4364) );
  MUX2X1 U4584 ( .B(mem[493]), .A(mem[526]), .S(n4493), .Y(n4368) );
  MUX2X1 U4585 ( .B(mem[427]), .A(mem[460]), .S(n4493), .Y(n4367) );
  MUX2X1 U4586 ( .B(mem[361]), .A(mem[394]), .S(n4493), .Y(n4371) );
  MUX2X1 U4587 ( .B(mem[295]), .A(mem[328]), .S(n4493), .Y(n4370) );
  MUX2X1 U4588 ( .B(n4369), .A(n4366), .S(n14), .Y(n4380) );
  MUX2X1 U4589 ( .B(mem[229]), .A(mem[262]), .S(n4493), .Y(n4374) );
  MUX2X1 U4590 ( .B(mem[163]), .A(mem[196]), .S(n4493), .Y(n4373) );
  MUX2X1 U4591 ( .B(mem[97]), .A(mem[130]), .S(n4493), .Y(n4377) );
  MUX2X1 U4592 ( .B(mem[31]), .A(mem[64]), .S(n4493), .Y(n4376) );
  MUX2X1 U4593 ( .B(n4375), .A(n4372), .S(n14), .Y(n4379) );
  MUX2X1 U4594 ( .B(n4378), .A(n4363), .S(n16), .Y(n4442) );
  MUX2X1 U4595 ( .B(mem[1022]), .A(mem[1055]), .S(n4493), .Y(n4383) );
  MUX2X1 U4596 ( .B(mem[956]), .A(mem[989]), .S(n4493), .Y(n4382) );
  MUX2X1 U4597 ( .B(mem[890]), .A(mem[923]), .S(n4493), .Y(n4386) );
  MUX2X1 U4598 ( .B(mem[824]), .A(mem[857]), .S(n4493), .Y(n4385) );
  MUX2X1 U4599 ( .B(n4384), .A(n4381), .S(n14), .Y(n4395) );
  MUX2X1 U4600 ( .B(mem[758]), .A(mem[791]), .S(n4494), .Y(n4389) );
  MUX2X1 U4601 ( .B(mem[692]), .A(mem[725]), .S(n4494), .Y(n4388) );
  MUX2X1 U4602 ( .B(mem[626]), .A(mem[659]), .S(n4494), .Y(n4392) );
  MUX2X1 U4603 ( .B(mem[560]), .A(mem[593]), .S(n4494), .Y(n4391) );
  MUX2X1 U4604 ( .B(n4390), .A(n4387), .S(n14), .Y(n4394) );
  MUX2X1 U4605 ( .B(mem[494]), .A(mem[527]), .S(n4494), .Y(n4398) );
  MUX2X1 U4606 ( .B(mem[428]), .A(mem[461]), .S(n4494), .Y(n4397) );
  MUX2X1 U4607 ( .B(mem[362]), .A(mem[395]), .S(n4494), .Y(n4401) );
  MUX2X1 U4608 ( .B(mem[296]), .A(mem[329]), .S(n4494), .Y(n4400) );
  MUX2X1 U4609 ( .B(n4399), .A(n4396), .S(n14), .Y(n4410) );
  MUX2X1 U4610 ( .B(mem[230]), .A(mem[263]), .S(n4494), .Y(n4404) );
  MUX2X1 U4611 ( .B(mem[164]), .A(mem[197]), .S(n4494), .Y(n4403) );
  MUX2X1 U4612 ( .B(mem[98]), .A(mem[131]), .S(n4494), .Y(n4407) );
  MUX2X1 U4613 ( .B(mem[32]), .A(mem[65]), .S(n4494), .Y(n4406) );
  MUX2X1 U4614 ( .B(n4405), .A(n4402), .S(n14), .Y(n4409) );
  MUX2X1 U4615 ( .B(n4408), .A(n4393), .S(n16), .Y(n4443) );
  OR2X1 U4616 ( .A(n4585), .B(wr_ptr[0]), .Y(sub_93_carry[1]) );
  XNOR2X1 U4617 ( .A(wr_ptr[0]), .B(n4585), .Y(fillcount[0]) );
  XOR2X1 U4618 ( .A(add_51_carry[4]), .B(wr_ptr[4]), .Y(n23) );
  XOR2X1 U4619 ( .A(add_57_carry[4]), .B(n16), .Y(n93) );
endmodule


module FIFO_DEPTH_P25_WIDTH41 ( clk, reset, data_in, put, get, data_out, 
        empty_bar, full_bar, fillcount );
  input [40:0] data_in;
  output [40:0] data_out;
  output [5:0] fillcount;
  input clk, reset, put, get;
  output empty_bar, full_bar;
  wire   n12, n13, n14, n15, n16, n5721, n5722, n20, n21, n22, n23, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n98, n99, n100,
         n101, n381, n383, n385, n387, n389, n391, n393, n395, n397, n399,
         n401, n403, n405, n407, n409, n411, n413, n415, n417, n419, n421,
         n423, n425, n427, n429, n431, n433, n435, n437, n439, n441, n443,
         n445, n447, n449, n451, n453, n455, n457, n459, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n17, n18, n19,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n97, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n382, n384, n386,
         n388, n390, n392, n394, n396, n398, n400, n402, n404, n406, n408,
         n410, n412, n414, n416, n418, n420, n422, n424, n426, n428, n430,
         n432, n434, n436, n438, n440, n442, n444, n446, n448, n450, n452,
         n454, n456, n458, n460, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720;
  wire   [4:0] wr_ptr;
  wire   [1311:0] mem;
  wire   [4:2] add_57_carry;
  wire   [4:2] add_51_carry;
  wire   [5:1] sub_93_carry;

  DFFPOSX1 wr_ptr_reg_0_ ( .D(n3163), .CLK(clk), .Q(wr_ptr[0]) );
  DFFPOSX1 rd_ptr_reg_4_ ( .D(n3162), .CLK(clk), .Q(n16) );
  DFFPOSX1 rd_ptr_reg_0_ ( .D(n3161), .CLK(clk), .Q(n12) );
  DFFPOSX1 rd_ptr_reg_1_ ( .D(n3160), .CLK(clk), .Q(n13) );
  DFFPOSX1 rd_ptr_reg_2_ ( .D(n3159), .CLK(clk), .Q(n14) );
  DFFPOSX1 rd_ptr_reg_3_ ( .D(n3158), .CLK(clk), .Q(n15) );
  DFFPOSX1 wr_ptr_reg_4_ ( .D(n3157), .CLK(clk), .Q(wr_ptr[4]) );
  DFFPOSX1 wr_ptr_reg_1_ ( .D(n3156), .CLK(clk), .Q(wr_ptr[1]) );
  DFFPOSX1 wr_ptr_reg_2_ ( .D(n3155), .CLK(clk), .Q(wr_ptr[2]) );
  DFFPOSX1 wr_ptr_reg_3_ ( .D(n3154), .CLK(clk), .Q(wr_ptr[3]) );
  DFFPOSX1 data_out_reg_40_ ( .D(n5715), .CLK(clk), .Q(data_out[40]) );
  DFFPOSX1 data_out_reg_39_ ( .D(n5714), .CLK(clk), .Q(data_out[39]) );
  DFFPOSX1 data_out_reg_38_ ( .D(n5713), .CLK(clk), .Q(data_out[38]) );
  DFFPOSX1 data_out_reg_37_ ( .D(n5712), .CLK(clk), .Q(data_out[37]) );
  DFFPOSX1 data_out_reg_36_ ( .D(n5711), .CLK(clk), .Q(data_out[36]) );
  DFFPOSX1 data_out_reg_35_ ( .D(n5710), .CLK(clk), .Q(data_out[35]) );
  DFFPOSX1 data_out_reg_34_ ( .D(n5709), .CLK(clk), .Q(data_out[34]) );
  DFFPOSX1 data_out_reg_33_ ( .D(n5708), .CLK(clk), .Q(data_out[33]) );
  DFFPOSX1 data_out_reg_32_ ( .D(n5707), .CLK(clk), .Q(data_out[32]) );
  DFFPOSX1 data_out_reg_31_ ( .D(n5706), .CLK(clk), .Q(data_out[31]) );
  DFFPOSX1 data_out_reg_30_ ( .D(n5705), .CLK(clk), .Q(data_out[30]) );
  DFFPOSX1 data_out_reg_29_ ( .D(n5704), .CLK(clk), .Q(data_out[29]) );
  DFFPOSX1 data_out_reg_28_ ( .D(n5703), .CLK(clk), .Q(data_out[28]) );
  DFFPOSX1 data_out_reg_27_ ( .D(n5702), .CLK(clk), .Q(data_out[27]) );
  DFFPOSX1 data_out_reg_26_ ( .D(n5701), .CLK(clk), .Q(data_out[26]) );
  DFFPOSX1 data_out_reg_25_ ( .D(n5700), .CLK(clk), .Q(data_out[25]) );
  DFFPOSX1 data_out_reg_24_ ( .D(n5699), .CLK(clk), .Q(data_out[24]) );
  DFFPOSX1 data_out_reg_23_ ( .D(n5698), .CLK(clk), .Q(data_out[23]) );
  DFFPOSX1 data_out_reg_22_ ( .D(n5697), .CLK(clk), .Q(data_out[22]) );
  DFFPOSX1 data_out_reg_21_ ( .D(n5696), .CLK(clk), .Q(data_out[21]) );
  DFFPOSX1 data_out_reg_20_ ( .D(n5695), .CLK(clk), .Q(data_out[20]) );
  DFFPOSX1 data_out_reg_19_ ( .D(n5694), .CLK(clk), .Q(data_out[19]) );
  DFFPOSX1 data_out_reg_18_ ( .D(n5693), .CLK(clk), .Q(data_out[18]) );
  DFFPOSX1 data_out_reg_17_ ( .D(n5692), .CLK(clk), .Q(data_out[17]) );
  DFFPOSX1 data_out_reg_16_ ( .D(n5691), .CLK(clk), .Q(data_out[16]) );
  DFFPOSX1 data_out_reg_15_ ( .D(n5690), .CLK(clk), .Q(data_out[15]) );
  DFFPOSX1 data_out_reg_14_ ( .D(n5689), .CLK(clk), .Q(data_out[14]) );
  DFFPOSX1 data_out_reg_13_ ( .D(n5688), .CLK(clk), .Q(data_out[13]) );
  DFFPOSX1 data_out_reg_12_ ( .D(n5687), .CLK(clk), .Q(data_out[12]) );
  DFFPOSX1 data_out_reg_11_ ( .D(n5686), .CLK(clk), .Q(data_out[11]) );
  DFFPOSX1 data_out_reg_10_ ( .D(n5685), .CLK(clk), .Q(data_out[10]) );
  DFFPOSX1 data_out_reg_9_ ( .D(n5684), .CLK(clk), .Q(data_out[9]) );
  DFFPOSX1 data_out_reg_8_ ( .D(n5683), .CLK(clk), .Q(data_out[8]) );
  DFFPOSX1 data_out_reg_7_ ( .D(n5682), .CLK(clk), .Q(data_out[7]) );
  DFFPOSX1 data_out_reg_6_ ( .D(n5681), .CLK(clk), .Q(data_out[6]) );
  DFFPOSX1 data_out_reg_5_ ( .D(n5680), .CLK(clk), .Q(data_out[5]) );
  DFFPOSX1 data_out_reg_4_ ( .D(n5679), .CLK(clk), .Q(data_out[4]) );
  DFFPOSX1 data_out_reg_3_ ( .D(n5678), .CLK(clk), .Q(data_out[3]) );
  DFFPOSX1 data_out_reg_2_ ( .D(n5677), .CLK(clk), .Q(data_out[2]) );
  DFFPOSX1 data_out_reg_1_ ( .D(n5676), .CLK(clk), .Q(data_out[1]) );
  DFFPOSX1 data_out_reg_0_ ( .D(n5675), .CLK(clk), .Q(data_out[0]) );
  DFFPOSX1 mem_reg_31__40_ ( .D(n3153), .CLK(clk), .Q(mem[1311]) );
  DFFPOSX1 mem_reg_31__39_ ( .D(n3152), .CLK(clk), .Q(mem[1310]) );
  DFFPOSX1 mem_reg_31__38_ ( .D(n3151), .CLK(clk), .Q(mem[1309]) );
  DFFPOSX1 mem_reg_31__37_ ( .D(n3150), .CLK(clk), .Q(mem[1308]) );
  DFFPOSX1 mem_reg_31__36_ ( .D(n3149), .CLK(clk), .Q(mem[1307]) );
  DFFPOSX1 mem_reg_31__35_ ( .D(n3148), .CLK(clk), .Q(mem[1306]) );
  DFFPOSX1 mem_reg_31__34_ ( .D(n3147), .CLK(clk), .Q(mem[1305]) );
  DFFPOSX1 mem_reg_31__33_ ( .D(n3146), .CLK(clk), .Q(mem[1304]) );
  DFFPOSX1 mem_reg_31__32_ ( .D(n3145), .CLK(clk), .Q(mem[1303]) );
  DFFPOSX1 mem_reg_31__31_ ( .D(n3144), .CLK(clk), .Q(mem[1302]) );
  DFFPOSX1 mem_reg_31__30_ ( .D(n3143), .CLK(clk), .Q(mem[1301]) );
  DFFPOSX1 mem_reg_31__29_ ( .D(n3142), .CLK(clk), .Q(mem[1300]) );
  DFFPOSX1 mem_reg_31__28_ ( .D(n3141), .CLK(clk), .Q(mem[1299]) );
  DFFPOSX1 mem_reg_31__27_ ( .D(n3140), .CLK(clk), .Q(mem[1298]) );
  DFFPOSX1 mem_reg_31__26_ ( .D(n3139), .CLK(clk), .Q(mem[1297]) );
  DFFPOSX1 mem_reg_31__25_ ( .D(n3138), .CLK(clk), .Q(mem[1296]) );
  DFFPOSX1 mem_reg_31__24_ ( .D(n3137), .CLK(clk), .Q(mem[1295]) );
  DFFPOSX1 mem_reg_31__23_ ( .D(n3136), .CLK(clk), .Q(mem[1294]) );
  DFFPOSX1 mem_reg_31__22_ ( .D(n3135), .CLK(clk), .Q(mem[1293]) );
  DFFPOSX1 mem_reg_31__21_ ( .D(n3134), .CLK(clk), .Q(mem[1292]) );
  DFFPOSX1 mem_reg_31__20_ ( .D(n3133), .CLK(clk), .Q(mem[1291]) );
  DFFPOSX1 mem_reg_31__19_ ( .D(n3132), .CLK(clk), .Q(mem[1290]) );
  DFFPOSX1 mem_reg_31__18_ ( .D(n3131), .CLK(clk), .Q(mem[1289]) );
  DFFPOSX1 mem_reg_31__17_ ( .D(n3130), .CLK(clk), .Q(mem[1288]) );
  DFFPOSX1 mem_reg_31__16_ ( .D(n3129), .CLK(clk), .Q(mem[1287]) );
  DFFPOSX1 mem_reg_31__15_ ( .D(n3128), .CLK(clk), .Q(mem[1286]) );
  DFFPOSX1 mem_reg_31__14_ ( .D(n3127), .CLK(clk), .Q(mem[1285]) );
  DFFPOSX1 mem_reg_31__13_ ( .D(n3126), .CLK(clk), .Q(mem[1284]) );
  DFFPOSX1 mem_reg_31__12_ ( .D(n3125), .CLK(clk), .Q(mem[1283]) );
  DFFPOSX1 mem_reg_31__11_ ( .D(n3124), .CLK(clk), .Q(mem[1282]) );
  DFFPOSX1 mem_reg_31__10_ ( .D(n3123), .CLK(clk), .Q(mem[1281]) );
  DFFPOSX1 mem_reg_31__9_ ( .D(n3122), .CLK(clk), .Q(mem[1280]) );
  DFFPOSX1 mem_reg_31__8_ ( .D(n3121), .CLK(clk), .Q(mem[1279]) );
  DFFPOSX1 mem_reg_31__7_ ( .D(n3120), .CLK(clk), .Q(mem[1278]) );
  DFFPOSX1 mem_reg_31__6_ ( .D(n3119), .CLK(clk), .Q(mem[1277]) );
  DFFPOSX1 mem_reg_31__5_ ( .D(n3118), .CLK(clk), .Q(mem[1276]) );
  DFFPOSX1 mem_reg_31__4_ ( .D(n3117), .CLK(clk), .Q(mem[1275]) );
  DFFPOSX1 mem_reg_31__3_ ( .D(n3116), .CLK(clk), .Q(mem[1274]) );
  DFFPOSX1 mem_reg_31__2_ ( .D(n3115), .CLK(clk), .Q(mem[1273]) );
  DFFPOSX1 mem_reg_31__1_ ( .D(n3114), .CLK(clk), .Q(mem[1272]) );
  DFFPOSX1 mem_reg_31__0_ ( .D(n3113), .CLK(clk), .Q(mem[1271]) );
  DFFPOSX1 mem_reg_30__40_ ( .D(n3112), .CLK(clk), .Q(mem[1270]) );
  DFFPOSX1 mem_reg_30__39_ ( .D(n3111), .CLK(clk), .Q(mem[1269]) );
  DFFPOSX1 mem_reg_30__38_ ( .D(n3110), .CLK(clk), .Q(mem[1268]) );
  DFFPOSX1 mem_reg_30__37_ ( .D(n3109), .CLK(clk), .Q(mem[1267]) );
  DFFPOSX1 mem_reg_30__36_ ( .D(n3108), .CLK(clk), .Q(mem[1266]) );
  DFFPOSX1 mem_reg_30__35_ ( .D(n3107), .CLK(clk), .Q(mem[1265]) );
  DFFPOSX1 mem_reg_30__34_ ( .D(n3106), .CLK(clk), .Q(mem[1264]) );
  DFFPOSX1 mem_reg_30__33_ ( .D(n3105), .CLK(clk), .Q(mem[1263]) );
  DFFPOSX1 mem_reg_30__32_ ( .D(n3104), .CLK(clk), .Q(mem[1262]) );
  DFFPOSX1 mem_reg_30__31_ ( .D(n3103), .CLK(clk), .Q(mem[1261]) );
  DFFPOSX1 mem_reg_30__30_ ( .D(n3102), .CLK(clk), .Q(mem[1260]) );
  DFFPOSX1 mem_reg_30__29_ ( .D(n3101), .CLK(clk), .Q(mem[1259]) );
  DFFPOSX1 mem_reg_30__28_ ( .D(n3100), .CLK(clk), .Q(mem[1258]) );
  DFFPOSX1 mem_reg_30__27_ ( .D(n3099), .CLK(clk), .Q(mem[1257]) );
  DFFPOSX1 mem_reg_30__26_ ( .D(n3098), .CLK(clk), .Q(mem[1256]) );
  DFFPOSX1 mem_reg_30__25_ ( .D(n3097), .CLK(clk), .Q(mem[1255]) );
  DFFPOSX1 mem_reg_30__24_ ( .D(n3096), .CLK(clk), .Q(mem[1254]) );
  DFFPOSX1 mem_reg_30__23_ ( .D(n3095), .CLK(clk), .Q(mem[1253]) );
  DFFPOSX1 mem_reg_30__22_ ( .D(n3094), .CLK(clk), .Q(mem[1252]) );
  DFFPOSX1 mem_reg_30__21_ ( .D(n3093), .CLK(clk), .Q(mem[1251]) );
  DFFPOSX1 mem_reg_30__20_ ( .D(n3092), .CLK(clk), .Q(mem[1250]) );
  DFFPOSX1 mem_reg_30__19_ ( .D(n3091), .CLK(clk), .Q(mem[1249]) );
  DFFPOSX1 mem_reg_30__18_ ( .D(n3090), .CLK(clk), .Q(mem[1248]) );
  DFFPOSX1 mem_reg_30__17_ ( .D(n3089), .CLK(clk), .Q(mem[1247]) );
  DFFPOSX1 mem_reg_30__16_ ( .D(n3088), .CLK(clk), .Q(mem[1246]) );
  DFFPOSX1 mem_reg_30__15_ ( .D(n3087), .CLK(clk), .Q(mem[1245]) );
  DFFPOSX1 mem_reg_30__14_ ( .D(n3086), .CLK(clk), .Q(mem[1244]) );
  DFFPOSX1 mem_reg_30__13_ ( .D(n3085), .CLK(clk), .Q(mem[1243]) );
  DFFPOSX1 mem_reg_30__12_ ( .D(n3084), .CLK(clk), .Q(mem[1242]) );
  DFFPOSX1 mem_reg_30__11_ ( .D(n3083), .CLK(clk), .Q(mem[1241]) );
  DFFPOSX1 mem_reg_30__10_ ( .D(n3082), .CLK(clk), .Q(mem[1240]) );
  DFFPOSX1 mem_reg_30__9_ ( .D(n3081), .CLK(clk), .Q(mem[1239]) );
  DFFPOSX1 mem_reg_30__8_ ( .D(n3080), .CLK(clk), .Q(mem[1238]) );
  DFFPOSX1 mem_reg_30__7_ ( .D(n3079), .CLK(clk), .Q(mem[1237]) );
  DFFPOSX1 mem_reg_30__6_ ( .D(n3078), .CLK(clk), .Q(mem[1236]) );
  DFFPOSX1 mem_reg_30__5_ ( .D(n3077), .CLK(clk), .Q(mem[1235]) );
  DFFPOSX1 mem_reg_30__4_ ( .D(n3076), .CLK(clk), .Q(mem[1234]) );
  DFFPOSX1 mem_reg_30__3_ ( .D(n3075), .CLK(clk), .Q(mem[1233]) );
  DFFPOSX1 mem_reg_30__2_ ( .D(n3074), .CLK(clk), .Q(mem[1232]) );
  DFFPOSX1 mem_reg_30__1_ ( .D(n3073), .CLK(clk), .Q(mem[1231]) );
  DFFPOSX1 mem_reg_30__0_ ( .D(n3072), .CLK(clk), .Q(mem[1230]) );
  DFFPOSX1 mem_reg_29__40_ ( .D(n3071), .CLK(clk), .Q(mem[1229]) );
  DFFPOSX1 mem_reg_29__39_ ( .D(n3070), .CLK(clk), .Q(mem[1228]) );
  DFFPOSX1 mem_reg_29__38_ ( .D(n3069), .CLK(clk), .Q(mem[1227]) );
  DFFPOSX1 mem_reg_29__37_ ( .D(n3068), .CLK(clk), .Q(mem[1226]) );
  DFFPOSX1 mem_reg_29__36_ ( .D(n3067), .CLK(clk), .Q(mem[1225]) );
  DFFPOSX1 mem_reg_29__35_ ( .D(n3066), .CLK(clk), .Q(mem[1224]) );
  DFFPOSX1 mem_reg_29__34_ ( .D(n3065), .CLK(clk), .Q(mem[1223]) );
  DFFPOSX1 mem_reg_29__33_ ( .D(n3064), .CLK(clk), .Q(mem[1222]) );
  DFFPOSX1 mem_reg_29__32_ ( .D(n3063), .CLK(clk), .Q(mem[1221]) );
  DFFPOSX1 mem_reg_29__31_ ( .D(n3062), .CLK(clk), .Q(mem[1220]) );
  DFFPOSX1 mem_reg_29__30_ ( .D(n3061), .CLK(clk), .Q(mem[1219]) );
  DFFPOSX1 mem_reg_29__29_ ( .D(n3060), .CLK(clk), .Q(mem[1218]) );
  DFFPOSX1 mem_reg_29__28_ ( .D(n3059), .CLK(clk), .Q(mem[1217]) );
  DFFPOSX1 mem_reg_29__27_ ( .D(n3058), .CLK(clk), .Q(mem[1216]) );
  DFFPOSX1 mem_reg_29__26_ ( .D(n3057), .CLK(clk), .Q(mem[1215]) );
  DFFPOSX1 mem_reg_29__25_ ( .D(n3056), .CLK(clk), .Q(mem[1214]) );
  DFFPOSX1 mem_reg_29__24_ ( .D(n3055), .CLK(clk), .Q(mem[1213]) );
  DFFPOSX1 mem_reg_29__23_ ( .D(n3054), .CLK(clk), .Q(mem[1212]) );
  DFFPOSX1 mem_reg_29__22_ ( .D(n3053), .CLK(clk), .Q(mem[1211]) );
  DFFPOSX1 mem_reg_29__21_ ( .D(n3052), .CLK(clk), .Q(mem[1210]) );
  DFFPOSX1 mem_reg_29__20_ ( .D(n3051), .CLK(clk), .Q(mem[1209]) );
  DFFPOSX1 mem_reg_29__19_ ( .D(n3050), .CLK(clk), .Q(mem[1208]) );
  DFFPOSX1 mem_reg_29__18_ ( .D(n3049), .CLK(clk), .Q(mem[1207]) );
  DFFPOSX1 mem_reg_29__17_ ( .D(n3048), .CLK(clk), .Q(mem[1206]) );
  DFFPOSX1 mem_reg_29__16_ ( .D(n3047), .CLK(clk), .Q(mem[1205]) );
  DFFPOSX1 mem_reg_29__15_ ( .D(n3046), .CLK(clk), .Q(mem[1204]) );
  DFFPOSX1 mem_reg_29__14_ ( .D(n3045), .CLK(clk), .Q(mem[1203]) );
  DFFPOSX1 mem_reg_29__13_ ( .D(n3044), .CLK(clk), .Q(mem[1202]) );
  DFFPOSX1 mem_reg_29__12_ ( .D(n3043), .CLK(clk), .Q(mem[1201]) );
  DFFPOSX1 mem_reg_29__11_ ( .D(n3042), .CLK(clk), .Q(mem[1200]) );
  DFFPOSX1 mem_reg_29__10_ ( .D(n3041), .CLK(clk), .Q(mem[1199]) );
  DFFPOSX1 mem_reg_29__9_ ( .D(n3040), .CLK(clk), .Q(mem[1198]) );
  DFFPOSX1 mem_reg_29__8_ ( .D(n3039), .CLK(clk), .Q(mem[1197]) );
  DFFPOSX1 mem_reg_29__7_ ( .D(n3038), .CLK(clk), .Q(mem[1196]) );
  DFFPOSX1 mem_reg_29__6_ ( .D(n3037), .CLK(clk), .Q(mem[1195]) );
  DFFPOSX1 mem_reg_29__5_ ( .D(n3036), .CLK(clk), .Q(mem[1194]) );
  DFFPOSX1 mem_reg_29__4_ ( .D(n3035), .CLK(clk), .Q(mem[1193]) );
  DFFPOSX1 mem_reg_29__3_ ( .D(n3034), .CLK(clk), .Q(mem[1192]) );
  DFFPOSX1 mem_reg_29__2_ ( .D(n3033), .CLK(clk), .Q(mem[1191]) );
  DFFPOSX1 mem_reg_29__1_ ( .D(n3032), .CLK(clk), .Q(mem[1190]) );
  DFFPOSX1 mem_reg_29__0_ ( .D(n3031), .CLK(clk), .Q(mem[1189]) );
  DFFPOSX1 mem_reg_28__40_ ( .D(n3030), .CLK(clk), .Q(mem[1188]) );
  DFFPOSX1 mem_reg_28__39_ ( .D(n3029), .CLK(clk), .Q(mem[1187]) );
  DFFPOSX1 mem_reg_28__38_ ( .D(n3028), .CLK(clk), .Q(mem[1186]) );
  DFFPOSX1 mem_reg_28__37_ ( .D(n3027), .CLK(clk), .Q(mem[1185]) );
  DFFPOSX1 mem_reg_28__36_ ( .D(n3026), .CLK(clk), .Q(mem[1184]) );
  DFFPOSX1 mem_reg_28__35_ ( .D(n3025), .CLK(clk), .Q(mem[1183]) );
  DFFPOSX1 mem_reg_28__34_ ( .D(n3024), .CLK(clk), .Q(mem[1182]) );
  DFFPOSX1 mem_reg_28__33_ ( .D(n3023), .CLK(clk), .Q(mem[1181]) );
  DFFPOSX1 mem_reg_28__32_ ( .D(n3022), .CLK(clk), .Q(mem[1180]) );
  DFFPOSX1 mem_reg_28__31_ ( .D(n3021), .CLK(clk), .Q(mem[1179]) );
  DFFPOSX1 mem_reg_28__30_ ( .D(n3020), .CLK(clk), .Q(mem[1178]) );
  DFFPOSX1 mem_reg_28__29_ ( .D(n3019), .CLK(clk), .Q(mem[1177]) );
  DFFPOSX1 mem_reg_28__28_ ( .D(n3018), .CLK(clk), .Q(mem[1176]) );
  DFFPOSX1 mem_reg_28__27_ ( .D(n3017), .CLK(clk), .Q(mem[1175]) );
  DFFPOSX1 mem_reg_28__26_ ( .D(n3016), .CLK(clk), .Q(mem[1174]) );
  DFFPOSX1 mem_reg_28__25_ ( .D(n3015), .CLK(clk), .Q(mem[1173]) );
  DFFPOSX1 mem_reg_28__24_ ( .D(n3014), .CLK(clk), .Q(mem[1172]) );
  DFFPOSX1 mem_reg_28__23_ ( .D(n3013), .CLK(clk), .Q(mem[1171]) );
  DFFPOSX1 mem_reg_28__22_ ( .D(n3012), .CLK(clk), .Q(mem[1170]) );
  DFFPOSX1 mem_reg_28__21_ ( .D(n3011), .CLK(clk), .Q(mem[1169]) );
  DFFPOSX1 mem_reg_28__20_ ( .D(n3010), .CLK(clk), .Q(mem[1168]) );
  DFFPOSX1 mem_reg_28__19_ ( .D(n3009), .CLK(clk), .Q(mem[1167]) );
  DFFPOSX1 mem_reg_28__18_ ( .D(n3008), .CLK(clk), .Q(mem[1166]) );
  DFFPOSX1 mem_reg_28__17_ ( .D(n3007), .CLK(clk), .Q(mem[1165]) );
  DFFPOSX1 mem_reg_28__16_ ( .D(n3006), .CLK(clk), .Q(mem[1164]) );
  DFFPOSX1 mem_reg_28__15_ ( .D(n3005), .CLK(clk), .Q(mem[1163]) );
  DFFPOSX1 mem_reg_28__14_ ( .D(n3004), .CLK(clk), .Q(mem[1162]) );
  DFFPOSX1 mem_reg_28__13_ ( .D(n3003), .CLK(clk), .Q(mem[1161]) );
  DFFPOSX1 mem_reg_28__12_ ( .D(n3002), .CLK(clk), .Q(mem[1160]) );
  DFFPOSX1 mem_reg_28__11_ ( .D(n3001), .CLK(clk), .Q(mem[1159]) );
  DFFPOSX1 mem_reg_28__10_ ( .D(n3000), .CLK(clk), .Q(mem[1158]) );
  DFFPOSX1 mem_reg_28__9_ ( .D(n2999), .CLK(clk), .Q(mem[1157]) );
  DFFPOSX1 mem_reg_28__8_ ( .D(n2998), .CLK(clk), .Q(mem[1156]) );
  DFFPOSX1 mem_reg_28__7_ ( .D(n2997), .CLK(clk), .Q(mem[1155]) );
  DFFPOSX1 mem_reg_28__6_ ( .D(n2996), .CLK(clk), .Q(mem[1154]) );
  DFFPOSX1 mem_reg_28__5_ ( .D(n2995), .CLK(clk), .Q(mem[1153]) );
  DFFPOSX1 mem_reg_28__4_ ( .D(n2994), .CLK(clk), .Q(mem[1152]) );
  DFFPOSX1 mem_reg_28__3_ ( .D(n2993), .CLK(clk), .Q(mem[1151]) );
  DFFPOSX1 mem_reg_28__2_ ( .D(n2992), .CLK(clk), .Q(mem[1150]) );
  DFFPOSX1 mem_reg_28__1_ ( .D(n2991), .CLK(clk), .Q(mem[1149]) );
  DFFPOSX1 mem_reg_28__0_ ( .D(n2990), .CLK(clk), .Q(mem[1148]) );
  DFFPOSX1 mem_reg_27__40_ ( .D(n2989), .CLK(clk), .Q(mem[1147]) );
  DFFPOSX1 mem_reg_27__39_ ( .D(n2988), .CLK(clk), .Q(mem[1146]) );
  DFFPOSX1 mem_reg_27__38_ ( .D(n2987), .CLK(clk), .Q(mem[1145]) );
  DFFPOSX1 mem_reg_27__37_ ( .D(n2986), .CLK(clk), .Q(mem[1144]) );
  DFFPOSX1 mem_reg_27__36_ ( .D(n2985), .CLK(clk), .Q(mem[1143]) );
  DFFPOSX1 mem_reg_27__35_ ( .D(n2984), .CLK(clk), .Q(mem[1142]) );
  DFFPOSX1 mem_reg_27__34_ ( .D(n2983), .CLK(clk), .Q(mem[1141]) );
  DFFPOSX1 mem_reg_27__33_ ( .D(n2982), .CLK(clk), .Q(mem[1140]) );
  DFFPOSX1 mem_reg_27__32_ ( .D(n2981), .CLK(clk), .Q(mem[1139]) );
  DFFPOSX1 mem_reg_27__31_ ( .D(n2980), .CLK(clk), .Q(mem[1138]) );
  DFFPOSX1 mem_reg_27__30_ ( .D(n2979), .CLK(clk), .Q(mem[1137]) );
  DFFPOSX1 mem_reg_27__29_ ( .D(n2978), .CLK(clk), .Q(mem[1136]) );
  DFFPOSX1 mem_reg_27__28_ ( .D(n2977), .CLK(clk), .Q(mem[1135]) );
  DFFPOSX1 mem_reg_27__27_ ( .D(n2976), .CLK(clk), .Q(mem[1134]) );
  DFFPOSX1 mem_reg_27__26_ ( .D(n2975), .CLK(clk), .Q(mem[1133]) );
  DFFPOSX1 mem_reg_27__25_ ( .D(n2974), .CLK(clk), .Q(mem[1132]) );
  DFFPOSX1 mem_reg_27__24_ ( .D(n2973), .CLK(clk), .Q(mem[1131]) );
  DFFPOSX1 mem_reg_27__23_ ( .D(n2972), .CLK(clk), .Q(mem[1130]) );
  DFFPOSX1 mem_reg_27__22_ ( .D(n2971), .CLK(clk), .Q(mem[1129]) );
  DFFPOSX1 mem_reg_27__21_ ( .D(n2970), .CLK(clk), .Q(mem[1128]) );
  DFFPOSX1 mem_reg_27__20_ ( .D(n2969), .CLK(clk), .Q(mem[1127]) );
  DFFPOSX1 mem_reg_27__19_ ( .D(n2968), .CLK(clk), .Q(mem[1126]) );
  DFFPOSX1 mem_reg_27__18_ ( .D(n2967), .CLK(clk), .Q(mem[1125]) );
  DFFPOSX1 mem_reg_27__17_ ( .D(n2966), .CLK(clk), .Q(mem[1124]) );
  DFFPOSX1 mem_reg_27__16_ ( .D(n2965), .CLK(clk), .Q(mem[1123]) );
  DFFPOSX1 mem_reg_27__15_ ( .D(n2964), .CLK(clk), .Q(mem[1122]) );
  DFFPOSX1 mem_reg_27__14_ ( .D(n2963), .CLK(clk), .Q(mem[1121]) );
  DFFPOSX1 mem_reg_27__13_ ( .D(n2962), .CLK(clk), .Q(mem[1120]) );
  DFFPOSX1 mem_reg_27__12_ ( .D(n2961), .CLK(clk), .Q(mem[1119]) );
  DFFPOSX1 mem_reg_27__11_ ( .D(n2960), .CLK(clk), .Q(mem[1118]) );
  DFFPOSX1 mem_reg_27__10_ ( .D(n2959), .CLK(clk), .Q(mem[1117]) );
  DFFPOSX1 mem_reg_27__9_ ( .D(n2958), .CLK(clk), .Q(mem[1116]) );
  DFFPOSX1 mem_reg_27__8_ ( .D(n2957), .CLK(clk), .Q(mem[1115]) );
  DFFPOSX1 mem_reg_27__7_ ( .D(n2956), .CLK(clk), .Q(mem[1114]) );
  DFFPOSX1 mem_reg_27__6_ ( .D(n2955), .CLK(clk), .Q(mem[1113]) );
  DFFPOSX1 mem_reg_27__5_ ( .D(n2954), .CLK(clk), .Q(mem[1112]) );
  DFFPOSX1 mem_reg_27__4_ ( .D(n2953), .CLK(clk), .Q(mem[1111]) );
  DFFPOSX1 mem_reg_27__3_ ( .D(n2952), .CLK(clk), .Q(mem[1110]) );
  DFFPOSX1 mem_reg_27__2_ ( .D(n2951), .CLK(clk), .Q(mem[1109]) );
  DFFPOSX1 mem_reg_27__1_ ( .D(n2950), .CLK(clk), .Q(mem[1108]) );
  DFFPOSX1 mem_reg_27__0_ ( .D(n2949), .CLK(clk), .Q(mem[1107]) );
  DFFPOSX1 mem_reg_26__40_ ( .D(n2948), .CLK(clk), .Q(mem[1106]) );
  DFFPOSX1 mem_reg_26__39_ ( .D(n2947), .CLK(clk), .Q(mem[1105]) );
  DFFPOSX1 mem_reg_26__38_ ( .D(n2946), .CLK(clk), .Q(mem[1104]) );
  DFFPOSX1 mem_reg_26__37_ ( .D(n2945), .CLK(clk), .Q(mem[1103]) );
  DFFPOSX1 mem_reg_26__36_ ( .D(n2944), .CLK(clk), .Q(mem[1102]) );
  DFFPOSX1 mem_reg_26__35_ ( .D(n2943), .CLK(clk), .Q(mem[1101]) );
  DFFPOSX1 mem_reg_26__34_ ( .D(n2942), .CLK(clk), .Q(mem[1100]) );
  DFFPOSX1 mem_reg_26__33_ ( .D(n2941), .CLK(clk), .Q(mem[1099]) );
  DFFPOSX1 mem_reg_26__32_ ( .D(n2940), .CLK(clk), .Q(mem[1098]) );
  DFFPOSX1 mem_reg_26__31_ ( .D(n2939), .CLK(clk), .Q(mem[1097]) );
  DFFPOSX1 mem_reg_26__30_ ( .D(n2938), .CLK(clk), .Q(mem[1096]) );
  DFFPOSX1 mem_reg_26__29_ ( .D(n2937), .CLK(clk), .Q(mem[1095]) );
  DFFPOSX1 mem_reg_26__28_ ( .D(n2936), .CLK(clk), .Q(mem[1094]) );
  DFFPOSX1 mem_reg_26__27_ ( .D(n2935), .CLK(clk), .Q(mem[1093]) );
  DFFPOSX1 mem_reg_26__26_ ( .D(n2934), .CLK(clk), .Q(mem[1092]) );
  DFFPOSX1 mem_reg_26__25_ ( .D(n2933), .CLK(clk), .Q(mem[1091]) );
  DFFPOSX1 mem_reg_26__24_ ( .D(n2932), .CLK(clk), .Q(mem[1090]) );
  DFFPOSX1 mem_reg_26__23_ ( .D(n2931), .CLK(clk), .Q(mem[1089]) );
  DFFPOSX1 mem_reg_26__22_ ( .D(n2930), .CLK(clk), .Q(mem[1088]) );
  DFFPOSX1 mem_reg_26__21_ ( .D(n2929), .CLK(clk), .Q(mem[1087]) );
  DFFPOSX1 mem_reg_26__20_ ( .D(n2928), .CLK(clk), .Q(mem[1086]) );
  DFFPOSX1 mem_reg_26__19_ ( .D(n2927), .CLK(clk), .Q(mem[1085]) );
  DFFPOSX1 mem_reg_26__18_ ( .D(n2926), .CLK(clk), .Q(mem[1084]) );
  DFFPOSX1 mem_reg_26__17_ ( .D(n2925), .CLK(clk), .Q(mem[1083]) );
  DFFPOSX1 mem_reg_26__16_ ( .D(n2924), .CLK(clk), .Q(mem[1082]) );
  DFFPOSX1 mem_reg_26__15_ ( .D(n2923), .CLK(clk), .Q(mem[1081]) );
  DFFPOSX1 mem_reg_26__14_ ( .D(n2922), .CLK(clk), .Q(mem[1080]) );
  DFFPOSX1 mem_reg_26__13_ ( .D(n2921), .CLK(clk), .Q(mem[1079]) );
  DFFPOSX1 mem_reg_26__12_ ( .D(n2920), .CLK(clk), .Q(mem[1078]) );
  DFFPOSX1 mem_reg_26__11_ ( .D(n2919), .CLK(clk), .Q(mem[1077]) );
  DFFPOSX1 mem_reg_26__10_ ( .D(n2918), .CLK(clk), .Q(mem[1076]) );
  DFFPOSX1 mem_reg_26__9_ ( .D(n2917), .CLK(clk), .Q(mem[1075]) );
  DFFPOSX1 mem_reg_26__8_ ( .D(n2916), .CLK(clk), .Q(mem[1074]) );
  DFFPOSX1 mem_reg_26__7_ ( .D(n2915), .CLK(clk), .Q(mem[1073]) );
  DFFPOSX1 mem_reg_26__6_ ( .D(n2914), .CLK(clk), .Q(mem[1072]) );
  DFFPOSX1 mem_reg_26__5_ ( .D(n2913), .CLK(clk), .Q(mem[1071]) );
  DFFPOSX1 mem_reg_26__4_ ( .D(n2912), .CLK(clk), .Q(mem[1070]) );
  DFFPOSX1 mem_reg_26__3_ ( .D(n2911), .CLK(clk), .Q(mem[1069]) );
  DFFPOSX1 mem_reg_26__2_ ( .D(n2910), .CLK(clk), .Q(mem[1068]) );
  DFFPOSX1 mem_reg_26__1_ ( .D(n2909), .CLK(clk), .Q(mem[1067]) );
  DFFPOSX1 mem_reg_26__0_ ( .D(n2908), .CLK(clk), .Q(mem[1066]) );
  DFFPOSX1 mem_reg_25__40_ ( .D(n2907), .CLK(clk), .Q(mem[1065]) );
  DFFPOSX1 mem_reg_25__39_ ( .D(n2906), .CLK(clk), .Q(mem[1064]) );
  DFFPOSX1 mem_reg_25__38_ ( .D(n2905), .CLK(clk), .Q(mem[1063]) );
  DFFPOSX1 mem_reg_25__37_ ( .D(n2904), .CLK(clk), .Q(mem[1062]) );
  DFFPOSX1 mem_reg_25__36_ ( .D(n2903), .CLK(clk), .Q(mem[1061]) );
  DFFPOSX1 mem_reg_25__35_ ( .D(n2902), .CLK(clk), .Q(mem[1060]) );
  DFFPOSX1 mem_reg_25__34_ ( .D(n2901), .CLK(clk), .Q(mem[1059]) );
  DFFPOSX1 mem_reg_25__33_ ( .D(n2900), .CLK(clk), .Q(mem[1058]) );
  DFFPOSX1 mem_reg_25__32_ ( .D(n2899), .CLK(clk), .Q(mem[1057]) );
  DFFPOSX1 mem_reg_25__31_ ( .D(n2898), .CLK(clk), .Q(mem[1056]) );
  DFFPOSX1 mem_reg_25__30_ ( .D(n2897), .CLK(clk), .Q(mem[1055]) );
  DFFPOSX1 mem_reg_25__29_ ( .D(n2896), .CLK(clk), .Q(mem[1054]) );
  DFFPOSX1 mem_reg_25__28_ ( .D(n2895), .CLK(clk), .Q(mem[1053]) );
  DFFPOSX1 mem_reg_25__27_ ( .D(n2894), .CLK(clk), .Q(mem[1052]) );
  DFFPOSX1 mem_reg_25__26_ ( .D(n2893), .CLK(clk), .Q(mem[1051]) );
  DFFPOSX1 mem_reg_25__25_ ( .D(n2892), .CLK(clk), .Q(mem[1050]) );
  DFFPOSX1 mem_reg_25__24_ ( .D(n2891), .CLK(clk), .Q(mem[1049]) );
  DFFPOSX1 mem_reg_25__23_ ( .D(n2890), .CLK(clk), .Q(mem[1048]) );
  DFFPOSX1 mem_reg_25__22_ ( .D(n2889), .CLK(clk), .Q(mem[1047]) );
  DFFPOSX1 mem_reg_25__21_ ( .D(n2888), .CLK(clk), .Q(mem[1046]) );
  DFFPOSX1 mem_reg_25__20_ ( .D(n2887), .CLK(clk), .Q(mem[1045]) );
  DFFPOSX1 mem_reg_25__19_ ( .D(n2886), .CLK(clk), .Q(mem[1044]) );
  DFFPOSX1 mem_reg_25__18_ ( .D(n2885), .CLK(clk), .Q(mem[1043]) );
  DFFPOSX1 mem_reg_25__17_ ( .D(n2884), .CLK(clk), .Q(mem[1042]) );
  DFFPOSX1 mem_reg_25__16_ ( .D(n2883), .CLK(clk), .Q(mem[1041]) );
  DFFPOSX1 mem_reg_25__15_ ( .D(n2882), .CLK(clk), .Q(mem[1040]) );
  DFFPOSX1 mem_reg_25__14_ ( .D(n2881), .CLK(clk), .Q(mem[1039]) );
  DFFPOSX1 mem_reg_25__13_ ( .D(n2880), .CLK(clk), .Q(mem[1038]) );
  DFFPOSX1 mem_reg_25__12_ ( .D(n2879), .CLK(clk), .Q(mem[1037]) );
  DFFPOSX1 mem_reg_25__11_ ( .D(n2878), .CLK(clk), .Q(mem[1036]) );
  DFFPOSX1 mem_reg_25__10_ ( .D(n2877), .CLK(clk), .Q(mem[1035]) );
  DFFPOSX1 mem_reg_25__9_ ( .D(n2876), .CLK(clk), .Q(mem[1034]) );
  DFFPOSX1 mem_reg_25__8_ ( .D(n2875), .CLK(clk), .Q(mem[1033]) );
  DFFPOSX1 mem_reg_25__7_ ( .D(n2874), .CLK(clk), .Q(mem[1032]) );
  DFFPOSX1 mem_reg_25__6_ ( .D(n2873), .CLK(clk), .Q(mem[1031]) );
  DFFPOSX1 mem_reg_25__5_ ( .D(n2872), .CLK(clk), .Q(mem[1030]) );
  DFFPOSX1 mem_reg_25__4_ ( .D(n2871), .CLK(clk), .Q(mem[1029]) );
  DFFPOSX1 mem_reg_25__3_ ( .D(n2870), .CLK(clk), .Q(mem[1028]) );
  DFFPOSX1 mem_reg_25__2_ ( .D(n2869), .CLK(clk), .Q(mem[1027]) );
  DFFPOSX1 mem_reg_25__1_ ( .D(n2868), .CLK(clk), .Q(mem[1026]) );
  DFFPOSX1 mem_reg_25__0_ ( .D(n2867), .CLK(clk), .Q(mem[1025]) );
  DFFPOSX1 mem_reg_24__40_ ( .D(n2866), .CLK(clk), .Q(mem[1024]) );
  DFFPOSX1 mem_reg_24__39_ ( .D(n2865), .CLK(clk), .Q(mem[1023]) );
  DFFPOSX1 mem_reg_24__38_ ( .D(n2864), .CLK(clk), .Q(mem[1022]) );
  DFFPOSX1 mem_reg_24__37_ ( .D(n2863), .CLK(clk), .Q(mem[1021]) );
  DFFPOSX1 mem_reg_24__36_ ( .D(n2862), .CLK(clk), .Q(mem[1020]) );
  DFFPOSX1 mem_reg_24__35_ ( .D(n2861), .CLK(clk), .Q(mem[1019]) );
  DFFPOSX1 mem_reg_24__34_ ( .D(n2860), .CLK(clk), .Q(mem[1018]) );
  DFFPOSX1 mem_reg_24__33_ ( .D(n2859), .CLK(clk), .Q(mem[1017]) );
  DFFPOSX1 mem_reg_24__32_ ( .D(n2858), .CLK(clk), .Q(mem[1016]) );
  DFFPOSX1 mem_reg_24__31_ ( .D(n2857), .CLK(clk), .Q(mem[1015]) );
  DFFPOSX1 mem_reg_24__30_ ( .D(n2856), .CLK(clk), .Q(mem[1014]) );
  DFFPOSX1 mem_reg_24__29_ ( .D(n2855), .CLK(clk), .Q(mem[1013]) );
  DFFPOSX1 mem_reg_24__28_ ( .D(n2854), .CLK(clk), .Q(mem[1012]) );
  DFFPOSX1 mem_reg_24__27_ ( .D(n2853), .CLK(clk), .Q(mem[1011]) );
  DFFPOSX1 mem_reg_24__26_ ( .D(n2852), .CLK(clk), .Q(mem[1010]) );
  DFFPOSX1 mem_reg_24__25_ ( .D(n2851), .CLK(clk), .Q(mem[1009]) );
  DFFPOSX1 mem_reg_24__24_ ( .D(n2850), .CLK(clk), .Q(mem[1008]) );
  DFFPOSX1 mem_reg_24__23_ ( .D(n2849), .CLK(clk), .Q(mem[1007]) );
  DFFPOSX1 mem_reg_24__22_ ( .D(n2848), .CLK(clk), .Q(mem[1006]) );
  DFFPOSX1 mem_reg_24__21_ ( .D(n2847), .CLK(clk), .Q(mem[1005]) );
  DFFPOSX1 mem_reg_24__20_ ( .D(n2846), .CLK(clk), .Q(mem[1004]) );
  DFFPOSX1 mem_reg_24__19_ ( .D(n2845), .CLK(clk), .Q(mem[1003]) );
  DFFPOSX1 mem_reg_24__18_ ( .D(n2844), .CLK(clk), .Q(mem[1002]) );
  DFFPOSX1 mem_reg_24__17_ ( .D(n2843), .CLK(clk), .Q(mem[1001]) );
  DFFPOSX1 mem_reg_24__16_ ( .D(n2842), .CLK(clk), .Q(mem[1000]) );
  DFFPOSX1 mem_reg_24__15_ ( .D(n2841), .CLK(clk), .Q(mem[999]) );
  DFFPOSX1 mem_reg_24__14_ ( .D(n2840), .CLK(clk), .Q(mem[998]) );
  DFFPOSX1 mem_reg_24__13_ ( .D(n2839), .CLK(clk), .Q(mem[997]) );
  DFFPOSX1 mem_reg_24__12_ ( .D(n2838), .CLK(clk), .Q(mem[996]) );
  DFFPOSX1 mem_reg_24__11_ ( .D(n2837), .CLK(clk), .Q(mem[995]) );
  DFFPOSX1 mem_reg_24__10_ ( .D(n2836), .CLK(clk), .Q(mem[994]) );
  DFFPOSX1 mem_reg_24__9_ ( .D(n2835), .CLK(clk), .Q(mem[993]) );
  DFFPOSX1 mem_reg_24__8_ ( .D(n2834), .CLK(clk), .Q(mem[992]) );
  DFFPOSX1 mem_reg_24__7_ ( .D(n2833), .CLK(clk), .Q(mem[991]) );
  DFFPOSX1 mem_reg_24__6_ ( .D(n2832), .CLK(clk), .Q(mem[990]) );
  DFFPOSX1 mem_reg_24__5_ ( .D(n2831), .CLK(clk), .Q(mem[989]) );
  DFFPOSX1 mem_reg_24__4_ ( .D(n2830), .CLK(clk), .Q(mem[988]) );
  DFFPOSX1 mem_reg_24__3_ ( .D(n2829), .CLK(clk), .Q(mem[987]) );
  DFFPOSX1 mem_reg_24__2_ ( .D(n2828), .CLK(clk), .Q(mem[986]) );
  DFFPOSX1 mem_reg_24__1_ ( .D(n2827), .CLK(clk), .Q(mem[985]) );
  DFFPOSX1 mem_reg_24__0_ ( .D(n2826), .CLK(clk), .Q(mem[984]) );
  DFFPOSX1 mem_reg_23__40_ ( .D(n2825), .CLK(clk), .Q(mem[983]) );
  DFFPOSX1 mem_reg_23__39_ ( .D(n2824), .CLK(clk), .Q(mem[982]) );
  DFFPOSX1 mem_reg_23__38_ ( .D(n2823), .CLK(clk), .Q(mem[981]) );
  DFFPOSX1 mem_reg_23__37_ ( .D(n2822), .CLK(clk), .Q(mem[980]) );
  DFFPOSX1 mem_reg_23__36_ ( .D(n2821), .CLK(clk), .Q(mem[979]) );
  DFFPOSX1 mem_reg_23__35_ ( .D(n2820), .CLK(clk), .Q(mem[978]) );
  DFFPOSX1 mem_reg_23__34_ ( .D(n2819), .CLK(clk), .Q(mem[977]) );
  DFFPOSX1 mem_reg_23__33_ ( .D(n2818), .CLK(clk), .Q(mem[976]) );
  DFFPOSX1 mem_reg_23__32_ ( .D(n2817), .CLK(clk), .Q(mem[975]) );
  DFFPOSX1 mem_reg_23__31_ ( .D(n2816), .CLK(clk), .Q(mem[974]) );
  DFFPOSX1 mem_reg_23__30_ ( .D(n2815), .CLK(clk), .Q(mem[973]) );
  DFFPOSX1 mem_reg_23__29_ ( .D(n2814), .CLK(clk), .Q(mem[972]) );
  DFFPOSX1 mem_reg_23__28_ ( .D(n2813), .CLK(clk), .Q(mem[971]) );
  DFFPOSX1 mem_reg_23__27_ ( .D(n2812), .CLK(clk), .Q(mem[970]) );
  DFFPOSX1 mem_reg_23__26_ ( .D(n2811), .CLK(clk), .Q(mem[969]) );
  DFFPOSX1 mem_reg_23__25_ ( .D(n2810), .CLK(clk), .Q(mem[968]) );
  DFFPOSX1 mem_reg_23__24_ ( .D(n2809), .CLK(clk), .Q(mem[967]) );
  DFFPOSX1 mem_reg_23__23_ ( .D(n2808), .CLK(clk), .Q(mem[966]) );
  DFFPOSX1 mem_reg_23__22_ ( .D(n2807), .CLK(clk), .Q(mem[965]) );
  DFFPOSX1 mem_reg_23__21_ ( .D(n2806), .CLK(clk), .Q(mem[964]) );
  DFFPOSX1 mem_reg_23__20_ ( .D(n2805), .CLK(clk), .Q(mem[963]) );
  DFFPOSX1 mem_reg_23__19_ ( .D(n2804), .CLK(clk), .Q(mem[962]) );
  DFFPOSX1 mem_reg_23__18_ ( .D(n2803), .CLK(clk), .Q(mem[961]) );
  DFFPOSX1 mem_reg_23__17_ ( .D(n2802), .CLK(clk), .Q(mem[960]) );
  DFFPOSX1 mem_reg_23__16_ ( .D(n2801), .CLK(clk), .Q(mem[959]) );
  DFFPOSX1 mem_reg_23__15_ ( .D(n2800), .CLK(clk), .Q(mem[958]) );
  DFFPOSX1 mem_reg_23__14_ ( .D(n2799), .CLK(clk), .Q(mem[957]) );
  DFFPOSX1 mem_reg_23__13_ ( .D(n2798), .CLK(clk), .Q(mem[956]) );
  DFFPOSX1 mem_reg_23__12_ ( .D(n2797), .CLK(clk), .Q(mem[955]) );
  DFFPOSX1 mem_reg_23__11_ ( .D(n2796), .CLK(clk), .Q(mem[954]) );
  DFFPOSX1 mem_reg_23__10_ ( .D(n2795), .CLK(clk), .Q(mem[953]) );
  DFFPOSX1 mem_reg_23__9_ ( .D(n2794), .CLK(clk), .Q(mem[952]) );
  DFFPOSX1 mem_reg_23__8_ ( .D(n2793), .CLK(clk), .Q(mem[951]) );
  DFFPOSX1 mem_reg_23__7_ ( .D(n2792), .CLK(clk), .Q(mem[950]) );
  DFFPOSX1 mem_reg_23__6_ ( .D(n2791), .CLK(clk), .Q(mem[949]) );
  DFFPOSX1 mem_reg_23__5_ ( .D(n2790), .CLK(clk), .Q(mem[948]) );
  DFFPOSX1 mem_reg_23__4_ ( .D(n2789), .CLK(clk), .Q(mem[947]) );
  DFFPOSX1 mem_reg_23__3_ ( .D(n2788), .CLK(clk), .Q(mem[946]) );
  DFFPOSX1 mem_reg_23__2_ ( .D(n2787), .CLK(clk), .Q(mem[945]) );
  DFFPOSX1 mem_reg_23__1_ ( .D(n2786), .CLK(clk), .Q(mem[944]) );
  DFFPOSX1 mem_reg_23__0_ ( .D(n2785), .CLK(clk), .Q(mem[943]) );
  DFFPOSX1 mem_reg_22__40_ ( .D(n2784), .CLK(clk), .Q(mem[942]) );
  DFFPOSX1 mem_reg_22__39_ ( .D(n2783), .CLK(clk), .Q(mem[941]) );
  DFFPOSX1 mem_reg_22__38_ ( .D(n2782), .CLK(clk), .Q(mem[940]) );
  DFFPOSX1 mem_reg_22__37_ ( .D(n2781), .CLK(clk), .Q(mem[939]) );
  DFFPOSX1 mem_reg_22__36_ ( .D(n2780), .CLK(clk), .Q(mem[938]) );
  DFFPOSX1 mem_reg_22__35_ ( .D(n2779), .CLK(clk), .Q(mem[937]) );
  DFFPOSX1 mem_reg_22__34_ ( .D(n2778), .CLK(clk), .Q(mem[936]) );
  DFFPOSX1 mem_reg_22__33_ ( .D(n2777), .CLK(clk), .Q(mem[935]) );
  DFFPOSX1 mem_reg_22__32_ ( .D(n2776), .CLK(clk), .Q(mem[934]) );
  DFFPOSX1 mem_reg_22__31_ ( .D(n2775), .CLK(clk), .Q(mem[933]) );
  DFFPOSX1 mem_reg_22__30_ ( .D(n2774), .CLK(clk), .Q(mem[932]) );
  DFFPOSX1 mem_reg_22__29_ ( .D(n2773), .CLK(clk), .Q(mem[931]) );
  DFFPOSX1 mem_reg_22__28_ ( .D(n2772), .CLK(clk), .Q(mem[930]) );
  DFFPOSX1 mem_reg_22__27_ ( .D(n2771), .CLK(clk), .Q(mem[929]) );
  DFFPOSX1 mem_reg_22__26_ ( .D(n2770), .CLK(clk), .Q(mem[928]) );
  DFFPOSX1 mem_reg_22__25_ ( .D(n2769), .CLK(clk), .Q(mem[927]) );
  DFFPOSX1 mem_reg_22__24_ ( .D(n2768), .CLK(clk), .Q(mem[926]) );
  DFFPOSX1 mem_reg_22__23_ ( .D(n2767), .CLK(clk), .Q(mem[925]) );
  DFFPOSX1 mem_reg_22__22_ ( .D(n2766), .CLK(clk), .Q(mem[924]) );
  DFFPOSX1 mem_reg_22__21_ ( .D(n2765), .CLK(clk), .Q(mem[923]) );
  DFFPOSX1 mem_reg_22__20_ ( .D(n2764), .CLK(clk), .Q(mem[922]) );
  DFFPOSX1 mem_reg_22__19_ ( .D(n2763), .CLK(clk), .Q(mem[921]) );
  DFFPOSX1 mem_reg_22__18_ ( .D(n2762), .CLK(clk), .Q(mem[920]) );
  DFFPOSX1 mem_reg_22__17_ ( .D(n2761), .CLK(clk), .Q(mem[919]) );
  DFFPOSX1 mem_reg_22__16_ ( .D(n2760), .CLK(clk), .Q(mem[918]) );
  DFFPOSX1 mem_reg_22__15_ ( .D(n2759), .CLK(clk), .Q(mem[917]) );
  DFFPOSX1 mem_reg_22__14_ ( .D(n2758), .CLK(clk), .Q(mem[916]) );
  DFFPOSX1 mem_reg_22__13_ ( .D(n2757), .CLK(clk), .Q(mem[915]) );
  DFFPOSX1 mem_reg_22__12_ ( .D(n2756), .CLK(clk), .Q(mem[914]) );
  DFFPOSX1 mem_reg_22__11_ ( .D(n2755), .CLK(clk), .Q(mem[913]) );
  DFFPOSX1 mem_reg_22__10_ ( .D(n2754), .CLK(clk), .Q(mem[912]) );
  DFFPOSX1 mem_reg_22__9_ ( .D(n2753), .CLK(clk), .Q(mem[911]) );
  DFFPOSX1 mem_reg_22__8_ ( .D(n2752), .CLK(clk), .Q(mem[910]) );
  DFFPOSX1 mem_reg_22__7_ ( .D(n2751), .CLK(clk), .Q(mem[909]) );
  DFFPOSX1 mem_reg_22__6_ ( .D(n2750), .CLK(clk), .Q(mem[908]) );
  DFFPOSX1 mem_reg_22__5_ ( .D(n2749), .CLK(clk), .Q(mem[907]) );
  DFFPOSX1 mem_reg_22__4_ ( .D(n2748), .CLK(clk), .Q(mem[906]) );
  DFFPOSX1 mem_reg_22__3_ ( .D(n2747), .CLK(clk), .Q(mem[905]) );
  DFFPOSX1 mem_reg_22__2_ ( .D(n2746), .CLK(clk), .Q(mem[904]) );
  DFFPOSX1 mem_reg_22__1_ ( .D(n2745), .CLK(clk), .Q(mem[903]) );
  DFFPOSX1 mem_reg_22__0_ ( .D(n2744), .CLK(clk), .Q(mem[902]) );
  DFFPOSX1 mem_reg_21__40_ ( .D(n2743), .CLK(clk), .Q(mem[901]) );
  DFFPOSX1 mem_reg_21__39_ ( .D(n2742), .CLK(clk), .Q(mem[900]) );
  DFFPOSX1 mem_reg_21__38_ ( .D(n2741), .CLK(clk), .Q(mem[899]) );
  DFFPOSX1 mem_reg_21__37_ ( .D(n2740), .CLK(clk), .Q(mem[898]) );
  DFFPOSX1 mem_reg_21__36_ ( .D(n2739), .CLK(clk), .Q(mem[897]) );
  DFFPOSX1 mem_reg_21__35_ ( .D(n2738), .CLK(clk), .Q(mem[896]) );
  DFFPOSX1 mem_reg_21__34_ ( .D(n2737), .CLK(clk), .Q(mem[895]) );
  DFFPOSX1 mem_reg_21__33_ ( .D(n2736), .CLK(clk), .Q(mem[894]) );
  DFFPOSX1 mem_reg_21__32_ ( .D(n2735), .CLK(clk), .Q(mem[893]) );
  DFFPOSX1 mem_reg_21__31_ ( .D(n2734), .CLK(clk), .Q(mem[892]) );
  DFFPOSX1 mem_reg_21__30_ ( .D(n2733), .CLK(clk), .Q(mem[891]) );
  DFFPOSX1 mem_reg_21__29_ ( .D(n2732), .CLK(clk), .Q(mem[890]) );
  DFFPOSX1 mem_reg_21__28_ ( .D(n2731), .CLK(clk), .Q(mem[889]) );
  DFFPOSX1 mem_reg_21__27_ ( .D(n2730), .CLK(clk), .Q(mem[888]) );
  DFFPOSX1 mem_reg_21__26_ ( .D(n2729), .CLK(clk), .Q(mem[887]) );
  DFFPOSX1 mem_reg_21__25_ ( .D(n2728), .CLK(clk), .Q(mem[886]) );
  DFFPOSX1 mem_reg_21__24_ ( .D(n2727), .CLK(clk), .Q(mem[885]) );
  DFFPOSX1 mem_reg_21__23_ ( .D(n2726), .CLK(clk), .Q(mem[884]) );
  DFFPOSX1 mem_reg_21__22_ ( .D(n2725), .CLK(clk), .Q(mem[883]) );
  DFFPOSX1 mem_reg_21__21_ ( .D(n2724), .CLK(clk), .Q(mem[882]) );
  DFFPOSX1 mem_reg_21__20_ ( .D(n2723), .CLK(clk), .Q(mem[881]) );
  DFFPOSX1 mem_reg_21__19_ ( .D(n2722), .CLK(clk), .Q(mem[880]) );
  DFFPOSX1 mem_reg_21__18_ ( .D(n2721), .CLK(clk), .Q(mem[879]) );
  DFFPOSX1 mem_reg_21__17_ ( .D(n2720), .CLK(clk), .Q(mem[878]) );
  DFFPOSX1 mem_reg_21__16_ ( .D(n2719), .CLK(clk), .Q(mem[877]) );
  DFFPOSX1 mem_reg_21__15_ ( .D(n2718), .CLK(clk), .Q(mem[876]) );
  DFFPOSX1 mem_reg_21__14_ ( .D(n2717), .CLK(clk), .Q(mem[875]) );
  DFFPOSX1 mem_reg_21__13_ ( .D(n2716), .CLK(clk), .Q(mem[874]) );
  DFFPOSX1 mem_reg_21__12_ ( .D(n2715), .CLK(clk), .Q(mem[873]) );
  DFFPOSX1 mem_reg_21__11_ ( .D(n2714), .CLK(clk), .Q(mem[872]) );
  DFFPOSX1 mem_reg_21__10_ ( .D(n2713), .CLK(clk), .Q(mem[871]) );
  DFFPOSX1 mem_reg_21__9_ ( .D(n2712), .CLK(clk), .Q(mem[870]) );
  DFFPOSX1 mem_reg_21__8_ ( .D(n2711), .CLK(clk), .Q(mem[869]) );
  DFFPOSX1 mem_reg_21__7_ ( .D(n2710), .CLK(clk), .Q(mem[868]) );
  DFFPOSX1 mem_reg_21__6_ ( .D(n2709), .CLK(clk), .Q(mem[867]) );
  DFFPOSX1 mem_reg_21__5_ ( .D(n2708), .CLK(clk), .Q(mem[866]) );
  DFFPOSX1 mem_reg_21__4_ ( .D(n2707), .CLK(clk), .Q(mem[865]) );
  DFFPOSX1 mem_reg_21__3_ ( .D(n2706), .CLK(clk), .Q(mem[864]) );
  DFFPOSX1 mem_reg_21__2_ ( .D(n2705), .CLK(clk), .Q(mem[863]) );
  DFFPOSX1 mem_reg_21__1_ ( .D(n2704), .CLK(clk), .Q(mem[862]) );
  DFFPOSX1 mem_reg_21__0_ ( .D(n2703), .CLK(clk), .Q(mem[861]) );
  DFFPOSX1 mem_reg_20__40_ ( .D(n2702), .CLK(clk), .Q(mem[860]) );
  DFFPOSX1 mem_reg_20__39_ ( .D(n2701), .CLK(clk), .Q(mem[859]) );
  DFFPOSX1 mem_reg_20__38_ ( .D(n2700), .CLK(clk), .Q(mem[858]) );
  DFFPOSX1 mem_reg_20__37_ ( .D(n2699), .CLK(clk), .Q(mem[857]) );
  DFFPOSX1 mem_reg_20__36_ ( .D(n2698), .CLK(clk), .Q(mem[856]) );
  DFFPOSX1 mem_reg_20__35_ ( .D(n2697), .CLK(clk), .Q(mem[855]) );
  DFFPOSX1 mem_reg_20__34_ ( .D(n2696), .CLK(clk), .Q(mem[854]) );
  DFFPOSX1 mem_reg_20__33_ ( .D(n2695), .CLK(clk), .Q(mem[853]) );
  DFFPOSX1 mem_reg_20__32_ ( .D(n2694), .CLK(clk), .Q(mem[852]) );
  DFFPOSX1 mem_reg_20__31_ ( .D(n2693), .CLK(clk), .Q(mem[851]) );
  DFFPOSX1 mem_reg_20__30_ ( .D(n2692), .CLK(clk), .Q(mem[850]) );
  DFFPOSX1 mem_reg_20__29_ ( .D(n2691), .CLK(clk), .Q(mem[849]) );
  DFFPOSX1 mem_reg_20__28_ ( .D(n2690), .CLK(clk), .Q(mem[848]) );
  DFFPOSX1 mem_reg_20__27_ ( .D(n2689), .CLK(clk), .Q(mem[847]) );
  DFFPOSX1 mem_reg_20__26_ ( .D(n2688), .CLK(clk), .Q(mem[846]) );
  DFFPOSX1 mem_reg_20__25_ ( .D(n2687), .CLK(clk), .Q(mem[845]) );
  DFFPOSX1 mem_reg_20__24_ ( .D(n2686), .CLK(clk), .Q(mem[844]) );
  DFFPOSX1 mem_reg_20__23_ ( .D(n2685), .CLK(clk), .Q(mem[843]) );
  DFFPOSX1 mem_reg_20__22_ ( .D(n2684), .CLK(clk), .Q(mem[842]) );
  DFFPOSX1 mem_reg_20__21_ ( .D(n2683), .CLK(clk), .Q(mem[841]) );
  DFFPOSX1 mem_reg_20__20_ ( .D(n2682), .CLK(clk), .Q(mem[840]) );
  DFFPOSX1 mem_reg_20__19_ ( .D(n2681), .CLK(clk), .Q(mem[839]) );
  DFFPOSX1 mem_reg_20__18_ ( .D(n2680), .CLK(clk), .Q(mem[838]) );
  DFFPOSX1 mem_reg_20__17_ ( .D(n2679), .CLK(clk), .Q(mem[837]) );
  DFFPOSX1 mem_reg_20__16_ ( .D(n2678), .CLK(clk), .Q(mem[836]) );
  DFFPOSX1 mem_reg_20__15_ ( .D(n2677), .CLK(clk), .Q(mem[835]) );
  DFFPOSX1 mem_reg_20__14_ ( .D(n2676), .CLK(clk), .Q(mem[834]) );
  DFFPOSX1 mem_reg_20__13_ ( .D(n2675), .CLK(clk), .Q(mem[833]) );
  DFFPOSX1 mem_reg_20__12_ ( .D(n2674), .CLK(clk), .Q(mem[832]) );
  DFFPOSX1 mem_reg_20__11_ ( .D(n2673), .CLK(clk), .Q(mem[831]) );
  DFFPOSX1 mem_reg_20__10_ ( .D(n2672), .CLK(clk), .Q(mem[830]) );
  DFFPOSX1 mem_reg_20__9_ ( .D(n2671), .CLK(clk), .Q(mem[829]) );
  DFFPOSX1 mem_reg_20__8_ ( .D(n2670), .CLK(clk), .Q(mem[828]) );
  DFFPOSX1 mem_reg_20__7_ ( .D(n2669), .CLK(clk), .Q(mem[827]) );
  DFFPOSX1 mem_reg_20__6_ ( .D(n2668), .CLK(clk), .Q(mem[826]) );
  DFFPOSX1 mem_reg_20__5_ ( .D(n2667), .CLK(clk), .Q(mem[825]) );
  DFFPOSX1 mem_reg_20__4_ ( .D(n2666), .CLK(clk), .Q(mem[824]) );
  DFFPOSX1 mem_reg_20__3_ ( .D(n2665), .CLK(clk), .Q(mem[823]) );
  DFFPOSX1 mem_reg_20__2_ ( .D(n2664), .CLK(clk), .Q(mem[822]) );
  DFFPOSX1 mem_reg_20__1_ ( .D(n2663), .CLK(clk), .Q(mem[821]) );
  DFFPOSX1 mem_reg_20__0_ ( .D(n2662), .CLK(clk), .Q(mem[820]) );
  DFFPOSX1 mem_reg_19__40_ ( .D(n2661), .CLK(clk), .Q(mem[819]) );
  DFFPOSX1 mem_reg_19__39_ ( .D(n2660), .CLK(clk), .Q(mem[818]) );
  DFFPOSX1 mem_reg_19__38_ ( .D(n2659), .CLK(clk), .Q(mem[817]) );
  DFFPOSX1 mem_reg_19__37_ ( .D(n2658), .CLK(clk), .Q(mem[816]) );
  DFFPOSX1 mem_reg_19__36_ ( .D(n2657), .CLK(clk), .Q(mem[815]) );
  DFFPOSX1 mem_reg_19__35_ ( .D(n2656), .CLK(clk), .Q(mem[814]) );
  DFFPOSX1 mem_reg_19__34_ ( .D(n2655), .CLK(clk), .Q(mem[813]) );
  DFFPOSX1 mem_reg_19__33_ ( .D(n2654), .CLK(clk), .Q(mem[812]) );
  DFFPOSX1 mem_reg_19__32_ ( .D(n2653), .CLK(clk), .Q(mem[811]) );
  DFFPOSX1 mem_reg_19__31_ ( .D(n2652), .CLK(clk), .Q(mem[810]) );
  DFFPOSX1 mem_reg_19__30_ ( .D(n2651), .CLK(clk), .Q(mem[809]) );
  DFFPOSX1 mem_reg_19__29_ ( .D(n2650), .CLK(clk), .Q(mem[808]) );
  DFFPOSX1 mem_reg_19__28_ ( .D(n2649), .CLK(clk), .Q(mem[807]) );
  DFFPOSX1 mem_reg_19__27_ ( .D(n2648), .CLK(clk), .Q(mem[806]) );
  DFFPOSX1 mem_reg_19__26_ ( .D(n2647), .CLK(clk), .Q(mem[805]) );
  DFFPOSX1 mem_reg_19__25_ ( .D(n2646), .CLK(clk), .Q(mem[804]) );
  DFFPOSX1 mem_reg_19__24_ ( .D(n2645), .CLK(clk), .Q(mem[803]) );
  DFFPOSX1 mem_reg_19__23_ ( .D(n2644), .CLK(clk), .Q(mem[802]) );
  DFFPOSX1 mem_reg_19__22_ ( .D(n2643), .CLK(clk), .Q(mem[801]) );
  DFFPOSX1 mem_reg_19__21_ ( .D(n2642), .CLK(clk), .Q(mem[800]) );
  DFFPOSX1 mem_reg_19__20_ ( .D(n2641), .CLK(clk), .Q(mem[799]) );
  DFFPOSX1 mem_reg_19__19_ ( .D(n2640), .CLK(clk), .Q(mem[798]) );
  DFFPOSX1 mem_reg_19__18_ ( .D(n2639), .CLK(clk), .Q(mem[797]) );
  DFFPOSX1 mem_reg_19__17_ ( .D(n2638), .CLK(clk), .Q(mem[796]) );
  DFFPOSX1 mem_reg_19__16_ ( .D(n2637), .CLK(clk), .Q(mem[795]) );
  DFFPOSX1 mem_reg_19__15_ ( .D(n2636), .CLK(clk), .Q(mem[794]) );
  DFFPOSX1 mem_reg_19__14_ ( .D(n2635), .CLK(clk), .Q(mem[793]) );
  DFFPOSX1 mem_reg_19__13_ ( .D(n2634), .CLK(clk), .Q(mem[792]) );
  DFFPOSX1 mem_reg_19__12_ ( .D(n2633), .CLK(clk), .Q(mem[791]) );
  DFFPOSX1 mem_reg_19__11_ ( .D(n2632), .CLK(clk), .Q(mem[790]) );
  DFFPOSX1 mem_reg_19__10_ ( .D(n2631), .CLK(clk), .Q(mem[789]) );
  DFFPOSX1 mem_reg_19__9_ ( .D(n2630), .CLK(clk), .Q(mem[788]) );
  DFFPOSX1 mem_reg_19__8_ ( .D(n2629), .CLK(clk), .Q(mem[787]) );
  DFFPOSX1 mem_reg_19__7_ ( .D(n2628), .CLK(clk), .Q(mem[786]) );
  DFFPOSX1 mem_reg_19__6_ ( .D(n2627), .CLK(clk), .Q(mem[785]) );
  DFFPOSX1 mem_reg_19__5_ ( .D(n2626), .CLK(clk), .Q(mem[784]) );
  DFFPOSX1 mem_reg_19__4_ ( .D(n2625), .CLK(clk), .Q(mem[783]) );
  DFFPOSX1 mem_reg_19__3_ ( .D(n2624), .CLK(clk), .Q(mem[782]) );
  DFFPOSX1 mem_reg_19__2_ ( .D(n2623), .CLK(clk), .Q(mem[781]) );
  DFFPOSX1 mem_reg_19__1_ ( .D(n2622), .CLK(clk), .Q(mem[780]) );
  DFFPOSX1 mem_reg_19__0_ ( .D(n2621), .CLK(clk), .Q(mem[779]) );
  DFFPOSX1 mem_reg_18__40_ ( .D(n2620), .CLK(clk), .Q(mem[778]) );
  DFFPOSX1 mem_reg_18__39_ ( .D(n2619), .CLK(clk), .Q(mem[777]) );
  DFFPOSX1 mem_reg_18__38_ ( .D(n2618), .CLK(clk), .Q(mem[776]) );
  DFFPOSX1 mem_reg_18__37_ ( .D(n2617), .CLK(clk), .Q(mem[775]) );
  DFFPOSX1 mem_reg_18__36_ ( .D(n2616), .CLK(clk), .Q(mem[774]) );
  DFFPOSX1 mem_reg_18__35_ ( .D(n2615), .CLK(clk), .Q(mem[773]) );
  DFFPOSX1 mem_reg_18__34_ ( .D(n2614), .CLK(clk), .Q(mem[772]) );
  DFFPOSX1 mem_reg_18__33_ ( .D(n2613), .CLK(clk), .Q(mem[771]) );
  DFFPOSX1 mem_reg_18__32_ ( .D(n2612), .CLK(clk), .Q(mem[770]) );
  DFFPOSX1 mem_reg_18__31_ ( .D(n2611), .CLK(clk), .Q(mem[769]) );
  DFFPOSX1 mem_reg_18__30_ ( .D(n2610), .CLK(clk), .Q(mem[768]) );
  DFFPOSX1 mem_reg_18__29_ ( .D(n2609), .CLK(clk), .Q(mem[767]) );
  DFFPOSX1 mem_reg_18__28_ ( .D(n2608), .CLK(clk), .Q(mem[766]) );
  DFFPOSX1 mem_reg_18__27_ ( .D(n2607), .CLK(clk), .Q(mem[765]) );
  DFFPOSX1 mem_reg_18__26_ ( .D(n2606), .CLK(clk), .Q(mem[764]) );
  DFFPOSX1 mem_reg_18__25_ ( .D(n2605), .CLK(clk), .Q(mem[763]) );
  DFFPOSX1 mem_reg_18__24_ ( .D(n2604), .CLK(clk), .Q(mem[762]) );
  DFFPOSX1 mem_reg_18__23_ ( .D(n2603), .CLK(clk), .Q(mem[761]) );
  DFFPOSX1 mem_reg_18__22_ ( .D(n2602), .CLK(clk), .Q(mem[760]) );
  DFFPOSX1 mem_reg_18__21_ ( .D(n2601), .CLK(clk), .Q(mem[759]) );
  DFFPOSX1 mem_reg_18__20_ ( .D(n2600), .CLK(clk), .Q(mem[758]) );
  DFFPOSX1 mem_reg_18__19_ ( .D(n2599), .CLK(clk), .Q(mem[757]) );
  DFFPOSX1 mem_reg_18__18_ ( .D(n2598), .CLK(clk), .Q(mem[756]) );
  DFFPOSX1 mem_reg_18__17_ ( .D(n2597), .CLK(clk), .Q(mem[755]) );
  DFFPOSX1 mem_reg_18__16_ ( .D(n2596), .CLK(clk), .Q(mem[754]) );
  DFFPOSX1 mem_reg_18__15_ ( .D(n2595), .CLK(clk), .Q(mem[753]) );
  DFFPOSX1 mem_reg_18__14_ ( .D(n2594), .CLK(clk), .Q(mem[752]) );
  DFFPOSX1 mem_reg_18__13_ ( .D(n2593), .CLK(clk), .Q(mem[751]) );
  DFFPOSX1 mem_reg_18__12_ ( .D(n2592), .CLK(clk), .Q(mem[750]) );
  DFFPOSX1 mem_reg_18__11_ ( .D(n2591), .CLK(clk), .Q(mem[749]) );
  DFFPOSX1 mem_reg_18__10_ ( .D(n2590), .CLK(clk), .Q(mem[748]) );
  DFFPOSX1 mem_reg_18__9_ ( .D(n2589), .CLK(clk), .Q(mem[747]) );
  DFFPOSX1 mem_reg_18__8_ ( .D(n2588), .CLK(clk), .Q(mem[746]) );
  DFFPOSX1 mem_reg_18__7_ ( .D(n2587), .CLK(clk), .Q(mem[745]) );
  DFFPOSX1 mem_reg_18__6_ ( .D(n2586), .CLK(clk), .Q(mem[744]) );
  DFFPOSX1 mem_reg_18__5_ ( .D(n2585), .CLK(clk), .Q(mem[743]) );
  DFFPOSX1 mem_reg_18__4_ ( .D(n2584), .CLK(clk), .Q(mem[742]) );
  DFFPOSX1 mem_reg_18__3_ ( .D(n2583), .CLK(clk), .Q(mem[741]) );
  DFFPOSX1 mem_reg_18__2_ ( .D(n2582), .CLK(clk), .Q(mem[740]) );
  DFFPOSX1 mem_reg_18__1_ ( .D(n2581), .CLK(clk), .Q(mem[739]) );
  DFFPOSX1 mem_reg_18__0_ ( .D(n2580), .CLK(clk), .Q(mem[738]) );
  DFFPOSX1 mem_reg_17__40_ ( .D(n2579), .CLK(clk), .Q(mem[737]) );
  DFFPOSX1 mem_reg_17__39_ ( .D(n2578), .CLK(clk), .Q(mem[736]) );
  DFFPOSX1 mem_reg_17__38_ ( .D(n2577), .CLK(clk), .Q(mem[735]) );
  DFFPOSX1 mem_reg_17__37_ ( .D(n2576), .CLK(clk), .Q(mem[734]) );
  DFFPOSX1 mem_reg_17__36_ ( .D(n2575), .CLK(clk), .Q(mem[733]) );
  DFFPOSX1 mem_reg_17__35_ ( .D(n2574), .CLK(clk), .Q(mem[732]) );
  DFFPOSX1 mem_reg_17__34_ ( .D(n2573), .CLK(clk), .Q(mem[731]) );
  DFFPOSX1 mem_reg_17__33_ ( .D(n2572), .CLK(clk), .Q(mem[730]) );
  DFFPOSX1 mem_reg_17__32_ ( .D(n2571), .CLK(clk), .Q(mem[729]) );
  DFFPOSX1 mem_reg_17__31_ ( .D(n2570), .CLK(clk), .Q(mem[728]) );
  DFFPOSX1 mem_reg_17__30_ ( .D(n2569), .CLK(clk), .Q(mem[727]) );
  DFFPOSX1 mem_reg_17__29_ ( .D(n2568), .CLK(clk), .Q(mem[726]) );
  DFFPOSX1 mem_reg_17__28_ ( .D(n2567), .CLK(clk), .Q(mem[725]) );
  DFFPOSX1 mem_reg_17__27_ ( .D(n2566), .CLK(clk), .Q(mem[724]) );
  DFFPOSX1 mem_reg_17__26_ ( .D(n2565), .CLK(clk), .Q(mem[723]) );
  DFFPOSX1 mem_reg_17__25_ ( .D(n2564), .CLK(clk), .Q(mem[722]) );
  DFFPOSX1 mem_reg_17__24_ ( .D(n2563), .CLK(clk), .Q(mem[721]) );
  DFFPOSX1 mem_reg_17__23_ ( .D(n2562), .CLK(clk), .Q(mem[720]) );
  DFFPOSX1 mem_reg_17__22_ ( .D(n2561), .CLK(clk), .Q(mem[719]) );
  DFFPOSX1 mem_reg_17__21_ ( .D(n2560), .CLK(clk), .Q(mem[718]) );
  DFFPOSX1 mem_reg_17__20_ ( .D(n2559), .CLK(clk), .Q(mem[717]) );
  DFFPOSX1 mem_reg_17__19_ ( .D(n2558), .CLK(clk), .Q(mem[716]) );
  DFFPOSX1 mem_reg_17__18_ ( .D(n2557), .CLK(clk), .Q(mem[715]) );
  DFFPOSX1 mem_reg_17__17_ ( .D(n2556), .CLK(clk), .Q(mem[714]) );
  DFFPOSX1 mem_reg_17__16_ ( .D(n2555), .CLK(clk), .Q(mem[713]) );
  DFFPOSX1 mem_reg_17__15_ ( .D(n2554), .CLK(clk), .Q(mem[712]) );
  DFFPOSX1 mem_reg_17__14_ ( .D(n2553), .CLK(clk), .Q(mem[711]) );
  DFFPOSX1 mem_reg_17__13_ ( .D(n2552), .CLK(clk), .Q(mem[710]) );
  DFFPOSX1 mem_reg_17__12_ ( .D(n2551), .CLK(clk), .Q(mem[709]) );
  DFFPOSX1 mem_reg_17__11_ ( .D(n2550), .CLK(clk), .Q(mem[708]) );
  DFFPOSX1 mem_reg_17__10_ ( .D(n2549), .CLK(clk), .Q(mem[707]) );
  DFFPOSX1 mem_reg_17__9_ ( .D(n2548), .CLK(clk), .Q(mem[706]) );
  DFFPOSX1 mem_reg_17__8_ ( .D(n2547), .CLK(clk), .Q(mem[705]) );
  DFFPOSX1 mem_reg_17__7_ ( .D(n2546), .CLK(clk), .Q(mem[704]) );
  DFFPOSX1 mem_reg_17__6_ ( .D(n2545), .CLK(clk), .Q(mem[703]) );
  DFFPOSX1 mem_reg_17__5_ ( .D(n2544), .CLK(clk), .Q(mem[702]) );
  DFFPOSX1 mem_reg_17__4_ ( .D(n2543), .CLK(clk), .Q(mem[701]) );
  DFFPOSX1 mem_reg_17__3_ ( .D(n2542), .CLK(clk), .Q(mem[700]) );
  DFFPOSX1 mem_reg_17__2_ ( .D(n2541), .CLK(clk), .Q(mem[699]) );
  DFFPOSX1 mem_reg_17__1_ ( .D(n2540), .CLK(clk), .Q(mem[698]) );
  DFFPOSX1 mem_reg_17__0_ ( .D(n2539), .CLK(clk), .Q(mem[697]) );
  DFFPOSX1 mem_reg_16__40_ ( .D(n2538), .CLK(clk), .Q(mem[696]) );
  DFFPOSX1 mem_reg_16__39_ ( .D(n2537), .CLK(clk), .Q(mem[695]) );
  DFFPOSX1 mem_reg_16__38_ ( .D(n2536), .CLK(clk), .Q(mem[694]) );
  DFFPOSX1 mem_reg_16__37_ ( .D(n2535), .CLK(clk), .Q(mem[693]) );
  DFFPOSX1 mem_reg_16__36_ ( .D(n2534), .CLK(clk), .Q(mem[692]) );
  DFFPOSX1 mem_reg_16__35_ ( .D(n2533), .CLK(clk), .Q(mem[691]) );
  DFFPOSX1 mem_reg_16__34_ ( .D(n2532), .CLK(clk), .Q(mem[690]) );
  DFFPOSX1 mem_reg_16__33_ ( .D(n2531), .CLK(clk), .Q(mem[689]) );
  DFFPOSX1 mem_reg_16__32_ ( .D(n2530), .CLK(clk), .Q(mem[688]) );
  DFFPOSX1 mem_reg_16__31_ ( .D(n2529), .CLK(clk), .Q(mem[687]) );
  DFFPOSX1 mem_reg_16__30_ ( .D(n2528), .CLK(clk), .Q(mem[686]) );
  DFFPOSX1 mem_reg_16__29_ ( .D(n2527), .CLK(clk), .Q(mem[685]) );
  DFFPOSX1 mem_reg_16__28_ ( .D(n2526), .CLK(clk), .Q(mem[684]) );
  DFFPOSX1 mem_reg_16__27_ ( .D(n2525), .CLK(clk), .Q(mem[683]) );
  DFFPOSX1 mem_reg_16__26_ ( .D(n2524), .CLK(clk), .Q(mem[682]) );
  DFFPOSX1 mem_reg_16__25_ ( .D(n2523), .CLK(clk), .Q(mem[681]) );
  DFFPOSX1 mem_reg_16__24_ ( .D(n2522), .CLK(clk), .Q(mem[680]) );
  DFFPOSX1 mem_reg_16__23_ ( .D(n2521), .CLK(clk), .Q(mem[679]) );
  DFFPOSX1 mem_reg_16__22_ ( .D(n2520), .CLK(clk), .Q(mem[678]) );
  DFFPOSX1 mem_reg_16__21_ ( .D(n2519), .CLK(clk), .Q(mem[677]) );
  DFFPOSX1 mem_reg_16__20_ ( .D(n2518), .CLK(clk), .Q(mem[676]) );
  DFFPOSX1 mem_reg_16__19_ ( .D(n2517), .CLK(clk), .Q(mem[675]) );
  DFFPOSX1 mem_reg_16__18_ ( .D(n2516), .CLK(clk), .Q(mem[674]) );
  DFFPOSX1 mem_reg_16__17_ ( .D(n2515), .CLK(clk), .Q(mem[673]) );
  DFFPOSX1 mem_reg_16__16_ ( .D(n2514), .CLK(clk), .Q(mem[672]) );
  DFFPOSX1 mem_reg_16__15_ ( .D(n2513), .CLK(clk), .Q(mem[671]) );
  DFFPOSX1 mem_reg_16__14_ ( .D(n2512), .CLK(clk), .Q(mem[670]) );
  DFFPOSX1 mem_reg_16__13_ ( .D(n2511), .CLK(clk), .Q(mem[669]) );
  DFFPOSX1 mem_reg_16__12_ ( .D(n2510), .CLK(clk), .Q(mem[668]) );
  DFFPOSX1 mem_reg_16__11_ ( .D(n2509), .CLK(clk), .Q(mem[667]) );
  DFFPOSX1 mem_reg_16__10_ ( .D(n2508), .CLK(clk), .Q(mem[666]) );
  DFFPOSX1 mem_reg_16__9_ ( .D(n2507), .CLK(clk), .Q(mem[665]) );
  DFFPOSX1 mem_reg_16__8_ ( .D(n2506), .CLK(clk), .Q(mem[664]) );
  DFFPOSX1 mem_reg_16__7_ ( .D(n2505), .CLK(clk), .Q(mem[663]) );
  DFFPOSX1 mem_reg_16__6_ ( .D(n2504), .CLK(clk), .Q(mem[662]) );
  DFFPOSX1 mem_reg_16__5_ ( .D(n2503), .CLK(clk), .Q(mem[661]) );
  DFFPOSX1 mem_reg_16__4_ ( .D(n2502), .CLK(clk), .Q(mem[660]) );
  DFFPOSX1 mem_reg_16__3_ ( .D(n2501), .CLK(clk), .Q(mem[659]) );
  DFFPOSX1 mem_reg_16__2_ ( .D(n2500), .CLK(clk), .Q(mem[658]) );
  DFFPOSX1 mem_reg_16__1_ ( .D(n2499), .CLK(clk), .Q(mem[657]) );
  DFFPOSX1 mem_reg_16__0_ ( .D(n2498), .CLK(clk), .Q(mem[656]) );
  DFFPOSX1 mem_reg_15__40_ ( .D(n2497), .CLK(clk), .Q(mem[655]) );
  DFFPOSX1 mem_reg_15__39_ ( .D(n2496), .CLK(clk), .Q(mem[654]) );
  DFFPOSX1 mem_reg_15__38_ ( .D(n2495), .CLK(clk), .Q(mem[653]) );
  DFFPOSX1 mem_reg_15__37_ ( .D(n2494), .CLK(clk), .Q(mem[652]) );
  DFFPOSX1 mem_reg_15__36_ ( .D(n2493), .CLK(clk), .Q(mem[651]) );
  DFFPOSX1 mem_reg_15__35_ ( .D(n2492), .CLK(clk), .Q(mem[650]) );
  DFFPOSX1 mem_reg_15__34_ ( .D(n2491), .CLK(clk), .Q(mem[649]) );
  DFFPOSX1 mem_reg_15__33_ ( .D(n2490), .CLK(clk), .Q(mem[648]) );
  DFFPOSX1 mem_reg_15__32_ ( .D(n2489), .CLK(clk), .Q(mem[647]) );
  DFFPOSX1 mem_reg_15__31_ ( .D(n2488), .CLK(clk), .Q(mem[646]) );
  DFFPOSX1 mem_reg_15__30_ ( .D(n2487), .CLK(clk), .Q(mem[645]) );
  DFFPOSX1 mem_reg_15__29_ ( .D(n2486), .CLK(clk), .Q(mem[644]) );
  DFFPOSX1 mem_reg_15__28_ ( .D(n2485), .CLK(clk), .Q(mem[643]) );
  DFFPOSX1 mem_reg_15__27_ ( .D(n2484), .CLK(clk), .Q(mem[642]) );
  DFFPOSX1 mem_reg_15__26_ ( .D(n2483), .CLK(clk), .Q(mem[641]) );
  DFFPOSX1 mem_reg_15__25_ ( .D(n2482), .CLK(clk), .Q(mem[640]) );
  DFFPOSX1 mem_reg_15__24_ ( .D(n2481), .CLK(clk), .Q(mem[639]) );
  DFFPOSX1 mem_reg_15__23_ ( .D(n2480), .CLK(clk), .Q(mem[638]) );
  DFFPOSX1 mem_reg_15__22_ ( .D(n2479), .CLK(clk), .Q(mem[637]) );
  DFFPOSX1 mem_reg_15__21_ ( .D(n2478), .CLK(clk), .Q(mem[636]) );
  DFFPOSX1 mem_reg_15__20_ ( .D(n2477), .CLK(clk), .Q(mem[635]) );
  DFFPOSX1 mem_reg_15__19_ ( .D(n2476), .CLK(clk), .Q(mem[634]) );
  DFFPOSX1 mem_reg_15__18_ ( .D(n2475), .CLK(clk), .Q(mem[633]) );
  DFFPOSX1 mem_reg_15__17_ ( .D(n2474), .CLK(clk), .Q(mem[632]) );
  DFFPOSX1 mem_reg_15__16_ ( .D(n2473), .CLK(clk), .Q(mem[631]) );
  DFFPOSX1 mem_reg_15__15_ ( .D(n2472), .CLK(clk), .Q(mem[630]) );
  DFFPOSX1 mem_reg_15__14_ ( .D(n2471), .CLK(clk), .Q(mem[629]) );
  DFFPOSX1 mem_reg_15__13_ ( .D(n2470), .CLK(clk), .Q(mem[628]) );
  DFFPOSX1 mem_reg_15__12_ ( .D(n2469), .CLK(clk), .Q(mem[627]) );
  DFFPOSX1 mem_reg_15__11_ ( .D(n2468), .CLK(clk), .Q(mem[626]) );
  DFFPOSX1 mem_reg_15__10_ ( .D(n2467), .CLK(clk), .Q(mem[625]) );
  DFFPOSX1 mem_reg_15__9_ ( .D(n2466), .CLK(clk), .Q(mem[624]) );
  DFFPOSX1 mem_reg_15__8_ ( .D(n2465), .CLK(clk), .Q(mem[623]) );
  DFFPOSX1 mem_reg_15__7_ ( .D(n2464), .CLK(clk), .Q(mem[622]) );
  DFFPOSX1 mem_reg_15__6_ ( .D(n2463), .CLK(clk), .Q(mem[621]) );
  DFFPOSX1 mem_reg_15__5_ ( .D(n2462), .CLK(clk), .Q(mem[620]) );
  DFFPOSX1 mem_reg_15__4_ ( .D(n2461), .CLK(clk), .Q(mem[619]) );
  DFFPOSX1 mem_reg_15__3_ ( .D(n2460), .CLK(clk), .Q(mem[618]) );
  DFFPOSX1 mem_reg_15__2_ ( .D(n2459), .CLK(clk), .Q(mem[617]) );
  DFFPOSX1 mem_reg_15__1_ ( .D(n2458), .CLK(clk), .Q(mem[616]) );
  DFFPOSX1 mem_reg_15__0_ ( .D(n2457), .CLK(clk), .Q(mem[615]) );
  DFFPOSX1 mem_reg_14__40_ ( .D(n2456), .CLK(clk), .Q(mem[614]) );
  DFFPOSX1 mem_reg_14__39_ ( .D(n2455), .CLK(clk), .Q(mem[613]) );
  DFFPOSX1 mem_reg_14__38_ ( .D(n2454), .CLK(clk), .Q(mem[612]) );
  DFFPOSX1 mem_reg_14__37_ ( .D(n2453), .CLK(clk), .Q(mem[611]) );
  DFFPOSX1 mem_reg_14__36_ ( .D(n2452), .CLK(clk), .Q(mem[610]) );
  DFFPOSX1 mem_reg_14__35_ ( .D(n2451), .CLK(clk), .Q(mem[609]) );
  DFFPOSX1 mem_reg_14__34_ ( .D(n2450), .CLK(clk), .Q(mem[608]) );
  DFFPOSX1 mem_reg_14__33_ ( .D(n2449), .CLK(clk), .Q(mem[607]) );
  DFFPOSX1 mem_reg_14__32_ ( .D(n2448), .CLK(clk), .Q(mem[606]) );
  DFFPOSX1 mem_reg_14__31_ ( .D(n2447), .CLK(clk), .Q(mem[605]) );
  DFFPOSX1 mem_reg_14__30_ ( .D(n2446), .CLK(clk), .Q(mem[604]) );
  DFFPOSX1 mem_reg_14__29_ ( .D(n2445), .CLK(clk), .Q(mem[603]) );
  DFFPOSX1 mem_reg_14__28_ ( .D(n2444), .CLK(clk), .Q(mem[602]) );
  DFFPOSX1 mem_reg_14__27_ ( .D(n2443), .CLK(clk), .Q(mem[601]) );
  DFFPOSX1 mem_reg_14__26_ ( .D(n2442), .CLK(clk), .Q(mem[600]) );
  DFFPOSX1 mem_reg_14__25_ ( .D(n2441), .CLK(clk), .Q(mem[599]) );
  DFFPOSX1 mem_reg_14__24_ ( .D(n2440), .CLK(clk), .Q(mem[598]) );
  DFFPOSX1 mem_reg_14__23_ ( .D(n2439), .CLK(clk), .Q(mem[597]) );
  DFFPOSX1 mem_reg_14__22_ ( .D(n2438), .CLK(clk), .Q(mem[596]) );
  DFFPOSX1 mem_reg_14__21_ ( .D(n2437), .CLK(clk), .Q(mem[595]) );
  DFFPOSX1 mem_reg_14__20_ ( .D(n2436), .CLK(clk), .Q(mem[594]) );
  DFFPOSX1 mem_reg_14__19_ ( .D(n2435), .CLK(clk), .Q(mem[593]) );
  DFFPOSX1 mem_reg_14__18_ ( .D(n2434), .CLK(clk), .Q(mem[592]) );
  DFFPOSX1 mem_reg_14__17_ ( .D(n2433), .CLK(clk), .Q(mem[591]) );
  DFFPOSX1 mem_reg_14__16_ ( .D(n2432), .CLK(clk), .Q(mem[590]) );
  DFFPOSX1 mem_reg_14__15_ ( .D(n2431), .CLK(clk), .Q(mem[589]) );
  DFFPOSX1 mem_reg_14__14_ ( .D(n2430), .CLK(clk), .Q(mem[588]) );
  DFFPOSX1 mem_reg_14__13_ ( .D(n2429), .CLK(clk), .Q(mem[587]) );
  DFFPOSX1 mem_reg_14__12_ ( .D(n2428), .CLK(clk), .Q(mem[586]) );
  DFFPOSX1 mem_reg_14__11_ ( .D(n2427), .CLK(clk), .Q(mem[585]) );
  DFFPOSX1 mem_reg_14__10_ ( .D(n2426), .CLK(clk), .Q(mem[584]) );
  DFFPOSX1 mem_reg_14__9_ ( .D(n2425), .CLK(clk), .Q(mem[583]) );
  DFFPOSX1 mem_reg_14__8_ ( .D(n2424), .CLK(clk), .Q(mem[582]) );
  DFFPOSX1 mem_reg_14__7_ ( .D(n2423), .CLK(clk), .Q(mem[581]) );
  DFFPOSX1 mem_reg_14__6_ ( .D(n2422), .CLK(clk), .Q(mem[580]) );
  DFFPOSX1 mem_reg_14__5_ ( .D(n2421), .CLK(clk), .Q(mem[579]) );
  DFFPOSX1 mem_reg_14__4_ ( .D(n2420), .CLK(clk), .Q(mem[578]) );
  DFFPOSX1 mem_reg_14__3_ ( .D(n2419), .CLK(clk), .Q(mem[577]) );
  DFFPOSX1 mem_reg_14__2_ ( .D(n2418), .CLK(clk), .Q(mem[576]) );
  DFFPOSX1 mem_reg_14__1_ ( .D(n2417), .CLK(clk), .Q(mem[575]) );
  DFFPOSX1 mem_reg_14__0_ ( .D(n2416), .CLK(clk), .Q(mem[574]) );
  DFFPOSX1 mem_reg_13__40_ ( .D(n2415), .CLK(clk), .Q(mem[573]) );
  DFFPOSX1 mem_reg_13__39_ ( .D(n2414), .CLK(clk), .Q(mem[572]) );
  DFFPOSX1 mem_reg_13__38_ ( .D(n2413), .CLK(clk), .Q(mem[571]) );
  DFFPOSX1 mem_reg_13__37_ ( .D(n2412), .CLK(clk), .Q(mem[570]) );
  DFFPOSX1 mem_reg_13__36_ ( .D(n2411), .CLK(clk), .Q(mem[569]) );
  DFFPOSX1 mem_reg_13__35_ ( .D(n2410), .CLK(clk), .Q(mem[568]) );
  DFFPOSX1 mem_reg_13__34_ ( .D(n2409), .CLK(clk), .Q(mem[567]) );
  DFFPOSX1 mem_reg_13__33_ ( .D(n2408), .CLK(clk), .Q(mem[566]) );
  DFFPOSX1 mem_reg_13__32_ ( .D(n2407), .CLK(clk), .Q(mem[565]) );
  DFFPOSX1 mem_reg_13__31_ ( .D(n2406), .CLK(clk), .Q(mem[564]) );
  DFFPOSX1 mem_reg_13__30_ ( .D(n2405), .CLK(clk), .Q(mem[563]) );
  DFFPOSX1 mem_reg_13__29_ ( .D(n2404), .CLK(clk), .Q(mem[562]) );
  DFFPOSX1 mem_reg_13__28_ ( .D(n2403), .CLK(clk), .Q(mem[561]) );
  DFFPOSX1 mem_reg_13__27_ ( .D(n2402), .CLK(clk), .Q(mem[560]) );
  DFFPOSX1 mem_reg_13__26_ ( .D(n2401), .CLK(clk), .Q(mem[559]) );
  DFFPOSX1 mem_reg_13__25_ ( .D(n2400), .CLK(clk), .Q(mem[558]) );
  DFFPOSX1 mem_reg_13__24_ ( .D(n2399), .CLK(clk), .Q(mem[557]) );
  DFFPOSX1 mem_reg_13__23_ ( .D(n2398), .CLK(clk), .Q(mem[556]) );
  DFFPOSX1 mem_reg_13__22_ ( .D(n2397), .CLK(clk), .Q(mem[555]) );
  DFFPOSX1 mem_reg_13__21_ ( .D(n2396), .CLK(clk), .Q(mem[554]) );
  DFFPOSX1 mem_reg_13__20_ ( .D(n2395), .CLK(clk), .Q(mem[553]) );
  DFFPOSX1 mem_reg_13__19_ ( .D(n2394), .CLK(clk), .Q(mem[552]) );
  DFFPOSX1 mem_reg_13__18_ ( .D(n2393), .CLK(clk), .Q(mem[551]) );
  DFFPOSX1 mem_reg_13__17_ ( .D(n2392), .CLK(clk), .Q(mem[550]) );
  DFFPOSX1 mem_reg_13__16_ ( .D(n2391), .CLK(clk), .Q(mem[549]) );
  DFFPOSX1 mem_reg_13__15_ ( .D(n2390), .CLK(clk), .Q(mem[548]) );
  DFFPOSX1 mem_reg_13__14_ ( .D(n2389), .CLK(clk), .Q(mem[547]) );
  DFFPOSX1 mem_reg_13__13_ ( .D(n2388), .CLK(clk), .Q(mem[546]) );
  DFFPOSX1 mem_reg_13__12_ ( .D(n2387), .CLK(clk), .Q(mem[545]) );
  DFFPOSX1 mem_reg_13__11_ ( .D(n2386), .CLK(clk), .Q(mem[544]) );
  DFFPOSX1 mem_reg_13__10_ ( .D(n2385), .CLK(clk), .Q(mem[543]) );
  DFFPOSX1 mem_reg_13__9_ ( .D(n2384), .CLK(clk), .Q(mem[542]) );
  DFFPOSX1 mem_reg_13__8_ ( .D(n2383), .CLK(clk), .Q(mem[541]) );
  DFFPOSX1 mem_reg_13__7_ ( .D(n2382), .CLK(clk), .Q(mem[540]) );
  DFFPOSX1 mem_reg_13__6_ ( .D(n2381), .CLK(clk), .Q(mem[539]) );
  DFFPOSX1 mem_reg_13__5_ ( .D(n2380), .CLK(clk), .Q(mem[538]) );
  DFFPOSX1 mem_reg_13__4_ ( .D(n2379), .CLK(clk), .Q(mem[537]) );
  DFFPOSX1 mem_reg_13__3_ ( .D(n2378), .CLK(clk), .Q(mem[536]) );
  DFFPOSX1 mem_reg_13__2_ ( .D(n2377), .CLK(clk), .Q(mem[535]) );
  DFFPOSX1 mem_reg_13__1_ ( .D(n2376), .CLK(clk), .Q(mem[534]) );
  DFFPOSX1 mem_reg_13__0_ ( .D(n2375), .CLK(clk), .Q(mem[533]) );
  DFFPOSX1 mem_reg_12__40_ ( .D(n2374), .CLK(clk), .Q(mem[532]) );
  DFFPOSX1 mem_reg_12__39_ ( .D(n2373), .CLK(clk), .Q(mem[531]) );
  DFFPOSX1 mem_reg_12__38_ ( .D(n2372), .CLK(clk), .Q(mem[530]) );
  DFFPOSX1 mem_reg_12__37_ ( .D(n2371), .CLK(clk), .Q(mem[529]) );
  DFFPOSX1 mem_reg_12__36_ ( .D(n2370), .CLK(clk), .Q(mem[528]) );
  DFFPOSX1 mem_reg_12__35_ ( .D(n2369), .CLK(clk), .Q(mem[527]) );
  DFFPOSX1 mem_reg_12__34_ ( .D(n2368), .CLK(clk), .Q(mem[526]) );
  DFFPOSX1 mem_reg_12__33_ ( .D(n2367), .CLK(clk), .Q(mem[525]) );
  DFFPOSX1 mem_reg_12__32_ ( .D(n2366), .CLK(clk), .Q(mem[524]) );
  DFFPOSX1 mem_reg_12__31_ ( .D(n2365), .CLK(clk), .Q(mem[523]) );
  DFFPOSX1 mem_reg_12__30_ ( .D(n2364), .CLK(clk), .Q(mem[522]) );
  DFFPOSX1 mem_reg_12__29_ ( .D(n2363), .CLK(clk), .Q(mem[521]) );
  DFFPOSX1 mem_reg_12__28_ ( .D(n2362), .CLK(clk), .Q(mem[520]) );
  DFFPOSX1 mem_reg_12__27_ ( .D(n2361), .CLK(clk), .Q(mem[519]) );
  DFFPOSX1 mem_reg_12__26_ ( .D(n2360), .CLK(clk), .Q(mem[518]) );
  DFFPOSX1 mem_reg_12__25_ ( .D(n2359), .CLK(clk), .Q(mem[517]) );
  DFFPOSX1 mem_reg_12__24_ ( .D(n2358), .CLK(clk), .Q(mem[516]) );
  DFFPOSX1 mem_reg_12__23_ ( .D(n2357), .CLK(clk), .Q(mem[515]) );
  DFFPOSX1 mem_reg_12__22_ ( .D(n2356), .CLK(clk), .Q(mem[514]) );
  DFFPOSX1 mem_reg_12__21_ ( .D(n2355), .CLK(clk), .Q(mem[513]) );
  DFFPOSX1 mem_reg_12__20_ ( .D(n2354), .CLK(clk), .Q(mem[512]) );
  DFFPOSX1 mem_reg_12__19_ ( .D(n2353), .CLK(clk), .Q(mem[511]) );
  DFFPOSX1 mem_reg_12__18_ ( .D(n2352), .CLK(clk), .Q(mem[510]) );
  DFFPOSX1 mem_reg_12__17_ ( .D(n2351), .CLK(clk), .Q(mem[509]) );
  DFFPOSX1 mem_reg_12__16_ ( .D(n2350), .CLK(clk), .Q(mem[508]) );
  DFFPOSX1 mem_reg_12__15_ ( .D(n2349), .CLK(clk), .Q(mem[507]) );
  DFFPOSX1 mem_reg_12__14_ ( .D(n2348), .CLK(clk), .Q(mem[506]) );
  DFFPOSX1 mem_reg_12__13_ ( .D(n2347), .CLK(clk), .Q(mem[505]) );
  DFFPOSX1 mem_reg_12__12_ ( .D(n2346), .CLK(clk), .Q(mem[504]) );
  DFFPOSX1 mem_reg_12__11_ ( .D(n2345), .CLK(clk), .Q(mem[503]) );
  DFFPOSX1 mem_reg_12__10_ ( .D(n2344), .CLK(clk), .Q(mem[502]) );
  DFFPOSX1 mem_reg_12__9_ ( .D(n2343), .CLK(clk), .Q(mem[501]) );
  DFFPOSX1 mem_reg_12__8_ ( .D(n2342), .CLK(clk), .Q(mem[500]) );
  DFFPOSX1 mem_reg_12__7_ ( .D(n2341), .CLK(clk), .Q(mem[499]) );
  DFFPOSX1 mem_reg_12__6_ ( .D(n2340), .CLK(clk), .Q(mem[498]) );
  DFFPOSX1 mem_reg_12__5_ ( .D(n2339), .CLK(clk), .Q(mem[497]) );
  DFFPOSX1 mem_reg_12__4_ ( .D(n2338), .CLK(clk), .Q(mem[496]) );
  DFFPOSX1 mem_reg_12__3_ ( .D(n2337), .CLK(clk), .Q(mem[495]) );
  DFFPOSX1 mem_reg_12__2_ ( .D(n2336), .CLK(clk), .Q(mem[494]) );
  DFFPOSX1 mem_reg_12__1_ ( .D(n2335), .CLK(clk), .Q(mem[493]) );
  DFFPOSX1 mem_reg_12__0_ ( .D(n2334), .CLK(clk), .Q(mem[492]) );
  DFFPOSX1 mem_reg_11__40_ ( .D(n2333), .CLK(clk), .Q(mem[491]) );
  DFFPOSX1 mem_reg_11__39_ ( .D(n2332), .CLK(clk), .Q(mem[490]) );
  DFFPOSX1 mem_reg_11__38_ ( .D(n2331), .CLK(clk), .Q(mem[489]) );
  DFFPOSX1 mem_reg_11__37_ ( .D(n2330), .CLK(clk), .Q(mem[488]) );
  DFFPOSX1 mem_reg_11__36_ ( .D(n2329), .CLK(clk), .Q(mem[487]) );
  DFFPOSX1 mem_reg_11__35_ ( .D(n2328), .CLK(clk), .Q(mem[486]) );
  DFFPOSX1 mem_reg_11__34_ ( .D(n2327), .CLK(clk), .Q(mem[485]) );
  DFFPOSX1 mem_reg_11__33_ ( .D(n2326), .CLK(clk), .Q(mem[484]) );
  DFFPOSX1 mem_reg_11__32_ ( .D(n2325), .CLK(clk), .Q(mem[483]) );
  DFFPOSX1 mem_reg_11__31_ ( .D(n2324), .CLK(clk), .Q(mem[482]) );
  DFFPOSX1 mem_reg_11__30_ ( .D(n2323), .CLK(clk), .Q(mem[481]) );
  DFFPOSX1 mem_reg_11__29_ ( .D(n2322), .CLK(clk), .Q(mem[480]) );
  DFFPOSX1 mem_reg_11__28_ ( .D(n2321), .CLK(clk), .Q(mem[479]) );
  DFFPOSX1 mem_reg_11__27_ ( .D(n2320), .CLK(clk), .Q(mem[478]) );
  DFFPOSX1 mem_reg_11__26_ ( .D(n2319), .CLK(clk), .Q(mem[477]) );
  DFFPOSX1 mem_reg_11__25_ ( .D(n2318), .CLK(clk), .Q(mem[476]) );
  DFFPOSX1 mem_reg_11__24_ ( .D(n2317), .CLK(clk), .Q(mem[475]) );
  DFFPOSX1 mem_reg_11__23_ ( .D(n2316), .CLK(clk), .Q(mem[474]) );
  DFFPOSX1 mem_reg_11__22_ ( .D(n2315), .CLK(clk), .Q(mem[473]) );
  DFFPOSX1 mem_reg_11__21_ ( .D(n2314), .CLK(clk), .Q(mem[472]) );
  DFFPOSX1 mem_reg_11__20_ ( .D(n2313), .CLK(clk), .Q(mem[471]) );
  DFFPOSX1 mem_reg_11__19_ ( .D(n2312), .CLK(clk), .Q(mem[470]) );
  DFFPOSX1 mem_reg_11__18_ ( .D(n2311), .CLK(clk), .Q(mem[469]) );
  DFFPOSX1 mem_reg_11__17_ ( .D(n2310), .CLK(clk), .Q(mem[468]) );
  DFFPOSX1 mem_reg_11__16_ ( .D(n2309), .CLK(clk), .Q(mem[467]) );
  DFFPOSX1 mem_reg_11__15_ ( .D(n2308), .CLK(clk), .Q(mem[466]) );
  DFFPOSX1 mem_reg_11__14_ ( .D(n2307), .CLK(clk), .Q(mem[465]) );
  DFFPOSX1 mem_reg_11__13_ ( .D(n2306), .CLK(clk), .Q(mem[464]) );
  DFFPOSX1 mem_reg_11__12_ ( .D(n2305), .CLK(clk), .Q(mem[463]) );
  DFFPOSX1 mem_reg_11__11_ ( .D(n2304), .CLK(clk), .Q(mem[462]) );
  DFFPOSX1 mem_reg_11__10_ ( .D(n2303), .CLK(clk), .Q(mem[461]) );
  DFFPOSX1 mem_reg_11__9_ ( .D(n2302), .CLK(clk), .Q(mem[460]) );
  DFFPOSX1 mem_reg_11__8_ ( .D(n2301), .CLK(clk), .Q(mem[459]) );
  DFFPOSX1 mem_reg_11__7_ ( .D(n2300), .CLK(clk), .Q(mem[458]) );
  DFFPOSX1 mem_reg_11__6_ ( .D(n2299), .CLK(clk), .Q(mem[457]) );
  DFFPOSX1 mem_reg_11__5_ ( .D(n2298), .CLK(clk), .Q(mem[456]) );
  DFFPOSX1 mem_reg_11__4_ ( .D(n2297), .CLK(clk), .Q(mem[455]) );
  DFFPOSX1 mem_reg_11__3_ ( .D(n2296), .CLK(clk), .Q(mem[454]) );
  DFFPOSX1 mem_reg_11__2_ ( .D(n2295), .CLK(clk), .Q(mem[453]) );
  DFFPOSX1 mem_reg_11__1_ ( .D(n2294), .CLK(clk), .Q(mem[452]) );
  DFFPOSX1 mem_reg_11__0_ ( .D(n2293), .CLK(clk), .Q(mem[451]) );
  DFFPOSX1 mem_reg_10__40_ ( .D(n2292), .CLK(clk), .Q(mem[450]) );
  DFFPOSX1 mem_reg_10__39_ ( .D(n2291), .CLK(clk), .Q(mem[449]) );
  DFFPOSX1 mem_reg_10__38_ ( .D(n2290), .CLK(clk), .Q(mem[448]) );
  DFFPOSX1 mem_reg_10__37_ ( .D(n2289), .CLK(clk), .Q(mem[447]) );
  DFFPOSX1 mem_reg_10__36_ ( .D(n2288), .CLK(clk), .Q(mem[446]) );
  DFFPOSX1 mem_reg_10__35_ ( .D(n2287), .CLK(clk), .Q(mem[445]) );
  DFFPOSX1 mem_reg_10__34_ ( .D(n2286), .CLK(clk), .Q(mem[444]) );
  DFFPOSX1 mem_reg_10__33_ ( .D(n2285), .CLK(clk), .Q(mem[443]) );
  DFFPOSX1 mem_reg_10__32_ ( .D(n2284), .CLK(clk), .Q(mem[442]) );
  DFFPOSX1 mem_reg_10__31_ ( .D(n2283), .CLK(clk), .Q(mem[441]) );
  DFFPOSX1 mem_reg_10__30_ ( .D(n2282), .CLK(clk), .Q(mem[440]) );
  DFFPOSX1 mem_reg_10__29_ ( .D(n2281), .CLK(clk), .Q(mem[439]) );
  DFFPOSX1 mem_reg_10__28_ ( .D(n2280), .CLK(clk), .Q(mem[438]) );
  DFFPOSX1 mem_reg_10__27_ ( .D(n2279), .CLK(clk), .Q(mem[437]) );
  DFFPOSX1 mem_reg_10__26_ ( .D(n2278), .CLK(clk), .Q(mem[436]) );
  DFFPOSX1 mem_reg_10__25_ ( .D(n2277), .CLK(clk), .Q(mem[435]) );
  DFFPOSX1 mem_reg_10__24_ ( .D(n2276), .CLK(clk), .Q(mem[434]) );
  DFFPOSX1 mem_reg_10__23_ ( .D(n2275), .CLK(clk), .Q(mem[433]) );
  DFFPOSX1 mem_reg_10__22_ ( .D(n2274), .CLK(clk), .Q(mem[432]) );
  DFFPOSX1 mem_reg_10__21_ ( .D(n2273), .CLK(clk), .Q(mem[431]) );
  DFFPOSX1 mem_reg_10__20_ ( .D(n2272), .CLK(clk), .Q(mem[430]) );
  DFFPOSX1 mem_reg_10__19_ ( .D(n2271), .CLK(clk), .Q(mem[429]) );
  DFFPOSX1 mem_reg_10__18_ ( .D(n2270), .CLK(clk), .Q(mem[428]) );
  DFFPOSX1 mem_reg_10__17_ ( .D(n2269), .CLK(clk), .Q(mem[427]) );
  DFFPOSX1 mem_reg_10__16_ ( .D(n2268), .CLK(clk), .Q(mem[426]) );
  DFFPOSX1 mem_reg_10__15_ ( .D(n2267), .CLK(clk), .Q(mem[425]) );
  DFFPOSX1 mem_reg_10__14_ ( .D(n2266), .CLK(clk), .Q(mem[424]) );
  DFFPOSX1 mem_reg_10__13_ ( .D(n2265), .CLK(clk), .Q(mem[423]) );
  DFFPOSX1 mem_reg_10__12_ ( .D(n2264), .CLK(clk), .Q(mem[422]) );
  DFFPOSX1 mem_reg_10__11_ ( .D(n2263), .CLK(clk), .Q(mem[421]) );
  DFFPOSX1 mem_reg_10__10_ ( .D(n2262), .CLK(clk), .Q(mem[420]) );
  DFFPOSX1 mem_reg_10__9_ ( .D(n2261), .CLK(clk), .Q(mem[419]) );
  DFFPOSX1 mem_reg_10__8_ ( .D(n2260), .CLK(clk), .Q(mem[418]) );
  DFFPOSX1 mem_reg_10__7_ ( .D(n2259), .CLK(clk), .Q(mem[417]) );
  DFFPOSX1 mem_reg_10__6_ ( .D(n2258), .CLK(clk), .Q(mem[416]) );
  DFFPOSX1 mem_reg_10__5_ ( .D(n2257), .CLK(clk), .Q(mem[415]) );
  DFFPOSX1 mem_reg_10__4_ ( .D(n2256), .CLK(clk), .Q(mem[414]) );
  DFFPOSX1 mem_reg_10__3_ ( .D(n2255), .CLK(clk), .Q(mem[413]) );
  DFFPOSX1 mem_reg_10__2_ ( .D(n2254), .CLK(clk), .Q(mem[412]) );
  DFFPOSX1 mem_reg_10__1_ ( .D(n2253), .CLK(clk), .Q(mem[411]) );
  DFFPOSX1 mem_reg_10__0_ ( .D(n2252), .CLK(clk), .Q(mem[410]) );
  DFFPOSX1 mem_reg_9__40_ ( .D(n2251), .CLK(clk), .Q(mem[409]) );
  DFFPOSX1 mem_reg_9__39_ ( .D(n2250), .CLK(clk), .Q(mem[408]) );
  DFFPOSX1 mem_reg_9__38_ ( .D(n2249), .CLK(clk), .Q(mem[407]) );
  DFFPOSX1 mem_reg_9__37_ ( .D(n2248), .CLK(clk), .Q(mem[406]) );
  DFFPOSX1 mem_reg_9__36_ ( .D(n2247), .CLK(clk), .Q(mem[405]) );
  DFFPOSX1 mem_reg_9__35_ ( .D(n2246), .CLK(clk), .Q(mem[404]) );
  DFFPOSX1 mem_reg_9__34_ ( .D(n2245), .CLK(clk), .Q(mem[403]) );
  DFFPOSX1 mem_reg_9__33_ ( .D(n2244), .CLK(clk), .Q(mem[402]) );
  DFFPOSX1 mem_reg_9__32_ ( .D(n2243), .CLK(clk), .Q(mem[401]) );
  DFFPOSX1 mem_reg_9__31_ ( .D(n2242), .CLK(clk), .Q(mem[400]) );
  DFFPOSX1 mem_reg_9__30_ ( .D(n2241), .CLK(clk), .Q(mem[399]) );
  DFFPOSX1 mem_reg_9__29_ ( .D(n2240), .CLK(clk), .Q(mem[398]) );
  DFFPOSX1 mem_reg_9__28_ ( .D(n2239), .CLK(clk), .Q(mem[397]) );
  DFFPOSX1 mem_reg_9__27_ ( .D(n2238), .CLK(clk), .Q(mem[396]) );
  DFFPOSX1 mem_reg_9__26_ ( .D(n2237), .CLK(clk), .Q(mem[395]) );
  DFFPOSX1 mem_reg_9__25_ ( .D(n2236), .CLK(clk), .Q(mem[394]) );
  DFFPOSX1 mem_reg_9__24_ ( .D(n2235), .CLK(clk), .Q(mem[393]) );
  DFFPOSX1 mem_reg_9__23_ ( .D(n2234), .CLK(clk), .Q(mem[392]) );
  DFFPOSX1 mem_reg_9__22_ ( .D(n2233), .CLK(clk), .Q(mem[391]) );
  DFFPOSX1 mem_reg_9__21_ ( .D(n2232), .CLK(clk), .Q(mem[390]) );
  DFFPOSX1 mem_reg_9__20_ ( .D(n2231), .CLK(clk), .Q(mem[389]) );
  DFFPOSX1 mem_reg_9__19_ ( .D(n2230), .CLK(clk), .Q(mem[388]) );
  DFFPOSX1 mem_reg_9__18_ ( .D(n2229), .CLK(clk), .Q(mem[387]) );
  DFFPOSX1 mem_reg_9__17_ ( .D(n2228), .CLK(clk), .Q(mem[386]) );
  DFFPOSX1 mem_reg_9__16_ ( .D(n2227), .CLK(clk), .Q(mem[385]) );
  DFFPOSX1 mem_reg_9__15_ ( .D(n2226), .CLK(clk), .Q(mem[384]) );
  DFFPOSX1 mem_reg_9__14_ ( .D(n2225), .CLK(clk), .Q(mem[383]) );
  DFFPOSX1 mem_reg_9__13_ ( .D(n2224), .CLK(clk), .Q(mem[382]) );
  DFFPOSX1 mem_reg_9__12_ ( .D(n2223), .CLK(clk), .Q(mem[381]) );
  DFFPOSX1 mem_reg_9__11_ ( .D(n2222), .CLK(clk), .Q(mem[380]) );
  DFFPOSX1 mem_reg_9__10_ ( .D(n2221), .CLK(clk), .Q(mem[379]) );
  DFFPOSX1 mem_reg_9__9_ ( .D(n2220), .CLK(clk), .Q(mem[378]) );
  DFFPOSX1 mem_reg_9__8_ ( .D(n2219), .CLK(clk), .Q(mem[377]) );
  DFFPOSX1 mem_reg_9__7_ ( .D(n2218), .CLK(clk), .Q(mem[376]) );
  DFFPOSX1 mem_reg_9__6_ ( .D(n2217), .CLK(clk), .Q(mem[375]) );
  DFFPOSX1 mem_reg_9__5_ ( .D(n2216), .CLK(clk), .Q(mem[374]) );
  DFFPOSX1 mem_reg_9__4_ ( .D(n2215), .CLK(clk), .Q(mem[373]) );
  DFFPOSX1 mem_reg_9__3_ ( .D(n2214), .CLK(clk), .Q(mem[372]) );
  DFFPOSX1 mem_reg_9__2_ ( .D(n2213), .CLK(clk), .Q(mem[371]) );
  DFFPOSX1 mem_reg_9__1_ ( .D(n2212), .CLK(clk), .Q(mem[370]) );
  DFFPOSX1 mem_reg_9__0_ ( .D(n2211), .CLK(clk), .Q(mem[369]) );
  DFFPOSX1 mem_reg_8__40_ ( .D(n2210), .CLK(clk), .Q(mem[368]) );
  DFFPOSX1 mem_reg_8__39_ ( .D(n2209), .CLK(clk), .Q(mem[367]) );
  DFFPOSX1 mem_reg_8__38_ ( .D(n2208), .CLK(clk), .Q(mem[366]) );
  DFFPOSX1 mem_reg_8__37_ ( .D(n2207), .CLK(clk), .Q(mem[365]) );
  DFFPOSX1 mem_reg_8__36_ ( .D(n2206), .CLK(clk), .Q(mem[364]) );
  DFFPOSX1 mem_reg_8__35_ ( .D(n2205), .CLK(clk), .Q(mem[363]) );
  DFFPOSX1 mem_reg_8__34_ ( .D(n2204), .CLK(clk), .Q(mem[362]) );
  DFFPOSX1 mem_reg_8__33_ ( .D(n2203), .CLK(clk), .Q(mem[361]) );
  DFFPOSX1 mem_reg_8__32_ ( .D(n2202), .CLK(clk), .Q(mem[360]) );
  DFFPOSX1 mem_reg_8__31_ ( .D(n2201), .CLK(clk), .Q(mem[359]) );
  DFFPOSX1 mem_reg_8__30_ ( .D(n2200), .CLK(clk), .Q(mem[358]) );
  DFFPOSX1 mem_reg_8__29_ ( .D(n2199), .CLK(clk), .Q(mem[357]) );
  DFFPOSX1 mem_reg_8__28_ ( .D(n2198), .CLK(clk), .Q(mem[356]) );
  DFFPOSX1 mem_reg_8__27_ ( .D(n2197), .CLK(clk), .Q(mem[355]) );
  DFFPOSX1 mem_reg_8__26_ ( .D(n2196), .CLK(clk), .Q(mem[354]) );
  DFFPOSX1 mem_reg_8__25_ ( .D(n2195), .CLK(clk), .Q(mem[353]) );
  DFFPOSX1 mem_reg_8__24_ ( .D(n2194), .CLK(clk), .Q(mem[352]) );
  DFFPOSX1 mem_reg_8__23_ ( .D(n2193), .CLK(clk), .Q(mem[351]) );
  DFFPOSX1 mem_reg_8__22_ ( .D(n2192), .CLK(clk), .Q(mem[350]) );
  DFFPOSX1 mem_reg_8__21_ ( .D(n2191), .CLK(clk), .Q(mem[349]) );
  DFFPOSX1 mem_reg_8__20_ ( .D(n2190), .CLK(clk), .Q(mem[348]) );
  DFFPOSX1 mem_reg_8__19_ ( .D(n2189), .CLK(clk), .Q(mem[347]) );
  DFFPOSX1 mem_reg_8__18_ ( .D(n2188), .CLK(clk), .Q(mem[346]) );
  DFFPOSX1 mem_reg_8__17_ ( .D(n2187), .CLK(clk), .Q(mem[345]) );
  DFFPOSX1 mem_reg_8__16_ ( .D(n2186), .CLK(clk), .Q(mem[344]) );
  DFFPOSX1 mem_reg_8__15_ ( .D(n2185), .CLK(clk), .Q(mem[343]) );
  DFFPOSX1 mem_reg_8__14_ ( .D(n2184), .CLK(clk), .Q(mem[342]) );
  DFFPOSX1 mem_reg_8__13_ ( .D(n2183), .CLK(clk), .Q(mem[341]) );
  DFFPOSX1 mem_reg_8__12_ ( .D(n2182), .CLK(clk), .Q(mem[340]) );
  DFFPOSX1 mem_reg_8__11_ ( .D(n2181), .CLK(clk), .Q(mem[339]) );
  DFFPOSX1 mem_reg_8__10_ ( .D(n2180), .CLK(clk), .Q(mem[338]) );
  DFFPOSX1 mem_reg_8__9_ ( .D(n2179), .CLK(clk), .Q(mem[337]) );
  DFFPOSX1 mem_reg_8__8_ ( .D(n2178), .CLK(clk), .Q(mem[336]) );
  DFFPOSX1 mem_reg_8__7_ ( .D(n2177), .CLK(clk), .Q(mem[335]) );
  DFFPOSX1 mem_reg_8__6_ ( .D(n2176), .CLK(clk), .Q(mem[334]) );
  DFFPOSX1 mem_reg_8__5_ ( .D(n2175), .CLK(clk), .Q(mem[333]) );
  DFFPOSX1 mem_reg_8__4_ ( .D(n2174), .CLK(clk), .Q(mem[332]) );
  DFFPOSX1 mem_reg_8__3_ ( .D(n2173), .CLK(clk), .Q(mem[331]) );
  DFFPOSX1 mem_reg_8__2_ ( .D(n2172), .CLK(clk), .Q(mem[330]) );
  DFFPOSX1 mem_reg_8__1_ ( .D(n2171), .CLK(clk), .Q(mem[329]) );
  DFFPOSX1 mem_reg_8__0_ ( .D(n2170), .CLK(clk), .Q(mem[328]) );
  DFFPOSX1 mem_reg_7__40_ ( .D(n2169), .CLK(clk), .Q(mem[327]) );
  DFFPOSX1 mem_reg_7__39_ ( .D(n2168), .CLK(clk), .Q(mem[326]) );
  DFFPOSX1 mem_reg_7__38_ ( .D(n2167), .CLK(clk), .Q(mem[325]) );
  DFFPOSX1 mem_reg_7__37_ ( .D(n2166), .CLK(clk), .Q(mem[324]) );
  DFFPOSX1 mem_reg_7__36_ ( .D(n2165), .CLK(clk), .Q(mem[323]) );
  DFFPOSX1 mem_reg_7__35_ ( .D(n2164), .CLK(clk), .Q(mem[322]) );
  DFFPOSX1 mem_reg_7__34_ ( .D(n2163), .CLK(clk), .Q(mem[321]) );
  DFFPOSX1 mem_reg_7__33_ ( .D(n2162), .CLK(clk), .Q(mem[320]) );
  DFFPOSX1 mem_reg_7__32_ ( .D(n2161), .CLK(clk), .Q(mem[319]) );
  DFFPOSX1 mem_reg_7__31_ ( .D(n2160), .CLK(clk), .Q(mem[318]) );
  DFFPOSX1 mem_reg_7__30_ ( .D(n2159), .CLK(clk), .Q(mem[317]) );
  DFFPOSX1 mem_reg_7__29_ ( .D(n2158), .CLK(clk), .Q(mem[316]) );
  DFFPOSX1 mem_reg_7__28_ ( .D(n2157), .CLK(clk), .Q(mem[315]) );
  DFFPOSX1 mem_reg_7__27_ ( .D(n2156), .CLK(clk), .Q(mem[314]) );
  DFFPOSX1 mem_reg_7__26_ ( .D(n2155), .CLK(clk), .Q(mem[313]) );
  DFFPOSX1 mem_reg_7__25_ ( .D(n2154), .CLK(clk), .Q(mem[312]) );
  DFFPOSX1 mem_reg_7__24_ ( .D(n2153), .CLK(clk), .Q(mem[311]) );
  DFFPOSX1 mem_reg_7__23_ ( .D(n2152), .CLK(clk), .Q(mem[310]) );
  DFFPOSX1 mem_reg_7__22_ ( .D(n2151), .CLK(clk), .Q(mem[309]) );
  DFFPOSX1 mem_reg_7__21_ ( .D(n2150), .CLK(clk), .Q(mem[308]) );
  DFFPOSX1 mem_reg_7__20_ ( .D(n2149), .CLK(clk), .Q(mem[307]) );
  DFFPOSX1 mem_reg_7__19_ ( .D(n2148), .CLK(clk), .Q(mem[306]) );
  DFFPOSX1 mem_reg_7__18_ ( .D(n2147), .CLK(clk), .Q(mem[305]) );
  DFFPOSX1 mem_reg_7__17_ ( .D(n2146), .CLK(clk), .Q(mem[304]) );
  DFFPOSX1 mem_reg_7__16_ ( .D(n2145), .CLK(clk), .Q(mem[303]) );
  DFFPOSX1 mem_reg_7__15_ ( .D(n2144), .CLK(clk), .Q(mem[302]) );
  DFFPOSX1 mem_reg_7__14_ ( .D(n2143), .CLK(clk), .Q(mem[301]) );
  DFFPOSX1 mem_reg_7__13_ ( .D(n2142), .CLK(clk), .Q(mem[300]) );
  DFFPOSX1 mem_reg_7__12_ ( .D(n2141), .CLK(clk), .Q(mem[299]) );
  DFFPOSX1 mem_reg_7__11_ ( .D(n2140), .CLK(clk), .Q(mem[298]) );
  DFFPOSX1 mem_reg_7__10_ ( .D(n2139), .CLK(clk), .Q(mem[297]) );
  DFFPOSX1 mem_reg_7__9_ ( .D(n2138), .CLK(clk), .Q(mem[296]) );
  DFFPOSX1 mem_reg_7__8_ ( .D(n2137), .CLK(clk), .Q(mem[295]) );
  DFFPOSX1 mem_reg_7__7_ ( .D(n2136), .CLK(clk), .Q(mem[294]) );
  DFFPOSX1 mem_reg_7__6_ ( .D(n2135), .CLK(clk), .Q(mem[293]) );
  DFFPOSX1 mem_reg_7__5_ ( .D(n2134), .CLK(clk), .Q(mem[292]) );
  DFFPOSX1 mem_reg_7__4_ ( .D(n2133), .CLK(clk), .Q(mem[291]) );
  DFFPOSX1 mem_reg_7__3_ ( .D(n2132), .CLK(clk), .Q(mem[290]) );
  DFFPOSX1 mem_reg_7__2_ ( .D(n2131), .CLK(clk), .Q(mem[289]) );
  DFFPOSX1 mem_reg_7__1_ ( .D(n2130), .CLK(clk), .Q(mem[288]) );
  DFFPOSX1 mem_reg_7__0_ ( .D(n2129), .CLK(clk), .Q(mem[287]) );
  DFFPOSX1 mem_reg_6__40_ ( .D(n2128), .CLK(clk), .Q(mem[286]) );
  DFFPOSX1 mem_reg_6__39_ ( .D(n2127), .CLK(clk), .Q(mem[285]) );
  DFFPOSX1 mem_reg_6__38_ ( .D(n2126), .CLK(clk), .Q(mem[284]) );
  DFFPOSX1 mem_reg_6__37_ ( .D(n2125), .CLK(clk), .Q(mem[283]) );
  DFFPOSX1 mem_reg_6__36_ ( .D(n2124), .CLK(clk), .Q(mem[282]) );
  DFFPOSX1 mem_reg_6__35_ ( .D(n2123), .CLK(clk), .Q(mem[281]) );
  DFFPOSX1 mem_reg_6__34_ ( .D(n2122), .CLK(clk), .Q(mem[280]) );
  DFFPOSX1 mem_reg_6__33_ ( .D(n2121), .CLK(clk), .Q(mem[279]) );
  DFFPOSX1 mem_reg_6__32_ ( .D(n2120), .CLK(clk), .Q(mem[278]) );
  DFFPOSX1 mem_reg_6__31_ ( .D(n2119), .CLK(clk), .Q(mem[277]) );
  DFFPOSX1 mem_reg_6__30_ ( .D(n2118), .CLK(clk), .Q(mem[276]) );
  DFFPOSX1 mem_reg_6__29_ ( .D(n2117), .CLK(clk), .Q(mem[275]) );
  DFFPOSX1 mem_reg_6__28_ ( .D(n2116), .CLK(clk), .Q(mem[274]) );
  DFFPOSX1 mem_reg_6__27_ ( .D(n2115), .CLK(clk), .Q(mem[273]) );
  DFFPOSX1 mem_reg_6__26_ ( .D(n2114), .CLK(clk), .Q(mem[272]) );
  DFFPOSX1 mem_reg_6__25_ ( .D(n2113), .CLK(clk), .Q(mem[271]) );
  DFFPOSX1 mem_reg_6__24_ ( .D(n2112), .CLK(clk), .Q(mem[270]) );
  DFFPOSX1 mem_reg_6__23_ ( .D(n2111), .CLK(clk), .Q(mem[269]) );
  DFFPOSX1 mem_reg_6__22_ ( .D(n2110), .CLK(clk), .Q(mem[268]) );
  DFFPOSX1 mem_reg_6__21_ ( .D(n2109), .CLK(clk), .Q(mem[267]) );
  DFFPOSX1 mem_reg_6__20_ ( .D(n2108), .CLK(clk), .Q(mem[266]) );
  DFFPOSX1 mem_reg_6__19_ ( .D(n2107), .CLK(clk), .Q(mem[265]) );
  DFFPOSX1 mem_reg_6__18_ ( .D(n2106), .CLK(clk), .Q(mem[264]) );
  DFFPOSX1 mem_reg_6__17_ ( .D(n2105), .CLK(clk), .Q(mem[263]) );
  DFFPOSX1 mem_reg_6__16_ ( .D(n2104), .CLK(clk), .Q(mem[262]) );
  DFFPOSX1 mem_reg_6__15_ ( .D(n2103), .CLK(clk), .Q(mem[261]) );
  DFFPOSX1 mem_reg_6__14_ ( .D(n2102), .CLK(clk), .Q(mem[260]) );
  DFFPOSX1 mem_reg_6__13_ ( .D(n2101), .CLK(clk), .Q(mem[259]) );
  DFFPOSX1 mem_reg_6__12_ ( .D(n2100), .CLK(clk), .Q(mem[258]) );
  DFFPOSX1 mem_reg_6__11_ ( .D(n2099), .CLK(clk), .Q(mem[257]) );
  DFFPOSX1 mem_reg_6__10_ ( .D(n2098), .CLK(clk), .Q(mem[256]) );
  DFFPOSX1 mem_reg_6__9_ ( .D(n2097), .CLK(clk), .Q(mem[255]) );
  DFFPOSX1 mem_reg_6__8_ ( .D(n2096), .CLK(clk), .Q(mem[254]) );
  DFFPOSX1 mem_reg_6__7_ ( .D(n2095), .CLK(clk), .Q(mem[253]) );
  DFFPOSX1 mem_reg_6__6_ ( .D(n2094), .CLK(clk), .Q(mem[252]) );
  DFFPOSX1 mem_reg_6__5_ ( .D(n2093), .CLK(clk), .Q(mem[251]) );
  DFFPOSX1 mem_reg_6__4_ ( .D(n2092), .CLK(clk), .Q(mem[250]) );
  DFFPOSX1 mem_reg_6__3_ ( .D(n2091), .CLK(clk), .Q(mem[249]) );
  DFFPOSX1 mem_reg_6__2_ ( .D(n2090), .CLK(clk), .Q(mem[248]) );
  DFFPOSX1 mem_reg_6__1_ ( .D(n2089), .CLK(clk), .Q(mem[247]) );
  DFFPOSX1 mem_reg_6__0_ ( .D(n2088), .CLK(clk), .Q(mem[246]) );
  DFFPOSX1 mem_reg_5__40_ ( .D(n2087), .CLK(clk), .Q(mem[245]) );
  DFFPOSX1 mem_reg_5__39_ ( .D(n2086), .CLK(clk), .Q(mem[244]) );
  DFFPOSX1 mem_reg_5__38_ ( .D(n2085), .CLK(clk), .Q(mem[243]) );
  DFFPOSX1 mem_reg_5__37_ ( .D(n2084), .CLK(clk), .Q(mem[242]) );
  DFFPOSX1 mem_reg_5__36_ ( .D(n2083), .CLK(clk), .Q(mem[241]) );
  DFFPOSX1 mem_reg_5__35_ ( .D(n2082), .CLK(clk), .Q(mem[240]) );
  DFFPOSX1 mem_reg_5__34_ ( .D(n2081), .CLK(clk), .Q(mem[239]) );
  DFFPOSX1 mem_reg_5__33_ ( .D(n2080), .CLK(clk), .Q(mem[238]) );
  DFFPOSX1 mem_reg_5__32_ ( .D(n2079), .CLK(clk), .Q(mem[237]) );
  DFFPOSX1 mem_reg_5__31_ ( .D(n2078), .CLK(clk), .Q(mem[236]) );
  DFFPOSX1 mem_reg_5__30_ ( .D(n2077), .CLK(clk), .Q(mem[235]) );
  DFFPOSX1 mem_reg_5__29_ ( .D(n2076), .CLK(clk), .Q(mem[234]) );
  DFFPOSX1 mem_reg_5__28_ ( .D(n2075), .CLK(clk), .Q(mem[233]) );
  DFFPOSX1 mem_reg_5__27_ ( .D(n2074), .CLK(clk), .Q(mem[232]) );
  DFFPOSX1 mem_reg_5__26_ ( .D(n2073), .CLK(clk), .Q(mem[231]) );
  DFFPOSX1 mem_reg_5__25_ ( .D(n2072), .CLK(clk), .Q(mem[230]) );
  DFFPOSX1 mem_reg_5__24_ ( .D(n2071), .CLK(clk), .Q(mem[229]) );
  DFFPOSX1 mem_reg_5__23_ ( .D(n2070), .CLK(clk), .Q(mem[228]) );
  DFFPOSX1 mem_reg_5__22_ ( .D(n2069), .CLK(clk), .Q(mem[227]) );
  DFFPOSX1 mem_reg_5__21_ ( .D(n2068), .CLK(clk), .Q(mem[226]) );
  DFFPOSX1 mem_reg_5__20_ ( .D(n2067), .CLK(clk), .Q(mem[225]) );
  DFFPOSX1 mem_reg_5__19_ ( .D(n2066), .CLK(clk), .Q(mem[224]) );
  DFFPOSX1 mem_reg_5__18_ ( .D(n2065), .CLK(clk), .Q(mem[223]) );
  DFFPOSX1 mem_reg_5__17_ ( .D(n2064), .CLK(clk), .Q(mem[222]) );
  DFFPOSX1 mem_reg_5__16_ ( .D(n2063), .CLK(clk), .Q(mem[221]) );
  DFFPOSX1 mem_reg_5__15_ ( .D(n2062), .CLK(clk), .Q(mem[220]) );
  DFFPOSX1 mem_reg_5__14_ ( .D(n2061), .CLK(clk), .Q(mem[219]) );
  DFFPOSX1 mem_reg_5__13_ ( .D(n2060), .CLK(clk), .Q(mem[218]) );
  DFFPOSX1 mem_reg_5__12_ ( .D(n2059), .CLK(clk), .Q(mem[217]) );
  DFFPOSX1 mem_reg_5__11_ ( .D(n2058), .CLK(clk), .Q(mem[216]) );
  DFFPOSX1 mem_reg_5__10_ ( .D(n2057), .CLK(clk), .Q(mem[215]) );
  DFFPOSX1 mem_reg_5__9_ ( .D(n2056), .CLK(clk), .Q(mem[214]) );
  DFFPOSX1 mem_reg_5__8_ ( .D(n2055), .CLK(clk), .Q(mem[213]) );
  DFFPOSX1 mem_reg_5__7_ ( .D(n2054), .CLK(clk), .Q(mem[212]) );
  DFFPOSX1 mem_reg_5__6_ ( .D(n2053), .CLK(clk), .Q(mem[211]) );
  DFFPOSX1 mem_reg_5__5_ ( .D(n2052), .CLK(clk), .Q(mem[210]) );
  DFFPOSX1 mem_reg_5__4_ ( .D(n2051), .CLK(clk), .Q(mem[209]) );
  DFFPOSX1 mem_reg_5__3_ ( .D(n2050), .CLK(clk), .Q(mem[208]) );
  DFFPOSX1 mem_reg_5__2_ ( .D(n2049), .CLK(clk), .Q(mem[207]) );
  DFFPOSX1 mem_reg_5__1_ ( .D(n2048), .CLK(clk), .Q(mem[206]) );
  DFFPOSX1 mem_reg_5__0_ ( .D(n2047), .CLK(clk), .Q(mem[205]) );
  DFFPOSX1 mem_reg_4__40_ ( .D(n2046), .CLK(clk), .Q(mem[204]) );
  DFFPOSX1 mem_reg_4__39_ ( .D(n2045), .CLK(clk), .Q(mem[203]) );
  DFFPOSX1 mem_reg_4__38_ ( .D(n2044), .CLK(clk), .Q(mem[202]) );
  DFFPOSX1 mem_reg_4__37_ ( .D(n2043), .CLK(clk), .Q(mem[201]) );
  DFFPOSX1 mem_reg_4__36_ ( .D(n2042), .CLK(clk), .Q(mem[200]) );
  DFFPOSX1 mem_reg_4__35_ ( .D(n2041), .CLK(clk), .Q(mem[199]) );
  DFFPOSX1 mem_reg_4__34_ ( .D(n2040), .CLK(clk), .Q(mem[198]) );
  DFFPOSX1 mem_reg_4__33_ ( .D(n2039), .CLK(clk), .Q(mem[197]) );
  DFFPOSX1 mem_reg_4__32_ ( .D(n2038), .CLK(clk), .Q(mem[196]) );
  DFFPOSX1 mem_reg_4__31_ ( .D(n2037), .CLK(clk), .Q(mem[195]) );
  DFFPOSX1 mem_reg_4__30_ ( .D(n2036), .CLK(clk), .Q(mem[194]) );
  DFFPOSX1 mem_reg_4__29_ ( .D(n2035), .CLK(clk), .Q(mem[193]) );
  DFFPOSX1 mem_reg_4__28_ ( .D(n2034), .CLK(clk), .Q(mem[192]) );
  DFFPOSX1 mem_reg_4__27_ ( .D(n2033), .CLK(clk), .Q(mem[191]) );
  DFFPOSX1 mem_reg_4__26_ ( .D(n2032), .CLK(clk), .Q(mem[190]) );
  DFFPOSX1 mem_reg_4__25_ ( .D(n2031), .CLK(clk), .Q(mem[189]) );
  DFFPOSX1 mem_reg_4__24_ ( .D(n2030), .CLK(clk), .Q(mem[188]) );
  DFFPOSX1 mem_reg_4__23_ ( .D(n2029), .CLK(clk), .Q(mem[187]) );
  DFFPOSX1 mem_reg_4__22_ ( .D(n2028), .CLK(clk), .Q(mem[186]) );
  DFFPOSX1 mem_reg_4__21_ ( .D(n2027), .CLK(clk), .Q(mem[185]) );
  DFFPOSX1 mem_reg_4__20_ ( .D(n2026), .CLK(clk), .Q(mem[184]) );
  DFFPOSX1 mem_reg_4__19_ ( .D(n2025), .CLK(clk), .Q(mem[183]) );
  DFFPOSX1 mem_reg_4__18_ ( .D(n2024), .CLK(clk), .Q(mem[182]) );
  DFFPOSX1 mem_reg_4__17_ ( .D(n2023), .CLK(clk), .Q(mem[181]) );
  DFFPOSX1 mem_reg_4__16_ ( .D(n2022), .CLK(clk), .Q(mem[180]) );
  DFFPOSX1 mem_reg_4__15_ ( .D(n2021), .CLK(clk), .Q(mem[179]) );
  DFFPOSX1 mem_reg_4__14_ ( .D(n2020), .CLK(clk), .Q(mem[178]) );
  DFFPOSX1 mem_reg_4__13_ ( .D(n2019), .CLK(clk), .Q(mem[177]) );
  DFFPOSX1 mem_reg_4__12_ ( .D(n2018), .CLK(clk), .Q(mem[176]) );
  DFFPOSX1 mem_reg_4__11_ ( .D(n2017), .CLK(clk), .Q(mem[175]) );
  DFFPOSX1 mem_reg_4__10_ ( .D(n2016), .CLK(clk), .Q(mem[174]) );
  DFFPOSX1 mem_reg_4__9_ ( .D(n2015), .CLK(clk), .Q(mem[173]) );
  DFFPOSX1 mem_reg_4__8_ ( .D(n2014), .CLK(clk), .Q(mem[172]) );
  DFFPOSX1 mem_reg_4__7_ ( .D(n2013), .CLK(clk), .Q(mem[171]) );
  DFFPOSX1 mem_reg_4__6_ ( .D(n2012), .CLK(clk), .Q(mem[170]) );
  DFFPOSX1 mem_reg_4__5_ ( .D(n2011), .CLK(clk), .Q(mem[169]) );
  DFFPOSX1 mem_reg_4__4_ ( .D(n2010), .CLK(clk), .Q(mem[168]) );
  DFFPOSX1 mem_reg_4__3_ ( .D(n2009), .CLK(clk), .Q(mem[167]) );
  DFFPOSX1 mem_reg_4__2_ ( .D(n2008), .CLK(clk), .Q(mem[166]) );
  DFFPOSX1 mem_reg_4__1_ ( .D(n2007), .CLK(clk), .Q(mem[165]) );
  DFFPOSX1 mem_reg_4__0_ ( .D(n2006), .CLK(clk), .Q(mem[164]) );
  DFFPOSX1 mem_reg_3__40_ ( .D(n2005), .CLK(clk), .Q(mem[163]) );
  DFFPOSX1 mem_reg_3__39_ ( .D(n2004), .CLK(clk), .Q(mem[162]) );
  DFFPOSX1 mem_reg_3__38_ ( .D(n2003), .CLK(clk), .Q(mem[161]) );
  DFFPOSX1 mem_reg_3__37_ ( .D(n2002), .CLK(clk), .Q(mem[160]) );
  DFFPOSX1 mem_reg_3__36_ ( .D(n2001), .CLK(clk), .Q(mem[159]) );
  DFFPOSX1 mem_reg_3__35_ ( .D(n2000), .CLK(clk), .Q(mem[158]) );
  DFFPOSX1 mem_reg_3__34_ ( .D(n1999), .CLK(clk), .Q(mem[157]) );
  DFFPOSX1 mem_reg_3__33_ ( .D(n1998), .CLK(clk), .Q(mem[156]) );
  DFFPOSX1 mem_reg_3__32_ ( .D(n1997), .CLK(clk), .Q(mem[155]) );
  DFFPOSX1 mem_reg_3__31_ ( .D(n1996), .CLK(clk), .Q(mem[154]) );
  DFFPOSX1 mem_reg_3__30_ ( .D(n1995), .CLK(clk), .Q(mem[153]) );
  DFFPOSX1 mem_reg_3__29_ ( .D(n1994), .CLK(clk), .Q(mem[152]) );
  DFFPOSX1 mem_reg_3__28_ ( .D(n1993), .CLK(clk), .Q(mem[151]) );
  DFFPOSX1 mem_reg_3__27_ ( .D(n1992), .CLK(clk), .Q(mem[150]) );
  DFFPOSX1 mem_reg_3__26_ ( .D(n1991), .CLK(clk), .Q(mem[149]) );
  DFFPOSX1 mem_reg_3__25_ ( .D(n1990), .CLK(clk), .Q(mem[148]) );
  DFFPOSX1 mem_reg_3__24_ ( .D(n1989), .CLK(clk), .Q(mem[147]) );
  DFFPOSX1 mem_reg_3__23_ ( .D(n1988), .CLK(clk), .Q(mem[146]) );
  DFFPOSX1 mem_reg_3__22_ ( .D(n1987), .CLK(clk), .Q(mem[145]) );
  DFFPOSX1 mem_reg_3__21_ ( .D(n1986), .CLK(clk), .Q(mem[144]) );
  DFFPOSX1 mem_reg_3__20_ ( .D(n1985), .CLK(clk), .Q(mem[143]) );
  DFFPOSX1 mem_reg_3__19_ ( .D(n1984), .CLK(clk), .Q(mem[142]) );
  DFFPOSX1 mem_reg_3__18_ ( .D(n1983), .CLK(clk), .Q(mem[141]) );
  DFFPOSX1 mem_reg_3__17_ ( .D(n1982), .CLK(clk), .Q(mem[140]) );
  DFFPOSX1 mem_reg_3__16_ ( .D(n1981), .CLK(clk), .Q(mem[139]) );
  DFFPOSX1 mem_reg_3__15_ ( .D(n1980), .CLK(clk), .Q(mem[138]) );
  DFFPOSX1 mem_reg_3__14_ ( .D(n1979), .CLK(clk), .Q(mem[137]) );
  DFFPOSX1 mem_reg_3__13_ ( .D(n1978), .CLK(clk), .Q(mem[136]) );
  DFFPOSX1 mem_reg_3__12_ ( .D(n1977), .CLK(clk), .Q(mem[135]) );
  DFFPOSX1 mem_reg_3__11_ ( .D(n1976), .CLK(clk), .Q(mem[134]) );
  DFFPOSX1 mem_reg_3__10_ ( .D(n1975), .CLK(clk), .Q(mem[133]) );
  DFFPOSX1 mem_reg_3__9_ ( .D(n1974), .CLK(clk), .Q(mem[132]) );
  DFFPOSX1 mem_reg_3__8_ ( .D(n1973), .CLK(clk), .Q(mem[131]) );
  DFFPOSX1 mem_reg_3__7_ ( .D(n1972), .CLK(clk), .Q(mem[130]) );
  DFFPOSX1 mem_reg_3__6_ ( .D(n1971), .CLK(clk), .Q(mem[129]) );
  DFFPOSX1 mem_reg_3__5_ ( .D(n1970), .CLK(clk), .Q(mem[128]) );
  DFFPOSX1 mem_reg_3__4_ ( .D(n1969), .CLK(clk), .Q(mem[127]) );
  DFFPOSX1 mem_reg_3__3_ ( .D(n1968), .CLK(clk), .Q(mem[126]) );
  DFFPOSX1 mem_reg_3__2_ ( .D(n1967), .CLK(clk), .Q(mem[125]) );
  DFFPOSX1 mem_reg_3__1_ ( .D(n1966), .CLK(clk), .Q(mem[124]) );
  DFFPOSX1 mem_reg_3__0_ ( .D(n1965), .CLK(clk), .Q(mem[123]) );
  DFFPOSX1 mem_reg_2__40_ ( .D(n1964), .CLK(clk), .Q(mem[122]) );
  DFFPOSX1 mem_reg_2__39_ ( .D(n1963), .CLK(clk), .Q(mem[121]) );
  DFFPOSX1 mem_reg_2__38_ ( .D(n1962), .CLK(clk), .Q(mem[120]) );
  DFFPOSX1 mem_reg_2__37_ ( .D(n1961), .CLK(clk), .Q(mem[119]) );
  DFFPOSX1 mem_reg_2__36_ ( .D(n1960), .CLK(clk), .Q(mem[118]) );
  DFFPOSX1 mem_reg_2__35_ ( .D(n1959), .CLK(clk), .Q(mem[117]) );
  DFFPOSX1 mem_reg_2__34_ ( .D(n1958), .CLK(clk), .Q(mem[116]) );
  DFFPOSX1 mem_reg_2__33_ ( .D(n1957), .CLK(clk), .Q(mem[115]) );
  DFFPOSX1 mem_reg_2__32_ ( .D(n1956), .CLK(clk), .Q(mem[114]) );
  DFFPOSX1 mem_reg_2__31_ ( .D(n1955), .CLK(clk), .Q(mem[113]) );
  DFFPOSX1 mem_reg_2__30_ ( .D(n1954), .CLK(clk), .Q(mem[112]) );
  DFFPOSX1 mem_reg_2__29_ ( .D(n1953), .CLK(clk), .Q(mem[111]) );
  DFFPOSX1 mem_reg_2__28_ ( .D(n1952), .CLK(clk), .Q(mem[110]) );
  DFFPOSX1 mem_reg_2__27_ ( .D(n1951), .CLK(clk), .Q(mem[109]) );
  DFFPOSX1 mem_reg_2__26_ ( .D(n1950), .CLK(clk), .Q(mem[108]) );
  DFFPOSX1 mem_reg_2__25_ ( .D(n1949), .CLK(clk), .Q(mem[107]) );
  DFFPOSX1 mem_reg_2__24_ ( .D(n1948), .CLK(clk), .Q(mem[106]) );
  DFFPOSX1 mem_reg_2__23_ ( .D(n1947), .CLK(clk), .Q(mem[105]) );
  DFFPOSX1 mem_reg_2__22_ ( .D(n1946), .CLK(clk), .Q(mem[104]) );
  DFFPOSX1 mem_reg_2__21_ ( .D(n1945), .CLK(clk), .Q(mem[103]) );
  DFFPOSX1 mem_reg_2__20_ ( .D(n1944), .CLK(clk), .Q(mem[102]) );
  DFFPOSX1 mem_reg_2__19_ ( .D(n1943), .CLK(clk), .Q(mem[101]) );
  DFFPOSX1 mem_reg_2__18_ ( .D(n1942), .CLK(clk), .Q(mem[100]) );
  DFFPOSX1 mem_reg_2__17_ ( .D(n1941), .CLK(clk), .Q(mem[99]) );
  DFFPOSX1 mem_reg_2__16_ ( .D(n1940), .CLK(clk), .Q(mem[98]) );
  DFFPOSX1 mem_reg_2__15_ ( .D(n1939), .CLK(clk), .Q(mem[97]) );
  DFFPOSX1 mem_reg_2__14_ ( .D(n1938), .CLK(clk), .Q(mem[96]) );
  DFFPOSX1 mem_reg_2__13_ ( .D(n1937), .CLK(clk), .Q(mem[95]) );
  DFFPOSX1 mem_reg_2__12_ ( .D(n1936), .CLK(clk), .Q(mem[94]) );
  DFFPOSX1 mem_reg_2__11_ ( .D(n1935), .CLK(clk), .Q(mem[93]) );
  DFFPOSX1 mem_reg_2__10_ ( .D(n1934), .CLK(clk), .Q(mem[92]) );
  DFFPOSX1 mem_reg_2__9_ ( .D(n1933), .CLK(clk), .Q(mem[91]) );
  DFFPOSX1 mem_reg_2__8_ ( .D(n1932), .CLK(clk), .Q(mem[90]) );
  DFFPOSX1 mem_reg_2__7_ ( .D(n1931), .CLK(clk), .Q(mem[89]) );
  DFFPOSX1 mem_reg_2__6_ ( .D(n1930), .CLK(clk), .Q(mem[88]) );
  DFFPOSX1 mem_reg_2__5_ ( .D(n1929), .CLK(clk), .Q(mem[87]) );
  DFFPOSX1 mem_reg_2__4_ ( .D(n1928), .CLK(clk), .Q(mem[86]) );
  DFFPOSX1 mem_reg_2__3_ ( .D(n1927), .CLK(clk), .Q(mem[85]) );
  DFFPOSX1 mem_reg_2__2_ ( .D(n1926), .CLK(clk), .Q(mem[84]) );
  DFFPOSX1 mem_reg_2__1_ ( .D(n1925), .CLK(clk), .Q(mem[83]) );
  DFFPOSX1 mem_reg_2__0_ ( .D(n1924), .CLK(clk), .Q(mem[82]) );
  DFFPOSX1 mem_reg_1__40_ ( .D(n1923), .CLK(clk), .Q(mem[81]) );
  DFFPOSX1 mem_reg_1__39_ ( .D(n1922), .CLK(clk), .Q(mem[80]) );
  DFFPOSX1 mem_reg_1__38_ ( .D(n1921), .CLK(clk), .Q(mem[79]) );
  DFFPOSX1 mem_reg_1__37_ ( .D(n1920), .CLK(clk), .Q(mem[78]) );
  DFFPOSX1 mem_reg_1__36_ ( .D(n1919), .CLK(clk), .Q(mem[77]) );
  DFFPOSX1 mem_reg_1__35_ ( .D(n1918), .CLK(clk), .Q(mem[76]) );
  DFFPOSX1 mem_reg_1__34_ ( .D(n1917), .CLK(clk), .Q(mem[75]) );
  DFFPOSX1 mem_reg_1__33_ ( .D(n1916), .CLK(clk), .Q(mem[74]) );
  DFFPOSX1 mem_reg_1__32_ ( .D(n1915), .CLK(clk), .Q(mem[73]) );
  DFFPOSX1 mem_reg_1__31_ ( .D(n1914), .CLK(clk), .Q(mem[72]) );
  DFFPOSX1 mem_reg_1__30_ ( .D(n1913), .CLK(clk), .Q(mem[71]) );
  DFFPOSX1 mem_reg_1__29_ ( .D(n1912), .CLK(clk), .Q(mem[70]) );
  DFFPOSX1 mem_reg_1__28_ ( .D(n1911), .CLK(clk), .Q(mem[69]) );
  DFFPOSX1 mem_reg_1__27_ ( .D(n1910), .CLK(clk), .Q(mem[68]) );
  DFFPOSX1 mem_reg_1__26_ ( .D(n1909), .CLK(clk), .Q(mem[67]) );
  DFFPOSX1 mem_reg_1__25_ ( .D(n1908), .CLK(clk), .Q(mem[66]) );
  DFFPOSX1 mem_reg_1__24_ ( .D(n1907), .CLK(clk), .Q(mem[65]) );
  DFFPOSX1 mem_reg_1__23_ ( .D(n1906), .CLK(clk), .Q(mem[64]) );
  DFFPOSX1 mem_reg_1__22_ ( .D(n1905), .CLK(clk), .Q(mem[63]) );
  DFFPOSX1 mem_reg_1__21_ ( .D(n1904), .CLK(clk), .Q(mem[62]) );
  DFFPOSX1 mem_reg_1__20_ ( .D(n1903), .CLK(clk), .Q(mem[61]) );
  DFFPOSX1 mem_reg_1__19_ ( .D(n1902), .CLK(clk), .Q(mem[60]) );
  DFFPOSX1 mem_reg_1__18_ ( .D(n1901), .CLK(clk), .Q(mem[59]) );
  DFFPOSX1 mem_reg_1__17_ ( .D(n1900), .CLK(clk), .Q(mem[58]) );
  DFFPOSX1 mem_reg_1__16_ ( .D(n1899), .CLK(clk), .Q(mem[57]) );
  DFFPOSX1 mem_reg_1__15_ ( .D(n1898), .CLK(clk), .Q(mem[56]) );
  DFFPOSX1 mem_reg_1__14_ ( .D(n1897), .CLK(clk), .Q(mem[55]) );
  DFFPOSX1 mem_reg_1__13_ ( .D(n1896), .CLK(clk), .Q(mem[54]) );
  DFFPOSX1 mem_reg_1__12_ ( .D(n1895), .CLK(clk), .Q(mem[53]) );
  DFFPOSX1 mem_reg_1__11_ ( .D(n1894), .CLK(clk), .Q(mem[52]) );
  DFFPOSX1 mem_reg_1__10_ ( .D(n1893), .CLK(clk), .Q(mem[51]) );
  DFFPOSX1 mem_reg_1__9_ ( .D(n1892), .CLK(clk), .Q(mem[50]) );
  DFFPOSX1 mem_reg_1__8_ ( .D(n1891), .CLK(clk), .Q(mem[49]) );
  DFFPOSX1 mem_reg_1__7_ ( .D(n1890), .CLK(clk), .Q(mem[48]) );
  DFFPOSX1 mem_reg_1__6_ ( .D(n1889), .CLK(clk), .Q(mem[47]) );
  DFFPOSX1 mem_reg_1__5_ ( .D(n1888), .CLK(clk), .Q(mem[46]) );
  DFFPOSX1 mem_reg_1__4_ ( .D(n1887), .CLK(clk), .Q(mem[45]) );
  DFFPOSX1 mem_reg_1__3_ ( .D(n1886), .CLK(clk), .Q(mem[44]) );
  DFFPOSX1 mem_reg_1__2_ ( .D(n1885), .CLK(clk), .Q(mem[43]) );
  DFFPOSX1 mem_reg_1__1_ ( .D(n1884), .CLK(clk), .Q(mem[42]) );
  DFFPOSX1 mem_reg_1__0_ ( .D(n1883), .CLK(clk), .Q(mem[41]) );
  DFFPOSX1 mem_reg_0__40_ ( .D(n1882), .CLK(clk), .Q(mem[40]) );
  DFFPOSX1 mem_reg_0__39_ ( .D(n1881), .CLK(clk), .Q(mem[39]) );
  DFFPOSX1 mem_reg_0__38_ ( .D(n1880), .CLK(clk), .Q(mem[38]) );
  DFFPOSX1 mem_reg_0__37_ ( .D(n1879), .CLK(clk), .Q(mem[37]) );
  DFFPOSX1 mem_reg_0__36_ ( .D(n1878), .CLK(clk), .Q(mem[36]) );
  DFFPOSX1 mem_reg_0__35_ ( .D(n1877), .CLK(clk), .Q(mem[35]) );
  DFFPOSX1 mem_reg_0__34_ ( .D(n1876), .CLK(clk), .Q(mem[34]) );
  DFFPOSX1 mem_reg_0__33_ ( .D(n1875), .CLK(clk), .Q(mem[33]) );
  DFFPOSX1 mem_reg_0__32_ ( .D(n1874), .CLK(clk), .Q(mem[32]) );
  DFFPOSX1 mem_reg_0__31_ ( .D(n1873), .CLK(clk), .Q(mem[31]) );
  DFFPOSX1 mem_reg_0__30_ ( .D(n1872), .CLK(clk), .Q(mem[30]) );
  DFFPOSX1 mem_reg_0__29_ ( .D(n1871), .CLK(clk), .Q(mem[29]) );
  DFFPOSX1 mem_reg_0__28_ ( .D(n1870), .CLK(clk), .Q(mem[28]) );
  DFFPOSX1 mem_reg_0__27_ ( .D(n1869), .CLK(clk), .Q(mem[27]) );
  DFFPOSX1 mem_reg_0__26_ ( .D(n1868), .CLK(clk), .Q(mem[26]) );
  DFFPOSX1 mem_reg_0__25_ ( .D(n1867), .CLK(clk), .Q(mem[25]) );
  DFFPOSX1 mem_reg_0__24_ ( .D(n1866), .CLK(clk), .Q(mem[24]) );
  DFFPOSX1 mem_reg_0__23_ ( .D(n1865), .CLK(clk), .Q(mem[23]) );
  DFFPOSX1 mem_reg_0__22_ ( .D(n1864), .CLK(clk), .Q(mem[22]) );
  DFFPOSX1 mem_reg_0__21_ ( .D(n1863), .CLK(clk), .Q(mem[21]) );
  DFFPOSX1 mem_reg_0__20_ ( .D(n1862), .CLK(clk), .Q(mem[20]) );
  DFFPOSX1 mem_reg_0__19_ ( .D(n1861), .CLK(clk), .Q(mem[19]) );
  DFFPOSX1 mem_reg_0__18_ ( .D(n1860), .CLK(clk), .Q(mem[18]) );
  DFFPOSX1 mem_reg_0__17_ ( .D(n1859), .CLK(clk), .Q(mem[17]) );
  DFFPOSX1 mem_reg_0__16_ ( .D(n1858), .CLK(clk), .Q(mem[16]) );
  DFFPOSX1 mem_reg_0__15_ ( .D(n1857), .CLK(clk), .Q(mem[15]) );
  DFFPOSX1 mem_reg_0__14_ ( .D(n1856), .CLK(clk), .Q(mem[14]) );
  DFFPOSX1 mem_reg_0__13_ ( .D(n1855), .CLK(clk), .Q(mem[13]) );
  DFFPOSX1 mem_reg_0__12_ ( .D(n1854), .CLK(clk), .Q(mem[12]) );
  DFFPOSX1 mem_reg_0__11_ ( .D(n1853), .CLK(clk), .Q(mem[11]) );
  DFFPOSX1 mem_reg_0__10_ ( .D(n1852), .CLK(clk), .Q(mem[10]) );
  DFFPOSX1 mem_reg_0__9_ ( .D(n1851), .CLK(clk), .Q(mem[9]) );
  DFFPOSX1 mem_reg_0__8_ ( .D(n1850), .CLK(clk), .Q(mem[8]) );
  DFFPOSX1 mem_reg_0__7_ ( .D(n1849), .CLK(clk), .Q(mem[7]) );
  DFFPOSX1 mem_reg_0__6_ ( .D(n1848), .CLK(clk), .Q(mem[6]) );
  DFFPOSX1 mem_reg_0__5_ ( .D(n1847), .CLK(clk), .Q(mem[5]) );
  DFFPOSX1 mem_reg_0__4_ ( .D(n1846), .CLK(clk), .Q(mem[4]) );
  DFFPOSX1 mem_reg_0__3_ ( .D(n1845), .CLK(clk), .Q(mem[3]) );
  DFFPOSX1 mem_reg_0__2_ ( .D(n1844), .CLK(clk), .Q(mem[2]) );
  DFFPOSX1 mem_reg_0__1_ ( .D(n1843), .CLK(clk), .Q(mem[1]) );
  DFFPOSX1 mem_reg_0__0_ ( .D(n1842), .CLK(clk), .Q(mem[0]) );
  OAI21X1 U91 ( .A(n5627), .B(n5668), .C(n4175), .Y(n1842) );
  OAI21X1 U93 ( .A(n5627), .B(n5667), .C(n4083), .Y(n1843) );
  OAI21X1 U95 ( .A(n5627), .B(n5666), .C(n3991), .Y(n1844) );
  OAI21X1 U97 ( .A(n5627), .B(n5665), .C(n3898), .Y(n1845) );
  OAI21X1 U99 ( .A(n5627), .B(n5664), .C(n4174), .Y(n1846) );
  OAI21X1 U101 ( .A(n5627), .B(n5663), .C(n3801), .Y(n1847) );
  OAI21X1 U103 ( .A(n5627), .B(n5662), .C(n3712), .Y(n1848) );
  OAI21X1 U105 ( .A(n5627), .B(n5661), .C(n3622), .Y(n1849) );
  OAI21X1 U107 ( .A(n5627), .B(n5660), .C(n3533), .Y(n1850) );
  OAI21X1 U109 ( .A(n5627), .B(n5659), .C(n3447), .Y(n1851) );
  OAI21X1 U111 ( .A(n5627), .B(n5658), .C(n4082), .Y(n1852) );
  OAI21X1 U113 ( .A(n5627), .B(n5657), .C(n3990), .Y(n1853) );
  OAI21X1 U115 ( .A(n5627), .B(n5656), .C(n3897), .Y(n1854) );
  OAI21X1 U117 ( .A(n5627), .B(n5655), .C(n3532), .Y(n1855) );
  OAI21X1 U119 ( .A(n5627), .B(n5654), .C(n3374), .Y(n1856) );
  OAI21X1 U121 ( .A(n5627), .B(n5653), .C(n3302), .Y(n1857) );
  OAI21X1 U123 ( .A(n5627), .B(n5652), .C(n3230), .Y(n1858) );
  OAI21X1 U125 ( .A(n5627), .B(n5651), .C(n450), .Y(n1859) );
  OAI21X1 U127 ( .A(n5627), .B(n5650), .C(n343), .Y(n1860) );
  OAI21X1 U129 ( .A(n5627), .B(n5649), .C(n3800), .Y(n1861) );
  OAI21X1 U131 ( .A(n5627), .B(n5648), .C(n3711), .Y(n1862) );
  OAI21X1 U133 ( .A(n5627), .B(n5647), .C(n3621), .Y(n1863) );
  OAI21X1 U135 ( .A(n5627), .B(n5646), .C(n271), .Y(n1864) );
  OAI21X1 U137 ( .A(n5627), .B(n5645), .C(n199), .Y(n1865) );
  OAI21X1 U139 ( .A(n5627), .B(n5644), .C(n127), .Y(n1866) );
  OAI21X1 U141 ( .A(n5627), .B(n5643), .C(n4173), .Y(n1867) );
  OAI21X1 U143 ( .A(n5627), .B(n5642), .C(n3531), .Y(n1868) );
  OAI21X1 U145 ( .A(n5627), .B(n5641), .C(n4081), .Y(n1869) );
  OAI21X1 U147 ( .A(n5627), .B(n5640), .C(n3989), .Y(n1870) );
  OAI21X1 U149 ( .A(n5627), .B(n5639), .C(n3896), .Y(n1871) );
  OAI21X1 U151 ( .A(n5627), .B(n5638), .C(n3446), .Y(n1872) );
  OAI21X1 U153 ( .A(n5627), .B(n5637), .C(n3373), .Y(n1873) );
  OAI21X1 U155 ( .A(n5627), .B(n5636), .C(n3301), .Y(n1874) );
  OAI21X1 U157 ( .A(n5627), .B(n5635), .C(n3229), .Y(n1875) );
  OAI21X1 U159 ( .A(n5627), .B(n5634), .C(n3799), .Y(n1876) );
  OAI21X1 U161 ( .A(n5627), .B(n5633), .C(n3710), .Y(n1877) );
  OAI21X1 U163 ( .A(n5627), .B(n5632), .C(n3620), .Y(n1878) );
  OAI21X1 U165 ( .A(n5627), .B(n5631), .C(n448), .Y(n1879) );
  OAI21X1 U167 ( .A(n5627), .B(n5630), .C(n342), .Y(n1880) );
  OAI21X1 U169 ( .A(n5627), .B(n5629), .C(n270), .Y(n1881) );
  OAI21X1 U171 ( .A(n5627), .B(n5628), .C(n3445), .Y(n1882) );
  OAI21X1 U173 ( .A(n3899), .B(n3806), .C(reset), .Y(n462) );
  OAI21X1 U174 ( .A(n5626), .B(n5668), .C(n4080), .Y(n1883) );
  OAI21X1 U176 ( .A(n5626), .B(n5667), .C(n4172), .Y(n1884) );
  OAI21X1 U178 ( .A(n5626), .B(n5666), .C(n3895), .Y(n1885) );
  OAI21X1 U180 ( .A(n5626), .B(n5665), .C(n3988), .Y(n1886) );
  OAI21X1 U182 ( .A(n5626), .B(n5664), .C(n4079), .Y(n1887) );
  OAI21X1 U184 ( .A(n5626), .B(n5663), .C(n3709), .Y(n1888) );
  OAI21X1 U186 ( .A(n5626), .B(n5662), .C(n3798), .Y(n1889) );
  OAI21X1 U188 ( .A(n5626), .B(n5661), .C(n3530), .Y(n1890) );
  OAI21X1 U190 ( .A(n5626), .B(n5660), .C(n3619), .Y(n1891) );
  OAI21X1 U192 ( .A(n5626), .B(n5659), .C(n3372), .Y(n1892) );
  OAI21X1 U194 ( .A(n5626), .B(n5658), .C(n4171), .Y(n1893) );
  OAI21X1 U196 ( .A(n5626), .B(n5657), .C(n3894), .Y(n1894) );
  OAI21X1 U198 ( .A(n5626), .B(n5656), .C(n3987), .Y(n1895) );
  OAI21X1 U200 ( .A(n5626), .B(n5655), .C(n3618), .Y(n1896) );
  OAI21X1 U202 ( .A(n5626), .B(n5654), .C(n3444), .Y(n1897) );
  OAI21X1 U204 ( .A(n5626), .B(n5653), .C(n3228), .Y(n1898) );
  OAI21X1 U206 ( .A(n5626), .B(n5652), .C(n3300), .Y(n1899) );
  OAI21X1 U208 ( .A(n5626), .B(n5651), .C(n341), .Y(n1900) );
  OAI21X1 U210 ( .A(n5626), .B(n5650), .C(n446), .Y(n1901) );
  OAI21X1 U212 ( .A(n5626), .B(n5649), .C(n3708), .Y(n1902) );
  OAI21X1 U214 ( .A(n5626), .B(n5648), .C(n3797), .Y(n1903) );
  OAI21X1 U216 ( .A(n5626), .B(n5647), .C(n3529), .Y(n1904) );
  OAI21X1 U218 ( .A(n5626), .B(n5646), .C(n198), .Y(n1905) );
  OAI21X1 U220 ( .A(n5626), .B(n5645), .C(n269), .Y(n1906) );
  OAI21X1 U222 ( .A(n5626), .B(n5644), .C(n126), .Y(n1907) );
  OAI21X1 U224 ( .A(n5626), .B(n5643), .C(n4078), .Y(n1908) );
  OAI21X1 U226 ( .A(n5626), .B(n5642), .C(n3617), .Y(n1909) );
  OAI21X1 U228 ( .A(n5626), .B(n5641), .C(n4170), .Y(n1910) );
  OAI21X1 U230 ( .A(n5626), .B(n5640), .C(n3893), .Y(n1911) );
  OAI21X1 U232 ( .A(n5626), .B(n5639), .C(n3986), .Y(n1912) );
  OAI21X1 U234 ( .A(n5626), .B(n5638), .C(n3371), .Y(n1913) );
  OAI21X1 U236 ( .A(n5626), .B(n5637), .C(n3443), .Y(n1914) );
  OAI21X1 U238 ( .A(n5626), .B(n5636), .C(n3227), .Y(n1915) );
  OAI21X1 U240 ( .A(n5626), .B(n5635), .C(n3299), .Y(n1916) );
  OAI21X1 U242 ( .A(n5626), .B(n5634), .C(n3707), .Y(n1917) );
  OAI21X1 U244 ( .A(n5626), .B(n5633), .C(n3796), .Y(n1918) );
  OAI21X1 U246 ( .A(n5626), .B(n5632), .C(n3528), .Y(n1919) );
  OAI21X1 U248 ( .A(n5626), .B(n5631), .C(n340), .Y(n1920) );
  OAI21X1 U250 ( .A(n5626), .B(n5630), .C(n444), .Y(n1921) );
  OAI21X1 U252 ( .A(n5626), .B(n5629), .C(n197), .Y(n1922) );
  OAI21X1 U254 ( .A(n5626), .B(n5628), .C(n3370), .Y(n1923) );
  OAI21X1 U256 ( .A(n3899), .B(n3714), .C(reset), .Y(n506) );
  OAI21X1 U257 ( .A(n5625), .B(n5668), .C(n3985), .Y(n1924) );
  OAI21X1 U259 ( .A(n5625), .B(n5667), .C(n3892), .Y(n1925) );
  OAI21X1 U261 ( .A(n5625), .B(n5666), .C(n4169), .Y(n1926) );
  OAI21X1 U263 ( .A(n5625), .B(n5665), .C(n4077), .Y(n1927) );
  OAI21X1 U265 ( .A(n5625), .B(n5664), .C(n3984), .Y(n1928) );
  OAI21X1 U267 ( .A(n5625), .B(n5663), .C(n3616), .Y(n1929) );
  OAI21X1 U269 ( .A(n5625), .B(n5662), .C(n3527), .Y(n1930) );
  OAI21X1 U271 ( .A(n5625), .B(n5661), .C(n3795), .Y(n1931) );
  OAI21X1 U273 ( .A(n5625), .B(n5660), .C(n3706), .Y(n1932) );
  OAI21X1 U275 ( .A(n5625), .B(n5659), .C(n3298), .Y(n1933) );
  OAI21X1 U277 ( .A(n5625), .B(n5658), .C(n3891), .Y(n1934) );
  OAI21X1 U279 ( .A(n5625), .B(n5657), .C(n4168), .Y(n1935) );
  OAI21X1 U281 ( .A(n5625), .B(n5656), .C(n4076), .Y(n1936) );
  OAI21X1 U283 ( .A(n5625), .B(n5655), .C(n3705), .Y(n1937) );
  OAI21X1 U285 ( .A(n5625), .B(n5654), .C(n3226), .Y(n1938) );
  OAI21X1 U287 ( .A(n5625), .B(n5653), .C(n3442), .Y(n1939) );
  OAI21X1 U289 ( .A(n5625), .B(n5652), .C(n3369), .Y(n1940) );
  OAI21X1 U291 ( .A(n5625), .B(n5651), .C(n268), .Y(n1941) );
  OAI21X1 U293 ( .A(n5625), .B(n5650), .C(n196), .Y(n1942) );
  OAI21X1 U295 ( .A(n5625), .B(n5649), .C(n3615), .Y(n1943) );
  OAI21X1 U297 ( .A(n5625), .B(n5648), .C(n3526), .Y(n1944) );
  OAI21X1 U299 ( .A(n5625), .B(n5647), .C(n3794), .Y(n1945) );
  OAI21X1 U301 ( .A(n5625), .B(n5646), .C(n442), .Y(n1946) );
  OAI21X1 U303 ( .A(n5625), .B(n5645), .C(n339), .Y(n1947) );
  OAI21X1 U305 ( .A(n5625), .B(n5644), .C(n125), .Y(n1948) );
  OAI21X1 U307 ( .A(n5625), .B(n5643), .C(n3983), .Y(n1949) );
  OAI21X1 U309 ( .A(n5625), .B(n5642), .C(n3704), .Y(n1950) );
  OAI21X1 U311 ( .A(n5625), .B(n5641), .C(n3890), .Y(n1951) );
  OAI21X1 U313 ( .A(n5625), .B(n5640), .C(n4167), .Y(n1952) );
  OAI21X1 U315 ( .A(n5625), .B(n5639), .C(n4075), .Y(n1953) );
  OAI21X1 U317 ( .A(n5625), .B(n5638), .C(n3297), .Y(n1954) );
  OAI21X1 U319 ( .A(n5625), .B(n5637), .C(n3225), .Y(n1955) );
  OAI21X1 U321 ( .A(n5625), .B(n5636), .C(n3441), .Y(n1956) );
  OAI21X1 U323 ( .A(n5625), .B(n5635), .C(n3368), .Y(n1957) );
  OAI21X1 U325 ( .A(n5625), .B(n5634), .C(n3614), .Y(n1958) );
  OAI21X1 U327 ( .A(n5625), .B(n5633), .C(n3525), .Y(n1959) );
  OAI21X1 U329 ( .A(n5625), .B(n5632), .C(n3793), .Y(n1960) );
  OAI21X1 U331 ( .A(n5625), .B(n5631), .C(n267), .Y(n1961) );
  OAI21X1 U333 ( .A(n5625), .B(n5630), .C(n195), .Y(n1962) );
  OAI21X1 U335 ( .A(n5625), .B(n5629), .C(n440), .Y(n1963) );
  OAI21X1 U337 ( .A(n5625), .B(n5628), .C(n3296), .Y(n1964) );
  OAI21X1 U339 ( .A(n3899), .B(n3624), .C(reset), .Y(n549) );
  OAI21X1 U340 ( .A(n5624), .B(n5668), .C(n3889), .Y(n1965) );
  OAI21X1 U342 ( .A(n5624), .B(n5667), .C(n3982), .Y(n1966) );
  OAI21X1 U344 ( .A(n5624), .B(n5666), .C(n4074), .Y(n1967) );
  OAI21X1 U346 ( .A(n5624), .B(n5665), .C(n4166), .Y(n1968) );
  OAI21X1 U348 ( .A(n5624), .B(n5664), .C(n3888), .Y(n1969) );
  OAI21X1 U350 ( .A(n5624), .B(n5663), .C(n3524), .Y(n1970) );
  OAI21X1 U352 ( .A(n5624), .B(n5662), .C(n3613), .Y(n1971) );
  OAI21X1 U354 ( .A(n5624), .B(n5661), .C(n3703), .Y(n1972) );
  OAI21X1 U356 ( .A(n5624), .B(n5660), .C(n3792), .Y(n1973) );
  OAI21X1 U358 ( .A(n5624), .B(n5659), .C(n3224), .Y(n1974) );
  OAI21X1 U360 ( .A(n5624), .B(n5658), .C(n3981), .Y(n1975) );
  OAI21X1 U362 ( .A(n5624), .B(n5657), .C(n4073), .Y(n1976) );
  OAI21X1 U364 ( .A(n5624), .B(n5656), .C(n4165), .Y(n1977) );
  OAI21X1 U366 ( .A(n5624), .B(n5655), .C(n3791), .Y(n1978) );
  OAI21X1 U368 ( .A(n5624), .B(n5654), .C(n3295), .Y(n1979) );
  OAI21X1 U370 ( .A(n5624), .B(n5653), .C(n3367), .Y(n1980) );
  OAI21X1 U372 ( .A(n5624), .B(n5652), .C(n3440), .Y(n1981) );
  OAI21X1 U374 ( .A(n5624), .B(n5651), .C(n194), .Y(n1982) );
  OAI21X1 U376 ( .A(n5624), .B(n5650), .C(n266), .Y(n1983) );
  OAI21X1 U378 ( .A(n5624), .B(n5649), .C(n3523), .Y(n1984) );
  OAI21X1 U380 ( .A(n5624), .B(n5648), .C(n3612), .Y(n1985) );
  OAI21X1 U382 ( .A(n5624), .B(n5647), .C(n3702), .Y(n1986) );
  OAI21X1 U384 ( .A(n5624), .B(n5646), .C(n338), .Y(n1987) );
  OAI21X1 U386 ( .A(n5624), .B(n5645), .C(n438), .Y(n1988) );
  OAI21X1 U388 ( .A(n5624), .B(n5644), .C(n124), .Y(n1989) );
  OAI21X1 U390 ( .A(n5624), .B(n5643), .C(n3887), .Y(n1990) );
  OAI21X1 U392 ( .A(n5624), .B(n5642), .C(n3790), .Y(n1991) );
  OAI21X1 U394 ( .A(n5624), .B(n5641), .C(n3980), .Y(n1992) );
  OAI21X1 U396 ( .A(n5624), .B(n5640), .C(n4072), .Y(n1993) );
  OAI21X1 U398 ( .A(n5624), .B(n5639), .C(n4164), .Y(n1994) );
  OAI21X1 U400 ( .A(n5624), .B(n5638), .C(n3223), .Y(n1995) );
  OAI21X1 U402 ( .A(n5624), .B(n5637), .C(n3294), .Y(n1996) );
  OAI21X1 U404 ( .A(n5624), .B(n5636), .C(n3366), .Y(n1997) );
  OAI21X1 U406 ( .A(n5624), .B(n5635), .C(n3439), .Y(n1998) );
  OAI21X1 U408 ( .A(n5624), .B(n5634), .C(n3522), .Y(n1999) );
  OAI21X1 U410 ( .A(n5624), .B(n5633), .C(n3611), .Y(n2000) );
  OAI21X1 U412 ( .A(n5624), .B(n5632), .C(n3701), .Y(n2001) );
  OAI21X1 U414 ( .A(n5624), .B(n5631), .C(n193), .Y(n2002) );
  OAI21X1 U416 ( .A(n5624), .B(n5630), .C(n265), .Y(n2003) );
  OAI21X1 U418 ( .A(n5624), .B(n5629), .C(n337), .Y(n2004) );
  OAI21X1 U420 ( .A(n5624), .B(n5628), .C(n3222), .Y(n2005) );
  OAI21X1 U422 ( .A(n3899), .B(n3535), .C(reset), .Y(n592) );
  OAI21X1 U423 ( .A(n5623), .B(n5668), .C(n3789), .Y(n2006) );
  OAI21X1 U425 ( .A(n5623), .B(n5667), .C(n3700), .Y(n2007) );
  OAI21X1 U427 ( .A(n5623), .B(n5666), .C(n3610), .Y(n2008) );
  OAI21X1 U429 ( .A(n5623), .B(n5665), .C(n3521), .Y(n2009) );
  OAI21X1 U431 ( .A(n5623), .B(n5664), .C(n3788), .Y(n2010) );
  OAI21X1 U433 ( .A(n5623), .B(n5663), .C(n4163), .Y(n2011) );
  OAI21X1 U435 ( .A(n5623), .B(n5662), .C(n4071), .Y(n2012) );
  OAI21X1 U437 ( .A(n5623), .B(n5661), .C(n3979), .Y(n2013) );
  OAI21X1 U439 ( .A(n5623), .B(n5660), .C(n3886), .Y(n2014) );
  OAI21X1 U441 ( .A(n5623), .B(n5659), .C(n436), .Y(n2015) );
  OAI21X1 U443 ( .A(n5623), .B(n5658), .C(n3699), .Y(n2016) );
  OAI21X1 U445 ( .A(n5623), .B(n5657), .C(n3609), .Y(n2017) );
  OAI21X1 U447 ( .A(n5623), .B(n5656), .C(n3520), .Y(n2018) );
  OAI21X1 U449 ( .A(n5623), .B(n5655), .C(n3885), .Y(n2019) );
  OAI21X1 U451 ( .A(n5623), .B(n5654), .C(n336), .Y(n2020) );
  OAI21X1 U453 ( .A(n5623), .B(n5653), .C(n264), .Y(n2021) );
  OAI21X1 U455 ( .A(n5623), .B(n5652), .C(n192), .Y(n2022) );
  OAI21X1 U457 ( .A(n5623), .B(n5651), .C(n3438), .Y(n2023) );
  OAI21X1 U459 ( .A(n5623), .B(n5650), .C(n3365), .Y(n2024) );
  OAI21X1 U461 ( .A(n5623), .B(n5649), .C(n4162), .Y(n2025) );
  OAI21X1 U463 ( .A(n5623), .B(n5648), .C(n4070), .Y(n2026) );
  OAI21X1 U465 ( .A(n5623), .B(n5647), .C(n3978), .Y(n2027) );
  OAI21X1 U467 ( .A(n5623), .B(n5646), .C(n3293), .Y(n2028) );
  OAI21X1 U469 ( .A(n5623), .B(n5645), .C(n3221), .Y(n2029) );
  OAI21X1 U471 ( .A(n5623), .B(n5644), .C(n123), .Y(n2030) );
  OAI21X1 U473 ( .A(n5623), .B(n5643), .C(n3787), .Y(n2031) );
  OAI21X1 U475 ( .A(n5623), .B(n5642), .C(n3884), .Y(n2032) );
  OAI21X1 U477 ( .A(n5623), .B(n5641), .C(n3698), .Y(n2033) );
  OAI21X1 U479 ( .A(n5623), .B(n5640), .C(n3608), .Y(n2034) );
  OAI21X1 U481 ( .A(n5623), .B(n5639), .C(n3519), .Y(n2035) );
  OAI21X1 U483 ( .A(n5623), .B(n5638), .C(n434), .Y(n2036) );
  OAI21X1 U485 ( .A(n5623), .B(n5637), .C(n335), .Y(n2037) );
  OAI21X1 U487 ( .A(n5623), .B(n5636), .C(n263), .Y(n2038) );
  OAI21X1 U489 ( .A(n5623), .B(n5635), .C(n191), .Y(n2039) );
  OAI21X1 U491 ( .A(n5623), .B(n5634), .C(n4161), .Y(n2040) );
  OAI21X1 U493 ( .A(n5623), .B(n5633), .C(n4069), .Y(n2041) );
  OAI21X1 U495 ( .A(n5623), .B(n5632), .C(n3977), .Y(n2042) );
  OAI21X1 U497 ( .A(n5623), .B(n5631), .C(n3437), .Y(n2043) );
  OAI21X1 U499 ( .A(n5623), .B(n5630), .C(n3364), .Y(n2044) );
  OAI21X1 U501 ( .A(n5623), .B(n5629), .C(n3292), .Y(n2045) );
  OAI21X1 U503 ( .A(n5623), .B(n5628), .C(n432), .Y(n2046) );
  OAI21X1 U505 ( .A(n3899), .B(n3534), .C(reset), .Y(n635) );
  OAI21X1 U506 ( .A(n5622), .B(n5668), .C(n3697), .Y(n2047) );
  OAI21X1 U508 ( .A(n5622), .B(n5667), .C(n3786), .Y(n2048) );
  OAI21X1 U510 ( .A(n5622), .B(n5666), .C(n3518), .Y(n2049) );
  OAI21X1 U512 ( .A(n5622), .B(n5665), .C(n3607), .Y(n2050) );
  OAI21X1 U514 ( .A(n5622), .B(n5664), .C(n3696), .Y(n2051) );
  OAI21X1 U516 ( .A(n5622), .B(n5663), .C(n4068), .Y(n2052) );
  OAI21X1 U518 ( .A(n5622), .B(n5662), .C(n4160), .Y(n2053) );
  OAI21X1 U520 ( .A(n5622), .B(n5661), .C(n3883), .Y(n2054) );
  OAI21X1 U522 ( .A(n5622), .B(n5660), .C(n3976), .Y(n2055) );
  OAI21X1 U524 ( .A(n5622), .B(n5659), .C(n334), .Y(n2056) );
  OAI21X1 U526 ( .A(n5622), .B(n5658), .C(n3785), .Y(n2057) );
  OAI21X1 U528 ( .A(n5622), .B(n5657), .C(n3517), .Y(n2058) );
  OAI21X1 U530 ( .A(n5622), .B(n5656), .C(n3606), .Y(n2059) );
  OAI21X1 U532 ( .A(n5622), .B(n5655), .C(n3975), .Y(n2060) );
  OAI21X1 U534 ( .A(n5622), .B(n5654), .C(n430), .Y(n2061) );
  OAI21X1 U536 ( .A(n5622), .B(n5653), .C(n190), .Y(n2062) );
  OAI21X1 U538 ( .A(n5622), .B(n5652), .C(n262), .Y(n2063) );
  OAI21X1 U540 ( .A(n5622), .B(n5651), .C(n3363), .Y(n2064) );
  OAI21X1 U542 ( .A(n5622), .B(n5650), .C(n3436), .Y(n2065) );
  OAI21X1 U544 ( .A(n5622), .B(n5649), .C(n4067), .Y(n2066) );
  OAI21X1 U546 ( .A(n5622), .B(n5648), .C(n4159), .Y(n2067) );
  OAI21X1 U548 ( .A(n5622), .B(n5647), .C(n3882), .Y(n2068) );
  OAI21X1 U550 ( .A(n5622), .B(n5646), .C(n3220), .Y(n2069) );
  OAI21X1 U552 ( .A(n5622), .B(n5645), .C(n3291), .Y(n2070) );
  OAI21X1 U554 ( .A(n5622), .B(n5644), .C(n122), .Y(n2071) );
  OAI21X1 U556 ( .A(n5622), .B(n5643), .C(n3695), .Y(n2072) );
  OAI21X1 U558 ( .A(n5622), .B(n5642), .C(n3974), .Y(n2073) );
  OAI21X1 U560 ( .A(n5622), .B(n5641), .C(n3784), .Y(n2074) );
  OAI21X1 U562 ( .A(n5622), .B(n5640), .C(n3516), .Y(n2075) );
  OAI21X1 U564 ( .A(n5622), .B(n5639), .C(n3605), .Y(n2076) );
  OAI21X1 U566 ( .A(n5622), .B(n5638), .C(n333), .Y(n2077) );
  OAI21X1 U568 ( .A(n5622), .B(n5637), .C(n428), .Y(n2078) );
  OAI21X1 U570 ( .A(n5622), .B(n5636), .C(n189), .Y(n2079) );
  OAI21X1 U572 ( .A(n5622), .B(n5635), .C(n261), .Y(n2080) );
  OAI21X1 U574 ( .A(n5622), .B(n5634), .C(n4066), .Y(n2081) );
  OAI21X1 U576 ( .A(n5622), .B(n5633), .C(n4158), .Y(n2082) );
  OAI21X1 U578 ( .A(n5622), .B(n5632), .C(n3881), .Y(n2083) );
  OAI21X1 U580 ( .A(n5622), .B(n5631), .C(n3362), .Y(n2084) );
  OAI21X1 U582 ( .A(n5622), .B(n5630), .C(n3435), .Y(n2085) );
  OAI21X1 U584 ( .A(n5622), .B(n5629), .C(n3219), .Y(n2086) );
  OAI21X1 U586 ( .A(n5622), .B(n5628), .C(n332), .Y(n2087) );
  OAI21X1 U588 ( .A(n3899), .B(n3623), .C(reset), .Y(n678) );
  OAI21X1 U589 ( .A(n5621), .B(n5668), .C(n3604), .Y(n2088) );
  OAI21X1 U591 ( .A(n5621), .B(n5667), .C(n3515), .Y(n2089) );
  OAI21X1 U593 ( .A(n5621), .B(n5666), .C(n3783), .Y(n2090) );
  OAI21X1 U595 ( .A(n5621), .B(n5665), .C(n3694), .Y(n2091) );
  OAI21X1 U597 ( .A(n5621), .B(n5664), .C(n3603), .Y(n2092) );
  OAI21X1 U599 ( .A(n5621), .B(n5663), .C(n3973), .Y(n2093) );
  OAI21X1 U601 ( .A(n5621), .B(n5662), .C(n3880), .Y(n2094) );
  OAI21X1 U603 ( .A(n5621), .B(n5661), .C(n4157), .Y(n2095) );
  OAI21X1 U605 ( .A(n5621), .B(n5660), .C(n4065), .Y(n2096) );
  OAI21X1 U607 ( .A(n5621), .B(n5659), .C(n260), .Y(n2097) );
  OAI21X1 U609 ( .A(n5621), .B(n5658), .C(n3514), .Y(n2098) );
  OAI21X1 U611 ( .A(n5621), .B(n5657), .C(n3782), .Y(n2099) );
  OAI21X1 U613 ( .A(n5621), .B(n5656), .C(n3693), .Y(n2100) );
  OAI21X1 U615 ( .A(n5621), .B(n5655), .C(n4064), .Y(n2101) );
  OAI21X1 U617 ( .A(n5621), .B(n5654), .C(n188), .Y(n2102) );
  OAI21X1 U619 ( .A(n5621), .B(n5653), .C(n426), .Y(n2103) );
  OAI21X1 U621 ( .A(n5621), .B(n5652), .C(n331), .Y(n2104) );
  OAI21X1 U623 ( .A(n5621), .B(n5651), .C(n3290), .Y(n2105) );
  OAI21X1 U625 ( .A(n5621), .B(n5650), .C(n3218), .Y(n2106) );
  OAI21X1 U627 ( .A(n5621), .B(n5649), .C(n3972), .Y(n2107) );
  OAI21X1 U629 ( .A(n5621), .B(n5648), .C(n3879), .Y(n2108) );
  OAI21X1 U631 ( .A(n5621), .B(n5647), .C(n4156), .Y(n2109) );
  OAI21X1 U633 ( .A(n5621), .B(n5646), .C(n3434), .Y(n2110) );
  OAI21X1 U635 ( .A(n5621), .B(n5645), .C(n3361), .Y(n2111) );
  OAI21X1 U637 ( .A(n5621), .B(n5644), .C(n121), .Y(n2112) );
  OAI21X1 U639 ( .A(n5621), .B(n5643), .C(n3602), .Y(n2113) );
  OAI21X1 U641 ( .A(n5621), .B(n5642), .C(n4063), .Y(n2114) );
  OAI21X1 U643 ( .A(n5621), .B(n5641), .C(n3513), .Y(n2115) );
  OAI21X1 U645 ( .A(n5621), .B(n5640), .C(n3781), .Y(n2116) );
  OAI21X1 U647 ( .A(n5621), .B(n5639), .C(n3692), .Y(n2117) );
  OAI21X1 U649 ( .A(n5621), .B(n5638), .C(n259), .Y(n2118) );
  OAI21X1 U651 ( .A(n5621), .B(n5637), .C(n187), .Y(n2119) );
  OAI21X1 U653 ( .A(n5621), .B(n5636), .C(n424), .Y(n2120) );
  OAI21X1 U655 ( .A(n5621), .B(n5635), .C(n330), .Y(n2121) );
  OAI21X1 U657 ( .A(n5621), .B(n5634), .C(n3971), .Y(n2122) );
  OAI21X1 U659 ( .A(n5621), .B(n5633), .C(n3878), .Y(n2123) );
  OAI21X1 U661 ( .A(n5621), .B(n5632), .C(n4155), .Y(n2124) );
  OAI21X1 U663 ( .A(n5621), .B(n5631), .C(n3289), .Y(n2125) );
  OAI21X1 U665 ( .A(n5621), .B(n5630), .C(n3217), .Y(n2126) );
  OAI21X1 U667 ( .A(n5621), .B(n5629), .C(n3433), .Y(n2127) );
  OAI21X1 U669 ( .A(n5621), .B(n5628), .C(n258), .Y(n2128) );
  OAI21X1 U671 ( .A(n3899), .B(n3713), .C(reset), .Y(n721) );
  OAI21X1 U672 ( .A(n5620), .B(n5668), .C(n3512), .Y(n2129) );
  OAI21X1 U674 ( .A(n5620), .B(n5667), .C(n3601), .Y(n2130) );
  OAI21X1 U676 ( .A(n5620), .B(n5666), .C(n3691), .Y(n2131) );
  OAI21X1 U678 ( .A(n5620), .B(n5665), .C(n3780), .Y(n2132) );
  OAI21X1 U680 ( .A(n5620), .B(n5664), .C(n3511), .Y(n2133) );
  OAI21X1 U682 ( .A(n5620), .B(n5663), .C(n3877), .Y(n2134) );
  OAI21X1 U684 ( .A(n5620), .B(n5662), .C(n3970), .Y(n2135) );
  OAI21X1 U686 ( .A(n5620), .B(n5661), .C(n4062), .Y(n2136) );
  OAI21X1 U688 ( .A(n5620), .B(n5660), .C(n4154), .Y(n2137) );
  OAI21X1 U690 ( .A(n5620), .B(n5659), .C(n186), .Y(n2138) );
  OAI21X1 U692 ( .A(n5620), .B(n5658), .C(n3600), .Y(n2139) );
  OAI21X1 U694 ( .A(n5620), .B(n5657), .C(n3690), .Y(n2140) );
  OAI21X1 U696 ( .A(n5620), .B(n5656), .C(n3779), .Y(n2141) );
  OAI21X1 U698 ( .A(n5620), .B(n5655), .C(n4153), .Y(n2142) );
  OAI21X1 U700 ( .A(n5620), .B(n5654), .C(n257), .Y(n2143) );
  OAI21X1 U702 ( .A(n5620), .B(n5653), .C(n329), .Y(n2144) );
  OAI21X1 U704 ( .A(n5620), .B(n5652), .C(n422), .Y(n2145) );
  OAI21X1 U706 ( .A(n5620), .B(n5651), .C(n3216), .Y(n2146) );
  OAI21X1 U708 ( .A(n5620), .B(n5650), .C(n3288), .Y(n2147) );
  OAI21X1 U710 ( .A(n5620), .B(n5649), .C(n3876), .Y(n2148) );
  OAI21X1 U712 ( .A(n5620), .B(n5648), .C(n3969), .Y(n2149) );
  OAI21X1 U714 ( .A(n5620), .B(n5647), .C(n4061), .Y(n2150) );
  OAI21X1 U716 ( .A(n5620), .B(n5646), .C(n3360), .Y(n2151) );
  OAI21X1 U718 ( .A(n5620), .B(n5645), .C(n3432), .Y(n2152) );
  OAI21X1 U720 ( .A(n5620), .B(n5644), .C(n120), .Y(n2153) );
  OAI21X1 U722 ( .A(n5620), .B(n5643), .C(n3510), .Y(n2154) );
  OAI21X1 U724 ( .A(n5620), .B(n5642), .C(n4152), .Y(n2155) );
  OAI21X1 U726 ( .A(n5620), .B(n5641), .C(n3599), .Y(n2156) );
  OAI21X1 U728 ( .A(n5620), .B(n5640), .C(n3689), .Y(n2157) );
  OAI21X1 U730 ( .A(n5620), .B(n5639), .C(n3778), .Y(n2158) );
  OAI21X1 U732 ( .A(n5620), .B(n5638), .C(n185), .Y(n2159) );
  OAI21X1 U734 ( .A(n5620), .B(n5637), .C(n256), .Y(n2160) );
  OAI21X1 U736 ( .A(n5620), .B(n5636), .C(n328), .Y(n2161) );
  OAI21X1 U738 ( .A(n5620), .B(n5635), .C(n420), .Y(n2162) );
  OAI21X1 U740 ( .A(n5620), .B(n5634), .C(n3875), .Y(n2163) );
  OAI21X1 U742 ( .A(n5620), .B(n5633), .C(n3968), .Y(n2164) );
  OAI21X1 U744 ( .A(n5620), .B(n5632), .C(n4060), .Y(n2165) );
  OAI21X1 U746 ( .A(n5620), .B(n5631), .C(n3215), .Y(n2166) );
  OAI21X1 U748 ( .A(n5620), .B(n5630), .C(n3287), .Y(n2167) );
  OAI21X1 U750 ( .A(n5620), .B(n5629), .C(n3359), .Y(n2168) );
  OAI21X1 U752 ( .A(n5620), .B(n5628), .C(n184), .Y(n2169) );
  OAI21X1 U754 ( .A(n3899), .B(n3805), .C(reset), .Y(n764) );
  NAND3X1 U755 ( .A(n5720), .B(n5717), .C(n1777), .Y(n463) );
  OAI21X1 U756 ( .A(n5619), .B(n5668), .C(n4151), .Y(n2170) );
  OAI21X1 U758 ( .A(n5619), .B(n5667), .C(n4059), .Y(n2171) );
  OAI21X1 U760 ( .A(n5619), .B(n5666), .C(n3967), .Y(n2172) );
  OAI21X1 U762 ( .A(n5619), .B(n5665), .C(n3874), .Y(n2173) );
  OAI21X1 U764 ( .A(n5619), .B(n5664), .C(n4150), .Y(n2174) );
  OAI21X1 U766 ( .A(n5619), .B(n5663), .C(n3777), .Y(n2175) );
  OAI21X1 U768 ( .A(n5619), .B(n5662), .C(n3688), .Y(n2176) );
  OAI21X1 U770 ( .A(n5619), .B(n5661), .C(n3598), .Y(n2177) );
  OAI21X1 U772 ( .A(n5619), .B(n5660), .C(n3509), .Y(n2178) );
  OAI21X1 U774 ( .A(n5619), .B(n5659), .C(n3431), .Y(n2179) );
  OAI21X1 U776 ( .A(n5619), .B(n5658), .C(n4058), .Y(n2180) );
  OAI21X1 U778 ( .A(n5619), .B(n5657), .C(n3966), .Y(n2181) );
  OAI21X1 U780 ( .A(n5619), .B(n5656), .C(n3873), .Y(n2182) );
  OAI21X1 U782 ( .A(n5619), .B(n5655), .C(n3508), .Y(n2183) );
  OAI21X1 U784 ( .A(n5619), .B(n5654), .C(n3358), .Y(n2184) );
  OAI21X1 U786 ( .A(n5619), .B(n5653), .C(n3286), .Y(n2185) );
  OAI21X1 U788 ( .A(n5619), .B(n5652), .C(n3214), .Y(n2186) );
  OAI21X1 U790 ( .A(n5619), .B(n5651), .C(n418), .Y(n2187) );
  OAI21X1 U792 ( .A(n5619), .B(n5650), .C(n327), .Y(n2188) );
  OAI21X1 U794 ( .A(n5619), .B(n5649), .C(n3776), .Y(n2189) );
  OAI21X1 U796 ( .A(n5619), .B(n5648), .C(n3687), .Y(n2190) );
  OAI21X1 U798 ( .A(n5619), .B(n5647), .C(n3597), .Y(n2191) );
  OAI21X1 U800 ( .A(n5619), .B(n5646), .C(n255), .Y(n2192) );
  OAI21X1 U802 ( .A(n5619), .B(n5645), .C(n183), .Y(n2193) );
  OAI21X1 U804 ( .A(n5619), .B(n5644), .C(n119), .Y(n2194) );
  OAI21X1 U806 ( .A(n5619), .B(n5643), .C(n4149), .Y(n2195) );
  OAI21X1 U808 ( .A(n5619), .B(n5642), .C(n3507), .Y(n2196) );
  OAI21X1 U810 ( .A(n5619), .B(n5641), .C(n4057), .Y(n2197) );
  OAI21X1 U812 ( .A(n5619), .B(n5640), .C(n3965), .Y(n2198) );
  OAI21X1 U814 ( .A(n5619), .B(n5639), .C(n3872), .Y(n2199) );
  OAI21X1 U816 ( .A(n5619), .B(n5638), .C(n3430), .Y(n2200) );
  OAI21X1 U818 ( .A(n5619), .B(n5637), .C(n3357), .Y(n2201) );
  OAI21X1 U820 ( .A(n5619), .B(n5636), .C(n3285), .Y(n2202) );
  OAI21X1 U822 ( .A(n5619), .B(n5635), .C(n3213), .Y(n2203) );
  OAI21X1 U824 ( .A(n5619), .B(n5634), .C(n3775), .Y(n2204) );
  OAI21X1 U826 ( .A(n5619), .B(n5633), .C(n3686), .Y(n2205) );
  OAI21X1 U828 ( .A(n5619), .B(n5632), .C(n3596), .Y(n2206) );
  OAI21X1 U830 ( .A(n5619), .B(n5631), .C(n416), .Y(n2207) );
  OAI21X1 U832 ( .A(n5619), .B(n5630), .C(n326), .Y(n2208) );
  OAI21X1 U834 ( .A(n5619), .B(n5629), .C(n254), .Y(n2209) );
  OAI21X1 U836 ( .A(n5619), .B(n5628), .C(n3429), .Y(n2210) );
  OAI21X1 U838 ( .A(n3806), .B(n4179), .C(reset), .Y(n807) );
  OAI21X1 U839 ( .A(n5618), .B(n5668), .C(n4056), .Y(n2211) );
  OAI21X1 U841 ( .A(n5618), .B(n5667), .C(n4148), .Y(n2212) );
  OAI21X1 U843 ( .A(n5618), .B(n5666), .C(n3871), .Y(n2213) );
  OAI21X1 U845 ( .A(n5618), .B(n5665), .C(n3964), .Y(n2214) );
  OAI21X1 U847 ( .A(n5618), .B(n5664), .C(n4055), .Y(n2215) );
  OAI21X1 U849 ( .A(n5618), .B(n5663), .C(n3685), .Y(n2216) );
  OAI21X1 U851 ( .A(n5618), .B(n5662), .C(n3774), .Y(n2217) );
  OAI21X1 U853 ( .A(n5618), .B(n5661), .C(n3506), .Y(n2218) );
  OAI21X1 U855 ( .A(n5618), .B(n5660), .C(n3595), .Y(n2219) );
  OAI21X1 U857 ( .A(n5618), .B(n5659), .C(n3356), .Y(n2220) );
  OAI21X1 U859 ( .A(n5618), .B(n5658), .C(n4147), .Y(n2221) );
  OAI21X1 U861 ( .A(n5618), .B(n5657), .C(n3870), .Y(n2222) );
  OAI21X1 U863 ( .A(n5618), .B(n5656), .C(n3963), .Y(n2223) );
  OAI21X1 U865 ( .A(n5618), .B(n5655), .C(n3594), .Y(n2224) );
  OAI21X1 U867 ( .A(n5618), .B(n5654), .C(n3428), .Y(n2225) );
  OAI21X1 U869 ( .A(n5618), .B(n5653), .C(n3212), .Y(n2226) );
  OAI21X1 U871 ( .A(n5618), .B(n5652), .C(n3284), .Y(n2227) );
  OAI21X1 U873 ( .A(n5618), .B(n5651), .C(n325), .Y(n2228) );
  OAI21X1 U875 ( .A(n5618), .B(n5650), .C(n414), .Y(n2229) );
  OAI21X1 U877 ( .A(n5618), .B(n5649), .C(n3684), .Y(n2230) );
  OAI21X1 U879 ( .A(n5618), .B(n5648), .C(n3773), .Y(n2231) );
  OAI21X1 U881 ( .A(n5618), .B(n5647), .C(n3505), .Y(n2232) );
  OAI21X1 U883 ( .A(n5618), .B(n5646), .C(n182), .Y(n2233) );
  OAI21X1 U885 ( .A(n5618), .B(n5645), .C(n253), .Y(n2234) );
  OAI21X1 U887 ( .A(n5618), .B(n5644), .C(n118), .Y(n2235) );
  OAI21X1 U889 ( .A(n5618), .B(n5643), .C(n4054), .Y(n2236) );
  OAI21X1 U891 ( .A(n5618), .B(n5642), .C(n3593), .Y(n2237) );
  OAI21X1 U893 ( .A(n5618), .B(n5641), .C(n4146), .Y(n2238) );
  OAI21X1 U895 ( .A(n5618), .B(n5640), .C(n3869), .Y(n2239) );
  OAI21X1 U897 ( .A(n5618), .B(n5639), .C(n3962), .Y(n2240) );
  OAI21X1 U899 ( .A(n5618), .B(n5638), .C(n3355), .Y(n2241) );
  OAI21X1 U901 ( .A(n5618), .B(n5637), .C(n3427), .Y(n2242) );
  OAI21X1 U903 ( .A(n5618), .B(n5636), .C(n3211), .Y(n2243) );
  OAI21X1 U905 ( .A(n5618), .B(n5635), .C(n3283), .Y(n2244) );
  OAI21X1 U907 ( .A(n5618), .B(n5634), .C(n3683), .Y(n2245) );
  OAI21X1 U909 ( .A(n5618), .B(n5633), .C(n3772), .Y(n2246) );
  OAI21X1 U911 ( .A(n5618), .B(n5632), .C(n3504), .Y(n2247) );
  OAI21X1 U913 ( .A(n5618), .B(n5631), .C(n324), .Y(n2248) );
  OAI21X1 U915 ( .A(n5618), .B(n5630), .C(n412), .Y(n2249) );
  OAI21X1 U917 ( .A(n5618), .B(n5629), .C(n181), .Y(n2250) );
  OAI21X1 U919 ( .A(n5618), .B(n5628), .C(n3354), .Y(n2251) );
  OAI21X1 U921 ( .A(n3714), .B(n4179), .C(reset), .Y(n850) );
  OAI21X1 U922 ( .A(n5617), .B(n5668), .C(n3961), .Y(n2252) );
  OAI21X1 U924 ( .A(n5617), .B(n5667), .C(n3868), .Y(n2253) );
  OAI21X1 U926 ( .A(n5617), .B(n5666), .C(n4145), .Y(n2254) );
  OAI21X1 U928 ( .A(n5617), .B(n5665), .C(n4053), .Y(n2255) );
  OAI21X1 U930 ( .A(n5617), .B(n5664), .C(n3960), .Y(n2256) );
  OAI21X1 U932 ( .A(n5617), .B(n5663), .C(n3592), .Y(n2257) );
  OAI21X1 U934 ( .A(n5617), .B(n5662), .C(n3503), .Y(n2258) );
  OAI21X1 U936 ( .A(n5617), .B(n5661), .C(n3771), .Y(n2259) );
  OAI21X1 U938 ( .A(n5617), .B(n5660), .C(n3682), .Y(n2260) );
  OAI21X1 U940 ( .A(n5617), .B(n5659), .C(n3282), .Y(n2261) );
  OAI21X1 U942 ( .A(n5617), .B(n5658), .C(n3867), .Y(n2262) );
  OAI21X1 U944 ( .A(n5617), .B(n5657), .C(n4144), .Y(n2263) );
  OAI21X1 U946 ( .A(n5617), .B(n5656), .C(n4052), .Y(n2264) );
  OAI21X1 U948 ( .A(n5617), .B(n5655), .C(n3681), .Y(n2265) );
  OAI21X1 U950 ( .A(n5617), .B(n5654), .C(n3210), .Y(n2266) );
  OAI21X1 U952 ( .A(n5617), .B(n5653), .C(n3426), .Y(n2267) );
  OAI21X1 U954 ( .A(n5617), .B(n5652), .C(n3353), .Y(n2268) );
  OAI21X1 U956 ( .A(n5617), .B(n5651), .C(n252), .Y(n2269) );
  OAI21X1 U958 ( .A(n5617), .B(n5650), .C(n180), .Y(n2270) );
  OAI21X1 U960 ( .A(n5617), .B(n5649), .C(n3591), .Y(n2271) );
  OAI21X1 U962 ( .A(n5617), .B(n5648), .C(n3502), .Y(n2272) );
  OAI21X1 U964 ( .A(n5617), .B(n5647), .C(n3770), .Y(n2273) );
  OAI21X1 U966 ( .A(n5617), .B(n5646), .C(n410), .Y(n2274) );
  OAI21X1 U968 ( .A(n5617), .B(n5645), .C(n323), .Y(n2275) );
  OAI21X1 U970 ( .A(n5617), .B(n5644), .C(n117), .Y(n2276) );
  OAI21X1 U972 ( .A(n5617), .B(n5643), .C(n3959), .Y(n2277) );
  OAI21X1 U974 ( .A(n5617), .B(n5642), .C(n3680), .Y(n2278) );
  OAI21X1 U976 ( .A(n5617), .B(n5641), .C(n3866), .Y(n2279) );
  OAI21X1 U978 ( .A(n5617), .B(n5640), .C(n4143), .Y(n2280) );
  OAI21X1 U980 ( .A(n5617), .B(n5639), .C(n4051), .Y(n2281) );
  OAI21X1 U982 ( .A(n5617), .B(n5638), .C(n3281), .Y(n2282) );
  OAI21X1 U984 ( .A(n5617), .B(n5637), .C(n3209), .Y(n2283) );
  OAI21X1 U986 ( .A(n5617), .B(n5636), .C(n3425), .Y(n2284) );
  OAI21X1 U988 ( .A(n5617), .B(n5635), .C(n3352), .Y(n2285) );
  OAI21X1 U990 ( .A(n5617), .B(n5634), .C(n3590), .Y(n2286) );
  OAI21X1 U992 ( .A(n5617), .B(n5633), .C(n3501), .Y(n2287) );
  OAI21X1 U994 ( .A(n5617), .B(n5632), .C(n3769), .Y(n2288) );
  OAI21X1 U996 ( .A(n5617), .B(n5631), .C(n251), .Y(n2289) );
  OAI21X1 U998 ( .A(n5617), .B(n5630), .C(n179), .Y(n2290) );
  OAI21X1 U1000 ( .A(n5617), .B(n5629), .C(n408), .Y(n2291) );
  OAI21X1 U1002 ( .A(n5617), .B(n5628), .C(n3280), .Y(n2292) );
  OAI21X1 U1004 ( .A(n3624), .B(n4179), .C(reset), .Y(n892) );
  OAI21X1 U1005 ( .A(n5616), .B(n5668), .C(n3865), .Y(n2293) );
  OAI21X1 U1007 ( .A(n5616), .B(n5667), .C(n3958), .Y(n2294) );
  OAI21X1 U1009 ( .A(n5616), .B(n5666), .C(n4050), .Y(n2295) );
  OAI21X1 U1011 ( .A(n5616), .B(n5665), .C(n4142), .Y(n2296) );
  OAI21X1 U1013 ( .A(n5616), .B(n5664), .C(n3864), .Y(n2297) );
  OAI21X1 U1015 ( .A(n5616), .B(n5663), .C(n3500), .Y(n2298) );
  OAI21X1 U1017 ( .A(n5616), .B(n5662), .C(n3589), .Y(n2299) );
  OAI21X1 U1019 ( .A(n5616), .B(n5661), .C(n3679), .Y(n2300) );
  OAI21X1 U1021 ( .A(n5616), .B(n5660), .C(n3768), .Y(n2301) );
  OAI21X1 U1023 ( .A(n5616), .B(n5659), .C(n3208), .Y(n2302) );
  OAI21X1 U1025 ( .A(n5616), .B(n5658), .C(n3957), .Y(n2303) );
  OAI21X1 U1027 ( .A(n5616), .B(n5657), .C(n4049), .Y(n2304) );
  OAI21X1 U1029 ( .A(n5616), .B(n5656), .C(n4141), .Y(n2305) );
  OAI21X1 U1031 ( .A(n5616), .B(n5655), .C(n3767), .Y(n2306) );
  OAI21X1 U1033 ( .A(n5616), .B(n5654), .C(n3279), .Y(n2307) );
  OAI21X1 U1035 ( .A(n5616), .B(n5653), .C(n3351), .Y(n2308) );
  OAI21X1 U1037 ( .A(n5616), .B(n5652), .C(n3424), .Y(n2309) );
  OAI21X1 U1039 ( .A(n5616), .B(n5651), .C(n178), .Y(n2310) );
  OAI21X1 U1041 ( .A(n5616), .B(n5650), .C(n250), .Y(n2311) );
  OAI21X1 U1043 ( .A(n5616), .B(n5649), .C(n3499), .Y(n2312) );
  OAI21X1 U1045 ( .A(n5616), .B(n5648), .C(n3588), .Y(n2313) );
  OAI21X1 U1047 ( .A(n5616), .B(n5647), .C(n3678), .Y(n2314) );
  OAI21X1 U1049 ( .A(n5616), .B(n5646), .C(n322), .Y(n2315) );
  OAI21X1 U1051 ( .A(n5616), .B(n5645), .C(n406), .Y(n2316) );
  OAI21X1 U1053 ( .A(n5616), .B(n5644), .C(n116), .Y(n2317) );
  OAI21X1 U1055 ( .A(n5616), .B(n5643), .C(n3863), .Y(n2318) );
  OAI21X1 U1057 ( .A(n5616), .B(n5642), .C(n3766), .Y(n2319) );
  OAI21X1 U1059 ( .A(n5616), .B(n5641), .C(n3956), .Y(n2320) );
  OAI21X1 U1061 ( .A(n5616), .B(n5640), .C(n4048), .Y(n2321) );
  OAI21X1 U1063 ( .A(n5616), .B(n5639), .C(n4140), .Y(n2322) );
  OAI21X1 U1065 ( .A(n5616), .B(n5638), .C(n3207), .Y(n2323) );
  OAI21X1 U1067 ( .A(n5616), .B(n5637), .C(n3278), .Y(n2324) );
  OAI21X1 U1069 ( .A(n5616), .B(n5636), .C(n3350), .Y(n2325) );
  OAI21X1 U1071 ( .A(n5616), .B(n5635), .C(n3423), .Y(n2326) );
  OAI21X1 U1073 ( .A(n5616), .B(n5634), .C(n3498), .Y(n2327) );
  OAI21X1 U1075 ( .A(n5616), .B(n5633), .C(n3587), .Y(n2328) );
  OAI21X1 U1077 ( .A(n5616), .B(n5632), .C(n3677), .Y(n2329) );
  OAI21X1 U1079 ( .A(n5616), .B(n5631), .C(n177), .Y(n2330) );
  OAI21X1 U1081 ( .A(n5616), .B(n5630), .C(n249), .Y(n2331) );
  OAI21X1 U1083 ( .A(n5616), .B(n5629), .C(n321), .Y(n2332) );
  OAI21X1 U1085 ( .A(n5616), .B(n5628), .C(n3206), .Y(n2333) );
  OAI21X1 U1087 ( .A(n3535), .B(n4179), .C(reset), .Y(n934) );
  OAI21X1 U1088 ( .A(n5615), .B(n5668), .C(n3765), .Y(n2334) );
  OAI21X1 U1090 ( .A(n5615), .B(n5667), .C(n3676), .Y(n2335) );
  OAI21X1 U1092 ( .A(n5615), .B(n5666), .C(n3586), .Y(n2336) );
  OAI21X1 U1094 ( .A(n5615), .B(n5665), .C(n3497), .Y(n2337) );
  OAI21X1 U1096 ( .A(n5615), .B(n5664), .C(n3764), .Y(n2338) );
  OAI21X1 U1098 ( .A(n5615), .B(n5663), .C(n4139), .Y(n2339) );
  OAI21X1 U1100 ( .A(n5615), .B(n5662), .C(n4047), .Y(n2340) );
  OAI21X1 U1102 ( .A(n5615), .B(n5661), .C(n3955), .Y(n2341) );
  OAI21X1 U1104 ( .A(n5615), .B(n5660), .C(n3862), .Y(n2342) );
  OAI21X1 U1106 ( .A(n5615), .B(n5659), .C(n404), .Y(n2343) );
  OAI21X1 U1108 ( .A(n5615), .B(n5658), .C(n3675), .Y(n2344) );
  OAI21X1 U1110 ( .A(n5615), .B(n5657), .C(n3585), .Y(n2345) );
  OAI21X1 U1112 ( .A(n5615), .B(n5656), .C(n3496), .Y(n2346) );
  OAI21X1 U1114 ( .A(n5615), .B(n5655), .C(n3861), .Y(n2347) );
  OAI21X1 U1116 ( .A(n5615), .B(n5654), .C(n320), .Y(n2348) );
  OAI21X1 U1118 ( .A(n5615), .B(n5653), .C(n248), .Y(n2349) );
  OAI21X1 U1120 ( .A(n5615), .B(n5652), .C(n176), .Y(n2350) );
  OAI21X1 U1122 ( .A(n5615), .B(n5651), .C(n3422), .Y(n2351) );
  OAI21X1 U1124 ( .A(n5615), .B(n5650), .C(n3349), .Y(n2352) );
  OAI21X1 U1126 ( .A(n5615), .B(n5649), .C(n4138), .Y(n2353) );
  OAI21X1 U1128 ( .A(n5615), .B(n5648), .C(n4046), .Y(n2354) );
  OAI21X1 U1130 ( .A(n5615), .B(n5647), .C(n3954), .Y(n2355) );
  OAI21X1 U1132 ( .A(n5615), .B(n5646), .C(n3277), .Y(n2356) );
  OAI21X1 U1134 ( .A(n5615), .B(n5645), .C(n3205), .Y(n2357) );
  OAI21X1 U1136 ( .A(n5615), .B(n5644), .C(n115), .Y(n2358) );
  OAI21X1 U1138 ( .A(n5615), .B(n5643), .C(n3763), .Y(n2359) );
  OAI21X1 U1140 ( .A(n5615), .B(n5642), .C(n3860), .Y(n2360) );
  OAI21X1 U1142 ( .A(n5615), .B(n5641), .C(n3674), .Y(n2361) );
  OAI21X1 U1144 ( .A(n5615), .B(n5640), .C(n3584), .Y(n2362) );
  OAI21X1 U1146 ( .A(n5615), .B(n5639), .C(n3495), .Y(n2363) );
  OAI21X1 U1148 ( .A(n5615), .B(n5638), .C(n402), .Y(n2364) );
  OAI21X1 U1150 ( .A(n5615), .B(n5637), .C(n319), .Y(n2365) );
  OAI21X1 U1152 ( .A(n5615), .B(n5636), .C(n247), .Y(n2366) );
  OAI21X1 U1154 ( .A(n5615), .B(n5635), .C(n175), .Y(n2367) );
  OAI21X1 U1156 ( .A(n5615), .B(n5634), .C(n4137), .Y(n2368) );
  OAI21X1 U1158 ( .A(n5615), .B(n5633), .C(n4045), .Y(n2369) );
  OAI21X1 U1160 ( .A(n5615), .B(n5632), .C(n3953), .Y(n2370) );
  OAI21X1 U1162 ( .A(n5615), .B(n5631), .C(n3421), .Y(n2371) );
  OAI21X1 U1164 ( .A(n5615), .B(n5630), .C(n3348), .Y(n2372) );
  OAI21X1 U1166 ( .A(n5615), .B(n5629), .C(n3276), .Y(n2373) );
  OAI21X1 U1168 ( .A(n5615), .B(n5628), .C(n400), .Y(n2374) );
  OAI21X1 U1170 ( .A(n3534), .B(n4179), .C(reset), .Y(n976) );
  OAI21X1 U1171 ( .A(n5614), .B(n5668), .C(n3673), .Y(n2375) );
  OAI21X1 U1173 ( .A(n5614), .B(n5667), .C(n3762), .Y(n2376) );
  OAI21X1 U1175 ( .A(n5614), .B(n5666), .C(n3494), .Y(n2377) );
  OAI21X1 U1177 ( .A(n5614), .B(n5665), .C(n3583), .Y(n2378) );
  OAI21X1 U1179 ( .A(n5614), .B(n5664), .C(n3672), .Y(n2379) );
  OAI21X1 U1181 ( .A(n5614), .B(n5663), .C(n4044), .Y(n2380) );
  OAI21X1 U1183 ( .A(n5614), .B(n5662), .C(n4136), .Y(n2381) );
  OAI21X1 U1185 ( .A(n5614), .B(n5661), .C(n3859), .Y(n2382) );
  OAI21X1 U1187 ( .A(n5614), .B(n5660), .C(n3952), .Y(n2383) );
  OAI21X1 U1189 ( .A(n5614), .B(n5659), .C(n318), .Y(n2384) );
  OAI21X1 U1191 ( .A(n5614), .B(n5658), .C(n3761), .Y(n2385) );
  OAI21X1 U1193 ( .A(n5614), .B(n5657), .C(n3493), .Y(n2386) );
  OAI21X1 U1195 ( .A(n5614), .B(n5656), .C(n3582), .Y(n2387) );
  OAI21X1 U1197 ( .A(n5614), .B(n5655), .C(n3951), .Y(n2388) );
  OAI21X1 U1199 ( .A(n5614), .B(n5654), .C(n398), .Y(n2389) );
  OAI21X1 U1201 ( .A(n5614), .B(n5653), .C(n174), .Y(n2390) );
  OAI21X1 U1203 ( .A(n5614), .B(n5652), .C(n246), .Y(n2391) );
  OAI21X1 U1205 ( .A(n5614), .B(n5651), .C(n3347), .Y(n2392) );
  OAI21X1 U1207 ( .A(n5614), .B(n5650), .C(n3420), .Y(n2393) );
  OAI21X1 U1209 ( .A(n5614), .B(n5649), .C(n4043), .Y(n2394) );
  OAI21X1 U1211 ( .A(n5614), .B(n5648), .C(n4135), .Y(n2395) );
  OAI21X1 U1213 ( .A(n5614), .B(n5647), .C(n3858), .Y(n2396) );
  OAI21X1 U1215 ( .A(n5614), .B(n5646), .C(n3204), .Y(n2397) );
  OAI21X1 U1217 ( .A(n5614), .B(n5645), .C(n3275), .Y(n2398) );
  OAI21X1 U1219 ( .A(n5614), .B(n5644), .C(n114), .Y(n2399) );
  OAI21X1 U1221 ( .A(n5614), .B(n5643), .C(n3671), .Y(n2400) );
  OAI21X1 U1223 ( .A(n5614), .B(n5642), .C(n3950), .Y(n2401) );
  OAI21X1 U1225 ( .A(n5614), .B(n5641), .C(n3760), .Y(n2402) );
  OAI21X1 U1227 ( .A(n5614), .B(n5640), .C(n3492), .Y(n2403) );
  OAI21X1 U1229 ( .A(n5614), .B(n5639), .C(n3581), .Y(n2404) );
  OAI21X1 U1231 ( .A(n5614), .B(n5638), .C(n317), .Y(n2405) );
  OAI21X1 U1233 ( .A(n5614), .B(n5637), .C(n396), .Y(n2406) );
  OAI21X1 U1235 ( .A(n5614), .B(n5636), .C(n173), .Y(n2407) );
  OAI21X1 U1237 ( .A(n5614), .B(n5635), .C(n245), .Y(n2408) );
  OAI21X1 U1239 ( .A(n5614), .B(n5634), .C(n4042), .Y(n2409) );
  OAI21X1 U1241 ( .A(n5614), .B(n5633), .C(n4134), .Y(n2410) );
  OAI21X1 U1243 ( .A(n5614), .B(n5632), .C(n3857), .Y(n2411) );
  OAI21X1 U1245 ( .A(n5614), .B(n5631), .C(n3346), .Y(n2412) );
  OAI21X1 U1247 ( .A(n5614), .B(n5630), .C(n3419), .Y(n2413) );
  OAI21X1 U1249 ( .A(n5614), .B(n5629), .C(n3203), .Y(n2414) );
  OAI21X1 U1251 ( .A(n5614), .B(n5628), .C(n316), .Y(n2415) );
  OAI21X1 U1253 ( .A(n3623), .B(n4179), .C(reset), .Y(n1018) );
  OAI21X1 U1254 ( .A(n5613), .B(n5668), .C(n3580), .Y(n2416) );
  OAI21X1 U1256 ( .A(n5613), .B(n5667), .C(n3491), .Y(n2417) );
  OAI21X1 U1258 ( .A(n5613), .B(n5666), .C(n3759), .Y(n2418) );
  OAI21X1 U1260 ( .A(n5613), .B(n5665), .C(n3670), .Y(n2419) );
  OAI21X1 U1262 ( .A(n5613), .B(n5664), .C(n3579), .Y(n2420) );
  OAI21X1 U1264 ( .A(n5613), .B(n5663), .C(n3949), .Y(n2421) );
  OAI21X1 U1266 ( .A(n5613), .B(n5662), .C(n3856), .Y(n2422) );
  OAI21X1 U1268 ( .A(n5613), .B(n5661), .C(n4133), .Y(n2423) );
  OAI21X1 U1270 ( .A(n5613), .B(n5660), .C(n4041), .Y(n2424) );
  OAI21X1 U1272 ( .A(n5613), .B(n5659), .C(n244), .Y(n2425) );
  OAI21X1 U1274 ( .A(n5613), .B(n5658), .C(n3490), .Y(n2426) );
  OAI21X1 U1276 ( .A(n5613), .B(n5657), .C(n3758), .Y(n2427) );
  OAI21X1 U1278 ( .A(n5613), .B(n5656), .C(n3669), .Y(n2428) );
  OAI21X1 U1280 ( .A(n5613), .B(n5655), .C(n4040), .Y(n2429) );
  OAI21X1 U1282 ( .A(n5613), .B(n5654), .C(n172), .Y(n2430) );
  OAI21X1 U1284 ( .A(n5613), .B(n5653), .C(n394), .Y(n2431) );
  OAI21X1 U1286 ( .A(n5613), .B(n5652), .C(n315), .Y(n2432) );
  OAI21X1 U1288 ( .A(n5613), .B(n5651), .C(n3274), .Y(n2433) );
  OAI21X1 U1290 ( .A(n5613), .B(n5650), .C(n3202), .Y(n2434) );
  OAI21X1 U1292 ( .A(n5613), .B(n5649), .C(n3948), .Y(n2435) );
  OAI21X1 U1294 ( .A(n5613), .B(n5648), .C(n3855), .Y(n2436) );
  OAI21X1 U1296 ( .A(n5613), .B(n5647), .C(n4132), .Y(n2437) );
  OAI21X1 U1298 ( .A(n5613), .B(n5646), .C(n3418), .Y(n2438) );
  OAI21X1 U1300 ( .A(n5613), .B(n5645), .C(n3345), .Y(n2439) );
  OAI21X1 U1302 ( .A(n5613), .B(n5644), .C(n113), .Y(n2440) );
  OAI21X1 U1304 ( .A(n5613), .B(n5643), .C(n3578), .Y(n2441) );
  OAI21X1 U1306 ( .A(n5613), .B(n5642), .C(n4039), .Y(n2442) );
  OAI21X1 U1308 ( .A(n5613), .B(n5641), .C(n3489), .Y(n2443) );
  OAI21X1 U1310 ( .A(n5613), .B(n5640), .C(n3757), .Y(n2444) );
  OAI21X1 U1312 ( .A(n5613), .B(n5639), .C(n3668), .Y(n2445) );
  OAI21X1 U1314 ( .A(n5613), .B(n5638), .C(n243), .Y(n2446) );
  OAI21X1 U1316 ( .A(n5613), .B(n5637), .C(n171), .Y(n2447) );
  OAI21X1 U1318 ( .A(n5613), .B(n5636), .C(n392), .Y(n2448) );
  OAI21X1 U1320 ( .A(n5613), .B(n5635), .C(n314), .Y(n2449) );
  OAI21X1 U1322 ( .A(n5613), .B(n5634), .C(n3947), .Y(n2450) );
  OAI21X1 U1324 ( .A(n5613), .B(n5633), .C(n3854), .Y(n2451) );
  OAI21X1 U1326 ( .A(n5613), .B(n5632), .C(n4131), .Y(n2452) );
  OAI21X1 U1328 ( .A(n5613), .B(n5631), .C(n3273), .Y(n2453) );
  OAI21X1 U1330 ( .A(n5613), .B(n5630), .C(n3201), .Y(n2454) );
  OAI21X1 U1332 ( .A(n5613), .B(n5629), .C(n3417), .Y(n2455) );
  OAI21X1 U1334 ( .A(n5613), .B(n5628), .C(n242), .Y(n2456) );
  OAI21X1 U1336 ( .A(n3713), .B(n4179), .C(reset), .Y(n1060) );
  OAI21X1 U1337 ( .A(n5612), .B(n5668), .C(n3488), .Y(n2457) );
  OAI21X1 U1339 ( .A(n5612), .B(n5667), .C(n3577), .Y(n2458) );
  OAI21X1 U1341 ( .A(n5612), .B(n5666), .C(n3667), .Y(n2459) );
  OAI21X1 U1343 ( .A(n5612), .B(n5665), .C(n3756), .Y(n2460) );
  OAI21X1 U1345 ( .A(n5612), .B(n5664), .C(n3487), .Y(n2461) );
  OAI21X1 U1347 ( .A(n5612), .B(n5663), .C(n3853), .Y(n2462) );
  OAI21X1 U1349 ( .A(n5612), .B(n5662), .C(n3946), .Y(n2463) );
  OAI21X1 U1351 ( .A(n5612), .B(n5661), .C(n4038), .Y(n2464) );
  OAI21X1 U1353 ( .A(n5612), .B(n5660), .C(n4130), .Y(n2465) );
  OAI21X1 U1355 ( .A(n5612), .B(n5659), .C(n170), .Y(n2466) );
  OAI21X1 U1357 ( .A(n5612), .B(n5658), .C(n3576), .Y(n2467) );
  OAI21X1 U1359 ( .A(n5612), .B(n5657), .C(n3666), .Y(n2468) );
  OAI21X1 U1361 ( .A(n5612), .B(n5656), .C(n3755), .Y(n2469) );
  OAI21X1 U1363 ( .A(n5612), .B(n5655), .C(n4129), .Y(n2470) );
  OAI21X1 U1365 ( .A(n5612), .B(n5654), .C(n241), .Y(n2471) );
  OAI21X1 U1367 ( .A(n5612), .B(n5653), .C(n313), .Y(n2472) );
  OAI21X1 U1369 ( .A(n5612), .B(n5652), .C(n390), .Y(n2473) );
  OAI21X1 U1371 ( .A(n5612), .B(n5651), .C(n3200), .Y(n2474) );
  OAI21X1 U1373 ( .A(n5612), .B(n5650), .C(n3272), .Y(n2475) );
  OAI21X1 U1375 ( .A(n5612), .B(n5649), .C(n3852), .Y(n2476) );
  OAI21X1 U1377 ( .A(n5612), .B(n5648), .C(n3945), .Y(n2477) );
  OAI21X1 U1379 ( .A(n5612), .B(n5647), .C(n4037), .Y(n2478) );
  OAI21X1 U1381 ( .A(n5612), .B(n5646), .C(n3344), .Y(n2479) );
  OAI21X1 U1383 ( .A(n5612), .B(n5645), .C(n3416), .Y(n2480) );
  OAI21X1 U1385 ( .A(n5612), .B(n5644), .C(n112), .Y(n2481) );
  OAI21X1 U1387 ( .A(n5612), .B(n5643), .C(n3486), .Y(n2482) );
  OAI21X1 U1389 ( .A(n5612), .B(n5642), .C(n4128), .Y(n2483) );
  OAI21X1 U1391 ( .A(n5612), .B(n5641), .C(n3575), .Y(n2484) );
  OAI21X1 U1393 ( .A(n5612), .B(n5640), .C(n3665), .Y(n2485) );
  OAI21X1 U1395 ( .A(n5612), .B(n5639), .C(n3754), .Y(n2486) );
  OAI21X1 U1397 ( .A(n5612), .B(n5638), .C(n169), .Y(n2487) );
  OAI21X1 U1399 ( .A(n5612), .B(n5637), .C(n240), .Y(n2488) );
  OAI21X1 U1401 ( .A(n5612), .B(n5636), .C(n312), .Y(n2489) );
  OAI21X1 U1403 ( .A(n5612), .B(n5635), .C(n388), .Y(n2490) );
  OAI21X1 U1405 ( .A(n5612), .B(n5634), .C(n3851), .Y(n2491) );
  OAI21X1 U1407 ( .A(n5612), .B(n5633), .C(n3944), .Y(n2492) );
  OAI21X1 U1409 ( .A(n5612), .B(n5632), .C(n4036), .Y(n2493) );
  OAI21X1 U1411 ( .A(n5612), .B(n5631), .C(n3199), .Y(n2494) );
  OAI21X1 U1413 ( .A(n5612), .B(n5630), .C(n3271), .Y(n2495) );
  OAI21X1 U1415 ( .A(n5612), .B(n5629), .C(n3343), .Y(n2496) );
  OAI21X1 U1417 ( .A(n5612), .B(n5628), .C(n168), .Y(n2497) );
  OAI21X1 U1419 ( .A(n3805), .B(n4179), .C(reset), .Y(n1102) );
  NAND3X1 U1420 ( .A(n1777), .B(n5717), .C(wr_ptr[3]), .Y(n808) );
  OAI21X1 U1421 ( .A(n5611), .B(n5668), .C(n3415), .Y(n2498) );
  OAI21X1 U1423 ( .A(n5611), .B(n5667), .C(n3342), .Y(n2499) );
  OAI21X1 U1425 ( .A(n5611), .B(n5666), .C(n3270), .Y(n2500) );
  OAI21X1 U1427 ( .A(n5611), .B(n5665), .C(n3198), .Y(n2501) );
  OAI21X1 U1429 ( .A(n5611), .B(n5664), .C(n3414), .Y(n2502) );
  OAI21X1 U1431 ( .A(n5611), .B(n5663), .C(n386), .Y(n2503) );
  OAI21X1 U1433 ( .A(n5611), .B(n5662), .C(n311), .Y(n2504) );
  OAI21X1 U1435 ( .A(n5611), .B(n5661), .C(n239), .Y(n2505) );
  OAI21X1 U1437 ( .A(n5611), .B(n5660), .C(n167), .Y(n2506) );
  OAI21X1 U1439 ( .A(n5611), .B(n5659), .C(n4127), .Y(n2507) );
  OAI21X1 U1441 ( .A(n5611), .B(n5658), .C(n3341), .Y(n2508) );
  OAI21X1 U1443 ( .A(n5611), .B(n5657), .C(n3269), .Y(n2509) );
  OAI21X1 U1445 ( .A(n5611), .B(n5656), .C(n3197), .Y(n2510) );
  OAI21X1 U1447 ( .A(n5611), .B(n5655), .C(n166), .Y(n2511) );
  OAI21X1 U1449 ( .A(n5611), .B(n5654), .C(n4035), .Y(n2512) );
  OAI21X1 U1451 ( .A(n5611), .B(n5653), .C(n3943), .Y(n2513) );
  OAI21X1 U1453 ( .A(n5611), .B(n5652), .C(n3850), .Y(n2514) );
  OAI21X1 U1455 ( .A(n5611), .B(n5651), .C(n3753), .Y(n2515) );
  OAI21X1 U1457 ( .A(n5611), .B(n5650), .C(n3664), .Y(n2516) );
  OAI21X1 U1459 ( .A(n5611), .B(n5649), .C(n384), .Y(n2517) );
  OAI21X1 U1461 ( .A(n5611), .B(n5648), .C(n310), .Y(n2518) );
  OAI21X1 U1463 ( .A(n5611), .B(n5647), .C(n238), .Y(n2519) );
  OAI21X1 U1465 ( .A(n5611), .B(n5646), .C(n3574), .Y(n2520) );
  OAI21X1 U1467 ( .A(n5611), .B(n5645), .C(n3485), .Y(n2521) );
  OAI21X1 U1469 ( .A(n5611), .B(n5644), .C(n111), .Y(n2522) );
  OAI21X1 U1471 ( .A(n5611), .B(n5643), .C(n3413), .Y(n2523) );
  OAI21X1 U1473 ( .A(n5611), .B(n5642), .C(n165), .Y(n2524) );
  OAI21X1 U1475 ( .A(n5611), .B(n5641), .C(n3340), .Y(n2525) );
  OAI21X1 U1477 ( .A(n5611), .B(n5640), .C(n3268), .Y(n2526) );
  OAI21X1 U1479 ( .A(n5611), .B(n5639), .C(n3196), .Y(n2527) );
  OAI21X1 U1481 ( .A(n5611), .B(n5638), .C(n4126), .Y(n2528) );
  OAI21X1 U1483 ( .A(n5611), .B(n5637), .C(n4034), .Y(n2529) );
  OAI21X1 U1485 ( .A(n5611), .B(n5636), .C(n3942), .Y(n2530) );
  OAI21X1 U1487 ( .A(n5611), .B(n5635), .C(n3849), .Y(n2531) );
  OAI21X1 U1489 ( .A(n5611), .B(n5634), .C(n382), .Y(n2532) );
  OAI21X1 U1491 ( .A(n5611), .B(n5633), .C(n309), .Y(n2533) );
  OAI21X1 U1493 ( .A(n5611), .B(n5632), .C(n237), .Y(n2534) );
  OAI21X1 U1495 ( .A(n5611), .B(n5631), .C(n3752), .Y(n2535) );
  OAI21X1 U1497 ( .A(n5611), .B(n5630), .C(n3663), .Y(n2536) );
  OAI21X1 U1499 ( .A(n5611), .B(n5629), .C(n3573), .Y(n2537) );
  OAI21X1 U1501 ( .A(n5611), .B(n5628), .C(n4125), .Y(n2538) );
  OAI21X1 U1503 ( .A(n3806), .B(n4085), .C(reset), .Y(n1144) );
  OAI21X1 U1504 ( .A(n5610), .B(n5668), .C(n3339), .Y(n2539) );
  OAI21X1 U1506 ( .A(n5610), .B(n5667), .C(n3412), .Y(n2540) );
  OAI21X1 U1508 ( .A(n5610), .B(n5666), .C(n3195), .Y(n2541) );
  OAI21X1 U1510 ( .A(n5610), .B(n5665), .C(n3267), .Y(n2542) );
  OAI21X1 U1512 ( .A(n5610), .B(n5664), .C(n3338), .Y(n2543) );
  OAI21X1 U1514 ( .A(n5610), .B(n5663), .C(n308), .Y(n2544) );
  OAI21X1 U1516 ( .A(n5610), .B(n5662), .C(n380), .Y(n2545) );
  OAI21X1 U1518 ( .A(n5610), .B(n5661), .C(n164), .Y(n2546) );
  OAI21X1 U1520 ( .A(n5610), .B(n5660), .C(n236), .Y(n2547) );
  OAI21X1 U1522 ( .A(n5610), .B(n5659), .C(n4033), .Y(n2548) );
  OAI21X1 U1524 ( .A(n5610), .B(n5658), .C(n3411), .Y(n2549) );
  OAI21X1 U1526 ( .A(n5610), .B(n5657), .C(n3194), .Y(n2550) );
  OAI21X1 U1528 ( .A(n5610), .B(n5656), .C(n3266), .Y(n2551) );
  OAI21X1 U1530 ( .A(n5610), .B(n5655), .C(n235), .Y(n2552) );
  OAI21X1 U1532 ( .A(n5610), .B(n5654), .C(n4124), .Y(n2553) );
  OAI21X1 U1534 ( .A(n5610), .B(n5653), .C(n3848), .Y(n2554) );
  OAI21X1 U1536 ( .A(n5610), .B(n5652), .C(n3941), .Y(n2555) );
  OAI21X1 U1538 ( .A(n5610), .B(n5651), .C(n3662), .Y(n2556) );
  OAI21X1 U1540 ( .A(n5610), .B(n5650), .C(n3751), .Y(n2557) );
  OAI21X1 U1542 ( .A(n5610), .B(n5649), .C(n307), .Y(n2558) );
  OAI21X1 U1544 ( .A(n5610), .B(n5648), .C(n379), .Y(n2559) );
  OAI21X1 U1546 ( .A(n5610), .B(n5647), .C(n163), .Y(n2560) );
  OAI21X1 U1548 ( .A(n5610), .B(n5646), .C(n3484), .Y(n2561) );
  OAI21X1 U1550 ( .A(n5610), .B(n5645), .C(n3572), .Y(n2562) );
  OAI21X1 U1552 ( .A(n5610), .B(n5644), .C(n110), .Y(n2563) );
  OAI21X1 U1554 ( .A(n5610), .B(n5643), .C(n3337), .Y(n2564) );
  OAI21X1 U1556 ( .A(n5610), .B(n5642), .C(n234), .Y(n2565) );
  OAI21X1 U1558 ( .A(n5610), .B(n5641), .C(n3410), .Y(n2566) );
  OAI21X1 U1560 ( .A(n5610), .B(n5640), .C(n3193), .Y(n2567) );
  OAI21X1 U1562 ( .A(n5610), .B(n5639), .C(n3265), .Y(n2568) );
  OAI21X1 U1564 ( .A(n5610), .B(n5638), .C(n4032), .Y(n2569) );
  OAI21X1 U1566 ( .A(n5610), .B(n5637), .C(n4123), .Y(n2570) );
  OAI21X1 U1568 ( .A(n5610), .B(n5636), .C(n3847), .Y(n2571) );
  OAI21X1 U1570 ( .A(n5610), .B(n5635), .C(n3940), .Y(n2572) );
  OAI21X1 U1572 ( .A(n5610), .B(n5634), .C(n306), .Y(n2573) );
  OAI21X1 U1574 ( .A(n5610), .B(n5633), .C(n378), .Y(n2574) );
  OAI21X1 U1576 ( .A(n5610), .B(n5632), .C(n162), .Y(n2575) );
  OAI21X1 U1578 ( .A(n5610), .B(n5631), .C(n3661), .Y(n2576) );
  OAI21X1 U1580 ( .A(n5610), .B(n5630), .C(n3750), .Y(n2577) );
  OAI21X1 U1582 ( .A(n5610), .B(n5629), .C(n3483), .Y(n2578) );
  OAI21X1 U1584 ( .A(n5610), .B(n5628), .C(n4031), .Y(n2579) );
  OAI21X1 U1586 ( .A(n3714), .B(n4085), .C(reset), .Y(n1187) );
  OAI21X1 U1587 ( .A(n5609), .B(n5668), .C(n3264), .Y(n2580) );
  OAI21X1 U1589 ( .A(n5609), .B(n5667), .C(n3192), .Y(n2581) );
  OAI21X1 U1591 ( .A(n5609), .B(n5666), .C(n3409), .Y(n2582) );
  OAI21X1 U1593 ( .A(n5609), .B(n5665), .C(n3336), .Y(n2583) );
  OAI21X1 U1595 ( .A(n5609), .B(n5664), .C(n3263), .Y(n2584) );
  OAI21X1 U1597 ( .A(n5609), .B(n5663), .C(n233), .Y(n2585) );
  OAI21X1 U1599 ( .A(n5609), .B(n5662), .C(n161), .Y(n2586) );
  OAI21X1 U1601 ( .A(n5609), .B(n5661), .C(n377), .Y(n2587) );
  OAI21X1 U1603 ( .A(n5609), .B(n5660), .C(n305), .Y(n2588) );
  OAI21X1 U1605 ( .A(n5609), .B(n5659), .C(n3939), .Y(n2589) );
  OAI21X1 U1607 ( .A(n5609), .B(n5658), .C(n3191), .Y(n2590) );
  OAI21X1 U1609 ( .A(n5609), .B(n5657), .C(n3408), .Y(n2591) );
  OAI21X1 U1611 ( .A(n5609), .B(n5656), .C(n3335), .Y(n2592) );
  OAI21X1 U1613 ( .A(n5609), .B(n5655), .C(n304), .Y(n2593) );
  OAI21X1 U1615 ( .A(n5609), .B(n5654), .C(n3846), .Y(n2594) );
  OAI21X1 U1617 ( .A(n5609), .B(n5653), .C(n4122), .Y(n2595) );
  OAI21X1 U1619 ( .A(n5609), .B(n5652), .C(n4030), .Y(n2596) );
  OAI21X1 U1621 ( .A(n5609), .B(n5651), .C(n3571), .Y(n2597) );
  OAI21X1 U1623 ( .A(n5609), .B(n5650), .C(n3482), .Y(n2598) );
  OAI21X1 U1625 ( .A(n5609), .B(n5649), .C(n232), .Y(n2599) );
  OAI21X1 U1627 ( .A(n5609), .B(n5648), .C(n160), .Y(n2600) );
  OAI21X1 U1629 ( .A(n5609), .B(n5647), .C(n376), .Y(n2601) );
  OAI21X1 U1631 ( .A(n5609), .B(n5646), .C(n3749), .Y(n2602) );
  OAI21X1 U1633 ( .A(n5609), .B(n5645), .C(n3660), .Y(n2603) );
  OAI21X1 U1635 ( .A(n5609), .B(n5644), .C(n109), .Y(n2604) );
  OAI21X1 U1637 ( .A(n5609), .B(n5643), .C(n3262), .Y(n2605) );
  OAI21X1 U1639 ( .A(n5609), .B(n5642), .C(n303), .Y(n2606) );
  OAI21X1 U1641 ( .A(n5609), .B(n5641), .C(n3190), .Y(n2607) );
  OAI21X1 U1643 ( .A(n5609), .B(n5640), .C(n3407), .Y(n2608) );
  OAI21X1 U1645 ( .A(n5609), .B(n5639), .C(n3334), .Y(n2609) );
  OAI21X1 U1647 ( .A(n5609), .B(n5638), .C(n3938), .Y(n2610) );
  OAI21X1 U1649 ( .A(n5609), .B(n5637), .C(n3845), .Y(n2611) );
  OAI21X1 U1651 ( .A(n5609), .B(n5636), .C(n4121), .Y(n2612) );
  OAI21X1 U1653 ( .A(n5609), .B(n5635), .C(n4029), .Y(n2613) );
  OAI21X1 U1655 ( .A(n5609), .B(n5634), .C(n231), .Y(n2614) );
  OAI21X1 U1657 ( .A(n5609), .B(n5633), .C(n159), .Y(n2615) );
  OAI21X1 U1659 ( .A(n5609), .B(n5632), .C(n375), .Y(n2616) );
  OAI21X1 U1661 ( .A(n5609), .B(n5631), .C(n3570), .Y(n2617) );
  OAI21X1 U1663 ( .A(n5609), .B(n5630), .C(n3481), .Y(n2618) );
  OAI21X1 U1665 ( .A(n5609), .B(n5629), .C(n3748), .Y(n2619) );
  OAI21X1 U1667 ( .A(n5609), .B(n5628), .C(n3937), .Y(n2620) );
  OAI21X1 U1669 ( .A(n3624), .B(n4085), .C(reset), .Y(n1229) );
  OAI21X1 U1670 ( .A(n5608), .B(n5668), .C(n3189), .Y(n2621) );
  OAI21X1 U1672 ( .A(n5608), .B(n5667), .C(n3261), .Y(n2622) );
  OAI21X1 U1674 ( .A(n5608), .B(n5666), .C(n3333), .Y(n2623) );
  OAI21X1 U1676 ( .A(n5608), .B(n5665), .C(n3406), .Y(n2624) );
  OAI21X1 U1678 ( .A(n5608), .B(n5664), .C(n3188), .Y(n2625) );
  OAI21X1 U1680 ( .A(n5608), .B(n5663), .C(n158), .Y(n2626) );
  OAI21X1 U1682 ( .A(n5608), .B(n5662), .C(n230), .Y(n2627) );
  OAI21X1 U1684 ( .A(n5608), .B(n5661), .C(n302), .Y(n2628) );
  OAI21X1 U1686 ( .A(n5608), .B(n5660), .C(n374), .Y(n2629) );
  OAI21X1 U1688 ( .A(n5608), .B(n5659), .C(n3844), .Y(n2630) );
  OAI21X1 U1690 ( .A(n5608), .B(n5658), .C(n3260), .Y(n2631) );
  OAI21X1 U1692 ( .A(n5608), .B(n5657), .C(n3332), .Y(n2632) );
  OAI21X1 U1694 ( .A(n5608), .B(n5656), .C(n3405), .Y(n2633) );
  OAI21X1 U1696 ( .A(n5608), .B(n5655), .C(n373), .Y(n2634) );
  OAI21X1 U1698 ( .A(n5608), .B(n5654), .C(n3936), .Y(n2635) );
  OAI21X1 U1700 ( .A(n5608), .B(n5653), .C(n4028), .Y(n2636) );
  OAI21X1 U1702 ( .A(n5608), .B(n5652), .C(n4120), .Y(n2637) );
  OAI21X1 U1704 ( .A(n5608), .B(n5651), .C(n3480), .Y(n2638) );
  OAI21X1 U1706 ( .A(n5608), .B(n5650), .C(n3569), .Y(n2639) );
  OAI21X1 U1708 ( .A(n5608), .B(n5649), .C(n157), .Y(n2640) );
  OAI21X1 U1710 ( .A(n5608), .B(n5648), .C(n229), .Y(n2641) );
  OAI21X1 U1712 ( .A(n5608), .B(n5647), .C(n301), .Y(n2642) );
  OAI21X1 U1714 ( .A(n5608), .B(n5646), .C(n3659), .Y(n2643) );
  OAI21X1 U1716 ( .A(n5608), .B(n5645), .C(n3747), .Y(n2644) );
  OAI21X1 U1718 ( .A(n5608), .B(n5644), .C(n108), .Y(n2645) );
  OAI21X1 U1720 ( .A(n5608), .B(n5643), .C(n3187), .Y(n2646) );
  OAI21X1 U1722 ( .A(n5608), .B(n5642), .C(n372), .Y(n2647) );
  OAI21X1 U1724 ( .A(n5608), .B(n5641), .C(n3259), .Y(n2648) );
  OAI21X1 U1726 ( .A(n5608), .B(n5640), .C(n3331), .Y(n2649) );
  OAI21X1 U1728 ( .A(n5608), .B(n5639), .C(n3404), .Y(n2650) );
  OAI21X1 U1730 ( .A(n5608), .B(n5638), .C(n3843), .Y(n2651) );
  OAI21X1 U1732 ( .A(n5608), .B(n5637), .C(n3935), .Y(n2652) );
  OAI21X1 U1734 ( .A(n5608), .B(n5636), .C(n4027), .Y(n2653) );
  OAI21X1 U1736 ( .A(n5608), .B(n5635), .C(n4119), .Y(n2654) );
  OAI21X1 U1738 ( .A(n5608), .B(n5634), .C(n156), .Y(n2655) );
  OAI21X1 U1740 ( .A(n5608), .B(n5633), .C(n228), .Y(n2656) );
  OAI21X1 U1742 ( .A(n5608), .B(n5632), .C(n300), .Y(n2657) );
  OAI21X1 U1744 ( .A(n5608), .B(n5631), .C(n3479), .Y(n2658) );
  OAI21X1 U1746 ( .A(n5608), .B(n5630), .C(n3568), .Y(n2659) );
  OAI21X1 U1748 ( .A(n5608), .B(n5629), .C(n3658), .Y(n2660) );
  OAI21X1 U1750 ( .A(n5608), .B(n5628), .C(n3842), .Y(n2661) );
  OAI21X1 U1752 ( .A(n3535), .B(n4085), .C(reset), .Y(n1271) );
  OAI21X1 U1753 ( .A(n5607), .B(n5668), .C(n4118), .Y(n2662) );
  OAI21X1 U1755 ( .A(n5607), .B(n5667), .C(n4026), .Y(n2663) );
  OAI21X1 U1757 ( .A(n5607), .B(n5666), .C(n3934), .Y(n2664) );
  OAI21X1 U1759 ( .A(n5607), .B(n5665), .C(n3841), .Y(n2665) );
  OAI21X1 U1761 ( .A(n5607), .B(n5664), .C(n4117), .Y(n2666) );
  OAI21X1 U1763 ( .A(n5607), .B(n5663), .C(n3746), .Y(n2667) );
  OAI21X1 U1765 ( .A(n5607), .B(n5662), .C(n3657), .Y(n2668) );
  OAI21X1 U1767 ( .A(n5607), .B(n5661), .C(n3567), .Y(n2669) );
  OAI21X1 U1769 ( .A(n5607), .B(n5660), .C(n3478), .Y(n2670) );
  OAI21X1 U1771 ( .A(n5607), .B(n5659), .C(n3403), .Y(n2671) );
  OAI21X1 U1773 ( .A(n5607), .B(n5658), .C(n4025), .Y(n2672) );
  OAI21X1 U1775 ( .A(n5607), .B(n5657), .C(n3933), .Y(n2673) );
  OAI21X1 U1777 ( .A(n5607), .B(n5656), .C(n3840), .Y(n2674) );
  OAI21X1 U1779 ( .A(n5607), .B(n5655), .C(n3477), .Y(n2675) );
  OAI21X1 U1781 ( .A(n5607), .B(n5654), .C(n3330), .Y(n2676) );
  OAI21X1 U1783 ( .A(n5607), .B(n5653), .C(n3258), .Y(n2677) );
  OAI21X1 U1785 ( .A(n5607), .B(n5652), .C(n3186), .Y(n2678) );
  OAI21X1 U1787 ( .A(n5607), .B(n5651), .C(n371), .Y(n2679) );
  OAI21X1 U1789 ( .A(n5607), .B(n5650), .C(n299), .Y(n2680) );
  OAI21X1 U1791 ( .A(n5607), .B(n5649), .C(n3745), .Y(n2681) );
  OAI21X1 U1793 ( .A(n5607), .B(n5648), .C(n3656), .Y(n2682) );
  OAI21X1 U1795 ( .A(n5607), .B(n5647), .C(n3566), .Y(n2683) );
  OAI21X1 U1797 ( .A(n5607), .B(n5646), .C(n227), .Y(n2684) );
  OAI21X1 U1799 ( .A(n5607), .B(n5645), .C(n155), .Y(n2685) );
  OAI21X1 U1801 ( .A(n5607), .B(n5644), .C(n107), .Y(n2686) );
  OAI21X1 U1803 ( .A(n5607), .B(n5643), .C(n4116), .Y(n2687) );
  OAI21X1 U1805 ( .A(n5607), .B(n5642), .C(n3476), .Y(n2688) );
  OAI21X1 U1807 ( .A(n5607), .B(n5641), .C(n4024), .Y(n2689) );
  OAI21X1 U1809 ( .A(n5607), .B(n5640), .C(n3932), .Y(n2690) );
  OAI21X1 U1811 ( .A(n5607), .B(n5639), .C(n3839), .Y(n2691) );
  OAI21X1 U1813 ( .A(n5607), .B(n5638), .C(n3402), .Y(n2692) );
  OAI21X1 U1815 ( .A(n5607), .B(n5637), .C(n3329), .Y(n2693) );
  OAI21X1 U1817 ( .A(n5607), .B(n5636), .C(n3257), .Y(n2694) );
  OAI21X1 U1819 ( .A(n5607), .B(n5635), .C(n3185), .Y(n2695) );
  OAI21X1 U1821 ( .A(n5607), .B(n5634), .C(n3744), .Y(n2696) );
  OAI21X1 U1823 ( .A(n5607), .B(n5633), .C(n3655), .Y(n2697) );
  OAI21X1 U1825 ( .A(n5607), .B(n5632), .C(n3565), .Y(n2698) );
  OAI21X1 U1827 ( .A(n5607), .B(n5631), .C(n370), .Y(n2699) );
  OAI21X1 U1829 ( .A(n5607), .B(n5630), .C(n298), .Y(n2700) );
  OAI21X1 U1831 ( .A(n5607), .B(n5629), .C(n226), .Y(n2701) );
  OAI21X1 U1833 ( .A(n5607), .B(n5628), .C(n3401), .Y(n2702) );
  OAI21X1 U1835 ( .A(n3534), .B(n4085), .C(reset), .Y(n1313) );
  OAI21X1 U1836 ( .A(n5606), .B(n5668), .C(n4023), .Y(n2703) );
  OAI21X1 U1838 ( .A(n5606), .B(n5667), .C(n4115), .Y(n2704) );
  OAI21X1 U1840 ( .A(n5606), .B(n5666), .C(n3838), .Y(n2705) );
  OAI21X1 U1842 ( .A(n5606), .B(n5665), .C(n3931), .Y(n2706) );
  OAI21X1 U1844 ( .A(n5606), .B(n5664), .C(n4022), .Y(n2707) );
  OAI21X1 U1846 ( .A(n5606), .B(n5663), .C(n3654), .Y(n2708) );
  OAI21X1 U1848 ( .A(n5606), .B(n5662), .C(n3743), .Y(n2709) );
  OAI21X1 U1850 ( .A(n5606), .B(n5661), .C(n3475), .Y(n2710) );
  OAI21X1 U1852 ( .A(n5606), .B(n5660), .C(n3564), .Y(n2711) );
  OAI21X1 U1854 ( .A(n5606), .B(n5659), .C(n3328), .Y(n2712) );
  OAI21X1 U1856 ( .A(n5606), .B(n5658), .C(n4114), .Y(n2713) );
  OAI21X1 U1858 ( .A(n5606), .B(n5657), .C(n3837), .Y(n2714) );
  OAI21X1 U1860 ( .A(n5606), .B(n5656), .C(n3930), .Y(n2715) );
  OAI21X1 U1862 ( .A(n5606), .B(n5655), .C(n3563), .Y(n2716) );
  OAI21X1 U1864 ( .A(n5606), .B(n5654), .C(n3400), .Y(n2717) );
  OAI21X1 U1866 ( .A(n5606), .B(n5653), .C(n3184), .Y(n2718) );
  OAI21X1 U1868 ( .A(n5606), .B(n5652), .C(n3256), .Y(n2719) );
  OAI21X1 U1870 ( .A(n5606), .B(n5651), .C(n297), .Y(n2720) );
  OAI21X1 U1872 ( .A(n5606), .B(n5650), .C(n369), .Y(n2721) );
  OAI21X1 U1874 ( .A(n5606), .B(n5649), .C(n3653), .Y(n2722) );
  OAI21X1 U1876 ( .A(n5606), .B(n5648), .C(n3742), .Y(n2723) );
  OAI21X1 U1878 ( .A(n5606), .B(n5647), .C(n3474), .Y(n2724) );
  OAI21X1 U1880 ( .A(n5606), .B(n5646), .C(n154), .Y(n2725) );
  OAI21X1 U1882 ( .A(n5606), .B(n5645), .C(n225), .Y(n2726) );
  OAI21X1 U1884 ( .A(n5606), .B(n5644), .C(n106), .Y(n2727) );
  OAI21X1 U1886 ( .A(n5606), .B(n5643), .C(n4021), .Y(n2728) );
  OAI21X1 U1888 ( .A(n5606), .B(n5642), .C(n3562), .Y(n2729) );
  OAI21X1 U1890 ( .A(n5606), .B(n5641), .C(n4113), .Y(n2730) );
  OAI21X1 U1892 ( .A(n5606), .B(n5640), .C(n3836), .Y(n2731) );
  OAI21X1 U1894 ( .A(n5606), .B(n5639), .C(n3929), .Y(n2732) );
  OAI21X1 U1896 ( .A(n5606), .B(n5638), .C(n3327), .Y(n2733) );
  OAI21X1 U1898 ( .A(n5606), .B(n5637), .C(n3399), .Y(n2734) );
  OAI21X1 U1900 ( .A(n5606), .B(n5636), .C(n3183), .Y(n2735) );
  OAI21X1 U1902 ( .A(n5606), .B(n5635), .C(n3255), .Y(n2736) );
  OAI21X1 U1904 ( .A(n5606), .B(n5634), .C(n3652), .Y(n2737) );
  OAI21X1 U1906 ( .A(n5606), .B(n5633), .C(n3741), .Y(n2738) );
  OAI21X1 U1908 ( .A(n5606), .B(n5632), .C(n3473), .Y(n2739) );
  OAI21X1 U1910 ( .A(n5606), .B(n5631), .C(n296), .Y(n2740) );
  OAI21X1 U1912 ( .A(n5606), .B(n5630), .C(n368), .Y(n2741) );
  OAI21X1 U1914 ( .A(n5606), .B(n5629), .C(n153), .Y(n2742) );
  OAI21X1 U1916 ( .A(n5606), .B(n5628), .C(n3326), .Y(n2743) );
  OAI21X1 U1918 ( .A(n3623), .B(n4085), .C(reset), .Y(n1355) );
  OAI21X1 U1919 ( .A(n5605), .B(n5668), .C(n3928), .Y(n2744) );
  OAI21X1 U1921 ( .A(n5605), .B(n5667), .C(n3835), .Y(n2745) );
  OAI21X1 U1923 ( .A(n5605), .B(n5666), .C(n4112), .Y(n2746) );
  OAI21X1 U1925 ( .A(n5605), .B(n5665), .C(n4020), .Y(n2747) );
  OAI21X1 U1927 ( .A(n5605), .B(n5664), .C(n3927), .Y(n2748) );
  OAI21X1 U1929 ( .A(n5605), .B(n5663), .C(n3561), .Y(n2749) );
  OAI21X1 U1931 ( .A(n5605), .B(n5662), .C(n3472), .Y(n2750) );
  OAI21X1 U1933 ( .A(n5605), .B(n5661), .C(n3740), .Y(n2751) );
  OAI21X1 U1935 ( .A(n5605), .B(n5660), .C(n3651), .Y(n2752) );
  OAI21X1 U1937 ( .A(n5605), .B(n5659), .C(n3254), .Y(n2753) );
  OAI21X1 U1939 ( .A(n5605), .B(n5658), .C(n3834), .Y(n2754) );
  OAI21X1 U1941 ( .A(n5605), .B(n5657), .C(n4111), .Y(n2755) );
  OAI21X1 U1943 ( .A(n5605), .B(n5656), .C(n4019), .Y(n2756) );
  OAI21X1 U1945 ( .A(n5605), .B(n5655), .C(n3650), .Y(n2757) );
  OAI21X1 U1947 ( .A(n5605), .B(n5654), .C(n3182), .Y(n2758) );
  OAI21X1 U1949 ( .A(n5605), .B(n5653), .C(n3398), .Y(n2759) );
  OAI21X1 U1951 ( .A(n5605), .B(n5652), .C(n3325), .Y(n2760) );
  OAI21X1 U1953 ( .A(n5605), .B(n5651), .C(n224), .Y(n2761) );
  OAI21X1 U1955 ( .A(n5605), .B(n5650), .C(n152), .Y(n2762) );
  OAI21X1 U1957 ( .A(n5605), .B(n5649), .C(n3560), .Y(n2763) );
  OAI21X1 U1959 ( .A(n5605), .B(n5648), .C(n3471), .Y(n2764) );
  OAI21X1 U1961 ( .A(n5605), .B(n5647), .C(n3739), .Y(n2765) );
  OAI21X1 U1963 ( .A(n5605), .B(n5646), .C(n367), .Y(n2766) );
  OAI21X1 U1965 ( .A(n5605), .B(n5645), .C(n295), .Y(n2767) );
  OAI21X1 U1967 ( .A(n5605), .B(n5644), .C(n105), .Y(n2768) );
  OAI21X1 U1969 ( .A(n5605), .B(n5643), .C(n3926), .Y(n2769) );
  OAI21X1 U1971 ( .A(n5605), .B(n5642), .C(n3649), .Y(n2770) );
  OAI21X1 U1973 ( .A(n5605), .B(n5641), .C(n3833), .Y(n2771) );
  OAI21X1 U1975 ( .A(n5605), .B(n5640), .C(n4110), .Y(n2772) );
  OAI21X1 U1977 ( .A(n5605), .B(n5639), .C(n4018), .Y(n2773) );
  OAI21X1 U1979 ( .A(n5605), .B(n5638), .C(n3253), .Y(n2774) );
  OAI21X1 U1981 ( .A(n5605), .B(n5637), .C(n3181), .Y(n2775) );
  OAI21X1 U1983 ( .A(n5605), .B(n5636), .C(n3397), .Y(n2776) );
  OAI21X1 U1985 ( .A(n5605), .B(n5635), .C(n3324), .Y(n2777) );
  OAI21X1 U1987 ( .A(n5605), .B(n5634), .C(n3559), .Y(n2778) );
  OAI21X1 U1989 ( .A(n5605), .B(n5633), .C(n3470), .Y(n2779) );
  OAI21X1 U1991 ( .A(n5605), .B(n5632), .C(n3738), .Y(n2780) );
  OAI21X1 U1993 ( .A(n5605), .B(n5631), .C(n223), .Y(n2781) );
  OAI21X1 U1995 ( .A(n5605), .B(n5630), .C(n151), .Y(n2782) );
  OAI21X1 U1997 ( .A(n5605), .B(n5629), .C(n366), .Y(n2783) );
  OAI21X1 U1999 ( .A(n5605), .B(n5628), .C(n3252), .Y(n2784) );
  OAI21X1 U2001 ( .A(n3713), .B(n4085), .C(reset), .Y(n1397) );
  OAI21X1 U2002 ( .A(n5604), .B(n5668), .C(n3832), .Y(n2785) );
  OAI21X1 U2004 ( .A(n5604), .B(n5667), .C(n3925), .Y(n2786) );
  OAI21X1 U2006 ( .A(n5604), .B(n5666), .C(n4017), .Y(n2787) );
  OAI21X1 U2008 ( .A(n5604), .B(n5665), .C(n4109), .Y(n2788) );
  OAI21X1 U2010 ( .A(n5604), .B(n5664), .C(n3831), .Y(n2789) );
  OAI21X1 U2012 ( .A(n5604), .B(n5663), .C(n3469), .Y(n2790) );
  OAI21X1 U2014 ( .A(n5604), .B(n5662), .C(n3558), .Y(n2791) );
  OAI21X1 U2016 ( .A(n5604), .B(n5661), .C(n3648), .Y(n2792) );
  OAI21X1 U2018 ( .A(n5604), .B(n5660), .C(n3737), .Y(n2793) );
  OAI21X1 U2020 ( .A(n5604), .B(n5659), .C(n3180), .Y(n2794) );
  OAI21X1 U2022 ( .A(n5604), .B(n5658), .C(n3924), .Y(n2795) );
  OAI21X1 U2024 ( .A(n5604), .B(n5657), .C(n4016), .Y(n2796) );
  OAI21X1 U2026 ( .A(n5604), .B(n5656), .C(n4108), .Y(n2797) );
  OAI21X1 U2028 ( .A(n5604), .B(n5655), .C(n3736), .Y(n2798) );
  OAI21X1 U2030 ( .A(n5604), .B(n5654), .C(n3251), .Y(n2799) );
  OAI21X1 U2032 ( .A(n5604), .B(n5653), .C(n3323), .Y(n2800) );
  OAI21X1 U2034 ( .A(n5604), .B(n5652), .C(n3396), .Y(n2801) );
  OAI21X1 U2036 ( .A(n5604), .B(n5651), .C(n150), .Y(n2802) );
  OAI21X1 U2038 ( .A(n5604), .B(n5650), .C(n222), .Y(n2803) );
  OAI21X1 U2040 ( .A(n5604), .B(n5649), .C(n3468), .Y(n2804) );
  OAI21X1 U2042 ( .A(n5604), .B(n5648), .C(n3557), .Y(n2805) );
  OAI21X1 U2044 ( .A(n5604), .B(n5647), .C(n3647), .Y(n2806) );
  OAI21X1 U2046 ( .A(n5604), .B(n5646), .C(n294), .Y(n2807) );
  OAI21X1 U2048 ( .A(n5604), .B(n5645), .C(n365), .Y(n2808) );
  OAI21X1 U2050 ( .A(n5604), .B(n5644), .C(n104), .Y(n2809) );
  OAI21X1 U2052 ( .A(n5604), .B(n5643), .C(n3830), .Y(n2810) );
  OAI21X1 U2054 ( .A(n5604), .B(n5642), .C(n3735), .Y(n2811) );
  OAI21X1 U2056 ( .A(n5604), .B(n5641), .C(n3923), .Y(n2812) );
  OAI21X1 U2058 ( .A(n5604), .B(n5640), .C(n4015), .Y(n2813) );
  OAI21X1 U2060 ( .A(n5604), .B(n5639), .C(n4107), .Y(n2814) );
  OAI21X1 U2062 ( .A(n5604), .B(n5638), .C(n3179), .Y(n2815) );
  OAI21X1 U2064 ( .A(n5604), .B(n5637), .C(n3250), .Y(n2816) );
  OAI21X1 U2066 ( .A(n5604), .B(n5636), .C(n3322), .Y(n2817) );
  OAI21X1 U2068 ( .A(n5604), .B(n5635), .C(n3395), .Y(n2818) );
  OAI21X1 U2070 ( .A(n5604), .B(n5634), .C(n3467), .Y(n2819) );
  OAI21X1 U2072 ( .A(n5604), .B(n5633), .C(n3556), .Y(n2820) );
  OAI21X1 U2074 ( .A(n5604), .B(n5632), .C(n3646), .Y(n2821) );
  OAI21X1 U2076 ( .A(n5604), .B(n5631), .C(n149), .Y(n2822) );
  OAI21X1 U2078 ( .A(n5604), .B(n5630), .C(n221), .Y(n2823) );
  OAI21X1 U2080 ( .A(n5604), .B(n5629), .C(n293), .Y(n2824) );
  OAI21X1 U2082 ( .A(n5604), .B(n5628), .C(n3178), .Y(n2825) );
  OAI21X1 U2084 ( .A(n3805), .B(n4085), .C(reset), .Y(n1439) );
  NAND3X1 U2085 ( .A(n1777), .B(n5720), .C(wr_ptr[4]), .Y(n1145) );
  OAI21X1 U2086 ( .A(n5603), .B(n5668), .C(n3734), .Y(n2826) );
  OAI21X1 U2088 ( .A(n5603), .B(n5667), .C(n3645), .Y(n2827) );
  OAI21X1 U2090 ( .A(n5603), .B(n5666), .C(n3555), .Y(n2828) );
  OAI21X1 U2092 ( .A(n5603), .B(n5665), .C(n3466), .Y(n2829) );
  OAI21X1 U2094 ( .A(n5603), .B(n5664), .C(n3733), .Y(n2830) );
  OAI21X1 U2096 ( .A(n5603), .B(n5663), .C(n4106), .Y(n2831) );
  OAI21X1 U2098 ( .A(n5603), .B(n5662), .C(n4014), .Y(n2832) );
  OAI21X1 U2100 ( .A(n5603), .B(n5661), .C(n3922), .Y(n2833) );
  OAI21X1 U2102 ( .A(n5603), .B(n5660), .C(n3829), .Y(n2834) );
  OAI21X1 U2104 ( .A(n5603), .B(n5659), .C(n364), .Y(n2835) );
  OAI21X1 U2106 ( .A(n5603), .B(n5658), .C(n3644), .Y(n2836) );
  OAI21X1 U2108 ( .A(n5603), .B(n5657), .C(n3554), .Y(n2837) );
  OAI21X1 U2110 ( .A(n5603), .B(n5656), .C(n3465), .Y(n2838) );
  OAI21X1 U2112 ( .A(n5603), .B(n5655), .C(n3828), .Y(n2839) );
  OAI21X1 U2114 ( .A(n5603), .B(n5654), .C(n292), .Y(n2840) );
  OAI21X1 U2116 ( .A(n5603), .B(n5653), .C(n220), .Y(n2841) );
  OAI21X1 U2118 ( .A(n5603), .B(n5652), .C(n148), .Y(n2842) );
  OAI21X1 U2120 ( .A(n5603), .B(n5651), .C(n3394), .Y(n2843) );
  OAI21X1 U2122 ( .A(n5603), .B(n5650), .C(n3321), .Y(n2844) );
  OAI21X1 U2124 ( .A(n5603), .B(n5649), .C(n4105), .Y(n2845) );
  OAI21X1 U2126 ( .A(n5603), .B(n5648), .C(n4013), .Y(n2846) );
  OAI21X1 U2128 ( .A(n5603), .B(n5647), .C(n3921), .Y(n2847) );
  OAI21X1 U2130 ( .A(n5603), .B(n5646), .C(n3249), .Y(n2848) );
  OAI21X1 U2132 ( .A(n5603), .B(n5645), .C(n3177), .Y(n2849) );
  OAI21X1 U2134 ( .A(n5603), .B(n5644), .C(n103), .Y(n2850) );
  OAI21X1 U2136 ( .A(n5603), .B(n5643), .C(n3732), .Y(n2851) );
  OAI21X1 U2138 ( .A(n5603), .B(n5642), .C(n3827), .Y(n2852) );
  OAI21X1 U2140 ( .A(n5603), .B(n5641), .C(n3643), .Y(n2853) );
  OAI21X1 U2142 ( .A(n5603), .B(n5640), .C(n3553), .Y(n2854) );
  OAI21X1 U2144 ( .A(n5603), .B(n5639), .C(n3464), .Y(n2855) );
  OAI21X1 U2146 ( .A(n5603), .B(n5638), .C(n363), .Y(n2856) );
  OAI21X1 U2148 ( .A(n5603), .B(n5637), .C(n291), .Y(n2857) );
  OAI21X1 U2150 ( .A(n5603), .B(n5636), .C(n219), .Y(n2858) );
  OAI21X1 U2152 ( .A(n5603), .B(n5635), .C(n147), .Y(n2859) );
  OAI21X1 U2154 ( .A(n5603), .B(n5634), .C(n4104), .Y(n2860) );
  OAI21X1 U2156 ( .A(n5603), .B(n5633), .C(n4012), .Y(n2861) );
  OAI21X1 U2158 ( .A(n5603), .B(n5632), .C(n3920), .Y(n2862) );
  OAI21X1 U2160 ( .A(n5603), .B(n5631), .C(n3393), .Y(n2863) );
  OAI21X1 U2162 ( .A(n5603), .B(n5630), .C(n3320), .Y(n2864) );
  OAI21X1 U2164 ( .A(n5603), .B(n5629), .C(n3248), .Y(n2865) );
  OAI21X1 U2166 ( .A(n5603), .B(n5628), .C(n362), .Y(n2866) );
  OAI21X1 U2168 ( .A(n3806), .B(n3992), .C(reset), .Y(n1481) );
  NAND3X1 U2169 ( .A(n5718), .B(n5719), .C(n5716), .Y(n464) );
  OAI21X1 U2170 ( .A(n5602), .B(n5668), .C(n3642), .Y(n2867) );
  OAI21X1 U2172 ( .A(n5602), .B(n5667), .C(n3731), .Y(n2868) );
  OAI21X1 U2174 ( .A(n5602), .B(n5666), .C(n3463), .Y(n2869) );
  OAI21X1 U2176 ( .A(n5602), .B(n5665), .C(n3552), .Y(n2870) );
  OAI21X1 U2178 ( .A(n5602), .B(n5664), .C(n3641), .Y(n2871) );
  OAI21X1 U2180 ( .A(n5602), .B(n5663), .C(n4011), .Y(n2872) );
  OAI21X1 U2182 ( .A(n5602), .B(n5662), .C(n4103), .Y(n2873) );
  OAI21X1 U2184 ( .A(n5602), .B(n5661), .C(n3826), .Y(n2874) );
  OAI21X1 U2186 ( .A(n5602), .B(n5660), .C(n3919), .Y(n2875) );
  OAI21X1 U2188 ( .A(n5602), .B(n5659), .C(n290), .Y(n2876) );
  OAI21X1 U2190 ( .A(n5602), .B(n5658), .C(n3730), .Y(n2877) );
  OAI21X1 U2192 ( .A(n5602), .B(n5657), .C(n3462), .Y(n2878) );
  OAI21X1 U2194 ( .A(n5602), .B(n5656), .C(n3551), .Y(n2879) );
  OAI21X1 U2196 ( .A(n5602), .B(n5655), .C(n3918), .Y(n2880) );
  OAI21X1 U2198 ( .A(n5602), .B(n5654), .C(n361), .Y(n2881) );
  OAI21X1 U2200 ( .A(n5602), .B(n5653), .C(n146), .Y(n2882) );
  OAI21X1 U2202 ( .A(n5602), .B(n5652), .C(n218), .Y(n2883) );
  OAI21X1 U2204 ( .A(n5602), .B(n5651), .C(n3319), .Y(n2884) );
  OAI21X1 U2206 ( .A(n5602), .B(n5650), .C(n3392), .Y(n2885) );
  OAI21X1 U2208 ( .A(n5602), .B(n5649), .C(n4010), .Y(n2886) );
  OAI21X1 U2210 ( .A(n5602), .B(n5648), .C(n4102), .Y(n2887) );
  OAI21X1 U2212 ( .A(n5602), .B(n5647), .C(n3825), .Y(n2888) );
  OAI21X1 U2214 ( .A(n5602), .B(n5646), .C(n3176), .Y(n2889) );
  OAI21X1 U2216 ( .A(n5602), .B(n5645), .C(n3247), .Y(n2890) );
  OAI21X1 U2218 ( .A(n5602), .B(n5644), .C(n102), .Y(n2891) );
  OAI21X1 U2220 ( .A(n5602), .B(n5643), .C(n3640), .Y(n2892) );
  OAI21X1 U2222 ( .A(n5602), .B(n5642), .C(n3917), .Y(n2893) );
  OAI21X1 U2224 ( .A(n5602), .B(n5641), .C(n3729), .Y(n2894) );
  OAI21X1 U2226 ( .A(n5602), .B(n5640), .C(n3461), .Y(n2895) );
  OAI21X1 U2228 ( .A(n5602), .B(n5639), .C(n3550), .Y(n2896) );
  OAI21X1 U2230 ( .A(n5602), .B(n5638), .C(n289), .Y(n2897) );
  OAI21X1 U2232 ( .A(n5602), .B(n5637), .C(n360), .Y(n2898) );
  OAI21X1 U2234 ( .A(n5602), .B(n5636), .C(n145), .Y(n2899) );
  OAI21X1 U2236 ( .A(n5602), .B(n5635), .C(n217), .Y(n2900) );
  OAI21X1 U2238 ( .A(n5602), .B(n5634), .C(n4009), .Y(n2901) );
  OAI21X1 U2240 ( .A(n5602), .B(n5633), .C(n4101), .Y(n2902) );
  OAI21X1 U2242 ( .A(n5602), .B(n5632), .C(n3824), .Y(n2903) );
  OAI21X1 U2244 ( .A(n5602), .B(n5631), .C(n3318), .Y(n2904) );
  OAI21X1 U2246 ( .A(n5602), .B(n5630), .C(n3391), .Y(n2905) );
  OAI21X1 U2248 ( .A(n5602), .B(n5629), .C(n3175), .Y(n2906) );
  OAI21X1 U2250 ( .A(n5602), .B(n5628), .C(n288), .Y(n2907) );
  OAI21X1 U2252 ( .A(n3714), .B(n3992), .C(reset), .Y(n1524) );
  NAND3X1 U2253 ( .A(n5718), .B(n5719), .C(wr_ptr[0]), .Y(n507) );
  OAI21X1 U2254 ( .A(n5601), .B(n5668), .C(n3549), .Y(n2908) );
  OAI21X1 U2256 ( .A(n5601), .B(n5667), .C(n3460), .Y(n2909) );
  OAI21X1 U2258 ( .A(n5601), .B(n5666), .C(n3728), .Y(n2910) );
  OAI21X1 U2260 ( .A(n5601), .B(n5665), .C(n3639), .Y(n2911) );
  OAI21X1 U2262 ( .A(n5601), .B(n5664), .C(n3548), .Y(n2912) );
  OAI21X1 U2264 ( .A(n5601), .B(n5663), .C(n3916), .Y(n2913) );
  OAI21X1 U2266 ( .A(n5601), .B(n5662), .C(n3823), .Y(n2914) );
  OAI21X1 U2268 ( .A(n5601), .B(n5661), .C(n4100), .Y(n2915) );
  OAI21X1 U2270 ( .A(n5601), .B(n5660), .C(n4008), .Y(n2916) );
  OAI21X1 U2272 ( .A(n5601), .B(n5659), .C(n216), .Y(n2917) );
  OAI21X1 U2274 ( .A(n5601), .B(n5658), .C(n3459), .Y(n2918) );
  OAI21X1 U2276 ( .A(n5601), .B(n5657), .C(n3727), .Y(n2919) );
  OAI21X1 U2278 ( .A(n5601), .B(n5656), .C(n3638), .Y(n2920) );
  OAI21X1 U2280 ( .A(n5601), .B(n5655), .C(n4007), .Y(n2921) );
  OAI21X1 U2282 ( .A(n5601), .B(n5654), .C(n144), .Y(n2922) );
  OAI21X1 U2284 ( .A(n5601), .B(n5653), .C(n359), .Y(n2923) );
  OAI21X1 U2286 ( .A(n5601), .B(n5652), .C(n287), .Y(n2924) );
  OAI21X1 U2288 ( .A(n5601), .B(n5651), .C(n3246), .Y(n2925) );
  OAI21X1 U2290 ( .A(n5601), .B(n5650), .C(n3174), .Y(n2926) );
  OAI21X1 U2292 ( .A(n5601), .B(n5649), .C(n3915), .Y(n2927) );
  OAI21X1 U2294 ( .A(n5601), .B(n5648), .C(n3822), .Y(n2928) );
  OAI21X1 U2296 ( .A(n5601), .B(n5647), .C(n4099), .Y(n2929) );
  OAI21X1 U2298 ( .A(n5601), .B(n5646), .C(n3390), .Y(n2930) );
  OAI21X1 U2300 ( .A(n5601), .B(n5645), .C(n3317), .Y(n2931) );
  OAI21X1 U2302 ( .A(n5601), .B(n5644), .C(n97), .Y(n2932) );
  OAI21X1 U2304 ( .A(n5601), .B(n5643), .C(n3547), .Y(n2933) );
  OAI21X1 U2306 ( .A(n5601), .B(n5642), .C(n4006), .Y(n2934) );
  OAI21X1 U2308 ( .A(n5601), .B(n5641), .C(n3458), .Y(n2935) );
  OAI21X1 U2310 ( .A(n5601), .B(n5640), .C(n3726), .Y(n2936) );
  OAI21X1 U2312 ( .A(n5601), .B(n5639), .C(n3637), .Y(n2937) );
  OAI21X1 U2314 ( .A(n5601), .B(n5638), .C(n215), .Y(n2938) );
  OAI21X1 U2316 ( .A(n5601), .B(n5637), .C(n143), .Y(n2939) );
  OAI21X1 U2318 ( .A(n5601), .B(n5636), .C(n358), .Y(n2940) );
  OAI21X1 U2320 ( .A(n5601), .B(n5635), .C(n286), .Y(n2941) );
  OAI21X1 U2322 ( .A(n5601), .B(n5634), .C(n3914), .Y(n2942) );
  OAI21X1 U2324 ( .A(n5601), .B(n5633), .C(n3821), .Y(n2943) );
  OAI21X1 U2326 ( .A(n5601), .B(n5632), .C(n4098), .Y(n2944) );
  OAI21X1 U2328 ( .A(n5601), .B(n5631), .C(n3245), .Y(n2945) );
  OAI21X1 U2330 ( .A(n5601), .B(n5630), .C(n3173), .Y(n2946) );
  OAI21X1 U2332 ( .A(n5601), .B(n5629), .C(n3389), .Y(n2947) );
  OAI21X1 U2334 ( .A(n5601), .B(n5628), .C(n214), .Y(n2948) );
  OAI21X1 U2336 ( .A(n3624), .B(n3992), .C(reset), .Y(n1566) );
  NAND3X1 U2337 ( .A(n5716), .B(n5719), .C(wr_ptr[1]), .Y(n550) );
  OAI21X1 U2338 ( .A(n5600), .B(n5668), .C(n3457), .Y(n2949) );
  OAI21X1 U2340 ( .A(n5600), .B(n5667), .C(n3546), .Y(n2950) );
  OAI21X1 U2342 ( .A(n5600), .B(n5666), .C(n3636), .Y(n2951) );
  OAI21X1 U2344 ( .A(n5600), .B(n5665), .C(n3725), .Y(n2952) );
  OAI21X1 U2346 ( .A(n5600), .B(n5664), .C(n3456), .Y(n2953) );
  OAI21X1 U2348 ( .A(n5600), .B(n5663), .C(n3820), .Y(n2954) );
  OAI21X1 U2350 ( .A(n5600), .B(n5662), .C(n3913), .Y(n2955) );
  OAI21X1 U2352 ( .A(n5600), .B(n5661), .C(n4005), .Y(n2956) );
  OAI21X1 U2354 ( .A(n5600), .B(n5660), .C(n4097), .Y(n2957) );
  OAI21X1 U2356 ( .A(n5600), .B(n5659), .C(n142), .Y(n2958) );
  OAI21X1 U2358 ( .A(n5600), .B(n5658), .C(n3545), .Y(n2959) );
  OAI21X1 U2360 ( .A(n5600), .B(n5657), .C(n3635), .Y(n2960) );
  OAI21X1 U2362 ( .A(n5600), .B(n5656), .C(n3724), .Y(n2961) );
  OAI21X1 U2364 ( .A(n5600), .B(n5655), .C(n4096), .Y(n2962) );
  OAI21X1 U2366 ( .A(n5600), .B(n5654), .C(n213), .Y(n2963) );
  OAI21X1 U2368 ( .A(n5600), .B(n5653), .C(n285), .Y(n2964) );
  OAI21X1 U2370 ( .A(n5600), .B(n5652), .C(n357), .Y(n2965) );
  OAI21X1 U2372 ( .A(n5600), .B(n5651), .C(n3172), .Y(n2966) );
  OAI21X1 U2374 ( .A(n5600), .B(n5650), .C(n3244), .Y(n2967) );
  OAI21X1 U2376 ( .A(n5600), .B(n5649), .C(n3819), .Y(n2968) );
  OAI21X1 U2378 ( .A(n5600), .B(n5648), .C(n3912), .Y(n2969) );
  OAI21X1 U2380 ( .A(n5600), .B(n5647), .C(n4004), .Y(n2970) );
  OAI21X1 U2382 ( .A(n5600), .B(n5646), .C(n3316), .Y(n2971) );
  OAI21X1 U2384 ( .A(n5600), .B(n5645), .C(n3388), .Y(n2972) );
  OAI21X1 U2386 ( .A(n5600), .B(n5644), .C(n55), .Y(n2973) );
  OAI21X1 U2388 ( .A(n5600), .B(n5643), .C(n3455), .Y(n2974) );
  OAI21X1 U2390 ( .A(n5600), .B(n5642), .C(n4095), .Y(n2975) );
  OAI21X1 U2392 ( .A(n5600), .B(n5641), .C(n3544), .Y(n2976) );
  OAI21X1 U2394 ( .A(n5600), .B(n5640), .C(n3634), .Y(n2977) );
  OAI21X1 U2396 ( .A(n5600), .B(n5639), .C(n3723), .Y(n2978) );
  OAI21X1 U2398 ( .A(n5600), .B(n5638), .C(n141), .Y(n2979) );
  OAI21X1 U2400 ( .A(n5600), .B(n5637), .C(n212), .Y(n2980) );
  OAI21X1 U2402 ( .A(n5600), .B(n5636), .C(n284), .Y(n2981) );
  OAI21X1 U2404 ( .A(n5600), .B(n5635), .C(n356), .Y(n2982) );
  OAI21X1 U2406 ( .A(n5600), .B(n5634), .C(n3818), .Y(n2983) );
  OAI21X1 U2408 ( .A(n5600), .B(n5633), .C(n3911), .Y(n2984) );
  OAI21X1 U2410 ( .A(n5600), .B(n5632), .C(n4003), .Y(n2985) );
  OAI21X1 U2412 ( .A(n5600), .B(n5631), .C(n3171), .Y(n2986) );
  OAI21X1 U2414 ( .A(n5600), .B(n5630), .C(n3243), .Y(n2987) );
  OAI21X1 U2416 ( .A(n5600), .B(n5629), .C(n3315), .Y(n2988) );
  OAI21X1 U2418 ( .A(n5600), .B(n5628), .C(n140), .Y(n2989) );
  OAI21X1 U2420 ( .A(n3535), .B(n3992), .C(reset), .Y(n1608) );
  NAND3X1 U2421 ( .A(wr_ptr[0]), .B(n5719), .C(wr_ptr[1]), .Y(n593) );
  OAI21X1 U2422 ( .A(n5599), .B(n5668), .C(n3387), .Y(n2990) );
  OAI21X1 U2424 ( .A(n5599), .B(n5667), .C(n3314), .Y(n2991) );
  OAI21X1 U2426 ( .A(n5599), .B(n5666), .C(n3242), .Y(n2992) );
  OAI21X1 U2428 ( .A(n5599), .B(n5665), .C(n3170), .Y(n2993) );
  OAI21X1 U2430 ( .A(n5599), .B(n5664), .C(n3386), .Y(n2994) );
  OAI21X1 U2432 ( .A(n5599), .B(n5663), .C(n355), .Y(n2995) );
  OAI21X1 U2434 ( .A(n5599), .B(n5662), .C(n283), .Y(n2996) );
  OAI21X1 U2436 ( .A(n5599), .B(n5661), .C(n211), .Y(n2997) );
  OAI21X1 U2438 ( .A(n5599), .B(n5660), .C(n139), .Y(n2998) );
  OAI21X1 U2440 ( .A(n5599), .B(n5659), .C(n4094), .Y(n2999) );
  OAI21X1 U2442 ( .A(n5599), .B(n5658), .C(n3313), .Y(n3000) );
  OAI21X1 U2444 ( .A(n5599), .B(n5657), .C(n3241), .Y(n3001) );
  OAI21X1 U2446 ( .A(n5599), .B(n5656), .C(n3169), .Y(n3002) );
  OAI21X1 U2448 ( .A(n5599), .B(n5655), .C(n138), .Y(n3003) );
  OAI21X1 U2450 ( .A(n5599), .B(n5654), .C(n4002), .Y(n3004) );
  OAI21X1 U2452 ( .A(n5599), .B(n5653), .C(n3910), .Y(n3005) );
  OAI21X1 U2454 ( .A(n5599), .B(n5652), .C(n3817), .Y(n3006) );
  OAI21X1 U2456 ( .A(n5599), .B(n5651), .C(n3722), .Y(n3007) );
  OAI21X1 U2458 ( .A(n5599), .B(n5650), .C(n3633), .Y(n3008) );
  OAI21X1 U2460 ( .A(n5599), .B(n5649), .C(n354), .Y(n3009) );
  OAI21X1 U2462 ( .A(n5599), .B(n5648), .C(n282), .Y(n3010) );
  OAI21X1 U2464 ( .A(n5599), .B(n5647), .C(n210), .Y(n3011) );
  OAI21X1 U2466 ( .A(n5599), .B(n5646), .C(n3543), .Y(n3012) );
  OAI21X1 U2468 ( .A(n5599), .B(n5645), .C(n3454), .Y(n3013) );
  OAI21X1 U2470 ( .A(n5599), .B(n5644), .C(n54), .Y(n3014) );
  OAI21X1 U2472 ( .A(n5599), .B(n5643), .C(n3385), .Y(n3015) );
  OAI21X1 U2474 ( .A(n5599), .B(n5642), .C(n137), .Y(n3016) );
  OAI21X1 U2476 ( .A(n5599), .B(n5641), .C(n3312), .Y(n3017) );
  OAI21X1 U2478 ( .A(n5599), .B(n5640), .C(n3240), .Y(n3018) );
  OAI21X1 U2480 ( .A(n5599), .B(n5639), .C(n3168), .Y(n3019) );
  OAI21X1 U2482 ( .A(n5599), .B(n5638), .C(n4093), .Y(n3020) );
  OAI21X1 U2484 ( .A(n5599), .B(n5637), .C(n4001), .Y(n3021) );
  OAI21X1 U2486 ( .A(n5599), .B(n5636), .C(n3909), .Y(n3022) );
  OAI21X1 U2488 ( .A(n5599), .B(n5635), .C(n3816), .Y(n3023) );
  OAI21X1 U2490 ( .A(n5599), .B(n5634), .C(n353), .Y(n3024) );
  OAI21X1 U2492 ( .A(n5599), .B(n5633), .C(n281), .Y(n3025) );
  OAI21X1 U2494 ( .A(n5599), .B(n5632), .C(n209), .Y(n3026) );
  OAI21X1 U2496 ( .A(n5599), .B(n5631), .C(n3721), .Y(n3027) );
  OAI21X1 U2498 ( .A(n5599), .B(n5630), .C(n3632), .Y(n3028) );
  OAI21X1 U2500 ( .A(n5599), .B(n5629), .C(n3542), .Y(n3029) );
  OAI21X1 U2502 ( .A(n5599), .B(n5628), .C(n4092), .Y(n3030) );
  OAI21X1 U2504 ( .A(n3534), .B(n3992), .C(reset), .Y(n1650) );
  NAND3X1 U2505 ( .A(n5716), .B(n5718), .C(wr_ptr[2]), .Y(n636) );
  OAI21X1 U2506 ( .A(n5598), .B(n5668), .C(n3311), .Y(n3031) );
  OAI21X1 U2508 ( .A(n5598), .B(n5667), .C(n3384), .Y(n3032) );
  OAI21X1 U2510 ( .A(n5598), .B(n5666), .C(n3167), .Y(n3033) );
  OAI21X1 U2512 ( .A(n5598), .B(n5665), .C(n3239), .Y(n3034) );
  OAI21X1 U2514 ( .A(n5598), .B(n5664), .C(n3310), .Y(n3035) );
  OAI21X1 U2516 ( .A(n5598), .B(n5663), .C(n280), .Y(n3036) );
  OAI21X1 U2518 ( .A(n5598), .B(n5662), .C(n352), .Y(n3037) );
  OAI21X1 U2520 ( .A(n5598), .B(n5661), .C(n136), .Y(n3038) );
  OAI21X1 U2522 ( .A(n5598), .B(n5660), .C(n208), .Y(n3039) );
  OAI21X1 U2524 ( .A(n5598), .B(n5659), .C(n4000), .Y(n3040) );
  OAI21X1 U2526 ( .A(n5598), .B(n5658), .C(n3383), .Y(n3041) );
  OAI21X1 U2528 ( .A(n5598), .B(n5657), .C(n3166), .Y(n3042) );
  OAI21X1 U2530 ( .A(n5598), .B(n5656), .C(n3238), .Y(n3043) );
  OAI21X1 U2532 ( .A(n5598), .B(n5655), .C(n207), .Y(n3044) );
  OAI21X1 U2534 ( .A(n5598), .B(n5654), .C(n4091), .Y(n3045) );
  OAI21X1 U2536 ( .A(n5598), .B(n5653), .C(n3815), .Y(n3046) );
  OAI21X1 U2538 ( .A(n5598), .B(n5652), .C(n3908), .Y(n3047) );
  OAI21X1 U2540 ( .A(n5598), .B(n5651), .C(n3631), .Y(n3048) );
  OAI21X1 U2542 ( .A(n5598), .B(n5650), .C(n3720), .Y(n3049) );
  OAI21X1 U2544 ( .A(n5598), .B(n5649), .C(n279), .Y(n3050) );
  OAI21X1 U2546 ( .A(n5598), .B(n5648), .C(n351), .Y(n3051) );
  OAI21X1 U2548 ( .A(n5598), .B(n5647), .C(n135), .Y(n3052) );
  OAI21X1 U2550 ( .A(n5598), .B(n5646), .C(n3453), .Y(n3053) );
  OAI21X1 U2552 ( .A(n5598), .B(n5645), .C(n3541), .Y(n3054) );
  OAI21X1 U2554 ( .A(n5598), .B(n5644), .C(n53), .Y(n3055) );
  OAI21X1 U2556 ( .A(n5598), .B(n5643), .C(n3309), .Y(n3056) );
  OAI21X1 U2558 ( .A(n5598), .B(n5642), .C(n206), .Y(n3057) );
  OAI21X1 U2560 ( .A(n5598), .B(n5641), .C(n3382), .Y(n3058) );
  OAI21X1 U2562 ( .A(n5598), .B(n5640), .C(n3165), .Y(n3059) );
  OAI21X1 U2564 ( .A(n5598), .B(n5639), .C(n3237), .Y(n3060) );
  OAI21X1 U2566 ( .A(n5598), .B(n5638), .C(n3999), .Y(n3061) );
  OAI21X1 U2568 ( .A(n5598), .B(n5637), .C(n4090), .Y(n3062) );
  OAI21X1 U2570 ( .A(n5598), .B(n5636), .C(n3814), .Y(n3063) );
  OAI21X1 U2572 ( .A(n5598), .B(n5635), .C(n3907), .Y(n3064) );
  OAI21X1 U2574 ( .A(n5598), .B(n5634), .C(n278), .Y(n3065) );
  OAI21X1 U2576 ( .A(n5598), .B(n5633), .C(n350), .Y(n3066) );
  OAI21X1 U2578 ( .A(n5598), .B(n5632), .C(n134), .Y(n3067) );
  OAI21X1 U2580 ( .A(n5598), .B(n5631), .C(n3630), .Y(n3068) );
  OAI21X1 U2582 ( .A(n5598), .B(n5630), .C(n3719), .Y(n3069) );
  OAI21X1 U2584 ( .A(n5598), .B(n5629), .C(n3452), .Y(n3070) );
  OAI21X1 U2586 ( .A(n5598), .B(n5628), .C(n3998), .Y(n3071) );
  OAI21X1 U2588 ( .A(n3623), .B(n3992), .C(reset), .Y(n1692) );
  NAND3X1 U2589 ( .A(wr_ptr[0]), .B(n5718), .C(wr_ptr[2]), .Y(n679) );
  OAI21X1 U2590 ( .A(n5597), .B(n5668), .C(n3236), .Y(n3072) );
  OAI21X1 U2592 ( .A(n5597), .B(n5667), .C(n3164), .Y(n3073) );
  OAI21X1 U2594 ( .A(n5597), .B(n5666), .C(n3381), .Y(n3074) );
  OAI21X1 U2596 ( .A(n5597), .B(n5665), .C(n3308), .Y(n3075) );
  OAI21X1 U2598 ( .A(n5597), .B(n5664), .C(n3235), .Y(n3076) );
  OAI21X1 U2600 ( .A(n5597), .B(n5663), .C(n205), .Y(n3077) );
  OAI21X1 U2602 ( .A(n5597), .B(n5662), .C(n133), .Y(n3078) );
  OAI21X1 U2604 ( .A(n5597), .B(n5661), .C(n349), .Y(n3079) );
  OAI21X1 U2606 ( .A(n5597), .B(n5660), .C(n277), .Y(n3080) );
  OAI21X1 U2608 ( .A(n5597), .B(n5659), .C(n3906), .Y(n3081) );
  OAI21X1 U2610 ( .A(n5597), .B(n5658), .C(n460), .Y(n3082) );
  OAI21X1 U2612 ( .A(n5597), .B(n5657), .C(n3380), .Y(n3083) );
  OAI21X1 U2614 ( .A(n5597), .B(n5656), .C(n3307), .Y(n3084) );
  OAI21X1 U2616 ( .A(n5597), .B(n5655), .C(n276), .Y(n3085) );
  OAI21X1 U2618 ( .A(n5597), .B(n5654), .C(n3813), .Y(n3086) );
  OAI21X1 U2620 ( .A(n5597), .B(n5653), .C(n4089), .Y(n3087) );
  OAI21X1 U2622 ( .A(n5597), .B(n5652), .C(n3997), .Y(n3088) );
  OAI21X1 U2624 ( .A(n5597), .B(n5651), .C(n3540), .Y(n3089) );
  OAI21X1 U2626 ( .A(n5597), .B(n5650), .C(n3451), .Y(n3090) );
  OAI21X1 U2628 ( .A(n5597), .B(n5649), .C(n204), .Y(n3091) );
  OAI21X1 U2630 ( .A(n5597), .B(n5648), .C(n132), .Y(n3092) );
  OAI21X1 U2632 ( .A(n5597), .B(n5647), .C(n348), .Y(n3093) );
  OAI21X1 U2634 ( .A(n5597), .B(n5646), .C(n3718), .Y(n3094) );
  OAI21X1 U2636 ( .A(n5597), .B(n5645), .C(n3629), .Y(n3095) );
  OAI21X1 U2638 ( .A(n5597), .B(n5644), .C(n52), .Y(n3096) );
  OAI21X1 U2640 ( .A(n5597), .B(n5643), .C(n3234), .Y(n3097) );
  OAI21X1 U2642 ( .A(n5597), .B(n5642), .C(n275), .Y(n3098) );
  OAI21X1 U2644 ( .A(n5597), .B(n5641), .C(n458), .Y(n3099) );
  OAI21X1 U2646 ( .A(n5597), .B(n5640), .C(n3379), .Y(n3100) );
  OAI21X1 U2648 ( .A(n5597), .B(n5639), .C(n3306), .Y(n3101) );
  OAI21X1 U2650 ( .A(n5597), .B(n5638), .C(n3905), .Y(n3102) );
  OAI21X1 U2652 ( .A(n5597), .B(n5637), .C(n3812), .Y(n3103) );
  OAI21X1 U2654 ( .A(n5597), .B(n5636), .C(n4088), .Y(n3104) );
  OAI21X1 U2656 ( .A(n5597), .B(n5635), .C(n3996), .Y(n3105) );
  OAI21X1 U2658 ( .A(n5597), .B(n5634), .C(n203), .Y(n3106) );
  OAI21X1 U2660 ( .A(n5597), .B(n5633), .C(n131), .Y(n3107) );
  OAI21X1 U2662 ( .A(n5597), .B(n5632), .C(n347), .Y(n3108) );
  OAI21X1 U2664 ( .A(n5597), .B(n5631), .C(n3539), .Y(n3109) );
  OAI21X1 U2666 ( .A(n5597), .B(n5630), .C(n3450), .Y(n3110) );
  OAI21X1 U2668 ( .A(n5597), .B(n5629), .C(n3717), .Y(n3111) );
  OAI21X1 U2670 ( .A(n5597), .B(n5628), .C(n3904), .Y(n3112) );
  OAI21X1 U2672 ( .A(n3713), .B(n3992), .C(reset), .Y(n1734) );
  NAND3X1 U2673 ( .A(wr_ptr[1]), .B(n5716), .C(wr_ptr[2]), .Y(n722) );
  OAI21X1 U2674 ( .A(n5596), .B(n5668), .C(n456), .Y(n3113) );
  OAI21X1 U2677 ( .A(n5596), .B(n5667), .C(n3233), .Y(n3114) );
  OAI21X1 U2680 ( .A(n5596), .B(n5666), .C(n3305), .Y(n3115) );
  OAI21X1 U2683 ( .A(n5596), .B(n5665), .C(n3378), .Y(n3116) );
  OAI21X1 U2686 ( .A(n5596), .B(n5664), .C(n454), .Y(n3117) );
  OAI21X1 U2689 ( .A(n5596), .B(n5663), .C(n130), .Y(n3118) );
  OAI21X1 U2692 ( .A(n5596), .B(n5662), .C(n202), .Y(n3119) );
  OAI21X1 U2695 ( .A(n5596), .B(n5661), .C(n274), .Y(n3120) );
  OAI21X1 U2698 ( .A(n5596), .B(n5660), .C(n346), .Y(n3121) );
  OAI21X1 U2701 ( .A(n5596), .B(n5659), .C(n3811), .Y(n3122) );
  OAI21X1 U2704 ( .A(n5596), .B(n5658), .C(n3232), .Y(n3123) );
  OAI21X1 U2707 ( .A(n5596), .B(n5657), .C(n3304), .Y(n3124) );
  OAI21X1 U2710 ( .A(n5596), .B(n5656), .C(n3377), .Y(n3125) );
  OAI21X1 U2713 ( .A(n5596), .B(n5655), .C(n345), .Y(n3126) );
  OAI21X1 U2716 ( .A(n5596), .B(n5654), .C(n3903), .Y(n3127) );
  OAI21X1 U2719 ( .A(n5596), .B(n5653), .C(n3995), .Y(n3128) );
  OAI21X1 U2722 ( .A(n5596), .B(n5652), .C(n4087), .Y(n3129) );
  OAI21X1 U2725 ( .A(n5596), .B(n5651), .C(n3449), .Y(n3130) );
  OAI21X1 U2728 ( .A(n5596), .B(n5650), .C(n3538), .Y(n3131) );
  OAI21X1 U2731 ( .A(n5596), .B(n5649), .C(n129), .Y(n3132) );
  OAI21X1 U2734 ( .A(n5596), .B(n5648), .C(n201), .Y(n3133) );
  OAI21X1 U2737 ( .A(n5596), .B(n5647), .C(n273), .Y(n3134) );
  OAI21X1 U2740 ( .A(n5596), .B(n5646), .C(n3628), .Y(n3135) );
  OAI21X1 U2743 ( .A(n5596), .B(n5645), .C(n3716), .Y(n3136) );
  OAI21X1 U2746 ( .A(n5596), .B(n5644), .C(n51), .Y(n3137) );
  OAI21X1 U2749 ( .A(n5596), .B(n5643), .C(n452), .Y(n3138) );
  OAI21X1 U2752 ( .A(n5596), .B(n5642), .C(n344), .Y(n3139) );
  OAI21X1 U2755 ( .A(n5596), .B(n5641), .C(n3231), .Y(n3140) );
  OAI21X1 U2758 ( .A(n5596), .B(n5640), .C(n3303), .Y(n3141) );
  OAI21X1 U2761 ( .A(n5596), .B(n5639), .C(n3376), .Y(n3142) );
  OAI21X1 U2764 ( .A(n5596), .B(n5638), .C(n3810), .Y(n3143) );
  OAI21X1 U2767 ( .A(n5596), .B(n5637), .C(n3902), .Y(n3144) );
  OAI21X1 U2770 ( .A(n5596), .B(n5636), .C(n3994), .Y(n3145) );
  OAI21X1 U2773 ( .A(n5596), .B(n5635), .C(n4086), .Y(n3146) );
  OAI21X1 U2776 ( .A(n5596), .B(n5634), .C(n128), .Y(n3147) );
  OAI21X1 U2779 ( .A(n5596), .B(n5633), .C(n200), .Y(n3148) );
  OAI21X1 U2782 ( .A(n5596), .B(n5632), .C(n272), .Y(n3149) );
  OAI21X1 U2785 ( .A(n5596), .B(n5631), .C(n3448), .Y(n3150) );
  OAI21X1 U2788 ( .A(n5596), .B(n5630), .C(n3537), .Y(n3151) );
  OAI21X1 U2791 ( .A(n5596), .B(n5629), .C(n3627), .Y(n3152) );
  OAI21X1 U2794 ( .A(n5596), .B(n5628), .C(n3809), .Y(n3153) );
  OAI21X1 U2797 ( .A(n3805), .B(n3992), .C(reset), .Y(n1776) );
  NAND3X1 U2798 ( .A(wr_ptr[3]), .B(n1777), .C(wr_ptr[4]), .Y(n1482) );
  NAND3X1 U2799 ( .A(wr_ptr[1]), .B(wr_ptr[0]), .C(wr_ptr[2]), .Y(n765) );
  OAI21X1 U2800 ( .A(n5720), .B(n4084), .C(n3626), .Y(n3154) );
  OAI21X1 U2802 ( .A(n5719), .B(n4084), .C(n3901), .Y(n3155) );
  OAI21X1 U2804 ( .A(n5718), .B(n4084), .C(n3808), .Y(n3156) );
  OAI21X1 U2806 ( .A(n5717), .B(n4084), .C(n3536), .Y(n3157) );
  OAI21X1 U2808 ( .A(n5670), .B(n4176), .C(n3993), .Y(n3158) );
  OAI21X1 U2810 ( .A(n5671), .B(n4176), .C(n3900), .Y(n3159) );
  OAI21X1 U2812 ( .A(n5672), .B(n4176), .C(n3807), .Y(n3160) );
  OAI21X1 U2814 ( .A(n5674), .B(n4176), .C(n3715), .Y(n3161) );
  OAI21X1 U2816 ( .A(n5669), .B(n4176), .C(n3625), .Y(n3162) );
  AOI22X1 U2818 ( .A(n56), .B(n1786), .C(data_out[40]), .D(n1784), .Y(n1791)
         );
  AOI22X1 U2819 ( .A(n57), .B(n1786), .C(data_out[39]), .D(n1784), .Y(n1792)
         );
  AOI22X1 U2820 ( .A(n58), .B(n1786), .C(data_out[38]), .D(n1784), .Y(n1793)
         );
  AOI22X1 U2821 ( .A(n59), .B(n1786), .C(data_out[37]), .D(n1784), .Y(n1794)
         );
  AOI22X1 U2822 ( .A(n60), .B(n1786), .C(data_out[36]), .D(n1784), .Y(n1795)
         );
  AOI22X1 U2823 ( .A(n61), .B(n1786), .C(data_out[35]), .D(n1784), .Y(n1796)
         );
  AOI22X1 U2824 ( .A(n62), .B(n1786), .C(data_out[34]), .D(n1784), .Y(n1797)
         );
  AOI22X1 U2825 ( .A(n63), .B(n1786), .C(data_out[33]), .D(n1784), .Y(n1798)
         );
  AOI22X1 U2826 ( .A(n64), .B(n1786), .C(data_out[32]), .D(n1784), .Y(n1799)
         );
  AOI22X1 U2827 ( .A(n65), .B(n1786), .C(data_out[31]), .D(n1784), .Y(n1800)
         );
  AOI22X1 U2828 ( .A(n66), .B(n1786), .C(data_out[30]), .D(n1784), .Y(n1801)
         );
  AOI22X1 U2829 ( .A(n67), .B(n1786), .C(data_out[29]), .D(n1784), .Y(n1802)
         );
  AOI22X1 U2830 ( .A(n68), .B(n1786), .C(data_out[28]), .D(n1784), .Y(n1803)
         );
  AOI22X1 U2831 ( .A(n69), .B(n1786), .C(data_out[27]), .D(n1784), .Y(n1804)
         );
  AOI22X1 U2832 ( .A(n70), .B(n1786), .C(data_out[26]), .D(n1784), .Y(n1805)
         );
  AOI22X1 U2833 ( .A(n71), .B(n1786), .C(data_out[25]), .D(n1784), .Y(n1806)
         );
  AOI22X1 U2834 ( .A(n72), .B(n1786), .C(data_out[24]), .D(n1784), .Y(n1807)
         );
  AOI22X1 U2835 ( .A(n73), .B(n1786), .C(data_out[23]), .D(n1784), .Y(n1808)
         );
  AOI22X1 U2836 ( .A(n74), .B(n1786), .C(data_out[22]), .D(n1784), .Y(n1809)
         );
  AOI22X1 U2837 ( .A(n75), .B(n1786), .C(data_out[21]), .D(n1784), .Y(n1810)
         );
  AOI22X1 U2838 ( .A(n76), .B(n1786), .C(data_out[20]), .D(n1784), .Y(n1811)
         );
  AOI22X1 U2839 ( .A(n77), .B(n1786), .C(data_out[19]), .D(n1784), .Y(n1812)
         );
  AOI22X1 U2840 ( .A(n78), .B(n1786), .C(data_out[18]), .D(n1784), .Y(n1813)
         );
  AOI22X1 U2841 ( .A(n79), .B(n1786), .C(data_out[17]), .D(n1784), .Y(n1814)
         );
  AOI22X1 U2842 ( .A(n80), .B(n1786), .C(data_out[16]), .D(n1784), .Y(n1815)
         );
  AOI22X1 U2843 ( .A(n81), .B(n1786), .C(data_out[15]), .D(n1784), .Y(n1816)
         );
  AOI22X1 U2844 ( .A(n82), .B(n1786), .C(data_out[14]), .D(n1784), .Y(n1817)
         );
  AOI22X1 U2845 ( .A(n83), .B(n1786), .C(data_out[13]), .D(n1784), .Y(n1818)
         );
  AOI22X1 U2846 ( .A(n84), .B(n1786), .C(data_out[12]), .D(n1784), .Y(n1819)
         );
  AOI22X1 U2847 ( .A(n85), .B(n1786), .C(data_out[11]), .D(n1784), .Y(n1820)
         );
  AOI22X1 U2848 ( .A(n86), .B(n1786), .C(data_out[10]), .D(n1784), .Y(n1821)
         );
  AOI22X1 U2849 ( .A(n87), .B(n1786), .C(data_out[9]), .D(n1784), .Y(n1822) );
  AOI22X1 U2850 ( .A(n88), .B(n1786), .C(data_out[8]), .D(n1784), .Y(n1823) );
  AOI22X1 U2851 ( .A(n89), .B(n1786), .C(data_out[7]), .D(n1784), .Y(n1824) );
  AOI22X1 U2852 ( .A(n90), .B(n1786), .C(data_out[6]), .D(n1784), .Y(n1825) );
  AOI22X1 U2853 ( .A(n91), .B(n1786), .C(data_out[5]), .D(n1784), .Y(n1826) );
  AOI22X1 U2854 ( .A(n92), .B(n1786), .C(data_out[4]), .D(n1784), .Y(n1827) );
  AOI22X1 U2855 ( .A(n93), .B(n1786), .C(data_out[3]), .D(n1784), .Y(n1828) );
  AOI22X1 U2856 ( .A(n94), .B(n1786), .C(data_out[2]), .D(n1784), .Y(n1829) );
  AOI22X1 U2857 ( .A(n95), .B(n1786), .C(data_out[1]), .D(n1784), .Y(n1830) );
  AOI22X1 U2858 ( .A(n96), .B(n1786), .C(data_out[0]), .D(n1784), .Y(n1831) );
  OAI21X1 U2861 ( .A(n5716), .B(n4084), .C(n3375), .Y(n3163) );
  NAND3X1 U2865 ( .A(n3804), .B(fillcount[5]), .C(n1835), .Y(n5722) );
  NOR3X1 U2866 ( .A(fillcount[2]), .B(fillcount[4]), .C(fillcount[3]), .Y(
        n1835) );
  NAND3X1 U2868 ( .A(n1836), .B(n1837), .C(n1838), .Y(n5721) );
  NOR3X1 U2869 ( .A(n1839), .B(n1840), .C(n1841), .Y(n1838) );
  XNOR2X1 U2870 ( .A(n5719), .B(n14), .Y(n1841) );
  XNOR2X1 U2871 ( .A(n5720), .B(n15), .Y(n1840) );
  XNOR2X1 U2872 ( .A(n5716), .B(n5673), .Y(n1839) );
  XNOR2X1 U2873 ( .A(n5572), .B(wr_ptr[1]), .Y(n1837) );
  XNOR2X1 U2874 ( .A(n16), .B(wr_ptr[4]), .Y(n1836) );
  HAX1 add_57_U1_1_1 ( .A(n5573), .B(n5673), .YC(add_57_carry[2]), .YS(n98) );
  HAX1 add_57_U1_1_2 ( .A(n14), .B(add_57_carry[2]), .YC(add_57_carry[3]), 
        .YS(n99) );
  HAX1 add_57_U1_1_3 ( .A(n15), .B(add_57_carry[3]), .YC(add_57_carry[4]), 
        .YS(n100) );
  HAX1 add_51_U1_1_1 ( .A(wr_ptr[1]), .B(wr_ptr[0]), .YC(add_51_carry[2]), 
        .YS(n20) );
  HAX1 add_51_U1_1_2 ( .A(wr_ptr[2]), .B(add_51_carry[2]), .YC(add_51_carry[3]), .YS(n21) );
  HAX1 add_51_U1_1_3 ( .A(wr_ptr[3]), .B(add_51_carry[3]), .YC(add_51_carry[4]), .YS(n22) );
  FAX1 sub_93_U2_1 ( .A(wr_ptr[1]), .B(n5672), .C(sub_93_carry[1]), .YC(
        sub_93_carry[2]), .YS(fillcount[1]) );
  FAX1 sub_93_U2_2 ( .A(wr_ptr[2]), .B(n5671), .C(sub_93_carry[2]), .YC(
        sub_93_carry[3]), .YS(fillcount[2]) );
  FAX1 sub_93_U2_3 ( .A(wr_ptr[3]), .B(n5670), .C(sub_93_carry[3]), .YC(
        sub_93_carry[4]), .YS(fillcount[3]) );
  FAX1 sub_93_U2_4 ( .A(wr_ptr[4]), .B(n5669), .C(sub_93_carry[4]), .YC(
        sub_93_carry[5]), .YS(fillcount[4]) );
  AND2X1 U3 ( .A(get), .B(empty_bar), .Y(n1832) );
  AND2X1 U4 ( .A(reset), .B(n3802), .Y(n1778) );
  AND2X1 U5 ( .A(reset), .B(n4177), .Y(n1784) );
  AND2X1 U6 ( .A(reset), .B(n4176), .Y(n1786) );
  AND2X1 U7 ( .A(put), .B(full_bar), .Y(n1777) );
  BUFX2 U8 ( .A(n1831), .Y(n1) );
  BUFX2 U9 ( .A(n1830), .Y(n2) );
  BUFX2 U10 ( .A(n1829), .Y(n3) );
  BUFX2 U11 ( .A(n1828), .Y(n4) );
  BUFX2 U12 ( .A(n1827), .Y(n5) );
  BUFX2 U13 ( .A(n1826), .Y(n6) );
  BUFX2 U14 ( .A(n1825), .Y(n7) );
  BUFX2 U15 ( .A(n1824), .Y(n8) );
  BUFX2 U16 ( .A(n1823), .Y(n9) );
  BUFX2 U17 ( .A(n1822), .Y(n10) );
  BUFX2 U18 ( .A(n1821), .Y(n11) );
  BUFX2 U19 ( .A(n1820), .Y(n17) );
  BUFX2 U20 ( .A(n1819), .Y(n18) );
  BUFX2 U21 ( .A(n1818), .Y(n19) );
  BUFX2 U22 ( .A(n1817), .Y(n24) );
  BUFX2 U23 ( .A(n1816), .Y(n25) );
  BUFX2 U24 ( .A(n1815), .Y(n26) );
  BUFX2 U25 ( .A(n1814), .Y(n27) );
  BUFX2 U26 ( .A(n1813), .Y(n28) );
  BUFX2 U27 ( .A(n1812), .Y(n29) );
  BUFX2 U28 ( .A(n1811), .Y(n30) );
  BUFX2 U29 ( .A(n1810), .Y(n31) );
  BUFX2 U30 ( .A(n1809), .Y(n32) );
  BUFX2 U31 ( .A(n1808), .Y(n33) );
  BUFX2 U32 ( .A(n1807), .Y(n34) );
  BUFX2 U33 ( .A(n1806), .Y(n35) );
  BUFX2 U34 ( .A(n1805), .Y(n36) );
  BUFX2 U35 ( .A(n1804), .Y(n37) );
  BUFX2 U36 ( .A(n1803), .Y(n38) );
  BUFX2 U37 ( .A(n1802), .Y(n39) );
  BUFX2 U38 ( .A(n1801), .Y(n40) );
  BUFX2 U39 ( .A(n1800), .Y(n41) );
  BUFX2 U40 ( .A(n1799), .Y(n42) );
  BUFX2 U41 ( .A(n1798), .Y(n43) );
  BUFX2 U42 ( .A(n1797), .Y(n44) );
  BUFX2 U43 ( .A(n1796), .Y(n45) );
  BUFX2 U44 ( .A(n1795), .Y(n46) );
  BUFX2 U45 ( .A(n1794), .Y(n47) );
  BUFX2 U46 ( .A(n1793), .Y(n48) );
  BUFX2 U47 ( .A(n1792), .Y(n49) );
  BUFX2 U48 ( .A(n1791), .Y(n50) );
  AND2X1 U49 ( .A(mem[1295]), .B(n5596), .Y(n1759) );
  INVX1 U50 ( .A(n1759), .Y(n51) );
  AND2X1 U51 ( .A(mem[1254]), .B(n5597), .Y(n1717) );
  INVX1 U52 ( .A(n1717), .Y(n52) );
  AND2X1 U53 ( .A(mem[1213]), .B(n5598), .Y(n1675) );
  INVX1 U54 ( .A(n1675), .Y(n53) );
  AND2X1 U55 ( .A(mem[1172]), .B(n5599), .Y(n1633) );
  INVX1 U56 ( .A(n1633), .Y(n54) );
  AND2X1 U57 ( .A(mem[1131]), .B(n5600), .Y(n1591) );
  INVX1 U58 ( .A(n1591), .Y(n55) );
  AND2X1 U59 ( .A(mem[1090]), .B(n5601), .Y(n1549) );
  INVX1 U60 ( .A(n1549), .Y(n97) );
  AND2X1 U61 ( .A(mem[1049]), .B(n5602), .Y(n1507) );
  INVX1 U62 ( .A(n1507), .Y(n102) );
  AND2X1 U63 ( .A(mem[1008]), .B(n5603), .Y(n1464) );
  INVX1 U64 ( .A(n1464), .Y(n103) );
  AND2X1 U65 ( .A(mem[967]), .B(n5604), .Y(n1422) );
  INVX1 U66 ( .A(n1422), .Y(n104) );
  AND2X1 U67 ( .A(mem[926]), .B(n5605), .Y(n1380) );
  INVX1 U68 ( .A(n1380), .Y(n105) );
  AND2X1 U69 ( .A(mem[885]), .B(n5606), .Y(n1338) );
  INVX1 U70 ( .A(n1338), .Y(n106) );
  AND2X1 U71 ( .A(mem[844]), .B(n5607), .Y(n1296) );
  INVX1 U72 ( .A(n1296), .Y(n107) );
  AND2X1 U73 ( .A(mem[803]), .B(n5608), .Y(n1254) );
  INVX1 U74 ( .A(n1254), .Y(n108) );
  AND2X1 U75 ( .A(mem[762]), .B(n5609), .Y(n1212) );
  INVX1 U76 ( .A(n1212), .Y(n109) );
  AND2X1 U77 ( .A(mem[721]), .B(n5610), .Y(n1170) );
  INVX1 U78 ( .A(n1170), .Y(n110) );
  AND2X1 U79 ( .A(mem[680]), .B(n5611), .Y(n1127) );
  INVX1 U80 ( .A(n1127), .Y(n111) );
  AND2X1 U81 ( .A(mem[639]), .B(n5612), .Y(n1085) );
  INVX1 U82 ( .A(n1085), .Y(n112) );
  AND2X1 U83 ( .A(mem[598]), .B(n5613), .Y(n1043) );
  INVX1 U84 ( .A(n1043), .Y(n113) );
  AND2X1 U85 ( .A(mem[557]), .B(n5614), .Y(n1001) );
  INVX1 U86 ( .A(n1001), .Y(n114) );
  AND2X1 U87 ( .A(mem[516]), .B(n5615), .Y(n959) );
  INVX1 U88 ( .A(n959), .Y(n115) );
  AND2X1 U89 ( .A(mem[475]), .B(n5616), .Y(n917) );
  INVX1 U90 ( .A(n917), .Y(n116) );
  AND2X1 U92 ( .A(mem[434]), .B(n5617), .Y(n875) );
  INVX1 U94 ( .A(n875), .Y(n117) );
  AND2X1 U96 ( .A(mem[393]), .B(n5618), .Y(n833) );
  INVX1 U98 ( .A(n833), .Y(n118) );
  AND2X1 U100 ( .A(mem[352]), .B(n5619), .Y(n790) );
  INVX1 U102 ( .A(n790), .Y(n119) );
  AND2X1 U104 ( .A(mem[311]), .B(n5620), .Y(n747) );
  INVX1 U106 ( .A(n747), .Y(n120) );
  AND2X1 U108 ( .A(mem[270]), .B(n5621), .Y(n704) );
  INVX1 U110 ( .A(n704), .Y(n121) );
  AND2X1 U112 ( .A(mem[229]), .B(n5622), .Y(n661) );
  INVX1 U114 ( .A(n661), .Y(n122) );
  AND2X1 U116 ( .A(mem[188]), .B(n5623), .Y(n618) );
  INVX1 U118 ( .A(n618), .Y(n123) );
  AND2X1 U120 ( .A(mem[147]), .B(n5624), .Y(n575) );
  INVX1 U122 ( .A(n575), .Y(n124) );
  AND2X1 U124 ( .A(mem[106]), .B(n5625), .Y(n532) );
  INVX1 U126 ( .A(n532), .Y(n125) );
  AND2X1 U128 ( .A(mem[65]), .B(n5626), .Y(n489) );
  INVX1 U130 ( .A(n489), .Y(n126) );
  AND2X1 U132 ( .A(mem[24]), .B(n5627), .Y(n429) );
  INVX1 U134 ( .A(n429), .Y(n127) );
  AND2X1 U136 ( .A(mem[1305]), .B(n5596), .Y(n1769) );
  INVX1 U138 ( .A(n1769), .Y(n128) );
  AND2X1 U140 ( .A(mem[1290]), .B(n5596), .Y(n1754) );
  INVX1 U142 ( .A(n1754), .Y(n129) );
  AND2X1 U144 ( .A(mem[1276]), .B(n5596), .Y(n1740) );
  INVX1 U146 ( .A(n1740), .Y(n130) );
  AND2X1 U148 ( .A(mem[1265]), .B(n5597), .Y(n1728) );
  INVX1 U150 ( .A(n1728), .Y(n131) );
  AND2X1 U152 ( .A(mem[1250]), .B(n5597), .Y(n1713) );
  INVX1 U154 ( .A(n1713), .Y(n132) );
  AND2X1 U156 ( .A(mem[1236]), .B(n5597), .Y(n1699) );
  INVX1 U158 ( .A(n1699), .Y(n133) );
  AND2X1 U160 ( .A(mem[1225]), .B(n5598), .Y(n1687) );
  INVX1 U162 ( .A(n1687), .Y(n134) );
  AND2X1 U164 ( .A(mem[1210]), .B(n5598), .Y(n1672) );
  INVX1 U166 ( .A(n1672), .Y(n135) );
  AND2X1 U168 ( .A(mem[1196]), .B(n5598), .Y(n1658) );
  INVX1 U170 ( .A(n1658), .Y(n136) );
  AND2X1 U172 ( .A(mem[1174]), .B(n5599), .Y(n1635) );
  INVX1 U175 ( .A(n1635), .Y(n137) );
  AND2X1 U177 ( .A(mem[1161]), .B(n5599), .Y(n1622) );
  INVX1 U179 ( .A(n1622), .Y(n138) );
  AND2X1 U181 ( .A(mem[1156]), .B(n5599), .Y(n1617) );
  INVX1 U183 ( .A(n1617), .Y(n139) );
  AND2X1 U185 ( .A(mem[1147]), .B(n5600), .Y(n1607) );
  INVX1 U187 ( .A(n1607), .Y(n140) );
  AND2X1 U189 ( .A(mem[1137]), .B(n5600), .Y(n1597) );
  INVX1 U191 ( .A(n1597), .Y(n141) );
  AND2X1 U193 ( .A(mem[1116]), .B(n5600), .Y(n1576) );
  INVX1 U195 ( .A(n1576), .Y(n142) );
  AND2X1 U197 ( .A(mem[1097]), .B(n5601), .Y(n1556) );
  INVX1 U199 ( .A(n1556), .Y(n143) );
  AND2X1 U201 ( .A(mem[1080]), .B(n5601), .Y(n1539) );
  INVX1 U203 ( .A(n1539), .Y(n144) );
  AND2X1 U205 ( .A(mem[1057]), .B(n5602), .Y(n1515) );
  INVX1 U207 ( .A(n1515), .Y(n145) );
  AND2X1 U209 ( .A(mem[1040]), .B(n5602), .Y(n1498) );
  INVX1 U211 ( .A(n1498), .Y(n146) );
  AND2X1 U213 ( .A(mem[1017]), .B(n5603), .Y(n1473) );
  INVX1 U215 ( .A(n1473), .Y(n147) );
  AND2X1 U217 ( .A(mem[1000]), .B(n5603), .Y(n1456) );
  INVX1 U219 ( .A(n1456), .Y(n148) );
  AND2X1 U221 ( .A(mem[980]), .B(n5604), .Y(n1435) );
  INVX1 U223 ( .A(n1435), .Y(n149) );
  AND2X1 U225 ( .A(mem[960]), .B(n5604), .Y(n1415) );
  INVX1 U227 ( .A(n1415), .Y(n150) );
  AND2X1 U229 ( .A(mem[940]), .B(n5605), .Y(n1394) );
  INVX1 U231 ( .A(n1394), .Y(n151) );
  AND2X1 U233 ( .A(mem[920]), .B(n5605), .Y(n1374) );
  INVX1 U235 ( .A(n1374), .Y(n152) );
  AND2X1 U237 ( .A(mem[900]), .B(n5606), .Y(n1353) );
  INVX1 U239 ( .A(n1353), .Y(n153) );
  AND2X1 U241 ( .A(mem[883]), .B(n5606), .Y(n1336) );
  INVX1 U243 ( .A(n1336), .Y(n154) );
  AND2X1 U245 ( .A(mem[843]), .B(n5607), .Y(n1295) );
  INVX1 U247 ( .A(n1295), .Y(n155) );
  AND2X1 U249 ( .A(mem[813]), .B(n5608), .Y(n1264) );
  INVX1 U251 ( .A(n1264), .Y(n156) );
  AND2X1 U253 ( .A(mem[798]), .B(n5608), .Y(n1249) );
  INVX1 U255 ( .A(n1249), .Y(n157) );
  AND2X1 U258 ( .A(mem[784]), .B(n5608), .Y(n1235) );
  INVX1 U260 ( .A(n1235), .Y(n158) );
  AND2X1 U262 ( .A(mem[773]), .B(n5609), .Y(n1223) );
  INVX1 U264 ( .A(n1223), .Y(n159) );
  AND2X1 U266 ( .A(mem[758]), .B(n5609), .Y(n1208) );
  INVX1 U268 ( .A(n1208), .Y(n160) );
  AND2X1 U270 ( .A(mem[744]), .B(n5609), .Y(n1194) );
  INVX1 U272 ( .A(n1194), .Y(n161) );
  AND2X1 U274 ( .A(mem[733]), .B(n5610), .Y(n1182) );
  INVX1 U276 ( .A(n1182), .Y(n162) );
  AND2X1 U278 ( .A(mem[718]), .B(n5610), .Y(n1167) );
  INVX1 U280 ( .A(n1167), .Y(n163) );
  AND2X1 U282 ( .A(mem[704]), .B(n5610), .Y(n1153) );
  INVX1 U284 ( .A(n1153), .Y(n164) );
  AND2X1 U286 ( .A(mem[682]), .B(n5611), .Y(n1129) );
  INVX1 U288 ( .A(n1129), .Y(n165) );
  AND2X1 U290 ( .A(mem[669]), .B(n5611), .Y(n1116) );
  INVX1 U292 ( .A(n1116), .Y(n166) );
  AND2X1 U294 ( .A(mem[664]), .B(n5611), .Y(n1111) );
  INVX1 U296 ( .A(n1111), .Y(n167) );
  AND2X1 U298 ( .A(mem[655]), .B(n5612), .Y(n1101) );
  INVX1 U300 ( .A(n1101), .Y(n168) );
  AND2X1 U302 ( .A(mem[645]), .B(n5612), .Y(n1091) );
  INVX1 U304 ( .A(n1091), .Y(n169) );
  AND2X1 U306 ( .A(mem[624]), .B(n5612), .Y(n1070) );
  INVX1 U308 ( .A(n1070), .Y(n170) );
  AND2X1 U310 ( .A(mem[605]), .B(n5613), .Y(n1050) );
  INVX1 U312 ( .A(n1050), .Y(n171) );
  AND2X1 U314 ( .A(mem[588]), .B(n5613), .Y(n1033) );
  INVX1 U316 ( .A(n1033), .Y(n172) );
  AND2X1 U318 ( .A(mem[565]), .B(n5614), .Y(n1009) );
  INVX1 U320 ( .A(n1009), .Y(n173) );
  AND2X1 U322 ( .A(mem[548]), .B(n5614), .Y(n992) );
  INVX1 U324 ( .A(n992), .Y(n174) );
  AND2X1 U326 ( .A(mem[525]), .B(n5615), .Y(n968) );
  INVX1 U328 ( .A(n968), .Y(n175) );
  AND2X1 U330 ( .A(mem[508]), .B(n5615), .Y(n951) );
  INVX1 U332 ( .A(n951), .Y(n176) );
  AND2X1 U334 ( .A(mem[488]), .B(n5616), .Y(n930) );
  INVX1 U336 ( .A(n930), .Y(n177) );
  AND2X1 U338 ( .A(mem[468]), .B(n5616), .Y(n910) );
  INVX1 U341 ( .A(n910), .Y(n178) );
  AND2X1 U343 ( .A(mem[448]), .B(n5617), .Y(n889) );
  INVX1 U345 ( .A(n889), .Y(n179) );
  AND2X1 U347 ( .A(mem[428]), .B(n5617), .Y(n869) );
  INVX1 U349 ( .A(n869), .Y(n180) );
  AND2X1 U351 ( .A(mem[408]), .B(n5618), .Y(n848) );
  INVX1 U353 ( .A(n848), .Y(n181) );
  AND2X1 U355 ( .A(mem[391]), .B(n5618), .Y(n831) );
  INVX1 U357 ( .A(n831), .Y(n182) );
  AND2X1 U359 ( .A(mem[351]), .B(n5619), .Y(n789) );
  INVX1 U361 ( .A(n789), .Y(n183) );
  AND2X1 U363 ( .A(mem[327]), .B(n5620), .Y(n763) );
  INVX1 U365 ( .A(n763), .Y(n184) );
  AND2X1 U367 ( .A(mem[317]), .B(n5620), .Y(n753) );
  INVX1 U369 ( .A(n753), .Y(n185) );
  AND2X1 U371 ( .A(mem[296]), .B(n5620), .Y(n732) );
  INVX1 U373 ( .A(n732), .Y(n186) );
  AND2X1 U375 ( .A(mem[277]), .B(n5621), .Y(n711) );
  INVX1 U377 ( .A(n711), .Y(n187) );
  AND2X1 U379 ( .A(mem[260]), .B(n5621), .Y(n694) );
  INVX1 U381 ( .A(n694), .Y(n188) );
  AND2X1 U383 ( .A(mem[237]), .B(n5622), .Y(n669) );
  INVX1 U385 ( .A(n669), .Y(n189) );
  AND2X1 U387 ( .A(mem[220]), .B(n5622), .Y(n652) );
  INVX1 U389 ( .A(n652), .Y(n190) );
  AND2X1 U391 ( .A(mem[197]), .B(n5623), .Y(n627) );
  INVX1 U393 ( .A(n627), .Y(n191) );
  AND2X1 U395 ( .A(mem[180]), .B(n5623), .Y(n610) );
  INVX1 U397 ( .A(n610), .Y(n192) );
  AND2X1 U399 ( .A(mem[160]), .B(n5624), .Y(n588) );
  INVX1 U401 ( .A(n588), .Y(n193) );
  AND2X1 U403 ( .A(mem[140]), .B(n5624), .Y(n568) );
  INVX1 U405 ( .A(n568), .Y(n194) );
  AND2X1 U407 ( .A(mem[120]), .B(n5625), .Y(n546) );
  INVX1 U409 ( .A(n546), .Y(n195) );
  AND2X1 U411 ( .A(mem[100]), .B(n5625), .Y(n526) );
  INVX1 U413 ( .A(n526), .Y(n196) );
  AND2X1 U415 ( .A(mem[80]), .B(n5626), .Y(n504) );
  INVX1 U417 ( .A(n504), .Y(n197) );
  AND2X1 U419 ( .A(mem[63]), .B(n5626), .Y(n487) );
  INVX1 U421 ( .A(n487), .Y(n198) );
  AND2X1 U424 ( .A(mem[23]), .B(n5627), .Y(n427) );
  INVX1 U426 ( .A(n427), .Y(n199) );
  AND2X1 U428 ( .A(mem[1306]), .B(n5596), .Y(n1770) );
  INVX1 U430 ( .A(n1770), .Y(n200) );
  AND2X1 U432 ( .A(mem[1291]), .B(n5596), .Y(n1755) );
  INVX1 U434 ( .A(n1755), .Y(n201) );
  AND2X1 U436 ( .A(mem[1277]), .B(n5596), .Y(n1741) );
  INVX1 U438 ( .A(n1741), .Y(n202) );
  AND2X1 U440 ( .A(mem[1264]), .B(n5597), .Y(n1727) );
  INVX1 U442 ( .A(n1727), .Y(n203) );
  AND2X1 U444 ( .A(mem[1249]), .B(n5597), .Y(n1712) );
  INVX1 U446 ( .A(n1712), .Y(n204) );
  AND2X1 U448 ( .A(mem[1235]), .B(n5597), .Y(n1698) );
  INVX1 U450 ( .A(n1698), .Y(n205) );
  AND2X1 U452 ( .A(mem[1215]), .B(n5598), .Y(n1677) );
  INVX1 U454 ( .A(n1677), .Y(n206) );
  AND2X1 U456 ( .A(mem[1202]), .B(n5598), .Y(n1664) );
  INVX1 U458 ( .A(n1664), .Y(n207) );
  AND2X1 U460 ( .A(mem[1197]), .B(n5598), .Y(n1659) );
  INVX1 U462 ( .A(n1659), .Y(n208) );
  AND2X1 U464 ( .A(mem[1184]), .B(n5599), .Y(n1645) );
  INVX1 U466 ( .A(n1645), .Y(n209) );
  AND2X1 U468 ( .A(mem[1169]), .B(n5599), .Y(n1630) );
  INVX1 U470 ( .A(n1630), .Y(n210) );
  AND2X1 U472 ( .A(mem[1155]), .B(n5599), .Y(n1616) );
  INVX1 U474 ( .A(n1616), .Y(n211) );
  AND2X1 U476 ( .A(mem[1138]), .B(n5600), .Y(n1598) );
  INVX1 U478 ( .A(n1598), .Y(n212) );
  AND2X1 U480 ( .A(mem[1121]), .B(n5600), .Y(n1581) );
  INVX1 U482 ( .A(n1581), .Y(n213) );
  AND2X1 U484 ( .A(mem[1106]), .B(n5601), .Y(n1565) );
  INVX1 U486 ( .A(n1565), .Y(n214) );
  AND2X1 U488 ( .A(mem[1096]), .B(n5601), .Y(n1555) );
  INVX1 U490 ( .A(n1555), .Y(n215) );
  AND2X1 U492 ( .A(mem[1075]), .B(n5601), .Y(n1534) );
  INVX1 U494 ( .A(n1534), .Y(n216) );
  AND2X1 U496 ( .A(mem[1058]), .B(n5602), .Y(n1516) );
  INVX1 U498 ( .A(n1516), .Y(n217) );
  AND2X1 U500 ( .A(mem[1041]), .B(n5602), .Y(n1499) );
  INVX1 U502 ( .A(n1499), .Y(n218) );
  AND2X1 U504 ( .A(mem[1016]), .B(n5603), .Y(n1472) );
  INVX1 U507 ( .A(n1472), .Y(n219) );
  AND2X1 U509 ( .A(mem[999]), .B(n5603), .Y(n1455) );
  INVX1 U511 ( .A(n1455), .Y(n220) );
  AND2X1 U513 ( .A(mem[981]), .B(n5604), .Y(n1436) );
  INVX1 U515 ( .A(n1436), .Y(n221) );
  AND2X1 U517 ( .A(mem[961]), .B(n5604), .Y(n1416) );
  INVX1 U519 ( .A(n1416), .Y(n222) );
  AND2X1 U521 ( .A(mem[939]), .B(n5605), .Y(n1393) );
  INVX1 U523 ( .A(n1393), .Y(n223) );
  AND2X1 U525 ( .A(mem[919]), .B(n5605), .Y(n1373) );
  INVX1 U527 ( .A(n1373), .Y(n224) );
  AND2X1 U529 ( .A(mem[884]), .B(n5606), .Y(n1337) );
  INVX1 U531 ( .A(n1337), .Y(n225) );
  AND2X1 U533 ( .A(mem[859]), .B(n5607), .Y(n1311) );
  INVX1 U535 ( .A(n1311), .Y(n226) );
  AND2X1 U537 ( .A(mem[842]), .B(n5607), .Y(n1294) );
  INVX1 U539 ( .A(n1294), .Y(n227) );
  AND2X1 U541 ( .A(mem[814]), .B(n5608), .Y(n1265) );
  INVX1 U543 ( .A(n1265), .Y(n228) );
  AND2X1 U545 ( .A(mem[799]), .B(n5608), .Y(n1250) );
  INVX1 U547 ( .A(n1250), .Y(n229) );
  AND2X1 U549 ( .A(mem[785]), .B(n5608), .Y(n1236) );
  INVX1 U551 ( .A(n1236), .Y(n230) );
  AND2X1 U553 ( .A(mem[772]), .B(n5609), .Y(n1222) );
  INVX1 U555 ( .A(n1222), .Y(n231) );
  AND2X1 U557 ( .A(mem[757]), .B(n5609), .Y(n1207) );
  INVX1 U559 ( .A(n1207), .Y(n232) );
  AND2X1 U561 ( .A(mem[743]), .B(n5609), .Y(n1193) );
  INVX1 U563 ( .A(n1193), .Y(n233) );
  AND2X1 U565 ( .A(mem[723]), .B(n5610), .Y(n1172) );
  INVX1 U567 ( .A(n1172), .Y(n234) );
  AND2X1 U569 ( .A(mem[710]), .B(n5610), .Y(n1159) );
  INVX1 U571 ( .A(n1159), .Y(n235) );
  AND2X1 U573 ( .A(mem[705]), .B(n5610), .Y(n1154) );
  INVX1 U575 ( .A(n1154), .Y(n236) );
  AND2X1 U577 ( .A(mem[692]), .B(n5611), .Y(n1139) );
  INVX1 U579 ( .A(n1139), .Y(n237) );
  AND2X1 U581 ( .A(mem[677]), .B(n5611), .Y(n1124) );
  INVX1 U583 ( .A(n1124), .Y(n238) );
  AND2X1 U585 ( .A(mem[663]), .B(n5611), .Y(n1110) );
  INVX1 U587 ( .A(n1110), .Y(n239) );
  AND2X1 U590 ( .A(mem[646]), .B(n5612), .Y(n1092) );
  INVX1 U592 ( .A(n1092), .Y(n240) );
  AND2X1 U594 ( .A(mem[629]), .B(n5612), .Y(n1075) );
  INVX1 U596 ( .A(n1075), .Y(n241) );
  AND2X1 U598 ( .A(mem[614]), .B(n5613), .Y(n1059) );
  INVX1 U600 ( .A(n1059), .Y(n242) );
  AND2X1 U602 ( .A(mem[604]), .B(n5613), .Y(n1049) );
  INVX1 U604 ( .A(n1049), .Y(n243) );
  AND2X1 U606 ( .A(mem[583]), .B(n5613), .Y(n1028) );
  INVX1 U608 ( .A(n1028), .Y(n244) );
  AND2X1 U610 ( .A(mem[566]), .B(n5614), .Y(n1010) );
  INVX1 U612 ( .A(n1010), .Y(n245) );
  AND2X1 U614 ( .A(mem[549]), .B(n5614), .Y(n993) );
  INVX1 U616 ( .A(n993), .Y(n246) );
  AND2X1 U618 ( .A(mem[524]), .B(n5615), .Y(n967) );
  INVX1 U620 ( .A(n967), .Y(n247) );
  AND2X1 U622 ( .A(mem[507]), .B(n5615), .Y(n950) );
  INVX1 U624 ( .A(n950), .Y(n248) );
  AND2X1 U626 ( .A(mem[489]), .B(n5616), .Y(n931) );
  INVX1 U628 ( .A(n931), .Y(n249) );
  AND2X1 U630 ( .A(mem[469]), .B(n5616), .Y(n911) );
  INVX1 U632 ( .A(n911), .Y(n250) );
  AND2X1 U634 ( .A(mem[447]), .B(n5617), .Y(n888) );
  INVX1 U636 ( .A(n888), .Y(n251) );
  AND2X1 U638 ( .A(mem[427]), .B(n5617), .Y(n868) );
  INVX1 U640 ( .A(n868), .Y(n252) );
  AND2X1 U642 ( .A(mem[392]), .B(n5618), .Y(n832) );
  INVX1 U644 ( .A(n832), .Y(n253) );
  AND2X1 U646 ( .A(mem[367]), .B(n5619), .Y(n805) );
  INVX1 U648 ( .A(n805), .Y(n254) );
  AND2X1 U650 ( .A(mem[350]), .B(n5619), .Y(n788) );
  INVX1 U652 ( .A(n788), .Y(n255) );
  AND2X1 U654 ( .A(mem[318]), .B(n5620), .Y(n754) );
  INVX1 U656 ( .A(n754), .Y(n256) );
  AND2X1 U658 ( .A(mem[301]), .B(n5620), .Y(n737) );
  INVX1 U660 ( .A(n737), .Y(n257) );
  AND2X1 U662 ( .A(mem[286]), .B(n5621), .Y(n720) );
  INVX1 U664 ( .A(n720), .Y(n258) );
  AND2X1 U666 ( .A(mem[276]), .B(n5621), .Y(n710) );
  INVX1 U668 ( .A(n710), .Y(n259) );
  AND2X1 U670 ( .A(mem[255]), .B(n5621), .Y(n689) );
  INVX1 U673 ( .A(n689), .Y(n260) );
  AND2X1 U675 ( .A(mem[238]), .B(n5622), .Y(n670) );
  INVX1 U677 ( .A(n670), .Y(n261) );
  AND2X1 U679 ( .A(mem[221]), .B(n5622), .Y(n653) );
  INVX1 U681 ( .A(n653), .Y(n262) );
  AND2X1 U683 ( .A(mem[196]), .B(n5623), .Y(n626) );
  INVX1 U685 ( .A(n626), .Y(n263) );
  AND2X1 U687 ( .A(mem[179]), .B(n5623), .Y(n609) );
  INVX1 U689 ( .A(n609), .Y(n264) );
  AND2X1 U691 ( .A(mem[161]), .B(n5624), .Y(n589) );
  INVX1 U693 ( .A(n589), .Y(n265) );
  AND2X1 U695 ( .A(mem[141]), .B(n5624), .Y(n569) );
  INVX1 U697 ( .A(n569), .Y(n266) );
  AND2X1 U699 ( .A(mem[119]), .B(n5625), .Y(n545) );
  INVX1 U701 ( .A(n545), .Y(n267) );
  AND2X1 U703 ( .A(mem[99]), .B(n5625), .Y(n525) );
  INVX1 U705 ( .A(n525), .Y(n268) );
  AND2X1 U707 ( .A(mem[64]), .B(n5626), .Y(n488) );
  INVX1 U709 ( .A(n488), .Y(n269) );
  AND2X1 U711 ( .A(mem[39]), .B(n5627), .Y(n459) );
  INVX1 U713 ( .A(n459), .Y(n270) );
  AND2X1 U715 ( .A(mem[22]), .B(n5627), .Y(n425) );
  INVX1 U717 ( .A(n425), .Y(n271) );
  AND2X1 U719 ( .A(mem[1307]), .B(n5596), .Y(n1771) );
  INVX1 U721 ( .A(n1771), .Y(n272) );
  AND2X1 U723 ( .A(mem[1292]), .B(n5596), .Y(n1756) );
  INVX1 U725 ( .A(n1756), .Y(n273) );
  AND2X1 U727 ( .A(mem[1278]), .B(n5596), .Y(n1742) );
  INVX1 U729 ( .A(n1742), .Y(n274) );
  AND2X1 U731 ( .A(mem[1256]), .B(n5597), .Y(n1719) );
  INVX1 U733 ( .A(n1719), .Y(n275) );
  AND2X1 U735 ( .A(mem[1243]), .B(n5597), .Y(n1706) );
  INVX1 U737 ( .A(n1706), .Y(n276) );
  AND2X1 U739 ( .A(mem[1238]), .B(n5597), .Y(n1701) );
  INVX1 U741 ( .A(n1701), .Y(n277) );
  AND2X1 U743 ( .A(mem[1223]), .B(n5598), .Y(n1685) );
  INVX1 U745 ( .A(n1685), .Y(n278) );
  AND2X1 U747 ( .A(mem[1208]), .B(n5598), .Y(n1670) );
  INVX1 U749 ( .A(n1670), .Y(n279) );
  AND2X1 U751 ( .A(mem[1194]), .B(n5598), .Y(n1656) );
  INVX1 U753 ( .A(n1656), .Y(n280) );
  AND2X1 U757 ( .A(mem[1183]), .B(n5599), .Y(n1644) );
  INVX1 U759 ( .A(n1644), .Y(n281) );
  AND2X1 U761 ( .A(mem[1168]), .B(n5599), .Y(n1629) );
  INVX1 U763 ( .A(n1629), .Y(n282) );
  AND2X1 U765 ( .A(mem[1154]), .B(n5599), .Y(n1615) );
  INVX1 U767 ( .A(n1615), .Y(n283) );
  AND2X1 U769 ( .A(mem[1139]), .B(n5600), .Y(n1599) );
  INVX1 U771 ( .A(n1599), .Y(n284) );
  AND2X1 U773 ( .A(mem[1122]), .B(n5600), .Y(n1582) );
  INVX1 U775 ( .A(n1582), .Y(n285) );
  AND2X1 U777 ( .A(mem[1099]), .B(n5601), .Y(n1558) );
  INVX1 U779 ( .A(n1558), .Y(n286) );
  AND2X1 U781 ( .A(mem[1082]), .B(n5601), .Y(n1541) );
  INVX1 U783 ( .A(n1541), .Y(n287) );
  AND2X1 U785 ( .A(mem[1065]), .B(n5602), .Y(n1523) );
  INVX1 U787 ( .A(n1523), .Y(n288) );
  AND2X1 U789 ( .A(mem[1055]), .B(n5602), .Y(n1513) );
  INVX1 U791 ( .A(n1513), .Y(n289) );
  AND2X1 U793 ( .A(mem[1034]), .B(n5602), .Y(n1492) );
  INVX1 U795 ( .A(n1492), .Y(n290) );
  AND2X1 U797 ( .A(mem[1015]), .B(n5603), .Y(n1471) );
  INVX1 U799 ( .A(n1471), .Y(n291) );
  AND2X1 U801 ( .A(mem[998]), .B(n5603), .Y(n1454) );
  INVX1 U803 ( .A(n1454), .Y(n292) );
  AND2X1 U805 ( .A(mem[982]), .B(n5604), .Y(n1437) );
  INVX1 U807 ( .A(n1437), .Y(n293) );
  AND2X1 U809 ( .A(mem[965]), .B(n5604), .Y(n1420) );
  INVX1 U811 ( .A(n1420), .Y(n294) );
  AND2X1 U813 ( .A(mem[925]), .B(n5605), .Y(n1379) );
  INVX1 U815 ( .A(n1379), .Y(n295) );
  AND2X1 U817 ( .A(mem[898]), .B(n5606), .Y(n1351) );
  INVX1 U819 ( .A(n1351), .Y(n296) );
  AND2X1 U821 ( .A(mem[878]), .B(n5606), .Y(n1331) );
  INVX1 U823 ( .A(n1331), .Y(n297) );
  AND2X1 U825 ( .A(mem[858]), .B(n5607), .Y(n1310) );
  INVX1 U827 ( .A(n1310), .Y(n298) );
  AND2X1 U829 ( .A(mem[838]), .B(n5607), .Y(n1290) );
  INVX1 U831 ( .A(n1290), .Y(n299) );
  AND2X1 U833 ( .A(mem[815]), .B(n5608), .Y(n1266) );
  INVX1 U835 ( .A(n1266), .Y(n300) );
  AND2X1 U837 ( .A(mem[800]), .B(n5608), .Y(n1251) );
  INVX1 U840 ( .A(n1251), .Y(n301) );
  AND2X1 U842 ( .A(mem[786]), .B(n5608), .Y(n1237) );
  INVX1 U844 ( .A(n1237), .Y(n302) );
  AND2X1 U846 ( .A(mem[764]), .B(n5609), .Y(n1214) );
  INVX1 U848 ( .A(n1214), .Y(n303) );
  AND2X1 U850 ( .A(mem[751]), .B(n5609), .Y(n1201) );
  INVX1 U852 ( .A(n1201), .Y(n304) );
  AND2X1 U854 ( .A(mem[746]), .B(n5609), .Y(n1196) );
  INVX1 U856 ( .A(n1196), .Y(n305) );
  AND2X1 U858 ( .A(mem[731]), .B(n5610), .Y(n1180) );
  INVX1 U860 ( .A(n1180), .Y(n306) );
  AND2X1 U862 ( .A(mem[716]), .B(n5610), .Y(n1165) );
  INVX1 U864 ( .A(n1165), .Y(n307) );
  AND2X1 U866 ( .A(mem[702]), .B(n5610), .Y(n1151) );
  INVX1 U868 ( .A(n1151), .Y(n308) );
  AND2X1 U870 ( .A(mem[691]), .B(n5611), .Y(n1138) );
  INVX1 U872 ( .A(n1138), .Y(n309) );
  AND2X1 U874 ( .A(mem[676]), .B(n5611), .Y(n1123) );
  INVX1 U876 ( .A(n1123), .Y(n310) );
  AND2X1 U878 ( .A(mem[662]), .B(n5611), .Y(n1109) );
  INVX1 U880 ( .A(n1109), .Y(n311) );
  AND2X1 U882 ( .A(mem[647]), .B(n5612), .Y(n1093) );
  INVX1 U884 ( .A(n1093), .Y(n312) );
  AND2X1 U886 ( .A(mem[630]), .B(n5612), .Y(n1076) );
  INVX1 U888 ( .A(n1076), .Y(n313) );
  AND2X1 U890 ( .A(mem[607]), .B(n5613), .Y(n1052) );
  INVX1 U892 ( .A(n1052), .Y(n314) );
  AND2X1 U894 ( .A(mem[590]), .B(n5613), .Y(n1035) );
  INVX1 U896 ( .A(n1035), .Y(n315) );
  AND2X1 U898 ( .A(mem[573]), .B(n5614), .Y(n1017) );
  INVX1 U900 ( .A(n1017), .Y(n316) );
  AND2X1 U902 ( .A(mem[563]), .B(n5614), .Y(n1007) );
  INVX1 U904 ( .A(n1007), .Y(n317) );
  AND2X1 U906 ( .A(mem[542]), .B(n5614), .Y(n986) );
  INVX1 U908 ( .A(n986), .Y(n318) );
  AND2X1 U910 ( .A(mem[523]), .B(n5615), .Y(n966) );
  INVX1 U912 ( .A(n966), .Y(n319) );
  AND2X1 U914 ( .A(mem[506]), .B(n5615), .Y(n949) );
  INVX1 U916 ( .A(n949), .Y(n320) );
  AND2X1 U918 ( .A(mem[490]), .B(n5616), .Y(n932) );
  INVX1 U920 ( .A(n932), .Y(n321) );
  AND2X1 U923 ( .A(mem[473]), .B(n5616), .Y(n915) );
  INVX1 U925 ( .A(n915), .Y(n322) );
  AND2X1 U927 ( .A(mem[433]), .B(n5617), .Y(n874) );
  INVX1 U929 ( .A(n874), .Y(n323) );
  AND2X1 U931 ( .A(mem[406]), .B(n5618), .Y(n846) );
  INVX1 U933 ( .A(n846), .Y(n324) );
  AND2X1 U935 ( .A(mem[386]), .B(n5618), .Y(n826) );
  INVX1 U937 ( .A(n826), .Y(n325) );
  AND2X1 U939 ( .A(mem[366]), .B(n5619), .Y(n804) );
  INVX1 U941 ( .A(n804), .Y(n326) );
  AND2X1 U943 ( .A(mem[346]), .B(n5619), .Y(n784) );
  INVX1 U945 ( .A(n784), .Y(n327) );
  AND2X1 U947 ( .A(mem[319]), .B(n5620), .Y(n755) );
  INVX1 U949 ( .A(n755), .Y(n328) );
  AND2X1 U951 ( .A(mem[302]), .B(n5620), .Y(n738) );
  INVX1 U953 ( .A(n738), .Y(n329) );
  AND2X1 U955 ( .A(mem[279]), .B(n5621), .Y(n713) );
  INVX1 U957 ( .A(n713), .Y(n330) );
  AND2X1 U959 ( .A(mem[262]), .B(n5621), .Y(n696) );
  INVX1 U961 ( .A(n696), .Y(n331) );
  AND2X1 U963 ( .A(mem[245]), .B(n5622), .Y(n677) );
  INVX1 U965 ( .A(n677), .Y(n332) );
  AND2X1 U967 ( .A(mem[235]), .B(n5622), .Y(n667) );
  INVX1 U969 ( .A(n667), .Y(n333) );
  AND2X1 U971 ( .A(mem[214]), .B(n5622), .Y(n646) );
  INVX1 U973 ( .A(n646), .Y(n334) );
  AND2X1 U975 ( .A(mem[195]), .B(n5623), .Y(n625) );
  INVX1 U977 ( .A(n625), .Y(n335) );
  AND2X1 U979 ( .A(mem[178]), .B(n5623), .Y(n608) );
  INVX1 U981 ( .A(n608), .Y(n336) );
  AND2X1 U983 ( .A(mem[162]), .B(n5624), .Y(n590) );
  INVX1 U985 ( .A(n590), .Y(n337) );
  AND2X1 U987 ( .A(mem[145]), .B(n5624), .Y(n573) );
  INVX1 U989 ( .A(n573), .Y(n338) );
  AND2X1 U991 ( .A(mem[105]), .B(n5625), .Y(n531) );
  INVX1 U993 ( .A(n531), .Y(n339) );
  AND2X1 U995 ( .A(mem[78]), .B(n5626), .Y(n502) );
  INVX1 U997 ( .A(n502), .Y(n340) );
  AND2X1 U999 ( .A(mem[58]), .B(n5626), .Y(n482) );
  INVX1 U1001 ( .A(n482), .Y(n341) );
  AND2X1 U1003 ( .A(mem[38]), .B(n5627), .Y(n457) );
  INVX1 U1006 ( .A(n457), .Y(n342) );
  AND2X1 U1008 ( .A(mem[18]), .B(n5627), .Y(n417) );
  INVX1 U1010 ( .A(n417), .Y(n343) );
  AND2X1 U1012 ( .A(mem[1297]), .B(n5596), .Y(n1761) );
  INVX1 U1014 ( .A(n1761), .Y(n344) );
  AND2X1 U1016 ( .A(mem[1284]), .B(n5596), .Y(n1748) );
  INVX1 U1018 ( .A(n1748), .Y(n345) );
  AND2X1 U1020 ( .A(mem[1279]), .B(n5596), .Y(n1743) );
  INVX1 U1022 ( .A(n1743), .Y(n346) );
  AND2X1 U1024 ( .A(mem[1266]), .B(n5597), .Y(n1729) );
  INVX1 U1026 ( .A(n1729), .Y(n347) );
  AND2X1 U1028 ( .A(mem[1251]), .B(n5597), .Y(n1714) );
  INVX1 U1030 ( .A(n1714), .Y(n348) );
  AND2X1 U1032 ( .A(mem[1237]), .B(n5597), .Y(n1700) );
  INVX1 U1034 ( .A(n1700), .Y(n349) );
  AND2X1 U1036 ( .A(mem[1224]), .B(n5598), .Y(n1686) );
  INVX1 U1038 ( .A(n1686), .Y(n350) );
  AND2X1 U1040 ( .A(mem[1209]), .B(n5598), .Y(n1671) );
  INVX1 U1042 ( .A(n1671), .Y(n351) );
  AND2X1 U1044 ( .A(mem[1195]), .B(n5598), .Y(n1657) );
  INVX1 U1046 ( .A(n1657), .Y(n352) );
  AND2X1 U1048 ( .A(mem[1182]), .B(n5599), .Y(n1643) );
  INVX1 U1050 ( .A(n1643), .Y(n353) );
  AND2X1 U1052 ( .A(mem[1167]), .B(n5599), .Y(n1628) );
  INVX1 U1054 ( .A(n1628), .Y(n354) );
  AND2X1 U1056 ( .A(mem[1153]), .B(n5599), .Y(n1614) );
  INVX1 U1058 ( .A(n1614), .Y(n355) );
  AND2X1 U1060 ( .A(mem[1140]), .B(n5600), .Y(n1600) );
  INVX1 U1062 ( .A(n1600), .Y(n356) );
  AND2X1 U1064 ( .A(mem[1123]), .B(n5600), .Y(n1583) );
  INVX1 U1066 ( .A(n1583), .Y(n357) );
  AND2X1 U1068 ( .A(mem[1098]), .B(n5601), .Y(n1557) );
  INVX1 U1070 ( .A(n1557), .Y(n358) );
  AND2X1 U1072 ( .A(mem[1081]), .B(n5601), .Y(n1540) );
  INVX1 U1074 ( .A(n1540), .Y(n359) );
  AND2X1 U1076 ( .A(mem[1056]), .B(n5602), .Y(n1514) );
  INVX1 U1078 ( .A(n1514), .Y(n360) );
  AND2X1 U1080 ( .A(mem[1039]), .B(n5602), .Y(n1497) );
  INVX1 U1082 ( .A(n1497), .Y(n361) );
  AND2X1 U1084 ( .A(mem[1024]), .B(n5603), .Y(n1480) );
  INVX1 U1086 ( .A(n1480), .Y(n362) );
  AND2X1 U1089 ( .A(mem[1014]), .B(n5603), .Y(n1470) );
  INVX1 U1091 ( .A(n1470), .Y(n363) );
  AND2X1 U1093 ( .A(mem[993]), .B(n5603), .Y(n1449) );
  INVX1 U1095 ( .A(n1449), .Y(n364) );
  AND2X1 U1097 ( .A(mem[966]), .B(n5604), .Y(n1421) );
  INVX1 U1099 ( .A(n1421), .Y(n365) );
  AND2X1 U1101 ( .A(mem[941]), .B(n5605), .Y(n1395) );
  INVX1 U1103 ( .A(n1395), .Y(n366) );
  AND2X1 U1105 ( .A(mem[924]), .B(n5605), .Y(n1378) );
  INVX1 U1107 ( .A(n1378), .Y(n367) );
  AND2X1 U1109 ( .A(mem[899]), .B(n5606), .Y(n1352) );
  INVX1 U1111 ( .A(n1352), .Y(n368) );
  AND2X1 U1113 ( .A(mem[879]), .B(n5606), .Y(n1332) );
  INVX1 U1115 ( .A(n1332), .Y(n369) );
  AND2X1 U1117 ( .A(mem[857]), .B(n5607), .Y(n1309) );
  INVX1 U1119 ( .A(n1309), .Y(n370) );
  AND2X1 U1121 ( .A(mem[837]), .B(n5607), .Y(n1289) );
  INVX1 U1123 ( .A(n1289), .Y(n371) );
  AND2X1 U1125 ( .A(mem[805]), .B(n5608), .Y(n1256) );
  INVX1 U1127 ( .A(n1256), .Y(n372) );
  AND2X1 U1129 ( .A(mem[792]), .B(n5608), .Y(n1243) );
  INVX1 U1131 ( .A(n1243), .Y(n373) );
  AND2X1 U1133 ( .A(mem[787]), .B(n5608), .Y(n1238) );
  INVX1 U1135 ( .A(n1238), .Y(n374) );
  AND2X1 U1137 ( .A(mem[774]), .B(n5609), .Y(n1224) );
  INVX1 U1139 ( .A(n1224), .Y(n375) );
  AND2X1 U1141 ( .A(mem[759]), .B(n5609), .Y(n1209) );
  INVX1 U1143 ( .A(n1209), .Y(n376) );
  AND2X1 U1145 ( .A(mem[745]), .B(n5609), .Y(n1195) );
  INVX1 U1147 ( .A(n1195), .Y(n377) );
  AND2X1 U1149 ( .A(mem[732]), .B(n5610), .Y(n1181) );
  INVX1 U1151 ( .A(n1181), .Y(n378) );
  AND2X1 U1153 ( .A(mem[717]), .B(n5610), .Y(n1166) );
  INVX1 U1155 ( .A(n1166), .Y(n379) );
  AND2X1 U1157 ( .A(mem[703]), .B(n5610), .Y(n1152) );
  INVX1 U1159 ( .A(n1152), .Y(n380) );
  AND2X1 U1161 ( .A(mem[690]), .B(n5611), .Y(n1137) );
  INVX1 U1163 ( .A(n1137), .Y(n382) );
  AND2X1 U1165 ( .A(mem[675]), .B(n5611), .Y(n1122) );
  INVX1 U1167 ( .A(n1122), .Y(n384) );
  AND2X1 U1169 ( .A(mem[661]), .B(n5611), .Y(n1108) );
  INVX1 U1172 ( .A(n1108), .Y(n386) );
  AND2X1 U1174 ( .A(mem[648]), .B(n5612), .Y(n1094) );
  INVX1 U1176 ( .A(n1094), .Y(n388) );
  AND2X1 U1178 ( .A(mem[631]), .B(n5612), .Y(n1077) );
  INVX1 U1180 ( .A(n1077), .Y(n390) );
  AND2X1 U1182 ( .A(mem[606]), .B(n5613), .Y(n1051) );
  INVX1 U1184 ( .A(n1051), .Y(n392) );
  AND2X1 U1186 ( .A(mem[589]), .B(n5613), .Y(n1034) );
  INVX1 U1188 ( .A(n1034), .Y(n394) );
  AND2X1 U1190 ( .A(mem[564]), .B(n5614), .Y(n1008) );
  INVX1 U1192 ( .A(n1008), .Y(n396) );
  AND2X1 U1194 ( .A(mem[547]), .B(n5614), .Y(n991) );
  INVX1 U1196 ( .A(n991), .Y(n398) );
  AND2X1 U1198 ( .A(mem[532]), .B(n5615), .Y(n975) );
  INVX1 U1200 ( .A(n975), .Y(n400) );
  AND2X1 U1202 ( .A(mem[522]), .B(n5615), .Y(n965) );
  INVX1 U1204 ( .A(n965), .Y(n402) );
  AND2X1 U1206 ( .A(mem[501]), .B(n5615), .Y(n944) );
  INVX1 U1208 ( .A(n944), .Y(n404) );
  AND2X1 U1210 ( .A(mem[474]), .B(n5616), .Y(n916) );
  INVX1 U1212 ( .A(n916), .Y(n406) );
  AND2X1 U1214 ( .A(mem[449]), .B(n5617), .Y(n890) );
  INVX1 U1216 ( .A(n890), .Y(n408) );
  AND2X1 U1218 ( .A(mem[432]), .B(n5617), .Y(n873) );
  INVX1 U1220 ( .A(n873), .Y(n410) );
  AND2X1 U1222 ( .A(mem[407]), .B(n5618), .Y(n847) );
  INVX1 U1224 ( .A(n847), .Y(n412) );
  AND2X1 U1226 ( .A(mem[387]), .B(n5618), .Y(n827) );
  INVX1 U1228 ( .A(n827), .Y(n414) );
  AND2X1 U1230 ( .A(mem[365]), .B(n5619), .Y(n803) );
  INVX1 U1232 ( .A(n803), .Y(n416) );
  AND2X1 U1234 ( .A(mem[345]), .B(n5619), .Y(n783) );
  INVX1 U1236 ( .A(n783), .Y(n418) );
  AND2X1 U1238 ( .A(mem[320]), .B(n5620), .Y(n756) );
  INVX1 U1240 ( .A(n756), .Y(n420) );
  AND2X1 U1242 ( .A(mem[303]), .B(n5620), .Y(n739) );
  INVX1 U1244 ( .A(n739), .Y(n422) );
  AND2X1 U1246 ( .A(mem[278]), .B(n5621), .Y(n712) );
  INVX1 U1248 ( .A(n712), .Y(n424) );
  AND2X1 U1250 ( .A(mem[261]), .B(n5621), .Y(n695) );
  INVX1 U1252 ( .A(n695), .Y(n426) );
  AND2X1 U1255 ( .A(mem[236]), .B(n5622), .Y(n668) );
  INVX1 U1257 ( .A(n668), .Y(n428) );
  AND2X1 U1259 ( .A(mem[219]), .B(n5622), .Y(n651) );
  INVX1 U1261 ( .A(n651), .Y(n430) );
  AND2X1 U1263 ( .A(mem[204]), .B(n5623), .Y(n634) );
  INVX1 U1265 ( .A(n634), .Y(n432) );
  AND2X1 U1267 ( .A(mem[194]), .B(n5623), .Y(n624) );
  INVX1 U1269 ( .A(n624), .Y(n434) );
  AND2X1 U1271 ( .A(mem[173]), .B(n5623), .Y(n603) );
  INVX1 U1273 ( .A(n603), .Y(n436) );
  AND2X1 U1275 ( .A(mem[146]), .B(n5624), .Y(n574) );
  INVX1 U1277 ( .A(n574), .Y(n438) );
  AND2X1 U1279 ( .A(mem[121]), .B(n5625), .Y(n547) );
  INVX1 U1281 ( .A(n547), .Y(n440) );
  AND2X1 U1283 ( .A(mem[104]), .B(n5625), .Y(n530) );
  INVX1 U1285 ( .A(n530), .Y(n442) );
  AND2X1 U1287 ( .A(mem[79]), .B(n5626), .Y(n503) );
  INVX1 U1289 ( .A(n503), .Y(n444) );
  AND2X1 U1291 ( .A(mem[59]), .B(n5626), .Y(n483) );
  INVX1 U1293 ( .A(n483), .Y(n446) );
  AND2X1 U1295 ( .A(mem[37]), .B(n5627), .Y(n455) );
  INVX1 U1297 ( .A(n455), .Y(n448) );
  AND2X1 U1299 ( .A(mem[17]), .B(n5627), .Y(n415) );
  INVX1 U1301 ( .A(n415), .Y(n450) );
  AND2X1 U1303 ( .A(mem[1296]), .B(n5596), .Y(n1760) );
  INVX1 U1305 ( .A(n1760), .Y(n452) );
  AND2X1 U1307 ( .A(mem[1275]), .B(n5596), .Y(n1739) );
  INVX1 U1309 ( .A(n1739), .Y(n454) );
  AND2X1 U1311 ( .A(mem[1271]), .B(n5596), .Y(n1735) );
  INVX1 U1313 ( .A(n1735), .Y(n456) );
  AND2X1 U1315 ( .A(mem[1257]), .B(n5597), .Y(n1720) );
  INVX1 U1317 ( .A(n1720), .Y(n458) );
  AND2X1 U1319 ( .A(mem[1240]), .B(n5597), .Y(n1703) );
  INVX1 U1321 ( .A(n1703), .Y(n460) );
  AND2X1 U1323 ( .A(mem[1231]), .B(n5597), .Y(n1694) );
  INVX1 U1325 ( .A(n1694), .Y(n3164) );
  AND2X1 U1327 ( .A(mem[1217]), .B(n5598), .Y(n1679) );
  INVX1 U1329 ( .A(n1679), .Y(n3165) );
  AND2X1 U1331 ( .A(mem[1200]), .B(n5598), .Y(n1662) );
  INVX1 U1333 ( .A(n1662), .Y(n3166) );
  AND2X1 U1335 ( .A(mem[1191]), .B(n5598), .Y(n1653) );
  INVX1 U1338 ( .A(n1653), .Y(n3167) );
  AND2X1 U1340 ( .A(mem[1177]), .B(n5599), .Y(n1638) );
  INVX1 U1342 ( .A(n1638), .Y(n3168) );
  AND2X1 U1344 ( .A(mem[1160]), .B(n5599), .Y(n1621) );
  INVX1 U1346 ( .A(n1621), .Y(n3169) );
  AND2X1 U1348 ( .A(mem[1151]), .B(n5599), .Y(n1612) );
  INVX1 U1350 ( .A(n1612), .Y(n3170) );
  AND2X1 U1352 ( .A(mem[1144]), .B(n5600), .Y(n1604) );
  INVX1 U1354 ( .A(n1604), .Y(n3171) );
  AND2X1 U1356 ( .A(mem[1124]), .B(n5600), .Y(n1584) );
  INVX1 U1358 ( .A(n1584), .Y(n3172) );
  AND2X1 U1360 ( .A(mem[1104]), .B(n5601), .Y(n1563) );
  INVX1 U1362 ( .A(n1563), .Y(n3173) );
  AND2X1 U1364 ( .A(mem[1084]), .B(n5601), .Y(n1543) );
  INVX1 U1366 ( .A(n1543), .Y(n3174) );
  AND2X1 U1368 ( .A(mem[1064]), .B(n5602), .Y(n1522) );
  INVX1 U1370 ( .A(n1522), .Y(n3175) );
  AND2X1 U1372 ( .A(mem[1047]), .B(n5602), .Y(n1505) );
  INVX1 U1374 ( .A(n1505), .Y(n3176) );
  AND2X1 U1376 ( .A(mem[1007]), .B(n5603), .Y(n1463) );
  INVX1 U1378 ( .A(n1463), .Y(n3177) );
  AND2X1 U1380 ( .A(mem[983]), .B(n5604), .Y(n1438) );
  INVX1 U1382 ( .A(n1438), .Y(n3178) );
  AND2X1 U1384 ( .A(mem[973]), .B(n5604), .Y(n1428) );
  INVX1 U1386 ( .A(n1428), .Y(n3179) );
  AND2X1 U1388 ( .A(mem[952]), .B(n5604), .Y(n1407) );
  INVX1 U1390 ( .A(n1407), .Y(n3180) );
  AND2X1 U1392 ( .A(mem[933]), .B(n5605), .Y(n1387) );
  INVX1 U1394 ( .A(n1387), .Y(n3181) );
  AND2X1 U1396 ( .A(mem[916]), .B(n5605), .Y(n1370) );
  INVX1 U1398 ( .A(n1370), .Y(n3182) );
  AND2X1 U1400 ( .A(mem[893]), .B(n5606), .Y(n1346) );
  INVX1 U1402 ( .A(n1346), .Y(n3183) );
  AND2X1 U1404 ( .A(mem[876]), .B(n5606), .Y(n1329) );
  INVX1 U1406 ( .A(n1329), .Y(n3184) );
  AND2X1 U1408 ( .A(mem[853]), .B(n5607), .Y(n1305) );
  INVX1 U1410 ( .A(n1305), .Y(n3185) );
  AND2X1 U1412 ( .A(mem[836]), .B(n5607), .Y(n1288) );
  INVX1 U1414 ( .A(n1288), .Y(n3186) );
  AND2X1 U1416 ( .A(mem[804]), .B(n5608), .Y(n1255) );
  INVX1 U1418 ( .A(n1255), .Y(n3187) );
  AND2X1 U1422 ( .A(mem[783]), .B(n5608), .Y(n1234) );
  INVX1 U1424 ( .A(n1234), .Y(n3188) );
  AND2X1 U1426 ( .A(mem[779]), .B(n5608), .Y(n1230) );
  INVX1 U1428 ( .A(n1230), .Y(n3189) );
  AND2X1 U1430 ( .A(mem[765]), .B(n5609), .Y(n1215) );
  INVX1 U1432 ( .A(n1215), .Y(n3190) );
  AND2X1 U1434 ( .A(mem[748]), .B(n5609), .Y(n1198) );
  INVX1 U1436 ( .A(n1198), .Y(n3191) );
  AND2X1 U1438 ( .A(mem[739]), .B(n5609), .Y(n1189) );
  INVX1 U1440 ( .A(n1189), .Y(n3192) );
  AND2X1 U1442 ( .A(mem[725]), .B(n5610), .Y(n1174) );
  INVX1 U1444 ( .A(n1174), .Y(n3193) );
  AND2X1 U1446 ( .A(mem[708]), .B(n5610), .Y(n1157) );
  INVX1 U1448 ( .A(n1157), .Y(n3194) );
  AND2X1 U1450 ( .A(mem[699]), .B(n5610), .Y(n1148) );
  INVX1 U1452 ( .A(n1148), .Y(n3195) );
  AND2X1 U1454 ( .A(mem[685]), .B(n5611), .Y(n1132) );
  INVX1 U1456 ( .A(n1132), .Y(n3196) );
  AND2X1 U1458 ( .A(mem[668]), .B(n5611), .Y(n1115) );
  INVX1 U1460 ( .A(n1115), .Y(n3197) );
  AND2X1 U1462 ( .A(mem[659]), .B(n5611), .Y(n1106) );
  INVX1 U1464 ( .A(n1106), .Y(n3198) );
  AND2X1 U1466 ( .A(mem[652]), .B(n5612), .Y(n1098) );
  INVX1 U1468 ( .A(n1098), .Y(n3199) );
  AND2X1 U1470 ( .A(mem[632]), .B(n5612), .Y(n1078) );
  INVX1 U1472 ( .A(n1078), .Y(n3200) );
  AND2X1 U1474 ( .A(mem[612]), .B(n5613), .Y(n1057) );
  INVX1 U1476 ( .A(n1057), .Y(n3201) );
  AND2X1 U1478 ( .A(mem[592]), .B(n5613), .Y(n1037) );
  INVX1 U1480 ( .A(n1037), .Y(n3202) );
  AND2X1 U1482 ( .A(mem[572]), .B(n5614), .Y(n1016) );
  INVX1 U1484 ( .A(n1016), .Y(n3203) );
  AND2X1 U1486 ( .A(mem[555]), .B(n5614), .Y(n999) );
  INVX1 U1488 ( .A(n999), .Y(n3204) );
  AND2X1 U1490 ( .A(mem[515]), .B(n5615), .Y(n958) );
  INVX1 U1492 ( .A(n958), .Y(n3205) );
  AND2X1 U1494 ( .A(mem[491]), .B(n5616), .Y(n933) );
  INVX1 U1496 ( .A(n933), .Y(n3206) );
  AND2X1 U1498 ( .A(mem[481]), .B(n5616), .Y(n923) );
  INVX1 U1500 ( .A(n923), .Y(n3207) );
  AND2X1 U1502 ( .A(mem[460]), .B(n5616), .Y(n902) );
  INVX1 U1505 ( .A(n902), .Y(n3208) );
  AND2X1 U1507 ( .A(mem[441]), .B(n5617), .Y(n882) );
  INVX1 U1509 ( .A(n882), .Y(n3209) );
  AND2X1 U1511 ( .A(mem[424]), .B(n5617), .Y(n865) );
  INVX1 U1513 ( .A(n865), .Y(n3210) );
  AND2X1 U1515 ( .A(mem[401]), .B(n5618), .Y(n841) );
  INVX1 U1517 ( .A(n841), .Y(n3211) );
  AND2X1 U1519 ( .A(mem[384]), .B(n5618), .Y(n824) );
  INVX1 U1521 ( .A(n824), .Y(n3212) );
  AND2X1 U1523 ( .A(mem[361]), .B(n5619), .Y(n799) );
  INVX1 U1525 ( .A(n799), .Y(n3213) );
  AND2X1 U1527 ( .A(mem[344]), .B(n5619), .Y(n782) );
  INVX1 U1529 ( .A(n782), .Y(n3214) );
  AND2X1 U1531 ( .A(mem[324]), .B(n5620), .Y(n760) );
  INVX1 U1533 ( .A(n760), .Y(n3215) );
  AND2X1 U1535 ( .A(mem[304]), .B(n5620), .Y(n740) );
  INVX1 U1537 ( .A(n740), .Y(n3216) );
  AND2X1 U1539 ( .A(mem[284]), .B(n5621), .Y(n718) );
  INVX1 U1541 ( .A(n718), .Y(n3217) );
  AND2X1 U1543 ( .A(mem[264]), .B(n5621), .Y(n698) );
  INVX1 U1545 ( .A(n698), .Y(n3218) );
  AND2X1 U1547 ( .A(mem[244]), .B(n5622), .Y(n676) );
  INVX1 U1549 ( .A(n676), .Y(n3219) );
  AND2X1 U1551 ( .A(mem[227]), .B(n5622), .Y(n659) );
  INVX1 U1553 ( .A(n659), .Y(n3220) );
  AND2X1 U1555 ( .A(mem[187]), .B(n5623), .Y(n617) );
  INVX1 U1557 ( .A(n617), .Y(n3221) );
  AND2X1 U1559 ( .A(mem[163]), .B(n5624), .Y(n591) );
  INVX1 U1561 ( .A(n591), .Y(n3222) );
  AND2X1 U1563 ( .A(mem[153]), .B(n5624), .Y(n581) );
  INVX1 U1565 ( .A(n581), .Y(n3223) );
  AND2X1 U1567 ( .A(mem[132]), .B(n5624), .Y(n560) );
  INVX1 U1569 ( .A(n560), .Y(n3224) );
  AND2X1 U1571 ( .A(mem[113]), .B(n5625), .Y(n539) );
  INVX1 U1573 ( .A(n539), .Y(n3225) );
  AND2X1 U1575 ( .A(mem[96]), .B(n5625), .Y(n522) );
  INVX1 U1577 ( .A(n522), .Y(n3226) );
  AND2X1 U1579 ( .A(mem[73]), .B(n5626), .Y(n497) );
  INVX1 U1581 ( .A(n497), .Y(n3227) );
  AND2X1 U1583 ( .A(mem[56]), .B(n5626), .Y(n480) );
  INVX1 U1585 ( .A(n480), .Y(n3228) );
  AND2X1 U1588 ( .A(mem[33]), .B(n5627), .Y(n447) );
  INVX1 U1590 ( .A(n447), .Y(n3229) );
  AND2X1 U1592 ( .A(mem[16]), .B(n5627), .Y(n413) );
  INVX1 U1594 ( .A(n413), .Y(n3230) );
  AND2X1 U1596 ( .A(mem[1298]), .B(n5596), .Y(n1762) );
  INVX1 U1598 ( .A(n1762), .Y(n3231) );
  AND2X1 U1600 ( .A(mem[1281]), .B(n5596), .Y(n1745) );
  INVX1 U1602 ( .A(n1745), .Y(n3232) );
  AND2X1 U1604 ( .A(mem[1272]), .B(n5596), .Y(n1736) );
  INVX1 U1606 ( .A(n1736), .Y(n3233) );
  AND2X1 U1608 ( .A(mem[1255]), .B(n5597), .Y(n1718) );
  INVX1 U1610 ( .A(n1718), .Y(n3234) );
  AND2X1 U1612 ( .A(mem[1234]), .B(n5597), .Y(n1697) );
  INVX1 U1614 ( .A(n1697), .Y(n3235) );
  AND2X1 U1616 ( .A(mem[1230]), .B(n5597), .Y(n1693) );
  INVX1 U1618 ( .A(n1693), .Y(n3236) );
  AND2X1 U1620 ( .A(mem[1218]), .B(n5598), .Y(n1680) );
  INVX1 U1622 ( .A(n1680), .Y(n3237) );
  AND2X1 U1624 ( .A(mem[1201]), .B(n5598), .Y(n1663) );
  INVX1 U1626 ( .A(n1663), .Y(n3238) );
  AND2X1 U1628 ( .A(mem[1192]), .B(n5598), .Y(n1654) );
  INVX1 U1630 ( .A(n1654), .Y(n3239) );
  AND2X1 U1632 ( .A(mem[1176]), .B(n5599), .Y(n1637) );
  INVX1 U1634 ( .A(n1637), .Y(n3240) );
  AND2X1 U1636 ( .A(mem[1159]), .B(n5599), .Y(n1620) );
  INVX1 U1638 ( .A(n1620), .Y(n3241) );
  AND2X1 U1640 ( .A(mem[1150]), .B(n5599), .Y(n1611) );
  INVX1 U1642 ( .A(n1611), .Y(n3242) );
  AND2X1 U1644 ( .A(mem[1145]), .B(n5600), .Y(n1605) );
  INVX1 U1646 ( .A(n1605), .Y(n3243) );
  AND2X1 U1648 ( .A(mem[1125]), .B(n5600), .Y(n1585) );
  INVX1 U1650 ( .A(n1585), .Y(n3244) );
  AND2X1 U1652 ( .A(mem[1103]), .B(n5601), .Y(n1562) );
  INVX1 U1654 ( .A(n1562), .Y(n3245) );
  AND2X1 U1656 ( .A(mem[1083]), .B(n5601), .Y(n1542) );
  INVX1 U1658 ( .A(n1542), .Y(n3246) );
  AND2X1 U1660 ( .A(mem[1048]), .B(n5602), .Y(n1506) );
  INVX1 U1662 ( .A(n1506), .Y(n3247) );
  AND2X1 U1664 ( .A(mem[1023]), .B(n5603), .Y(n1479) );
  INVX1 U1666 ( .A(n1479), .Y(n3248) );
  AND2X1 U1668 ( .A(mem[1006]), .B(n5603), .Y(n1462) );
  INVX1 U1671 ( .A(n1462), .Y(n3249) );
  AND2X1 U1673 ( .A(mem[974]), .B(n5604), .Y(n1429) );
  INVX1 U1675 ( .A(n1429), .Y(n3250) );
  AND2X1 U1677 ( .A(mem[957]), .B(n5604), .Y(n1412) );
  INVX1 U1679 ( .A(n1412), .Y(n3251) );
  AND2X1 U1681 ( .A(mem[942]), .B(n5605), .Y(n1396) );
  INVX1 U1683 ( .A(n1396), .Y(n3252) );
  AND2X1 U1685 ( .A(mem[932]), .B(n5605), .Y(n1386) );
  INVX1 U1687 ( .A(n1386), .Y(n3253) );
  AND2X1 U1689 ( .A(mem[911]), .B(n5605), .Y(n1365) );
  INVX1 U1691 ( .A(n1365), .Y(n3254) );
  AND2X1 U1693 ( .A(mem[894]), .B(n5606), .Y(n1347) );
  INVX1 U1695 ( .A(n1347), .Y(n3255) );
  AND2X1 U1697 ( .A(mem[877]), .B(n5606), .Y(n1330) );
  INVX1 U1699 ( .A(n1330), .Y(n3256) );
  AND2X1 U1701 ( .A(mem[852]), .B(n5607), .Y(n1304) );
  INVX1 U1703 ( .A(n1304), .Y(n3257) );
  AND2X1 U1705 ( .A(mem[835]), .B(n5607), .Y(n1287) );
  INVX1 U1707 ( .A(n1287), .Y(n3258) );
  AND2X1 U1709 ( .A(mem[806]), .B(n5608), .Y(n1257) );
  INVX1 U1711 ( .A(n1257), .Y(n3259) );
  AND2X1 U1713 ( .A(mem[789]), .B(n5608), .Y(n1240) );
  INVX1 U1715 ( .A(n1240), .Y(n3260) );
  AND2X1 U1717 ( .A(mem[780]), .B(n5608), .Y(n1231) );
  INVX1 U1719 ( .A(n1231), .Y(n3261) );
  AND2X1 U1721 ( .A(mem[763]), .B(n5609), .Y(n1213) );
  INVX1 U1723 ( .A(n1213), .Y(n3262) );
  AND2X1 U1725 ( .A(mem[742]), .B(n5609), .Y(n1192) );
  INVX1 U1727 ( .A(n1192), .Y(n3263) );
  AND2X1 U1729 ( .A(mem[738]), .B(n5609), .Y(n1188) );
  INVX1 U1731 ( .A(n1188), .Y(n3264) );
  AND2X1 U1733 ( .A(mem[726]), .B(n5610), .Y(n1175) );
  INVX1 U1735 ( .A(n1175), .Y(n3265) );
  AND2X1 U1737 ( .A(mem[709]), .B(n5610), .Y(n1158) );
  INVX1 U1739 ( .A(n1158), .Y(n3266) );
  AND2X1 U1741 ( .A(mem[700]), .B(n5610), .Y(n1149) );
  INVX1 U1743 ( .A(n1149), .Y(n3267) );
  AND2X1 U1745 ( .A(mem[684]), .B(n5611), .Y(n1131) );
  INVX1 U1747 ( .A(n1131), .Y(n3268) );
  AND2X1 U1749 ( .A(mem[667]), .B(n5611), .Y(n1114) );
  INVX1 U1751 ( .A(n1114), .Y(n3269) );
  AND2X1 U1754 ( .A(mem[658]), .B(n5611), .Y(n1105) );
  INVX1 U1756 ( .A(n1105), .Y(n3270) );
  AND2X1 U1758 ( .A(mem[653]), .B(n5612), .Y(n1099) );
  INVX1 U1760 ( .A(n1099), .Y(n3271) );
  AND2X1 U1762 ( .A(mem[633]), .B(n5612), .Y(n1079) );
  INVX1 U1764 ( .A(n1079), .Y(n3272) );
  AND2X1 U1766 ( .A(mem[611]), .B(n5613), .Y(n1056) );
  INVX1 U1768 ( .A(n1056), .Y(n3273) );
  AND2X1 U1770 ( .A(mem[591]), .B(n5613), .Y(n1036) );
  INVX1 U1772 ( .A(n1036), .Y(n3274) );
  AND2X1 U1774 ( .A(mem[556]), .B(n5614), .Y(n1000) );
  INVX1 U1776 ( .A(n1000), .Y(n3275) );
  AND2X1 U1778 ( .A(mem[531]), .B(n5615), .Y(n974) );
  INVX1 U1780 ( .A(n974), .Y(n3276) );
  AND2X1 U1782 ( .A(mem[514]), .B(n5615), .Y(n957) );
  INVX1 U1784 ( .A(n957), .Y(n3277) );
  AND2X1 U1786 ( .A(mem[482]), .B(n5616), .Y(n924) );
  INVX1 U1788 ( .A(n924), .Y(n3278) );
  AND2X1 U1790 ( .A(mem[465]), .B(n5616), .Y(n907) );
  INVX1 U1792 ( .A(n907), .Y(n3279) );
  AND2X1 U1794 ( .A(mem[450]), .B(n5617), .Y(n891) );
  INVX1 U1796 ( .A(n891), .Y(n3280) );
  AND2X1 U1798 ( .A(mem[440]), .B(n5617), .Y(n881) );
  INVX1 U1800 ( .A(n881), .Y(n3281) );
  AND2X1 U1802 ( .A(mem[419]), .B(n5617), .Y(n860) );
  INVX1 U1804 ( .A(n860), .Y(n3282) );
  AND2X1 U1806 ( .A(mem[402]), .B(n5618), .Y(n842) );
  INVX1 U1808 ( .A(n842), .Y(n3283) );
  AND2X1 U1810 ( .A(mem[385]), .B(n5618), .Y(n825) );
  INVX1 U1812 ( .A(n825), .Y(n3284) );
  AND2X1 U1814 ( .A(mem[360]), .B(n5619), .Y(n798) );
  INVX1 U1816 ( .A(n798), .Y(n3285) );
  AND2X1 U1818 ( .A(mem[343]), .B(n5619), .Y(n781) );
  INVX1 U1820 ( .A(n781), .Y(n3286) );
  AND2X1 U1822 ( .A(mem[325]), .B(n5620), .Y(n761) );
  INVX1 U1824 ( .A(n761), .Y(n3287) );
  AND2X1 U1826 ( .A(mem[305]), .B(n5620), .Y(n741) );
  INVX1 U1828 ( .A(n741), .Y(n3288) );
  AND2X1 U1830 ( .A(mem[283]), .B(n5621), .Y(n717) );
  INVX1 U1832 ( .A(n717), .Y(n3289) );
  AND2X1 U1834 ( .A(mem[263]), .B(n5621), .Y(n697) );
  INVX1 U1837 ( .A(n697), .Y(n3290) );
  AND2X1 U1839 ( .A(mem[228]), .B(n5622), .Y(n660) );
  INVX1 U1841 ( .A(n660), .Y(n3291) );
  AND2X1 U1843 ( .A(mem[203]), .B(n5623), .Y(n633) );
  INVX1 U1845 ( .A(n633), .Y(n3292) );
  AND2X1 U1847 ( .A(mem[186]), .B(n5623), .Y(n616) );
  INVX1 U1849 ( .A(n616), .Y(n3293) );
  AND2X1 U1851 ( .A(mem[154]), .B(n5624), .Y(n582) );
  INVX1 U1853 ( .A(n582), .Y(n3294) );
  AND2X1 U1855 ( .A(mem[137]), .B(n5624), .Y(n565) );
  INVX1 U1857 ( .A(n565), .Y(n3295) );
  AND2X1 U1859 ( .A(mem[122]), .B(n5625), .Y(n548) );
  INVX1 U1861 ( .A(n548), .Y(n3296) );
  AND2X1 U1863 ( .A(mem[112]), .B(n5625), .Y(n538) );
  INVX1 U1865 ( .A(n538), .Y(n3297) );
  AND2X1 U1867 ( .A(mem[91]), .B(n5625), .Y(n517) );
  INVX1 U1869 ( .A(n517), .Y(n3298) );
  AND2X1 U1871 ( .A(mem[74]), .B(n5626), .Y(n498) );
  INVX1 U1873 ( .A(n498), .Y(n3299) );
  AND2X1 U1875 ( .A(mem[57]), .B(n5626), .Y(n481) );
  INVX1 U1877 ( .A(n481), .Y(n3300) );
  AND2X1 U1879 ( .A(mem[32]), .B(n5627), .Y(n445) );
  INVX1 U1881 ( .A(n445), .Y(n3301) );
  AND2X1 U1883 ( .A(mem[15]), .B(n5627), .Y(n411) );
  INVX1 U1885 ( .A(n411), .Y(n3302) );
  AND2X1 U1887 ( .A(mem[1299]), .B(n5596), .Y(n1763) );
  INVX1 U1889 ( .A(n1763), .Y(n3303) );
  AND2X1 U1891 ( .A(mem[1282]), .B(n5596), .Y(n1746) );
  INVX1 U1893 ( .A(n1746), .Y(n3304) );
  AND2X1 U1895 ( .A(mem[1273]), .B(n5596), .Y(n1737) );
  INVX1 U1897 ( .A(n1737), .Y(n3305) );
  AND2X1 U1899 ( .A(mem[1259]), .B(n5597), .Y(n1722) );
  INVX1 U1901 ( .A(n1722), .Y(n3306) );
  AND2X1 U1903 ( .A(mem[1242]), .B(n5597), .Y(n1705) );
  INVX1 U1905 ( .A(n1705), .Y(n3307) );
  AND2X1 U1907 ( .A(mem[1233]), .B(n5597), .Y(n1696) );
  INVX1 U1909 ( .A(n1696), .Y(n3308) );
  AND2X1 U1911 ( .A(mem[1214]), .B(n5598), .Y(n1676) );
  INVX1 U1913 ( .A(n1676), .Y(n3309) );
  AND2X1 U1915 ( .A(mem[1193]), .B(n5598), .Y(n1655) );
  INVX1 U1917 ( .A(n1655), .Y(n3310) );
  AND2X1 U1920 ( .A(mem[1189]), .B(n5598), .Y(n1651) );
  INVX1 U1922 ( .A(n1651), .Y(n3311) );
  AND2X1 U1924 ( .A(mem[1175]), .B(n5599), .Y(n1636) );
  INVX1 U1926 ( .A(n1636), .Y(n3312) );
  AND2X1 U1928 ( .A(mem[1158]), .B(n5599), .Y(n1619) );
  INVX1 U1930 ( .A(n1619), .Y(n3313) );
  AND2X1 U1932 ( .A(mem[1149]), .B(n5599), .Y(n1610) );
  INVX1 U1934 ( .A(n1610), .Y(n3314) );
  AND2X1 U1936 ( .A(mem[1146]), .B(n5600), .Y(n1606) );
  INVX1 U1938 ( .A(n1606), .Y(n3315) );
  AND2X1 U1940 ( .A(mem[1129]), .B(n5600), .Y(n1589) );
  INVX1 U1942 ( .A(n1589), .Y(n3316) );
  AND2X1 U1944 ( .A(mem[1089]), .B(n5601), .Y(n1548) );
  INVX1 U1946 ( .A(n1548), .Y(n3317) );
  AND2X1 U1948 ( .A(mem[1062]), .B(n5602), .Y(n1520) );
  INVX1 U1950 ( .A(n1520), .Y(n3318) );
  AND2X1 U1952 ( .A(mem[1042]), .B(n5602), .Y(n1500) );
  INVX1 U1954 ( .A(n1500), .Y(n3319) );
  AND2X1 U1956 ( .A(mem[1022]), .B(n5603), .Y(n1478) );
  INVX1 U1958 ( .A(n1478), .Y(n3320) );
  AND2X1 U1960 ( .A(mem[1002]), .B(n5603), .Y(n1458) );
  INVX1 U1962 ( .A(n1458), .Y(n3321) );
  AND2X1 U1964 ( .A(mem[975]), .B(n5604), .Y(n1430) );
  INVX1 U1966 ( .A(n1430), .Y(n3322) );
  AND2X1 U1968 ( .A(mem[958]), .B(n5604), .Y(n1413) );
  INVX1 U1970 ( .A(n1413), .Y(n3323) );
  AND2X1 U1972 ( .A(mem[935]), .B(n5605), .Y(n1389) );
  INVX1 U1974 ( .A(n1389), .Y(n3324) );
  AND2X1 U1976 ( .A(mem[918]), .B(n5605), .Y(n1372) );
  INVX1 U1978 ( .A(n1372), .Y(n3325) );
  AND2X1 U1980 ( .A(mem[901]), .B(n5606), .Y(n1354) );
  INVX1 U1982 ( .A(n1354), .Y(n3326) );
  AND2X1 U1984 ( .A(mem[891]), .B(n5606), .Y(n1344) );
  INVX1 U1986 ( .A(n1344), .Y(n3327) );
  AND2X1 U1988 ( .A(mem[870]), .B(n5606), .Y(n1323) );
  INVX1 U1990 ( .A(n1323), .Y(n3328) );
  AND2X1 U1992 ( .A(mem[851]), .B(n5607), .Y(n1303) );
  INVX1 U1994 ( .A(n1303), .Y(n3329) );
  AND2X1 U1996 ( .A(mem[834]), .B(n5607), .Y(n1286) );
  INVX1 U1998 ( .A(n1286), .Y(n3330) );
  AND2X1 U2000 ( .A(mem[807]), .B(n5608), .Y(n1258) );
  INVX1 U2003 ( .A(n1258), .Y(n3331) );
  AND2X1 U2005 ( .A(mem[790]), .B(n5608), .Y(n1241) );
  INVX1 U2007 ( .A(n1241), .Y(n3332) );
  AND2X1 U2009 ( .A(mem[781]), .B(n5608), .Y(n1232) );
  INVX1 U2011 ( .A(n1232), .Y(n3333) );
  AND2X1 U2013 ( .A(mem[767]), .B(n5609), .Y(n1217) );
  INVX1 U2015 ( .A(n1217), .Y(n3334) );
  AND2X1 U2017 ( .A(mem[750]), .B(n5609), .Y(n1200) );
  INVX1 U2019 ( .A(n1200), .Y(n3335) );
  AND2X1 U2021 ( .A(mem[741]), .B(n5609), .Y(n1191) );
  INVX1 U2023 ( .A(n1191), .Y(n3336) );
  AND2X1 U2025 ( .A(mem[722]), .B(n5610), .Y(n1171) );
  INVX1 U2027 ( .A(n1171), .Y(n3337) );
  AND2X1 U2029 ( .A(mem[701]), .B(n5610), .Y(n1150) );
  INVX1 U2031 ( .A(n1150), .Y(n3338) );
  AND2X1 U2033 ( .A(mem[697]), .B(n5610), .Y(n1146) );
  INVX1 U2035 ( .A(n1146), .Y(n3339) );
  AND2X1 U2037 ( .A(mem[683]), .B(n5611), .Y(n1130) );
  INVX1 U2039 ( .A(n1130), .Y(n3340) );
  AND2X1 U2041 ( .A(mem[666]), .B(n5611), .Y(n1113) );
  INVX1 U2043 ( .A(n1113), .Y(n3341) );
  AND2X1 U2045 ( .A(mem[657]), .B(n5611), .Y(n1104) );
  INVX1 U2047 ( .A(n1104), .Y(n3342) );
  AND2X1 U2049 ( .A(mem[654]), .B(n5612), .Y(n1100) );
  INVX1 U2051 ( .A(n1100), .Y(n3343) );
  AND2X1 U2053 ( .A(mem[637]), .B(n5612), .Y(n1083) );
  INVX1 U2055 ( .A(n1083), .Y(n3344) );
  AND2X1 U2057 ( .A(mem[597]), .B(n5613), .Y(n1042) );
  INVX1 U2059 ( .A(n1042), .Y(n3345) );
  AND2X1 U2061 ( .A(mem[570]), .B(n5614), .Y(n1014) );
  INVX1 U2063 ( .A(n1014), .Y(n3346) );
  AND2X1 U2065 ( .A(mem[550]), .B(n5614), .Y(n994) );
  INVX1 U2067 ( .A(n994), .Y(n3347) );
  AND2X1 U2069 ( .A(mem[530]), .B(n5615), .Y(n973) );
  INVX1 U2071 ( .A(n973), .Y(n3348) );
  AND2X1 U2073 ( .A(mem[510]), .B(n5615), .Y(n953) );
  INVX1 U2075 ( .A(n953), .Y(n3349) );
  AND2X1 U2077 ( .A(mem[483]), .B(n5616), .Y(n925) );
  INVX1 U2079 ( .A(n925), .Y(n3350) );
  AND2X1 U2081 ( .A(mem[466]), .B(n5616), .Y(n908) );
  INVX1 U2083 ( .A(n908), .Y(n3351) );
  AND2X1 U2087 ( .A(mem[443]), .B(n5617), .Y(n884) );
  INVX1 U2089 ( .A(n884), .Y(n3352) );
  AND2X1 U2091 ( .A(mem[426]), .B(n5617), .Y(n867) );
  INVX1 U2093 ( .A(n867), .Y(n3353) );
  AND2X1 U2095 ( .A(mem[409]), .B(n5618), .Y(n849) );
  INVX1 U2097 ( .A(n849), .Y(n3354) );
  AND2X1 U2099 ( .A(mem[399]), .B(n5618), .Y(n839) );
  INVX1 U2101 ( .A(n839), .Y(n3355) );
  AND2X1 U2103 ( .A(mem[378]), .B(n5618), .Y(n818) );
  INVX1 U2105 ( .A(n818), .Y(n3356) );
  AND2X1 U2107 ( .A(mem[359]), .B(n5619), .Y(n797) );
  INVX1 U2109 ( .A(n797), .Y(n3357) );
  AND2X1 U2111 ( .A(mem[342]), .B(n5619), .Y(n780) );
  INVX1 U2113 ( .A(n780), .Y(n3358) );
  AND2X1 U2115 ( .A(mem[326]), .B(n5620), .Y(n762) );
  INVX1 U2117 ( .A(n762), .Y(n3359) );
  AND2X1 U2119 ( .A(mem[309]), .B(n5620), .Y(n745) );
  INVX1 U2121 ( .A(n745), .Y(n3360) );
  AND2X1 U2123 ( .A(mem[269]), .B(n5621), .Y(n703) );
  INVX1 U2125 ( .A(n703), .Y(n3361) );
  AND2X1 U2127 ( .A(mem[242]), .B(n5622), .Y(n674) );
  INVX1 U2129 ( .A(n674), .Y(n3362) );
  AND2X1 U2131 ( .A(mem[222]), .B(n5622), .Y(n654) );
  INVX1 U2133 ( .A(n654), .Y(n3363) );
  AND2X1 U2135 ( .A(mem[202]), .B(n5623), .Y(n632) );
  INVX1 U2137 ( .A(n632), .Y(n3364) );
  AND2X1 U2139 ( .A(mem[182]), .B(n5623), .Y(n612) );
  INVX1 U2141 ( .A(n612), .Y(n3365) );
  AND2X1 U2143 ( .A(mem[155]), .B(n5624), .Y(n583) );
  INVX1 U2145 ( .A(n583), .Y(n3366) );
  AND2X1 U2147 ( .A(mem[138]), .B(n5624), .Y(n566) );
  INVX1 U2149 ( .A(n566), .Y(n3367) );
  AND2X1 U2151 ( .A(mem[115]), .B(n5625), .Y(n541) );
  INVX1 U2153 ( .A(n541), .Y(n3368) );
  AND2X1 U2155 ( .A(mem[98]), .B(n5625), .Y(n524) );
  INVX1 U2157 ( .A(n524), .Y(n3369) );
  AND2X1 U2159 ( .A(mem[81]), .B(n5626), .Y(n505) );
  INVX1 U2161 ( .A(n505), .Y(n3370) );
  AND2X1 U2163 ( .A(mem[71]), .B(n5626), .Y(n495) );
  INVX1 U2165 ( .A(n495), .Y(n3371) );
  AND2X1 U2167 ( .A(mem[50]), .B(n5626), .Y(n474) );
  INVX1 U2171 ( .A(n474), .Y(n3372) );
  AND2X1 U2173 ( .A(mem[31]), .B(n5627), .Y(n443) );
  INVX1 U2175 ( .A(n443), .Y(n3373) );
  AND2X1 U2177 ( .A(mem[14]), .B(n5627), .Y(n409) );
  INVX1 U2179 ( .A(n409), .Y(n3374) );
  AND2X1 U2181 ( .A(n5716), .B(n1780), .Y(n1833) );
  INVX1 U2183 ( .A(n1833), .Y(n3375) );
  AND2X1 U2185 ( .A(mem[1300]), .B(n5596), .Y(n1764) );
  INVX1 U2187 ( .A(n1764), .Y(n3376) );
  AND2X1 U2189 ( .A(mem[1283]), .B(n5596), .Y(n1747) );
  INVX1 U2191 ( .A(n1747), .Y(n3377) );
  AND2X1 U2193 ( .A(mem[1274]), .B(n5596), .Y(n1738) );
  INVX1 U2195 ( .A(n1738), .Y(n3378) );
  AND2X1 U2197 ( .A(mem[1258]), .B(n5597), .Y(n1721) );
  INVX1 U2199 ( .A(n1721), .Y(n3379) );
  AND2X1 U2201 ( .A(mem[1241]), .B(n5597), .Y(n1704) );
  INVX1 U2203 ( .A(n1704), .Y(n3380) );
  AND2X1 U2205 ( .A(mem[1232]), .B(n5597), .Y(n1695) );
  INVX1 U2207 ( .A(n1695), .Y(n3381) );
  AND2X1 U2209 ( .A(mem[1216]), .B(n5598), .Y(n1678) );
  INVX1 U2211 ( .A(n1678), .Y(n3382) );
  AND2X1 U2213 ( .A(mem[1199]), .B(n5598), .Y(n1661) );
  INVX1 U2215 ( .A(n1661), .Y(n3383) );
  AND2X1 U2217 ( .A(mem[1190]), .B(n5598), .Y(n1652) );
  INVX1 U2219 ( .A(n1652), .Y(n3384) );
  AND2X1 U2221 ( .A(mem[1173]), .B(n5599), .Y(n1634) );
  INVX1 U2223 ( .A(n1634), .Y(n3385) );
  AND2X1 U2225 ( .A(mem[1152]), .B(n5599), .Y(n1613) );
  INVX1 U2227 ( .A(n1613), .Y(n3386) );
  AND2X1 U2229 ( .A(mem[1148]), .B(n5599), .Y(n1609) );
  INVX1 U2231 ( .A(n1609), .Y(n3387) );
  AND2X1 U2233 ( .A(mem[1130]), .B(n5600), .Y(n1590) );
  INVX1 U2235 ( .A(n1590), .Y(n3388) );
  AND2X1 U2237 ( .A(mem[1105]), .B(n5601), .Y(n1564) );
  INVX1 U2239 ( .A(n1564), .Y(n3389) );
  AND2X1 U2241 ( .A(mem[1088]), .B(n5601), .Y(n1547) );
  INVX1 U2243 ( .A(n1547), .Y(n3390) );
  AND2X1 U2245 ( .A(mem[1063]), .B(n5602), .Y(n1521) );
  INVX1 U2247 ( .A(n1521), .Y(n3391) );
  AND2X1 U2249 ( .A(mem[1043]), .B(n5602), .Y(n1501) );
  INVX1 U2251 ( .A(n1501), .Y(n3392) );
  AND2X1 U2255 ( .A(mem[1021]), .B(n5603), .Y(n1477) );
  INVX1 U2257 ( .A(n1477), .Y(n3393) );
  AND2X1 U2259 ( .A(mem[1001]), .B(n5603), .Y(n1457) );
  INVX1 U2261 ( .A(n1457), .Y(n3394) );
  AND2X1 U2263 ( .A(mem[976]), .B(n5604), .Y(n1431) );
  INVX1 U2265 ( .A(n1431), .Y(n3395) );
  AND2X1 U2267 ( .A(mem[959]), .B(n5604), .Y(n1414) );
  INVX1 U2269 ( .A(n1414), .Y(n3396) );
  AND2X1 U2271 ( .A(mem[934]), .B(n5605), .Y(n1388) );
  INVX1 U2273 ( .A(n1388), .Y(n3397) );
  AND2X1 U2275 ( .A(mem[917]), .B(n5605), .Y(n1371) );
  INVX1 U2277 ( .A(n1371), .Y(n3398) );
  AND2X1 U2279 ( .A(mem[892]), .B(n5606), .Y(n1345) );
  INVX1 U2281 ( .A(n1345), .Y(n3399) );
  AND2X1 U2283 ( .A(mem[875]), .B(n5606), .Y(n1328) );
  INVX1 U2285 ( .A(n1328), .Y(n3400) );
  AND2X1 U2287 ( .A(mem[860]), .B(n5607), .Y(n1312) );
  INVX1 U2289 ( .A(n1312), .Y(n3401) );
  AND2X1 U2291 ( .A(mem[850]), .B(n5607), .Y(n1302) );
  INVX1 U2293 ( .A(n1302), .Y(n3402) );
  AND2X1 U2295 ( .A(mem[829]), .B(n5607), .Y(n1281) );
  INVX1 U2297 ( .A(n1281), .Y(n3403) );
  AND2X1 U2299 ( .A(mem[808]), .B(n5608), .Y(n1259) );
  INVX1 U2301 ( .A(n1259), .Y(n3404) );
  AND2X1 U2303 ( .A(mem[791]), .B(n5608), .Y(n1242) );
  INVX1 U2305 ( .A(n1242), .Y(n3405) );
  AND2X1 U2307 ( .A(mem[782]), .B(n5608), .Y(n1233) );
  INVX1 U2309 ( .A(n1233), .Y(n3406) );
  AND2X1 U2311 ( .A(mem[766]), .B(n5609), .Y(n1216) );
  INVX1 U2313 ( .A(n1216), .Y(n3407) );
  AND2X1 U2315 ( .A(mem[749]), .B(n5609), .Y(n1199) );
  INVX1 U2317 ( .A(n1199), .Y(n3408) );
  AND2X1 U2319 ( .A(mem[740]), .B(n5609), .Y(n1190) );
  INVX1 U2321 ( .A(n1190), .Y(n3409) );
  AND2X1 U2323 ( .A(mem[724]), .B(n5610), .Y(n1173) );
  INVX1 U2325 ( .A(n1173), .Y(n3410) );
  AND2X1 U2327 ( .A(mem[707]), .B(n5610), .Y(n1156) );
  INVX1 U2329 ( .A(n1156), .Y(n3411) );
  AND2X1 U2331 ( .A(mem[698]), .B(n5610), .Y(n1147) );
  INVX1 U2333 ( .A(n1147), .Y(n3412) );
  AND2X1 U2335 ( .A(mem[681]), .B(n5611), .Y(n1128) );
  INVX1 U2339 ( .A(n1128), .Y(n3413) );
  AND2X1 U2341 ( .A(mem[660]), .B(n5611), .Y(n1107) );
  INVX1 U2343 ( .A(n1107), .Y(n3414) );
  AND2X1 U2345 ( .A(mem[656]), .B(n5611), .Y(n1103) );
  INVX1 U2347 ( .A(n1103), .Y(n3415) );
  AND2X1 U2349 ( .A(mem[638]), .B(n5612), .Y(n1084) );
  INVX1 U2351 ( .A(n1084), .Y(n3416) );
  AND2X1 U2353 ( .A(mem[613]), .B(n5613), .Y(n1058) );
  INVX1 U2355 ( .A(n1058), .Y(n3417) );
  AND2X1 U2357 ( .A(mem[596]), .B(n5613), .Y(n1041) );
  INVX1 U2359 ( .A(n1041), .Y(n3418) );
  AND2X1 U2361 ( .A(mem[571]), .B(n5614), .Y(n1015) );
  INVX1 U2363 ( .A(n1015), .Y(n3419) );
  AND2X1 U2365 ( .A(mem[551]), .B(n5614), .Y(n995) );
  INVX1 U2367 ( .A(n995), .Y(n3420) );
  AND2X1 U2369 ( .A(mem[529]), .B(n5615), .Y(n972) );
  INVX1 U2371 ( .A(n972), .Y(n3421) );
  AND2X1 U2373 ( .A(mem[509]), .B(n5615), .Y(n952) );
  INVX1 U2375 ( .A(n952), .Y(n3422) );
  AND2X1 U2377 ( .A(mem[484]), .B(n5616), .Y(n926) );
  INVX1 U2379 ( .A(n926), .Y(n3423) );
  AND2X1 U2381 ( .A(mem[467]), .B(n5616), .Y(n909) );
  INVX1 U2383 ( .A(n909), .Y(n3424) );
  AND2X1 U2385 ( .A(mem[442]), .B(n5617), .Y(n883) );
  INVX1 U2387 ( .A(n883), .Y(n3425) );
  AND2X1 U2389 ( .A(mem[425]), .B(n5617), .Y(n866) );
  INVX1 U2391 ( .A(n866), .Y(n3426) );
  AND2X1 U2393 ( .A(mem[400]), .B(n5618), .Y(n840) );
  INVX1 U2395 ( .A(n840), .Y(n3427) );
  AND2X1 U2397 ( .A(mem[383]), .B(n5618), .Y(n823) );
  INVX1 U2399 ( .A(n823), .Y(n3428) );
  AND2X1 U2401 ( .A(mem[368]), .B(n5619), .Y(n806) );
  INVX1 U2403 ( .A(n806), .Y(n3429) );
  AND2X1 U2405 ( .A(mem[358]), .B(n5619), .Y(n796) );
  INVX1 U2407 ( .A(n796), .Y(n3430) );
  AND2X1 U2409 ( .A(mem[337]), .B(n5619), .Y(n775) );
  INVX1 U2411 ( .A(n775), .Y(n3431) );
  AND2X1 U2413 ( .A(mem[310]), .B(n5620), .Y(n746) );
  INVX1 U2415 ( .A(n746), .Y(n3432) );
  AND2X1 U2417 ( .A(mem[285]), .B(n5621), .Y(n719) );
  INVX1 U2419 ( .A(n719), .Y(n3433) );
  AND2X1 U2423 ( .A(mem[268]), .B(n5621), .Y(n702) );
  INVX1 U2425 ( .A(n702), .Y(n3434) );
  AND2X1 U2427 ( .A(mem[243]), .B(n5622), .Y(n675) );
  INVX1 U2429 ( .A(n675), .Y(n3435) );
  AND2X1 U2431 ( .A(mem[223]), .B(n5622), .Y(n655) );
  INVX1 U2433 ( .A(n655), .Y(n3436) );
  AND2X1 U2435 ( .A(mem[201]), .B(n5623), .Y(n631) );
  INVX1 U2437 ( .A(n631), .Y(n3437) );
  AND2X1 U2439 ( .A(mem[181]), .B(n5623), .Y(n611) );
  INVX1 U2441 ( .A(n611), .Y(n3438) );
  AND2X1 U2443 ( .A(mem[156]), .B(n5624), .Y(n584) );
  INVX1 U2445 ( .A(n584), .Y(n3439) );
  AND2X1 U2447 ( .A(mem[139]), .B(n5624), .Y(n567) );
  INVX1 U2449 ( .A(n567), .Y(n3440) );
  AND2X1 U2451 ( .A(mem[114]), .B(n5625), .Y(n540) );
  INVX1 U2453 ( .A(n540), .Y(n3441) );
  AND2X1 U2455 ( .A(mem[97]), .B(n5625), .Y(n523) );
  INVX1 U2457 ( .A(n523), .Y(n3442) );
  AND2X1 U2459 ( .A(mem[72]), .B(n5626), .Y(n496) );
  INVX1 U2461 ( .A(n496), .Y(n3443) );
  AND2X1 U2463 ( .A(mem[55]), .B(n5626), .Y(n479) );
  INVX1 U2465 ( .A(n479), .Y(n3444) );
  AND2X1 U2467 ( .A(mem[40]), .B(n5627), .Y(n461) );
  INVX1 U2469 ( .A(n461), .Y(n3445) );
  AND2X1 U2471 ( .A(mem[30]), .B(n5627), .Y(n441) );
  INVX1 U2473 ( .A(n441), .Y(n3446) );
  AND2X1 U2475 ( .A(mem[9]), .B(n5627), .Y(n399) );
  INVX1 U2477 ( .A(n399), .Y(n3447) );
  AND2X1 U2479 ( .A(mem[1308]), .B(n5596), .Y(n1772) );
  INVX1 U2481 ( .A(n1772), .Y(n3448) );
  AND2X1 U2483 ( .A(mem[1288]), .B(n5596), .Y(n1752) );
  INVX1 U2485 ( .A(n1752), .Y(n3449) );
  AND2X1 U2487 ( .A(mem[1268]), .B(n5597), .Y(n1731) );
  INVX1 U2489 ( .A(n1731), .Y(n3450) );
  AND2X1 U2491 ( .A(mem[1248]), .B(n5597), .Y(n1711) );
  INVX1 U2493 ( .A(n1711), .Y(n3451) );
  AND2X1 U2495 ( .A(mem[1228]), .B(n5598), .Y(n1690) );
  INVX1 U2497 ( .A(n1690), .Y(n3452) );
  AND2X1 U2499 ( .A(mem[1211]), .B(n5598), .Y(n1673) );
  INVX1 U2501 ( .A(n1673), .Y(n3453) );
  AND2X1 U2503 ( .A(mem[1171]), .B(n5599), .Y(n1632) );
  INVX1 U2507 ( .A(n1632), .Y(n3454) );
  AND2X1 U2509 ( .A(mem[1132]), .B(n5600), .Y(n1592) );
  INVX1 U2511 ( .A(n1592), .Y(n3455) );
  AND2X1 U2513 ( .A(mem[1111]), .B(n5600), .Y(n1571) );
  INVX1 U2515 ( .A(n1571), .Y(n3456) );
  AND2X1 U2517 ( .A(mem[1107]), .B(n5600), .Y(n1567) );
  INVX1 U2519 ( .A(n1567), .Y(n3457) );
  AND2X1 U2521 ( .A(mem[1093]), .B(n5601), .Y(n1552) );
  INVX1 U2523 ( .A(n1552), .Y(n3458) );
  AND2X1 U2525 ( .A(mem[1076]), .B(n5601), .Y(n1535) );
  INVX1 U2527 ( .A(n1535), .Y(n3459) );
  AND2X1 U2529 ( .A(mem[1067]), .B(n5601), .Y(n1526) );
  INVX1 U2531 ( .A(n1526), .Y(n3460) );
  AND2X1 U2533 ( .A(mem[1053]), .B(n5602), .Y(n1511) );
  INVX1 U2535 ( .A(n1511), .Y(n3461) );
  AND2X1 U2537 ( .A(mem[1036]), .B(n5602), .Y(n1494) );
  INVX1 U2539 ( .A(n1494), .Y(n3462) );
  AND2X1 U2541 ( .A(mem[1027]), .B(n5602), .Y(n1485) );
  INVX1 U2543 ( .A(n1485), .Y(n3463) );
  AND2X1 U2545 ( .A(mem[1013]), .B(n5603), .Y(n1469) );
  INVX1 U2547 ( .A(n1469), .Y(n3464) );
  AND2X1 U2549 ( .A(mem[996]), .B(n5603), .Y(n1452) );
  INVX1 U2551 ( .A(n1452), .Y(n3465) );
  AND2X1 U2553 ( .A(mem[987]), .B(n5603), .Y(n1443) );
  INVX1 U2555 ( .A(n1443), .Y(n3466) );
  AND2X1 U2557 ( .A(mem[977]), .B(n5604), .Y(n1432) );
  INVX1 U2559 ( .A(n1432), .Y(n3467) );
  AND2X1 U2561 ( .A(mem[962]), .B(n5604), .Y(n1417) );
  INVX1 U2563 ( .A(n1417), .Y(n3468) );
  AND2X1 U2565 ( .A(mem[948]), .B(n5604), .Y(n1403) );
  INVX1 U2567 ( .A(n1403), .Y(n3469) );
  AND2X1 U2569 ( .A(mem[937]), .B(n5605), .Y(n1391) );
  INVX1 U2571 ( .A(n1391), .Y(n3470) );
  AND2X1 U2573 ( .A(mem[922]), .B(n5605), .Y(n1376) );
  INVX1 U2575 ( .A(n1376), .Y(n3471) );
  AND2X1 U2577 ( .A(mem[908]), .B(n5605), .Y(n1362) );
  INVX1 U2579 ( .A(n1362), .Y(n3472) );
  AND2X1 U2581 ( .A(mem[897]), .B(n5606), .Y(n1350) );
  INVX1 U2583 ( .A(n1350), .Y(n3473) );
  AND2X1 U2585 ( .A(mem[882]), .B(n5606), .Y(n1335) );
  INVX1 U2587 ( .A(n1335), .Y(n3474) );
  AND2X1 U2591 ( .A(mem[868]), .B(n5606), .Y(n1321) );
  INVX1 U2593 ( .A(n1321), .Y(n3475) );
  AND2X1 U2595 ( .A(mem[846]), .B(n5607), .Y(n1298) );
  INVX1 U2597 ( .A(n1298), .Y(n3476) );
  AND2X1 U2599 ( .A(mem[833]), .B(n5607), .Y(n1285) );
  INVX1 U2601 ( .A(n1285), .Y(n3477) );
  AND2X1 U2603 ( .A(mem[828]), .B(n5607), .Y(n1280) );
  INVX1 U2605 ( .A(n1280), .Y(n3478) );
  AND2X1 U2607 ( .A(mem[816]), .B(n5608), .Y(n1267) );
  INVX1 U2609 ( .A(n1267), .Y(n3479) );
  AND2X1 U2611 ( .A(mem[796]), .B(n5608), .Y(n1247) );
  INVX1 U2613 ( .A(n1247), .Y(n3480) );
  AND2X1 U2615 ( .A(mem[776]), .B(n5609), .Y(n1226) );
  INVX1 U2617 ( .A(n1226), .Y(n3481) );
  AND2X1 U2619 ( .A(mem[756]), .B(n5609), .Y(n1206) );
  INVX1 U2621 ( .A(n1206), .Y(n3482) );
  AND2X1 U2623 ( .A(mem[736]), .B(n5610), .Y(n1185) );
  INVX1 U2625 ( .A(n1185), .Y(n3483) );
  AND2X1 U2627 ( .A(mem[719]), .B(n5610), .Y(n1168) );
  INVX1 U2629 ( .A(n1168), .Y(n3484) );
  AND2X1 U2631 ( .A(mem[679]), .B(n5611), .Y(n1126) );
  INVX1 U2633 ( .A(n1126), .Y(n3485) );
  AND2X1 U2635 ( .A(mem[640]), .B(n5612), .Y(n1086) );
  INVX1 U2637 ( .A(n1086), .Y(n3486) );
  AND2X1 U2639 ( .A(mem[619]), .B(n5612), .Y(n1065) );
  INVX1 U2641 ( .A(n1065), .Y(n3487) );
  AND2X1 U2643 ( .A(mem[615]), .B(n5612), .Y(n1061) );
  INVX1 U2645 ( .A(n1061), .Y(n3488) );
  AND2X1 U2647 ( .A(mem[601]), .B(n5613), .Y(n1046) );
  INVX1 U2649 ( .A(n1046), .Y(n3489) );
  AND2X1 U2651 ( .A(mem[584]), .B(n5613), .Y(n1029) );
  INVX1 U2653 ( .A(n1029), .Y(n3490) );
  AND2X1 U2655 ( .A(mem[575]), .B(n5613), .Y(n1020) );
  INVX1 U2657 ( .A(n1020), .Y(n3491) );
  AND2X1 U2659 ( .A(mem[561]), .B(n5614), .Y(n1005) );
  INVX1 U2661 ( .A(n1005), .Y(n3492) );
  AND2X1 U2663 ( .A(mem[544]), .B(n5614), .Y(n988) );
  INVX1 U2665 ( .A(n988), .Y(n3493) );
  AND2X1 U2667 ( .A(mem[535]), .B(n5614), .Y(n979) );
  INVX1 U2669 ( .A(n979), .Y(n3494) );
  AND2X1 U2671 ( .A(mem[521]), .B(n5615), .Y(n964) );
  INVX1 U2675 ( .A(n964), .Y(n3495) );
  AND2X1 U2676 ( .A(mem[504]), .B(n5615), .Y(n947) );
  INVX1 U2678 ( .A(n947), .Y(n3496) );
  AND2X1 U2679 ( .A(mem[495]), .B(n5615), .Y(n938) );
  INVX1 U2681 ( .A(n938), .Y(n3497) );
  AND2X1 U2682 ( .A(mem[485]), .B(n5616), .Y(n927) );
  INVX1 U2684 ( .A(n927), .Y(n3498) );
  AND2X1 U2685 ( .A(mem[470]), .B(n5616), .Y(n912) );
  INVX1 U2687 ( .A(n912), .Y(n3499) );
  AND2X1 U2688 ( .A(mem[456]), .B(n5616), .Y(n898) );
  INVX1 U2690 ( .A(n898), .Y(n3500) );
  AND2X1 U2691 ( .A(mem[445]), .B(n5617), .Y(n886) );
  INVX1 U2693 ( .A(n886), .Y(n3501) );
  AND2X1 U2694 ( .A(mem[430]), .B(n5617), .Y(n871) );
  INVX1 U2696 ( .A(n871), .Y(n3502) );
  AND2X1 U2697 ( .A(mem[416]), .B(n5617), .Y(n857) );
  INVX1 U2699 ( .A(n857), .Y(n3503) );
  AND2X1 U2700 ( .A(mem[405]), .B(n5618), .Y(n845) );
  INVX1 U2702 ( .A(n845), .Y(n3504) );
  AND2X1 U2703 ( .A(mem[390]), .B(n5618), .Y(n830) );
  INVX1 U2705 ( .A(n830), .Y(n3505) );
  AND2X1 U2706 ( .A(mem[376]), .B(n5618), .Y(n816) );
  INVX1 U2708 ( .A(n816), .Y(n3506) );
  AND2X1 U2709 ( .A(mem[354]), .B(n5619), .Y(n792) );
  INVX1 U2711 ( .A(n792), .Y(n3507) );
  AND2X1 U2712 ( .A(mem[341]), .B(n5619), .Y(n779) );
  INVX1 U2714 ( .A(n779), .Y(n3508) );
  AND2X1 U2715 ( .A(mem[336]), .B(n5619), .Y(n774) );
  INVX1 U2717 ( .A(n774), .Y(n3509) );
  AND2X1 U2718 ( .A(mem[312]), .B(n5620), .Y(n748) );
  INVX1 U2720 ( .A(n748), .Y(n3510) );
  AND2X1 U2721 ( .A(mem[291]), .B(n5620), .Y(n727) );
  INVX1 U2723 ( .A(n727), .Y(n3511) );
  AND2X1 U2724 ( .A(mem[287]), .B(n5620), .Y(n723) );
  INVX1 U2726 ( .A(n723), .Y(n3512) );
  AND2X1 U2727 ( .A(mem[273]), .B(n5621), .Y(n707) );
  INVX1 U2729 ( .A(n707), .Y(n3513) );
  AND2X1 U2730 ( .A(mem[256]), .B(n5621), .Y(n690) );
  INVX1 U2732 ( .A(n690), .Y(n3514) );
  AND2X1 U2733 ( .A(mem[247]), .B(n5621), .Y(n681) );
  INVX1 U2735 ( .A(n681), .Y(n3515) );
  AND2X1 U2736 ( .A(mem[233]), .B(n5622), .Y(n665) );
  INVX1 U2738 ( .A(n665), .Y(n3516) );
  AND2X1 U2739 ( .A(mem[216]), .B(n5622), .Y(n648) );
  INVX1 U2741 ( .A(n648), .Y(n3517) );
  AND2X1 U2742 ( .A(mem[207]), .B(n5622), .Y(n639) );
  INVX1 U2744 ( .A(n639), .Y(n3518) );
  AND2X1 U2745 ( .A(mem[193]), .B(n5623), .Y(n623) );
  INVX1 U2747 ( .A(n623), .Y(n3519) );
  AND2X1 U2748 ( .A(mem[176]), .B(n5623), .Y(n606) );
  INVX1 U2750 ( .A(n606), .Y(n3520) );
  AND2X1 U2751 ( .A(mem[167]), .B(n5623), .Y(n597) );
  INVX1 U2753 ( .A(n597), .Y(n3521) );
  AND2X1 U2754 ( .A(mem[157]), .B(n5624), .Y(n585) );
  INVX1 U2756 ( .A(n585), .Y(n3522) );
  AND2X1 U2757 ( .A(mem[142]), .B(n5624), .Y(n570) );
  INVX1 U2759 ( .A(n570), .Y(n3523) );
  AND2X1 U2760 ( .A(mem[128]), .B(n5624), .Y(n556) );
  INVX1 U2762 ( .A(n556), .Y(n3524) );
  AND2X1 U2763 ( .A(mem[117]), .B(n5625), .Y(n543) );
  INVX1 U2765 ( .A(n543), .Y(n3525) );
  AND2X1 U2766 ( .A(mem[102]), .B(n5625), .Y(n528) );
  INVX1 U2768 ( .A(n528), .Y(n3526) );
  AND2X1 U2769 ( .A(mem[88]), .B(n5625), .Y(n514) );
  INVX1 U2771 ( .A(n514), .Y(n3527) );
  AND2X1 U2772 ( .A(mem[77]), .B(n5626), .Y(n501) );
  INVX1 U2774 ( .A(n501), .Y(n3528) );
  AND2X1 U2775 ( .A(mem[62]), .B(n5626), .Y(n486) );
  INVX1 U2777 ( .A(n486), .Y(n3529) );
  AND2X1 U2778 ( .A(mem[48]), .B(n5626), .Y(n472) );
  INVX1 U2780 ( .A(n472), .Y(n3530) );
  AND2X1 U2781 ( .A(mem[26]), .B(n5627), .Y(n433) );
  INVX1 U2783 ( .A(n433), .Y(n3531) );
  AND2X1 U2784 ( .A(mem[13]), .B(n5627), .Y(n407) );
  INVX1 U2786 ( .A(n407), .Y(n3532) );
  AND2X1 U2787 ( .A(mem[8]), .B(n5627), .Y(n397) );
  INVX1 U2789 ( .A(n397), .Y(n3533) );
  BUFX2 U2790 ( .A(n636), .Y(n3534) );
  BUFX2 U2792 ( .A(n593), .Y(n3535) );
  AND2X1 U2793 ( .A(n23), .B(n1780), .Y(n1783) );
  INVX1 U2795 ( .A(n1783), .Y(n3536) );
  AND2X1 U2796 ( .A(mem[1309]), .B(n5596), .Y(n1773) );
  INVX1 U2801 ( .A(n1773), .Y(n3537) );
  AND2X1 U2803 ( .A(mem[1289]), .B(n5596), .Y(n1753) );
  INVX1 U2805 ( .A(n1753), .Y(n3538) );
  AND2X1 U2807 ( .A(mem[1267]), .B(n5597), .Y(n1730) );
  INVX1 U2809 ( .A(n1730), .Y(n3539) );
  AND2X1 U2811 ( .A(mem[1247]), .B(n5597), .Y(n1710) );
  INVX1 U2813 ( .A(n1710), .Y(n3540) );
  AND2X1 U2815 ( .A(mem[1212]), .B(n5598), .Y(n1674) );
  INVX1 U2817 ( .A(n1674), .Y(n3541) );
  AND2X1 U2859 ( .A(mem[1187]), .B(n5599), .Y(n1648) );
  INVX1 U2860 ( .A(n1648), .Y(n3542) );
  AND2X1 U2862 ( .A(mem[1170]), .B(n5599), .Y(n1631) );
  INVX1 U2863 ( .A(n1631), .Y(n3543) );
  AND2X1 U2864 ( .A(mem[1134]), .B(n5600), .Y(n1594) );
  INVX1 U2867 ( .A(n1594), .Y(n3544) );
  AND2X1 U2875 ( .A(mem[1117]), .B(n5600), .Y(n1577) );
  INVX1 U2876 ( .A(n1577), .Y(n3545) );
  AND2X1 U2877 ( .A(mem[1108]), .B(n5600), .Y(n1568) );
  INVX1 U2878 ( .A(n1568), .Y(n3546) );
  AND2X1 U2879 ( .A(mem[1091]), .B(n5601), .Y(n1550) );
  INVX1 U2880 ( .A(n1550), .Y(n3547) );
  AND2X1 U2881 ( .A(mem[1070]), .B(n5601), .Y(n1529) );
  INVX1 U2882 ( .A(n1529), .Y(n3548) );
  AND2X1 U2883 ( .A(mem[1066]), .B(n5601), .Y(n1525) );
  INVX1 U2884 ( .A(n1525), .Y(n3549) );
  AND2X1 U2885 ( .A(mem[1054]), .B(n5602), .Y(n1512) );
  INVX1 U2886 ( .A(n1512), .Y(n3550) );
  AND2X1 U2887 ( .A(mem[1037]), .B(n5602), .Y(n1495) );
  INVX1 U2888 ( .A(n1495), .Y(n3551) );
  AND2X1 U2889 ( .A(mem[1028]), .B(n5602), .Y(n1486) );
  INVX1 U2890 ( .A(n1486), .Y(n3552) );
  AND2X1 U2891 ( .A(mem[1012]), .B(n5603), .Y(n1468) );
  INVX1 U2892 ( .A(n1468), .Y(n3553) );
  AND2X1 U2893 ( .A(mem[995]), .B(n5603), .Y(n1451) );
  INVX1 U2894 ( .A(n1451), .Y(n3554) );
  AND2X1 U2895 ( .A(mem[986]), .B(n5603), .Y(n1442) );
  INVX1 U2896 ( .A(n1442), .Y(n3555) );
  AND2X1 U2897 ( .A(mem[978]), .B(n5604), .Y(n1433) );
  INVX1 U2898 ( .A(n1433), .Y(n3556) );
  AND2X1 U2899 ( .A(mem[963]), .B(n5604), .Y(n1418) );
  INVX1 U2900 ( .A(n1418), .Y(n3557) );
  AND2X1 U2901 ( .A(mem[949]), .B(n5604), .Y(n1404) );
  INVX1 U2902 ( .A(n1404), .Y(n3558) );
  AND2X1 U2903 ( .A(mem[936]), .B(n5605), .Y(n1390) );
  INVX1 U2904 ( .A(n1390), .Y(n3559) );
  AND2X1 U2905 ( .A(mem[921]), .B(n5605), .Y(n1375) );
  INVX1 U2906 ( .A(n1375), .Y(n3560) );
  AND2X1 U2907 ( .A(mem[907]), .B(n5605), .Y(n1361) );
  INVX1 U2908 ( .A(n1361), .Y(n3561) );
  AND2X1 U2909 ( .A(mem[887]), .B(n5606), .Y(n1340) );
  INVX1 U2910 ( .A(n1340), .Y(n3562) );
  AND2X1 U2911 ( .A(mem[874]), .B(n5606), .Y(n1327) );
  INVX1 U2912 ( .A(n1327), .Y(n3563) );
  AND2X1 U2913 ( .A(mem[869]), .B(n5606), .Y(n1322) );
  INVX1 U2914 ( .A(n1322), .Y(n3564) );
  AND2X1 U2915 ( .A(mem[856]), .B(n5607), .Y(n1308) );
  INVX1 U2916 ( .A(n1308), .Y(n3565) );
  AND2X1 U2917 ( .A(mem[841]), .B(n5607), .Y(n1293) );
  INVX1 U2918 ( .A(n1293), .Y(n3566) );
  AND2X1 U2919 ( .A(mem[827]), .B(n5607), .Y(n1279) );
  INVX1 U2920 ( .A(n1279), .Y(n3567) );
  AND2X1 U2921 ( .A(mem[817]), .B(n5608), .Y(n1268) );
  INVX1 U2922 ( .A(n1268), .Y(n3568) );
  AND2X1 U2923 ( .A(mem[797]), .B(n5608), .Y(n1248) );
  INVX1 U2924 ( .A(n1248), .Y(n3569) );
  AND2X1 U2925 ( .A(mem[775]), .B(n5609), .Y(n1225) );
  INVX1 U2926 ( .A(n1225), .Y(n3570) );
  AND2X1 U2927 ( .A(mem[755]), .B(n5609), .Y(n1205) );
  INVX1 U2928 ( .A(n1205), .Y(n3571) );
  AND2X1 U2929 ( .A(mem[720]), .B(n5610), .Y(n1169) );
  INVX1 U2930 ( .A(n1169), .Y(n3572) );
  AND2X1 U2931 ( .A(mem[695]), .B(n5611), .Y(n1142) );
  INVX1 U2932 ( .A(n1142), .Y(n3573) );
  AND2X1 U2933 ( .A(mem[678]), .B(n5611), .Y(n1125) );
  INVX1 U2934 ( .A(n1125), .Y(n3574) );
  AND2X1 U2935 ( .A(mem[642]), .B(n5612), .Y(n1088) );
  INVX1 U2936 ( .A(n1088), .Y(n3575) );
  AND2X1 U2937 ( .A(mem[625]), .B(n5612), .Y(n1071) );
  INVX1 U2938 ( .A(n1071), .Y(n3576) );
  AND2X1 U2939 ( .A(mem[616]), .B(n5612), .Y(n1062) );
  INVX1 U2940 ( .A(n1062), .Y(n3577) );
  AND2X1 U2941 ( .A(mem[599]), .B(n5613), .Y(n1044) );
  INVX1 U2942 ( .A(n1044), .Y(n3578) );
  AND2X1 U2943 ( .A(mem[578]), .B(n5613), .Y(n1023) );
  INVX1 U2944 ( .A(n1023), .Y(n3579) );
  AND2X1 U2945 ( .A(mem[574]), .B(n5613), .Y(n1019) );
  INVX1 U2946 ( .A(n1019), .Y(n3580) );
  AND2X1 U2947 ( .A(mem[562]), .B(n5614), .Y(n1006) );
  INVX1 U2948 ( .A(n1006), .Y(n3581) );
  AND2X1 U2949 ( .A(mem[545]), .B(n5614), .Y(n989) );
  INVX1 U2950 ( .A(n989), .Y(n3582) );
  AND2X1 U2951 ( .A(mem[536]), .B(n5614), .Y(n980) );
  INVX1 U2952 ( .A(n980), .Y(n3583) );
  AND2X1 U2953 ( .A(mem[520]), .B(n5615), .Y(n963) );
  INVX1 U2954 ( .A(n963), .Y(n3584) );
  AND2X1 U2955 ( .A(mem[503]), .B(n5615), .Y(n946) );
  INVX1 U2956 ( .A(n946), .Y(n3585) );
  AND2X1 U2957 ( .A(mem[494]), .B(n5615), .Y(n937) );
  INVX1 U2958 ( .A(n937), .Y(n3586) );
  AND2X1 U2959 ( .A(mem[486]), .B(n5616), .Y(n928) );
  INVX1 U2960 ( .A(n928), .Y(n3587) );
  AND2X1 U2961 ( .A(mem[471]), .B(n5616), .Y(n913) );
  INVX1 U2962 ( .A(n913), .Y(n3588) );
  AND2X1 U2963 ( .A(mem[457]), .B(n5616), .Y(n899) );
  INVX1 U2964 ( .A(n899), .Y(n3589) );
  AND2X1 U2965 ( .A(mem[444]), .B(n5617), .Y(n885) );
  INVX1 U2966 ( .A(n885), .Y(n3590) );
  AND2X1 U2967 ( .A(mem[429]), .B(n5617), .Y(n870) );
  INVX1 U2968 ( .A(n870), .Y(n3591) );
  AND2X1 U2969 ( .A(mem[415]), .B(n5617), .Y(n856) );
  INVX1 U2970 ( .A(n856), .Y(n3592) );
  AND2X1 U2971 ( .A(mem[395]), .B(n5618), .Y(n835) );
  INVX1 U2972 ( .A(n835), .Y(n3593) );
  AND2X1 U2973 ( .A(mem[382]), .B(n5618), .Y(n822) );
  INVX1 U2974 ( .A(n822), .Y(n3594) );
  AND2X1 U2975 ( .A(mem[377]), .B(n5618), .Y(n817) );
  INVX1 U2976 ( .A(n817), .Y(n3595) );
  AND2X1 U2977 ( .A(mem[364]), .B(n5619), .Y(n802) );
  INVX1 U2978 ( .A(n802), .Y(n3596) );
  AND2X1 U2979 ( .A(mem[349]), .B(n5619), .Y(n787) );
  INVX1 U2980 ( .A(n787), .Y(n3597) );
  AND2X1 U2981 ( .A(mem[335]), .B(n5619), .Y(n773) );
  INVX1 U2982 ( .A(n773), .Y(n3598) );
  AND2X1 U2983 ( .A(mem[314]), .B(n5620), .Y(n750) );
  INVX1 U2984 ( .A(n750), .Y(n3599) );
  AND2X1 U2985 ( .A(mem[297]), .B(n5620), .Y(n733) );
  INVX1 U2986 ( .A(n733), .Y(n3600) );
  AND2X1 U2987 ( .A(mem[288]), .B(n5620), .Y(n724) );
  INVX1 U2988 ( .A(n724), .Y(n3601) );
  AND2X1 U2989 ( .A(mem[271]), .B(n5621), .Y(n705) );
  INVX1 U2990 ( .A(n705), .Y(n3602) );
  AND2X1 U2991 ( .A(mem[250]), .B(n5621), .Y(n684) );
  INVX1 U2992 ( .A(n684), .Y(n3603) );
  AND2X1 U2993 ( .A(mem[246]), .B(n5621), .Y(n680) );
  INVX1 U2994 ( .A(n680), .Y(n3604) );
  AND2X1 U2995 ( .A(mem[234]), .B(n5622), .Y(n666) );
  INVX1 U2996 ( .A(n666), .Y(n3605) );
  AND2X1 U2997 ( .A(mem[217]), .B(n5622), .Y(n649) );
  INVX1 U2998 ( .A(n649), .Y(n3606) );
  AND2X1 U2999 ( .A(mem[208]), .B(n5622), .Y(n640) );
  INVX1 U3000 ( .A(n640), .Y(n3607) );
  AND2X1 U3001 ( .A(mem[192]), .B(n5623), .Y(n622) );
  INVX1 U3002 ( .A(n622), .Y(n3608) );
  AND2X1 U3003 ( .A(mem[175]), .B(n5623), .Y(n605) );
  INVX1 U3004 ( .A(n605), .Y(n3609) );
  AND2X1 U3005 ( .A(mem[166]), .B(n5623), .Y(n596) );
  INVX1 U3006 ( .A(n596), .Y(n3610) );
  AND2X1 U3007 ( .A(mem[158]), .B(n5624), .Y(n586) );
  INVX1 U3008 ( .A(n586), .Y(n3611) );
  AND2X1 U3009 ( .A(mem[143]), .B(n5624), .Y(n571) );
  INVX1 U3010 ( .A(n571), .Y(n3612) );
  AND2X1 U3011 ( .A(mem[129]), .B(n5624), .Y(n557) );
  INVX1 U3012 ( .A(n557), .Y(n3613) );
  AND2X1 U3013 ( .A(mem[116]), .B(n5625), .Y(n542) );
  INVX1 U3014 ( .A(n542), .Y(n3614) );
  AND2X1 U3015 ( .A(mem[101]), .B(n5625), .Y(n527) );
  INVX1 U3016 ( .A(n527), .Y(n3615) );
  AND2X1 U3017 ( .A(mem[87]), .B(n5625), .Y(n513) );
  INVX1 U3018 ( .A(n513), .Y(n3616) );
  AND2X1 U3019 ( .A(mem[67]), .B(n5626), .Y(n491) );
  INVX1 U3020 ( .A(n491), .Y(n3617) );
  AND2X1 U3021 ( .A(mem[54]), .B(n5626), .Y(n478) );
  INVX1 U3022 ( .A(n478), .Y(n3618) );
  AND2X1 U3023 ( .A(mem[49]), .B(n5626), .Y(n473) );
  INVX1 U3024 ( .A(n473), .Y(n3619) );
  AND2X1 U3025 ( .A(mem[36]), .B(n5627), .Y(n453) );
  INVX1 U3026 ( .A(n453), .Y(n3620) );
  AND2X1 U3027 ( .A(mem[21]), .B(n5627), .Y(n423) );
  INVX1 U3028 ( .A(n423), .Y(n3621) );
  AND2X1 U3029 ( .A(mem[7]), .B(n5627), .Y(n395) );
  INVX1 U3030 ( .A(n395), .Y(n3622) );
  BUFX2 U3031 ( .A(n679), .Y(n3623) );
  BUFX2 U3032 ( .A(n550), .Y(n3624) );
  AND2X1 U3033 ( .A(n101), .B(n1786), .Y(n1790) );
  INVX1 U3034 ( .A(n1790), .Y(n3625) );
  AND2X1 U3035 ( .A(n22), .B(n1780), .Y(n1779) );
  INVX1 U3036 ( .A(n1779), .Y(n3626) );
  AND2X1 U3037 ( .A(mem[1310]), .B(n5596), .Y(n1774) );
  INVX1 U3038 ( .A(n1774), .Y(n3627) );
  AND2X1 U3039 ( .A(mem[1293]), .B(n5596), .Y(n1757) );
  INVX1 U3040 ( .A(n1757), .Y(n3628) );
  AND2X1 U3041 ( .A(mem[1253]), .B(n5597), .Y(n1716) );
  INVX1 U3042 ( .A(n1716), .Y(n3629) );
  AND2X1 U3043 ( .A(mem[1226]), .B(n5598), .Y(n1688) );
  INVX1 U3044 ( .A(n1688), .Y(n3630) );
  AND2X1 U3045 ( .A(mem[1206]), .B(n5598), .Y(n1668) );
  INVX1 U3046 ( .A(n1668), .Y(n3631) );
  AND2X1 U3047 ( .A(mem[1186]), .B(n5599), .Y(n1647) );
  INVX1 U3048 ( .A(n1647), .Y(n3632) );
  AND2X1 U3049 ( .A(mem[1166]), .B(n5599), .Y(n1627) );
  INVX1 U3050 ( .A(n1627), .Y(n3633) );
  AND2X1 U3051 ( .A(mem[1135]), .B(n5600), .Y(n1595) );
  INVX1 U3052 ( .A(n1595), .Y(n3634) );
  AND2X1 U3053 ( .A(mem[1118]), .B(n5600), .Y(n1578) );
  INVX1 U3054 ( .A(n1578), .Y(n3635) );
  AND2X1 U3055 ( .A(mem[1109]), .B(n5600), .Y(n1569) );
  INVX1 U3056 ( .A(n1569), .Y(n3636) );
  AND2X1 U3057 ( .A(mem[1095]), .B(n5601), .Y(n1554) );
  INVX1 U3058 ( .A(n1554), .Y(n3637) );
  AND2X1 U3059 ( .A(mem[1078]), .B(n5601), .Y(n1537) );
  INVX1 U3060 ( .A(n1537), .Y(n3638) );
  AND2X1 U3061 ( .A(mem[1069]), .B(n5601), .Y(n1528) );
  INVX1 U3062 ( .A(n1528), .Y(n3639) );
  AND2X1 U3063 ( .A(mem[1050]), .B(n5602), .Y(n1508) );
  INVX1 U3064 ( .A(n1508), .Y(n3640) );
  AND2X1 U3065 ( .A(mem[1029]), .B(n5602), .Y(n1487) );
  INVX1 U3066 ( .A(n1487), .Y(n3641) );
  AND2X1 U3067 ( .A(mem[1025]), .B(n5602), .Y(n1483) );
  INVX1 U3068 ( .A(n1483), .Y(n3642) );
  AND2X1 U3069 ( .A(mem[1011]), .B(n5603), .Y(n1467) );
  INVX1 U3070 ( .A(n1467), .Y(n3643) );
  AND2X1 U3071 ( .A(mem[994]), .B(n5603), .Y(n1450) );
  INVX1 U3072 ( .A(n1450), .Y(n3644) );
  AND2X1 U3073 ( .A(mem[985]), .B(n5603), .Y(n1441) );
  INVX1 U3074 ( .A(n1441), .Y(n3645) );
  AND2X1 U3075 ( .A(mem[979]), .B(n5604), .Y(n1434) );
  INVX1 U3076 ( .A(n1434), .Y(n3646) );
  AND2X1 U3077 ( .A(mem[964]), .B(n5604), .Y(n1419) );
  INVX1 U3078 ( .A(n1419), .Y(n3647) );
  AND2X1 U3079 ( .A(mem[950]), .B(n5604), .Y(n1405) );
  INVX1 U3080 ( .A(n1405), .Y(n3648) );
  AND2X1 U3081 ( .A(mem[928]), .B(n5605), .Y(n1382) );
  INVX1 U3082 ( .A(n1382), .Y(n3649) );
  AND2X1 U3083 ( .A(mem[915]), .B(n5605), .Y(n1369) );
  INVX1 U3084 ( .A(n1369), .Y(n3650) );
  AND2X1 U3085 ( .A(mem[910]), .B(n5605), .Y(n1364) );
  INVX1 U3086 ( .A(n1364), .Y(n3651) );
  AND2X1 U3087 ( .A(mem[895]), .B(n5606), .Y(n1348) );
  INVX1 U3088 ( .A(n1348), .Y(n3652) );
  AND2X1 U3089 ( .A(mem[880]), .B(n5606), .Y(n1333) );
  INVX1 U3090 ( .A(n1333), .Y(n3653) );
  AND2X1 U3091 ( .A(mem[866]), .B(n5606), .Y(n1319) );
  INVX1 U3092 ( .A(n1319), .Y(n3654) );
  AND2X1 U3093 ( .A(mem[855]), .B(n5607), .Y(n1307) );
  INVX1 U3094 ( .A(n1307), .Y(n3655) );
  AND2X1 U3095 ( .A(mem[840]), .B(n5607), .Y(n1292) );
  INVX1 U3096 ( .A(n1292), .Y(n3656) );
  AND2X1 U3097 ( .A(mem[826]), .B(n5607), .Y(n1278) );
  INVX1 U3098 ( .A(n1278), .Y(n3657) );
  AND2X1 U3099 ( .A(mem[818]), .B(n5608), .Y(n1269) );
  INVX1 U3100 ( .A(n1269), .Y(n3658) );
  AND2X1 U3101 ( .A(mem[801]), .B(n5608), .Y(n1252) );
  INVX1 U3102 ( .A(n1252), .Y(n3659) );
  AND2X1 U3103 ( .A(mem[761]), .B(n5609), .Y(n1211) );
  INVX1 U3104 ( .A(n1211), .Y(n3660) );
  AND2X1 U3105 ( .A(mem[734]), .B(n5610), .Y(n1183) );
  INVX1 U3106 ( .A(n1183), .Y(n3661) );
  AND2X1 U3107 ( .A(mem[714]), .B(n5610), .Y(n1163) );
  INVX1 U3108 ( .A(n1163), .Y(n3662) );
  AND2X1 U3109 ( .A(mem[694]), .B(n5611), .Y(n1141) );
  INVX1 U3110 ( .A(n1141), .Y(n3663) );
  AND2X1 U3111 ( .A(mem[674]), .B(n5611), .Y(n1121) );
  INVX1 U3112 ( .A(n1121), .Y(n3664) );
  AND2X1 U3113 ( .A(mem[643]), .B(n5612), .Y(n1089) );
  INVX1 U3114 ( .A(n1089), .Y(n3665) );
  AND2X1 U3115 ( .A(mem[626]), .B(n5612), .Y(n1072) );
  INVX1 U3116 ( .A(n1072), .Y(n3666) );
  AND2X1 U3117 ( .A(mem[617]), .B(n5612), .Y(n1063) );
  INVX1 U3118 ( .A(n1063), .Y(n3667) );
  AND2X1 U3119 ( .A(mem[603]), .B(n5613), .Y(n1048) );
  INVX1 U3120 ( .A(n1048), .Y(n3668) );
  AND2X1 U3121 ( .A(mem[586]), .B(n5613), .Y(n1031) );
  INVX1 U3122 ( .A(n1031), .Y(n3669) );
  AND2X1 U3123 ( .A(mem[577]), .B(n5613), .Y(n1022) );
  INVX1 U3124 ( .A(n1022), .Y(n3670) );
  AND2X1 U3125 ( .A(mem[558]), .B(n5614), .Y(n1002) );
  INVX1 U3126 ( .A(n1002), .Y(n3671) );
  AND2X1 U3127 ( .A(mem[537]), .B(n5614), .Y(n981) );
  INVX1 U3128 ( .A(n981), .Y(n3672) );
  AND2X1 U3129 ( .A(mem[533]), .B(n5614), .Y(n977) );
  INVX1 U3130 ( .A(n977), .Y(n3673) );
  AND2X1 U3131 ( .A(mem[519]), .B(n5615), .Y(n962) );
  INVX1 U3132 ( .A(n962), .Y(n3674) );
  AND2X1 U3133 ( .A(mem[502]), .B(n5615), .Y(n945) );
  INVX1 U3134 ( .A(n945), .Y(n3675) );
  AND2X1 U3135 ( .A(mem[493]), .B(n5615), .Y(n936) );
  INVX1 U3136 ( .A(n936), .Y(n3676) );
  AND2X1 U3137 ( .A(mem[487]), .B(n5616), .Y(n929) );
  INVX1 U3138 ( .A(n929), .Y(n3677) );
  AND2X1 U3139 ( .A(mem[472]), .B(n5616), .Y(n914) );
  INVX1 U3140 ( .A(n914), .Y(n3678) );
  AND2X1 U3141 ( .A(mem[458]), .B(n5616), .Y(n900) );
  INVX1 U3142 ( .A(n900), .Y(n3679) );
  AND2X1 U3143 ( .A(mem[436]), .B(n5617), .Y(n877) );
  INVX1 U3144 ( .A(n877), .Y(n3680) );
  AND2X1 U3145 ( .A(mem[423]), .B(n5617), .Y(n864) );
  INVX1 U3146 ( .A(n864), .Y(n3681) );
  AND2X1 U3147 ( .A(mem[418]), .B(n5617), .Y(n859) );
  INVX1 U3148 ( .A(n859), .Y(n3682) );
  AND2X1 U3149 ( .A(mem[403]), .B(n5618), .Y(n843) );
  INVX1 U3150 ( .A(n843), .Y(n3683) );
  AND2X1 U3151 ( .A(mem[388]), .B(n5618), .Y(n828) );
  INVX1 U3152 ( .A(n828), .Y(n3684) );
  AND2X1 U3153 ( .A(mem[374]), .B(n5618), .Y(n814) );
  INVX1 U3154 ( .A(n814), .Y(n3685) );
  AND2X1 U3155 ( .A(mem[363]), .B(n5619), .Y(n801) );
  INVX1 U3156 ( .A(n801), .Y(n3686) );
  AND2X1 U3157 ( .A(mem[348]), .B(n5619), .Y(n786) );
  INVX1 U3158 ( .A(n786), .Y(n3687) );
  AND2X1 U3159 ( .A(mem[334]), .B(n5619), .Y(n772) );
  INVX1 U3160 ( .A(n772), .Y(n3688) );
  AND2X1 U3161 ( .A(mem[315]), .B(n5620), .Y(n751) );
  INVX1 U3162 ( .A(n751), .Y(n3689) );
  AND2X1 U3163 ( .A(mem[298]), .B(n5620), .Y(n734) );
  INVX1 U3164 ( .A(n734), .Y(n3690) );
  AND2X1 U3165 ( .A(mem[289]), .B(n5620), .Y(n725) );
  INVX1 U3166 ( .A(n725), .Y(n3691) );
  AND2X1 U3167 ( .A(mem[275]), .B(n5621), .Y(n709) );
  INVX1 U3168 ( .A(n709), .Y(n3692) );
  AND2X1 U3169 ( .A(mem[258]), .B(n5621), .Y(n692) );
  INVX1 U3170 ( .A(n692), .Y(n3693) );
  AND2X1 U3171 ( .A(mem[249]), .B(n5621), .Y(n683) );
  INVX1 U3172 ( .A(n683), .Y(n3694) );
  AND2X1 U3173 ( .A(mem[230]), .B(n5622), .Y(n662) );
  INVX1 U3174 ( .A(n662), .Y(n3695) );
  AND2X1 U3175 ( .A(mem[209]), .B(n5622), .Y(n641) );
  INVX1 U3176 ( .A(n641), .Y(n3696) );
  AND2X1 U3177 ( .A(mem[205]), .B(n5622), .Y(n637) );
  INVX1 U3178 ( .A(n637), .Y(n3697) );
  AND2X1 U3179 ( .A(mem[191]), .B(n5623), .Y(n621) );
  INVX1 U3180 ( .A(n621), .Y(n3698) );
  AND2X1 U3181 ( .A(mem[174]), .B(n5623), .Y(n604) );
  INVX1 U3182 ( .A(n604), .Y(n3699) );
  AND2X1 U3183 ( .A(mem[165]), .B(n5623), .Y(n595) );
  INVX1 U3184 ( .A(n595), .Y(n3700) );
  AND2X1 U3185 ( .A(mem[159]), .B(n5624), .Y(n587) );
  INVX1 U3186 ( .A(n587), .Y(n3701) );
  AND2X1 U3187 ( .A(mem[144]), .B(n5624), .Y(n572) );
  INVX1 U3188 ( .A(n572), .Y(n3702) );
  AND2X1 U3189 ( .A(mem[130]), .B(n5624), .Y(n558) );
  INVX1 U3190 ( .A(n558), .Y(n3703) );
  AND2X1 U3191 ( .A(mem[108]), .B(n5625), .Y(n534) );
  INVX1 U3192 ( .A(n534), .Y(n3704) );
  AND2X1 U3193 ( .A(mem[95]), .B(n5625), .Y(n521) );
  INVX1 U3194 ( .A(n521), .Y(n3705) );
  AND2X1 U3195 ( .A(mem[90]), .B(n5625), .Y(n516) );
  INVX1 U3196 ( .A(n516), .Y(n3706) );
  AND2X1 U3197 ( .A(mem[75]), .B(n5626), .Y(n499) );
  INVX1 U3198 ( .A(n499), .Y(n3707) );
  AND2X1 U3199 ( .A(mem[60]), .B(n5626), .Y(n484) );
  INVX1 U3200 ( .A(n484), .Y(n3708) );
  AND2X1 U3201 ( .A(mem[46]), .B(n5626), .Y(n470) );
  INVX1 U3202 ( .A(n470), .Y(n3709) );
  AND2X1 U3203 ( .A(mem[35]), .B(n5627), .Y(n451) );
  INVX1 U3204 ( .A(n451), .Y(n3710) );
  AND2X1 U3205 ( .A(mem[20]), .B(n5627), .Y(n421) );
  INVX1 U3206 ( .A(n421), .Y(n3711) );
  AND2X1 U3207 ( .A(mem[6]), .B(n5627), .Y(n393) );
  INVX1 U3208 ( .A(n393), .Y(n3712) );
  BUFX2 U3209 ( .A(n722), .Y(n3713) );
  BUFX2 U3210 ( .A(n507), .Y(n3714) );
  AND2X1 U3211 ( .A(n5674), .B(n1786), .Y(n1789) );
  INVX1 U3212 ( .A(n1789), .Y(n3715) );
  AND2X1 U3213 ( .A(mem[1294]), .B(n5596), .Y(n1758) );
  INVX1 U3214 ( .A(n1758), .Y(n3716) );
  AND2X1 U3215 ( .A(mem[1269]), .B(n5597), .Y(n1732) );
  INVX1 U3216 ( .A(n1732), .Y(n3717) );
  AND2X1 U3217 ( .A(mem[1252]), .B(n5597), .Y(n1715) );
  INVX1 U3218 ( .A(n1715), .Y(n3718) );
  AND2X1 U3219 ( .A(mem[1227]), .B(n5598), .Y(n1689) );
  INVX1 U3220 ( .A(n1689), .Y(n3719) );
  AND2X1 U3221 ( .A(mem[1207]), .B(n5598), .Y(n1669) );
  INVX1 U3222 ( .A(n1669), .Y(n3720) );
  AND2X1 U3223 ( .A(mem[1185]), .B(n5599), .Y(n1646) );
  INVX1 U3224 ( .A(n1646), .Y(n3721) );
  AND2X1 U3225 ( .A(mem[1165]), .B(n5599), .Y(n1626) );
  INVX1 U3226 ( .A(n1626), .Y(n3722) );
  AND2X1 U3227 ( .A(mem[1136]), .B(n5600), .Y(n1596) );
  INVX1 U3228 ( .A(n1596), .Y(n3723) );
  AND2X1 U3229 ( .A(mem[1119]), .B(n5600), .Y(n1579) );
  INVX1 U3230 ( .A(n1579), .Y(n3724) );
  AND2X1 U3231 ( .A(mem[1110]), .B(n5600), .Y(n1570) );
  INVX1 U3232 ( .A(n1570), .Y(n3725) );
  AND2X1 U3233 ( .A(mem[1094]), .B(n5601), .Y(n1553) );
  INVX1 U3234 ( .A(n1553), .Y(n3726) );
  AND2X1 U3235 ( .A(mem[1077]), .B(n5601), .Y(n1536) );
  INVX1 U3236 ( .A(n1536), .Y(n3727) );
  AND2X1 U3237 ( .A(mem[1068]), .B(n5601), .Y(n1527) );
  INVX1 U3238 ( .A(n1527), .Y(n3728) );
  AND2X1 U3239 ( .A(mem[1052]), .B(n5602), .Y(n1510) );
  INVX1 U3240 ( .A(n1510), .Y(n3729) );
  AND2X1 U3241 ( .A(mem[1035]), .B(n5602), .Y(n1493) );
  INVX1 U3242 ( .A(n1493), .Y(n3730) );
  AND2X1 U3243 ( .A(mem[1026]), .B(n5602), .Y(n1484) );
  INVX1 U3244 ( .A(n1484), .Y(n3731) );
  AND2X1 U3245 ( .A(mem[1009]), .B(n5603), .Y(n1465) );
  INVX1 U3246 ( .A(n1465), .Y(n3732) );
  AND2X1 U3247 ( .A(mem[988]), .B(n5603), .Y(n1444) );
  INVX1 U3248 ( .A(n1444), .Y(n3733) );
  AND2X1 U3249 ( .A(mem[984]), .B(n5603), .Y(n1440) );
  INVX1 U3250 ( .A(n1440), .Y(n3734) );
  AND2X1 U3251 ( .A(mem[969]), .B(n5604), .Y(n1424) );
  INVX1 U3252 ( .A(n1424), .Y(n3735) );
  AND2X1 U3253 ( .A(mem[956]), .B(n5604), .Y(n1411) );
  INVX1 U3254 ( .A(n1411), .Y(n3736) );
  AND2X1 U3255 ( .A(mem[951]), .B(n5604), .Y(n1406) );
  INVX1 U3256 ( .A(n1406), .Y(n3737) );
  AND2X1 U3257 ( .A(mem[938]), .B(n5605), .Y(n1392) );
  INVX1 U3258 ( .A(n1392), .Y(n3738) );
  AND2X1 U3259 ( .A(mem[923]), .B(n5605), .Y(n1377) );
  INVX1 U3260 ( .A(n1377), .Y(n3739) );
  AND2X1 U3261 ( .A(mem[909]), .B(n5605), .Y(n1363) );
  INVX1 U3262 ( .A(n1363), .Y(n3740) );
  AND2X1 U3263 ( .A(mem[896]), .B(n5606), .Y(n1349) );
  INVX1 U3264 ( .A(n1349), .Y(n3741) );
  AND2X1 U3265 ( .A(mem[881]), .B(n5606), .Y(n1334) );
  INVX1 U3266 ( .A(n1334), .Y(n3742) );
  AND2X1 U3267 ( .A(mem[867]), .B(n5606), .Y(n1320) );
  INVX1 U3268 ( .A(n1320), .Y(n3743) );
  AND2X1 U3269 ( .A(mem[854]), .B(n5607), .Y(n1306) );
  INVX1 U3270 ( .A(n1306), .Y(n3744) );
  AND2X1 U3271 ( .A(mem[839]), .B(n5607), .Y(n1291) );
  INVX1 U3272 ( .A(n1291), .Y(n3745) );
  AND2X1 U3273 ( .A(mem[825]), .B(n5607), .Y(n1277) );
  INVX1 U3274 ( .A(n1277), .Y(n3746) );
  AND2X1 U3275 ( .A(mem[802]), .B(n5608), .Y(n1253) );
  INVX1 U3276 ( .A(n1253), .Y(n3747) );
  AND2X1 U3277 ( .A(mem[777]), .B(n5609), .Y(n1227) );
  INVX1 U3278 ( .A(n1227), .Y(n3748) );
  AND2X1 U3279 ( .A(mem[760]), .B(n5609), .Y(n1210) );
  INVX1 U3280 ( .A(n1210), .Y(n3749) );
  AND2X1 U3281 ( .A(mem[735]), .B(n5610), .Y(n1184) );
  INVX1 U3282 ( .A(n1184), .Y(n3750) );
  AND2X1 U3283 ( .A(mem[715]), .B(n5610), .Y(n1164) );
  INVX1 U3284 ( .A(n1164), .Y(n3751) );
  AND2X1 U3285 ( .A(mem[693]), .B(n5611), .Y(n1140) );
  INVX1 U3286 ( .A(n1140), .Y(n3752) );
  AND2X1 U3287 ( .A(mem[673]), .B(n5611), .Y(n1120) );
  INVX1 U3288 ( .A(n1120), .Y(n3753) );
  AND2X1 U3289 ( .A(mem[644]), .B(n5612), .Y(n1090) );
  INVX1 U3290 ( .A(n1090), .Y(n3754) );
  AND2X1 U3291 ( .A(mem[627]), .B(n5612), .Y(n1073) );
  INVX1 U3292 ( .A(n1073), .Y(n3755) );
  AND2X1 U3293 ( .A(mem[618]), .B(n5612), .Y(n1064) );
  INVX1 U3294 ( .A(n1064), .Y(n3756) );
  AND2X1 U3295 ( .A(mem[602]), .B(n5613), .Y(n1047) );
  INVX1 U3296 ( .A(n1047), .Y(n3757) );
  AND2X1 U3297 ( .A(mem[585]), .B(n5613), .Y(n1030) );
  INVX1 U3298 ( .A(n1030), .Y(n3758) );
  AND2X1 U3299 ( .A(mem[576]), .B(n5613), .Y(n1021) );
  INVX1 U3300 ( .A(n1021), .Y(n3759) );
  AND2X1 U3301 ( .A(mem[560]), .B(n5614), .Y(n1004) );
  INVX1 U3302 ( .A(n1004), .Y(n3760) );
  AND2X1 U3303 ( .A(mem[543]), .B(n5614), .Y(n987) );
  INVX1 U3304 ( .A(n987), .Y(n3761) );
  AND2X1 U3305 ( .A(mem[534]), .B(n5614), .Y(n978) );
  INVX1 U3306 ( .A(n978), .Y(n3762) );
  AND2X1 U3307 ( .A(mem[517]), .B(n5615), .Y(n960) );
  INVX1 U3308 ( .A(n960), .Y(n3763) );
  AND2X1 U3309 ( .A(mem[496]), .B(n5615), .Y(n939) );
  INVX1 U3310 ( .A(n939), .Y(n3764) );
  AND2X1 U3311 ( .A(mem[492]), .B(n5615), .Y(n935) );
  INVX1 U3312 ( .A(n935), .Y(n3765) );
  AND2X1 U3313 ( .A(mem[477]), .B(n5616), .Y(n919) );
  INVX1 U3314 ( .A(n919), .Y(n3766) );
  AND2X1 U3315 ( .A(mem[464]), .B(n5616), .Y(n906) );
  INVX1 U3316 ( .A(n906), .Y(n3767) );
  AND2X1 U3317 ( .A(mem[459]), .B(n5616), .Y(n901) );
  INVX1 U3318 ( .A(n901), .Y(n3768) );
  AND2X1 U3319 ( .A(mem[446]), .B(n5617), .Y(n887) );
  INVX1 U3320 ( .A(n887), .Y(n3769) );
  AND2X1 U3321 ( .A(mem[431]), .B(n5617), .Y(n872) );
  INVX1 U3322 ( .A(n872), .Y(n3770) );
  AND2X1 U3323 ( .A(mem[417]), .B(n5617), .Y(n858) );
  INVX1 U3324 ( .A(n858), .Y(n3771) );
  AND2X1 U3325 ( .A(mem[404]), .B(n5618), .Y(n844) );
  INVX1 U3326 ( .A(n844), .Y(n3772) );
  AND2X1 U3327 ( .A(mem[389]), .B(n5618), .Y(n829) );
  INVX1 U3328 ( .A(n829), .Y(n3773) );
  AND2X1 U3329 ( .A(mem[375]), .B(n5618), .Y(n815) );
  INVX1 U3330 ( .A(n815), .Y(n3774) );
  AND2X1 U3331 ( .A(mem[362]), .B(n5619), .Y(n800) );
  INVX1 U3332 ( .A(n800), .Y(n3775) );
  AND2X1 U3333 ( .A(mem[347]), .B(n5619), .Y(n785) );
  INVX1 U3334 ( .A(n785), .Y(n3776) );
  AND2X1 U3335 ( .A(mem[333]), .B(n5619), .Y(n771) );
  INVX1 U3336 ( .A(n771), .Y(n3777) );
  AND2X1 U3337 ( .A(mem[316]), .B(n5620), .Y(n752) );
  INVX1 U3338 ( .A(n752), .Y(n3778) );
  AND2X1 U3339 ( .A(mem[299]), .B(n5620), .Y(n735) );
  INVX1 U3340 ( .A(n735), .Y(n3779) );
  AND2X1 U3341 ( .A(mem[290]), .B(n5620), .Y(n726) );
  INVX1 U3342 ( .A(n726), .Y(n3780) );
  AND2X1 U3343 ( .A(mem[274]), .B(n5621), .Y(n708) );
  INVX1 U3344 ( .A(n708), .Y(n3781) );
  AND2X1 U3345 ( .A(mem[257]), .B(n5621), .Y(n691) );
  INVX1 U3346 ( .A(n691), .Y(n3782) );
  AND2X1 U3347 ( .A(mem[248]), .B(n5621), .Y(n682) );
  INVX1 U3348 ( .A(n682), .Y(n3783) );
  AND2X1 U3349 ( .A(mem[232]), .B(n5622), .Y(n664) );
  INVX1 U3350 ( .A(n664), .Y(n3784) );
  AND2X1 U3351 ( .A(mem[215]), .B(n5622), .Y(n647) );
  INVX1 U3352 ( .A(n647), .Y(n3785) );
  AND2X1 U3353 ( .A(mem[206]), .B(n5622), .Y(n638) );
  INVX1 U3354 ( .A(n638), .Y(n3786) );
  AND2X1 U3355 ( .A(mem[189]), .B(n5623), .Y(n619) );
  INVX1 U3356 ( .A(n619), .Y(n3787) );
  AND2X1 U3357 ( .A(mem[168]), .B(n5623), .Y(n598) );
  INVX1 U3358 ( .A(n598), .Y(n3788) );
  AND2X1 U3359 ( .A(mem[164]), .B(n5623), .Y(n594) );
  INVX1 U3360 ( .A(n594), .Y(n3789) );
  AND2X1 U3361 ( .A(mem[149]), .B(n5624), .Y(n577) );
  INVX1 U3362 ( .A(n577), .Y(n3790) );
  AND2X1 U3363 ( .A(mem[136]), .B(n5624), .Y(n564) );
  INVX1 U3364 ( .A(n564), .Y(n3791) );
  AND2X1 U3365 ( .A(mem[131]), .B(n5624), .Y(n559) );
  INVX1 U3366 ( .A(n559), .Y(n3792) );
  AND2X1 U3367 ( .A(mem[118]), .B(n5625), .Y(n544) );
  INVX1 U3368 ( .A(n544), .Y(n3793) );
  AND2X1 U3369 ( .A(mem[103]), .B(n5625), .Y(n529) );
  INVX1 U3370 ( .A(n529), .Y(n3794) );
  AND2X1 U3371 ( .A(mem[89]), .B(n5625), .Y(n515) );
  INVX1 U3372 ( .A(n515), .Y(n3795) );
  AND2X1 U3373 ( .A(mem[76]), .B(n5626), .Y(n500) );
  INVX1 U3374 ( .A(n500), .Y(n3796) );
  AND2X1 U3375 ( .A(mem[61]), .B(n5626), .Y(n485) );
  INVX1 U3376 ( .A(n485), .Y(n3797) );
  AND2X1 U3377 ( .A(mem[47]), .B(n5626), .Y(n471) );
  INVX1 U3378 ( .A(n471), .Y(n3798) );
  AND2X1 U3379 ( .A(mem[34]), .B(n5627), .Y(n449) );
  INVX1 U3380 ( .A(n449), .Y(n3799) );
  AND2X1 U3381 ( .A(mem[19]), .B(n5627), .Y(n419) );
  INVX1 U3382 ( .A(n419), .Y(n3800) );
  AND2X1 U3383 ( .A(mem[5]), .B(n5627), .Y(n391) );
  INVX1 U3384 ( .A(n391), .Y(n3801) );
  INVX1 U3385 ( .A(n1777), .Y(n3802) );
  BUFX2 U3386 ( .A(n5722), .Y(full_bar) );
  OR2X1 U3387 ( .A(fillcount[1]), .B(fillcount[0]), .Y(n1834) );
  INVX1 U3388 ( .A(n1834), .Y(n3804) );
  BUFX2 U3389 ( .A(n765), .Y(n3805) );
  BUFX2 U3390 ( .A(n464), .Y(n3806) );
  AND2X1 U3391 ( .A(n98), .B(n1786), .Y(n1788) );
  INVX1 U3392 ( .A(n1788), .Y(n3807) );
  AND2X1 U3393 ( .A(n20), .B(n1780), .Y(n1782) );
  INVX1 U3394 ( .A(n1782), .Y(n3808) );
  AND2X1 U3395 ( .A(mem[1311]), .B(n5596), .Y(n1775) );
  INVX1 U3396 ( .A(n1775), .Y(n3809) );
  AND2X1 U3397 ( .A(mem[1301]), .B(n5596), .Y(n1765) );
  INVX1 U3398 ( .A(n1765), .Y(n3810) );
  AND2X1 U3399 ( .A(mem[1280]), .B(n5596), .Y(n1744) );
  INVX1 U3400 ( .A(n1744), .Y(n3811) );
  AND2X1 U3401 ( .A(mem[1261]), .B(n5597), .Y(n1724) );
  INVX1 U3402 ( .A(n1724), .Y(n3812) );
  AND2X1 U3403 ( .A(mem[1244]), .B(n5597), .Y(n1707) );
  INVX1 U3404 ( .A(n1707), .Y(n3813) );
  AND2X1 U3405 ( .A(mem[1221]), .B(n5598), .Y(n1683) );
  INVX1 U3406 ( .A(n1683), .Y(n3814) );
  AND2X1 U3407 ( .A(mem[1204]), .B(n5598), .Y(n1666) );
  INVX1 U3408 ( .A(n1666), .Y(n3815) );
  AND2X1 U3409 ( .A(mem[1181]), .B(n5599), .Y(n1642) );
  INVX1 U3410 ( .A(n1642), .Y(n3816) );
  AND2X1 U3411 ( .A(mem[1164]), .B(n5599), .Y(n1625) );
  INVX1 U3412 ( .A(n1625), .Y(n3817) );
  AND2X1 U3413 ( .A(mem[1141]), .B(n5600), .Y(n1601) );
  INVX1 U3414 ( .A(n1601), .Y(n3818) );
  AND2X1 U3415 ( .A(mem[1126]), .B(n5600), .Y(n1586) );
  INVX1 U3416 ( .A(n1586), .Y(n3819) );
  AND2X1 U3417 ( .A(mem[1112]), .B(n5600), .Y(n1572) );
  INVX1 U3418 ( .A(n1572), .Y(n3820) );
  AND2X1 U3419 ( .A(mem[1101]), .B(n5601), .Y(n1560) );
  INVX1 U3420 ( .A(n1560), .Y(n3821) );
  AND2X1 U3421 ( .A(mem[1086]), .B(n5601), .Y(n1545) );
  INVX1 U3422 ( .A(n1545), .Y(n3822) );
  AND2X1 U3423 ( .A(mem[1072]), .B(n5601), .Y(n1531) );
  INVX1 U3424 ( .A(n1531), .Y(n3823) );
  AND2X1 U3425 ( .A(mem[1061]), .B(n5602), .Y(n1519) );
  INVX1 U3426 ( .A(n1519), .Y(n3824) );
  AND2X1 U3427 ( .A(mem[1046]), .B(n5602), .Y(n1504) );
  INVX1 U3428 ( .A(n1504), .Y(n3825) );
  AND2X1 U3429 ( .A(mem[1032]), .B(n5602), .Y(n1490) );
  INVX1 U3430 ( .A(n1490), .Y(n3826) );
  AND2X1 U3431 ( .A(mem[1010]), .B(n5603), .Y(n1466) );
  INVX1 U3432 ( .A(n1466), .Y(n3827) );
  AND2X1 U3433 ( .A(mem[997]), .B(n5603), .Y(n1453) );
  INVX1 U3434 ( .A(n1453), .Y(n3828) );
  AND2X1 U3435 ( .A(mem[992]), .B(n5603), .Y(n1448) );
  INVX1 U3436 ( .A(n1448), .Y(n3829) );
  AND2X1 U3437 ( .A(mem[968]), .B(n5604), .Y(n1423) );
  INVX1 U3438 ( .A(n1423), .Y(n3830) );
  AND2X1 U3439 ( .A(mem[947]), .B(n5604), .Y(n1402) );
  INVX1 U3440 ( .A(n1402), .Y(n3831) );
  AND2X1 U3441 ( .A(mem[943]), .B(n5604), .Y(n1398) );
  INVX1 U3442 ( .A(n1398), .Y(n3832) );
  AND2X1 U3443 ( .A(mem[929]), .B(n5605), .Y(n1383) );
  INVX1 U3444 ( .A(n1383), .Y(n3833) );
  AND2X1 U3445 ( .A(mem[912]), .B(n5605), .Y(n1366) );
  INVX1 U3446 ( .A(n1366), .Y(n3834) );
  AND2X1 U3447 ( .A(mem[903]), .B(n5605), .Y(n1357) );
  INVX1 U3448 ( .A(n1357), .Y(n3835) );
  AND2X1 U3449 ( .A(mem[889]), .B(n5606), .Y(n1342) );
  INVX1 U3450 ( .A(n1342), .Y(n3836) );
  AND2X1 U3451 ( .A(mem[872]), .B(n5606), .Y(n1325) );
  INVX1 U3452 ( .A(n1325), .Y(n3837) );
  AND2X1 U3453 ( .A(mem[863]), .B(n5606), .Y(n1316) );
  INVX1 U3454 ( .A(n1316), .Y(n3838) );
  AND2X1 U3455 ( .A(mem[849]), .B(n5607), .Y(n1301) );
  INVX1 U3456 ( .A(n1301), .Y(n3839) );
  AND2X1 U3457 ( .A(mem[832]), .B(n5607), .Y(n1284) );
  INVX1 U3458 ( .A(n1284), .Y(n3840) );
  AND2X1 U3459 ( .A(mem[823]), .B(n5607), .Y(n1275) );
  INVX1 U3460 ( .A(n1275), .Y(n3841) );
  AND2X1 U3461 ( .A(mem[819]), .B(n5608), .Y(n1270) );
  INVX1 U3462 ( .A(n1270), .Y(n3842) );
  AND2X1 U3463 ( .A(mem[809]), .B(n5608), .Y(n1260) );
  INVX1 U3464 ( .A(n1260), .Y(n3843) );
  AND2X1 U3465 ( .A(mem[788]), .B(n5608), .Y(n1239) );
  INVX1 U3466 ( .A(n1239), .Y(n3844) );
  AND2X1 U3467 ( .A(mem[769]), .B(n5609), .Y(n1219) );
  INVX1 U3468 ( .A(n1219), .Y(n3845) );
  AND2X1 U3469 ( .A(mem[752]), .B(n5609), .Y(n1202) );
  INVX1 U3470 ( .A(n1202), .Y(n3846) );
  AND2X1 U3471 ( .A(mem[729]), .B(n5610), .Y(n1178) );
  INVX1 U3472 ( .A(n1178), .Y(n3847) );
  AND2X1 U3473 ( .A(mem[712]), .B(n5610), .Y(n1161) );
  INVX1 U3474 ( .A(n1161), .Y(n3848) );
  AND2X1 U3475 ( .A(mem[689]), .B(n5611), .Y(n1136) );
  INVX1 U3476 ( .A(n1136), .Y(n3849) );
  AND2X1 U3477 ( .A(mem[672]), .B(n5611), .Y(n1119) );
  INVX1 U3478 ( .A(n1119), .Y(n3850) );
  AND2X1 U3479 ( .A(mem[649]), .B(n5612), .Y(n1095) );
  INVX1 U3480 ( .A(n1095), .Y(n3851) );
  AND2X1 U3481 ( .A(mem[634]), .B(n5612), .Y(n1080) );
  INVX1 U3482 ( .A(n1080), .Y(n3852) );
  AND2X1 U3483 ( .A(mem[620]), .B(n5612), .Y(n1066) );
  INVX1 U3484 ( .A(n1066), .Y(n3853) );
  AND2X1 U3485 ( .A(mem[609]), .B(n5613), .Y(n1054) );
  INVX1 U3486 ( .A(n1054), .Y(n3854) );
  AND2X1 U3487 ( .A(mem[594]), .B(n5613), .Y(n1039) );
  INVX1 U3488 ( .A(n1039), .Y(n3855) );
  AND2X1 U3489 ( .A(mem[580]), .B(n5613), .Y(n1025) );
  INVX1 U3490 ( .A(n1025), .Y(n3856) );
  AND2X1 U3491 ( .A(mem[569]), .B(n5614), .Y(n1013) );
  INVX1 U3492 ( .A(n1013), .Y(n3857) );
  AND2X1 U3493 ( .A(mem[554]), .B(n5614), .Y(n998) );
  INVX1 U3494 ( .A(n998), .Y(n3858) );
  AND2X1 U3495 ( .A(mem[540]), .B(n5614), .Y(n984) );
  INVX1 U3496 ( .A(n984), .Y(n3859) );
  AND2X1 U3497 ( .A(mem[518]), .B(n5615), .Y(n961) );
  INVX1 U3498 ( .A(n961), .Y(n3860) );
  AND2X1 U3499 ( .A(mem[505]), .B(n5615), .Y(n948) );
  INVX1 U3500 ( .A(n948), .Y(n3861) );
  AND2X1 U3501 ( .A(mem[500]), .B(n5615), .Y(n943) );
  INVX1 U3502 ( .A(n943), .Y(n3862) );
  AND2X1 U3503 ( .A(mem[476]), .B(n5616), .Y(n918) );
  INVX1 U3504 ( .A(n918), .Y(n3863) );
  AND2X1 U3505 ( .A(mem[455]), .B(n5616), .Y(n897) );
  INVX1 U3506 ( .A(n897), .Y(n3864) );
  AND2X1 U3507 ( .A(mem[451]), .B(n5616), .Y(n893) );
  INVX1 U3508 ( .A(n893), .Y(n3865) );
  AND2X1 U3509 ( .A(mem[437]), .B(n5617), .Y(n878) );
  INVX1 U3510 ( .A(n878), .Y(n3866) );
  AND2X1 U3511 ( .A(mem[420]), .B(n5617), .Y(n861) );
  INVX1 U3512 ( .A(n861), .Y(n3867) );
  AND2X1 U3513 ( .A(mem[411]), .B(n5617), .Y(n852) );
  INVX1 U3514 ( .A(n852), .Y(n3868) );
  AND2X1 U3515 ( .A(mem[397]), .B(n5618), .Y(n837) );
  INVX1 U3516 ( .A(n837), .Y(n3869) );
  AND2X1 U3517 ( .A(mem[380]), .B(n5618), .Y(n820) );
  INVX1 U3518 ( .A(n820), .Y(n3870) );
  AND2X1 U3519 ( .A(mem[371]), .B(n5618), .Y(n811) );
  INVX1 U3520 ( .A(n811), .Y(n3871) );
  AND2X1 U3521 ( .A(mem[357]), .B(n5619), .Y(n795) );
  INVX1 U3522 ( .A(n795), .Y(n3872) );
  AND2X1 U3523 ( .A(mem[340]), .B(n5619), .Y(n778) );
  INVX1 U3524 ( .A(n778), .Y(n3873) );
  AND2X1 U3525 ( .A(mem[331]), .B(n5619), .Y(n769) );
  INVX1 U3526 ( .A(n769), .Y(n3874) );
  AND2X1 U3527 ( .A(mem[321]), .B(n5620), .Y(n757) );
  INVX1 U3528 ( .A(n757), .Y(n3875) );
  AND2X1 U3529 ( .A(mem[306]), .B(n5620), .Y(n742) );
  INVX1 U3530 ( .A(n742), .Y(n3876) );
  AND2X1 U3531 ( .A(mem[292]), .B(n5620), .Y(n728) );
  INVX1 U3532 ( .A(n728), .Y(n3877) );
  AND2X1 U3533 ( .A(mem[281]), .B(n5621), .Y(n715) );
  INVX1 U3534 ( .A(n715), .Y(n3878) );
  AND2X1 U3535 ( .A(mem[266]), .B(n5621), .Y(n700) );
  INVX1 U3536 ( .A(n700), .Y(n3879) );
  AND2X1 U3537 ( .A(mem[252]), .B(n5621), .Y(n686) );
  INVX1 U3538 ( .A(n686), .Y(n3880) );
  AND2X1 U3539 ( .A(mem[241]), .B(n5622), .Y(n673) );
  INVX1 U3540 ( .A(n673), .Y(n3881) );
  AND2X1 U3541 ( .A(mem[226]), .B(n5622), .Y(n658) );
  INVX1 U3542 ( .A(n658), .Y(n3882) );
  AND2X1 U3543 ( .A(mem[212]), .B(n5622), .Y(n644) );
  INVX1 U3544 ( .A(n644), .Y(n3883) );
  AND2X1 U3545 ( .A(mem[190]), .B(n5623), .Y(n620) );
  INVX1 U3546 ( .A(n620), .Y(n3884) );
  AND2X1 U3547 ( .A(mem[177]), .B(n5623), .Y(n607) );
  INVX1 U3548 ( .A(n607), .Y(n3885) );
  AND2X1 U3549 ( .A(mem[172]), .B(n5623), .Y(n602) );
  INVX1 U3550 ( .A(n602), .Y(n3886) );
  AND2X1 U3551 ( .A(mem[148]), .B(n5624), .Y(n576) );
  INVX1 U3552 ( .A(n576), .Y(n3887) );
  AND2X1 U3553 ( .A(mem[127]), .B(n5624), .Y(n555) );
  INVX1 U3554 ( .A(n555), .Y(n3888) );
  AND2X1 U3555 ( .A(mem[123]), .B(n5624), .Y(n551) );
  INVX1 U3556 ( .A(n551), .Y(n3889) );
  AND2X1 U3557 ( .A(mem[109]), .B(n5625), .Y(n535) );
  INVX1 U3558 ( .A(n535), .Y(n3890) );
  AND2X1 U3559 ( .A(mem[92]), .B(n5625), .Y(n518) );
  INVX1 U3560 ( .A(n518), .Y(n3891) );
  AND2X1 U3561 ( .A(mem[83]), .B(n5625), .Y(n509) );
  INVX1 U3562 ( .A(n509), .Y(n3892) );
  AND2X1 U3563 ( .A(mem[69]), .B(n5626), .Y(n493) );
  INVX1 U3564 ( .A(n493), .Y(n3893) );
  AND2X1 U3565 ( .A(mem[52]), .B(n5626), .Y(n476) );
  INVX1 U3566 ( .A(n476), .Y(n3894) );
  AND2X1 U3567 ( .A(mem[43]), .B(n5626), .Y(n467) );
  INVX1 U3568 ( .A(n467), .Y(n3895) );
  AND2X1 U3569 ( .A(mem[29]), .B(n5627), .Y(n439) );
  INVX1 U3570 ( .A(n439), .Y(n3896) );
  AND2X1 U3571 ( .A(mem[12]), .B(n5627), .Y(n405) );
  INVX1 U3572 ( .A(n405), .Y(n3897) );
  AND2X1 U3573 ( .A(mem[3]), .B(n5627), .Y(n387) );
  INVX1 U3574 ( .A(n387), .Y(n3898) );
  BUFX2 U3575 ( .A(n463), .Y(n3899) );
  AND2X1 U3576 ( .A(n99), .B(n1786), .Y(n1787) );
  INVX1 U3577 ( .A(n1787), .Y(n3900) );
  AND2X1 U3578 ( .A(n21), .B(n1780), .Y(n1781) );
  INVX1 U3579 ( .A(n1781), .Y(n3901) );
  AND2X1 U3580 ( .A(reset), .B(n4084), .Y(n1780) );
  AND2X1 U3581 ( .A(mem[1302]), .B(n5596), .Y(n1766) );
  INVX1 U3582 ( .A(n1766), .Y(n3902) );
  AND2X1 U3583 ( .A(mem[1285]), .B(n5596), .Y(n1749) );
  INVX1 U3584 ( .A(n1749), .Y(n3903) );
  AND2X1 U3585 ( .A(mem[1270]), .B(n5597), .Y(n1733) );
  INVX1 U3586 ( .A(n1733), .Y(n3904) );
  AND2X1 U3587 ( .A(mem[1260]), .B(n5597), .Y(n1723) );
  INVX1 U3588 ( .A(n1723), .Y(n3905) );
  AND2X1 U3589 ( .A(mem[1239]), .B(n5597), .Y(n1702) );
  INVX1 U3590 ( .A(n1702), .Y(n3906) );
  AND2X1 U3591 ( .A(mem[1222]), .B(n5598), .Y(n1684) );
  INVX1 U3592 ( .A(n1684), .Y(n3907) );
  AND2X1 U3593 ( .A(mem[1205]), .B(n5598), .Y(n1667) );
  INVX1 U3594 ( .A(n1667), .Y(n3908) );
  AND2X1 U3595 ( .A(mem[1180]), .B(n5599), .Y(n1641) );
  INVX1 U3596 ( .A(n1641), .Y(n3909) );
  AND2X1 U3597 ( .A(mem[1163]), .B(n5599), .Y(n1624) );
  INVX1 U3598 ( .A(n1624), .Y(n3910) );
  AND2X1 U3599 ( .A(mem[1142]), .B(n5600), .Y(n1602) );
  INVX1 U3600 ( .A(n1602), .Y(n3911) );
  AND2X1 U3601 ( .A(mem[1127]), .B(n5600), .Y(n1587) );
  INVX1 U3602 ( .A(n1587), .Y(n3912) );
  AND2X1 U3603 ( .A(mem[1113]), .B(n5600), .Y(n1573) );
  INVX1 U3604 ( .A(n1573), .Y(n3913) );
  AND2X1 U3605 ( .A(mem[1100]), .B(n5601), .Y(n1559) );
  INVX1 U3606 ( .A(n1559), .Y(n3914) );
  AND2X1 U3607 ( .A(mem[1085]), .B(n5601), .Y(n1544) );
  INVX1 U3608 ( .A(n1544), .Y(n3915) );
  AND2X1 U3609 ( .A(mem[1071]), .B(n5601), .Y(n1530) );
  INVX1 U3610 ( .A(n1530), .Y(n3916) );
  AND2X1 U3611 ( .A(mem[1051]), .B(n5602), .Y(n1509) );
  INVX1 U3612 ( .A(n1509), .Y(n3917) );
  AND2X1 U3613 ( .A(mem[1038]), .B(n5602), .Y(n1496) );
  INVX1 U3614 ( .A(n1496), .Y(n3918) );
  AND2X1 U3615 ( .A(mem[1033]), .B(n5602), .Y(n1491) );
  INVX1 U3616 ( .A(n1491), .Y(n3919) );
  AND2X1 U3617 ( .A(mem[1020]), .B(n5603), .Y(n1476) );
  INVX1 U3618 ( .A(n1476), .Y(n3920) );
  AND2X1 U3619 ( .A(mem[1005]), .B(n5603), .Y(n1461) );
  INVX1 U3620 ( .A(n1461), .Y(n3921) );
  AND2X1 U3621 ( .A(mem[991]), .B(n5603), .Y(n1447) );
  INVX1 U3622 ( .A(n1447), .Y(n3922) );
  AND2X1 U3623 ( .A(mem[970]), .B(n5604), .Y(n1425) );
  INVX1 U3624 ( .A(n1425), .Y(n3923) );
  AND2X1 U3625 ( .A(mem[953]), .B(n5604), .Y(n1408) );
  INVX1 U3626 ( .A(n1408), .Y(n3924) );
  AND2X1 U3627 ( .A(mem[944]), .B(n5604), .Y(n1399) );
  INVX1 U3628 ( .A(n1399), .Y(n3925) );
  AND2X1 U3629 ( .A(mem[927]), .B(n5605), .Y(n1381) );
  INVX1 U3630 ( .A(n1381), .Y(n3926) );
  AND2X1 U3631 ( .A(mem[906]), .B(n5605), .Y(n1360) );
  INVX1 U3632 ( .A(n1360), .Y(n3927) );
  AND2X1 U3633 ( .A(mem[902]), .B(n5605), .Y(n1356) );
  INVX1 U3634 ( .A(n1356), .Y(n3928) );
  AND2X1 U3635 ( .A(mem[890]), .B(n5606), .Y(n1343) );
  INVX1 U3636 ( .A(n1343), .Y(n3929) );
  AND2X1 U3637 ( .A(mem[873]), .B(n5606), .Y(n1326) );
  INVX1 U3638 ( .A(n1326), .Y(n3930) );
  AND2X1 U3639 ( .A(mem[864]), .B(n5606), .Y(n1317) );
  INVX1 U3640 ( .A(n1317), .Y(n3931) );
  AND2X1 U3641 ( .A(mem[848]), .B(n5607), .Y(n1300) );
  INVX1 U3642 ( .A(n1300), .Y(n3932) );
  AND2X1 U3643 ( .A(mem[831]), .B(n5607), .Y(n1283) );
  INVX1 U3644 ( .A(n1283), .Y(n3933) );
  AND2X1 U3645 ( .A(mem[822]), .B(n5607), .Y(n1274) );
  INVX1 U3646 ( .A(n1274), .Y(n3934) );
  AND2X1 U3647 ( .A(mem[810]), .B(n5608), .Y(n1261) );
  INVX1 U3648 ( .A(n1261), .Y(n3935) );
  AND2X1 U3649 ( .A(mem[793]), .B(n5608), .Y(n1244) );
  INVX1 U3650 ( .A(n1244), .Y(n3936) );
  AND2X1 U3651 ( .A(mem[778]), .B(n5609), .Y(n1228) );
  INVX1 U3652 ( .A(n1228), .Y(n3937) );
  AND2X1 U3653 ( .A(mem[768]), .B(n5609), .Y(n1218) );
  INVX1 U3654 ( .A(n1218), .Y(n3938) );
  AND2X1 U3655 ( .A(mem[747]), .B(n5609), .Y(n1197) );
  INVX1 U3656 ( .A(n1197), .Y(n3939) );
  AND2X1 U3657 ( .A(mem[730]), .B(n5610), .Y(n1179) );
  INVX1 U3658 ( .A(n1179), .Y(n3940) );
  AND2X1 U3659 ( .A(mem[713]), .B(n5610), .Y(n1162) );
  INVX1 U3660 ( .A(n1162), .Y(n3941) );
  AND2X1 U3661 ( .A(mem[688]), .B(n5611), .Y(n1135) );
  INVX1 U3662 ( .A(n1135), .Y(n3942) );
  AND2X1 U3663 ( .A(mem[671]), .B(n5611), .Y(n1118) );
  INVX1 U3664 ( .A(n1118), .Y(n3943) );
  AND2X1 U3665 ( .A(mem[650]), .B(n5612), .Y(n1096) );
  INVX1 U3666 ( .A(n1096), .Y(n3944) );
  AND2X1 U3667 ( .A(mem[635]), .B(n5612), .Y(n1081) );
  INVX1 U3668 ( .A(n1081), .Y(n3945) );
  AND2X1 U3669 ( .A(mem[621]), .B(n5612), .Y(n1067) );
  INVX1 U3670 ( .A(n1067), .Y(n3946) );
  AND2X1 U3671 ( .A(mem[608]), .B(n5613), .Y(n1053) );
  INVX1 U3672 ( .A(n1053), .Y(n3947) );
  AND2X1 U3673 ( .A(mem[593]), .B(n5613), .Y(n1038) );
  INVX1 U3674 ( .A(n1038), .Y(n3948) );
  AND2X1 U3675 ( .A(mem[579]), .B(n5613), .Y(n1024) );
  INVX1 U3676 ( .A(n1024), .Y(n3949) );
  AND2X1 U3677 ( .A(mem[559]), .B(n5614), .Y(n1003) );
  INVX1 U3678 ( .A(n1003), .Y(n3950) );
  AND2X1 U3679 ( .A(mem[546]), .B(n5614), .Y(n990) );
  INVX1 U3680 ( .A(n990), .Y(n3951) );
  AND2X1 U3681 ( .A(mem[541]), .B(n5614), .Y(n985) );
  INVX1 U3682 ( .A(n985), .Y(n3952) );
  AND2X1 U3683 ( .A(mem[528]), .B(n5615), .Y(n971) );
  INVX1 U3684 ( .A(n971), .Y(n3953) );
  AND2X1 U3685 ( .A(mem[513]), .B(n5615), .Y(n956) );
  INVX1 U3686 ( .A(n956), .Y(n3954) );
  AND2X1 U3687 ( .A(mem[499]), .B(n5615), .Y(n942) );
  INVX1 U3688 ( .A(n942), .Y(n3955) );
  AND2X1 U3689 ( .A(mem[478]), .B(n5616), .Y(n920) );
  INVX1 U3690 ( .A(n920), .Y(n3956) );
  AND2X1 U3691 ( .A(mem[461]), .B(n5616), .Y(n903) );
  INVX1 U3692 ( .A(n903), .Y(n3957) );
  AND2X1 U3693 ( .A(mem[452]), .B(n5616), .Y(n894) );
  INVX1 U3694 ( .A(n894), .Y(n3958) );
  AND2X1 U3695 ( .A(mem[435]), .B(n5617), .Y(n876) );
  INVX1 U3696 ( .A(n876), .Y(n3959) );
  AND2X1 U3697 ( .A(mem[414]), .B(n5617), .Y(n855) );
  INVX1 U3698 ( .A(n855), .Y(n3960) );
  AND2X1 U3699 ( .A(mem[410]), .B(n5617), .Y(n851) );
  INVX1 U3700 ( .A(n851), .Y(n3961) );
  AND2X1 U3701 ( .A(mem[398]), .B(n5618), .Y(n838) );
  INVX1 U3702 ( .A(n838), .Y(n3962) );
  AND2X1 U3703 ( .A(mem[381]), .B(n5618), .Y(n821) );
  INVX1 U3704 ( .A(n821), .Y(n3963) );
  AND2X1 U3705 ( .A(mem[372]), .B(n5618), .Y(n812) );
  INVX1 U3706 ( .A(n812), .Y(n3964) );
  AND2X1 U3707 ( .A(mem[356]), .B(n5619), .Y(n794) );
  INVX1 U3708 ( .A(n794), .Y(n3965) );
  AND2X1 U3709 ( .A(mem[339]), .B(n5619), .Y(n777) );
  INVX1 U3710 ( .A(n777), .Y(n3966) );
  AND2X1 U3711 ( .A(mem[330]), .B(n5619), .Y(n768) );
  INVX1 U3712 ( .A(n768), .Y(n3967) );
  AND2X1 U3713 ( .A(mem[322]), .B(n5620), .Y(n758) );
  INVX1 U3714 ( .A(n758), .Y(n3968) );
  AND2X1 U3715 ( .A(mem[307]), .B(n5620), .Y(n743) );
  INVX1 U3716 ( .A(n743), .Y(n3969) );
  AND2X1 U3717 ( .A(mem[293]), .B(n5620), .Y(n729) );
  INVX1 U3718 ( .A(n729), .Y(n3970) );
  AND2X1 U3719 ( .A(mem[280]), .B(n5621), .Y(n714) );
  INVX1 U3720 ( .A(n714), .Y(n3971) );
  AND2X1 U3721 ( .A(mem[265]), .B(n5621), .Y(n699) );
  INVX1 U3722 ( .A(n699), .Y(n3972) );
  AND2X1 U3723 ( .A(mem[251]), .B(n5621), .Y(n685) );
  INVX1 U3724 ( .A(n685), .Y(n3973) );
  AND2X1 U3725 ( .A(mem[231]), .B(n5622), .Y(n663) );
  INVX1 U3726 ( .A(n663), .Y(n3974) );
  AND2X1 U3727 ( .A(mem[218]), .B(n5622), .Y(n650) );
  INVX1 U3728 ( .A(n650), .Y(n3975) );
  AND2X1 U3729 ( .A(mem[213]), .B(n5622), .Y(n645) );
  INVX1 U3730 ( .A(n645), .Y(n3976) );
  AND2X1 U3731 ( .A(mem[200]), .B(n5623), .Y(n630) );
  INVX1 U3732 ( .A(n630), .Y(n3977) );
  AND2X1 U3733 ( .A(mem[185]), .B(n5623), .Y(n615) );
  INVX1 U3734 ( .A(n615), .Y(n3978) );
  AND2X1 U3735 ( .A(mem[171]), .B(n5623), .Y(n601) );
  INVX1 U3736 ( .A(n601), .Y(n3979) );
  AND2X1 U3737 ( .A(mem[150]), .B(n5624), .Y(n578) );
  INVX1 U3738 ( .A(n578), .Y(n3980) );
  AND2X1 U3739 ( .A(mem[133]), .B(n5624), .Y(n561) );
  INVX1 U3740 ( .A(n561), .Y(n3981) );
  AND2X1 U3741 ( .A(mem[124]), .B(n5624), .Y(n552) );
  INVX1 U3742 ( .A(n552), .Y(n3982) );
  AND2X1 U3743 ( .A(mem[107]), .B(n5625), .Y(n533) );
  INVX1 U3744 ( .A(n533), .Y(n3983) );
  AND2X1 U3745 ( .A(mem[86]), .B(n5625), .Y(n512) );
  INVX1 U3746 ( .A(n512), .Y(n3984) );
  AND2X1 U3747 ( .A(mem[82]), .B(n5625), .Y(n508) );
  INVX1 U3748 ( .A(n508), .Y(n3985) );
  AND2X1 U3749 ( .A(mem[70]), .B(n5626), .Y(n494) );
  INVX1 U3750 ( .A(n494), .Y(n3986) );
  AND2X1 U3751 ( .A(mem[53]), .B(n5626), .Y(n477) );
  INVX1 U3752 ( .A(n477), .Y(n3987) );
  AND2X1 U3753 ( .A(mem[44]), .B(n5626), .Y(n468) );
  INVX1 U3754 ( .A(n468), .Y(n3988) );
  AND2X1 U3755 ( .A(mem[28]), .B(n5627), .Y(n437) );
  INVX1 U3756 ( .A(n437), .Y(n3989) );
  AND2X1 U3757 ( .A(mem[11]), .B(n5627), .Y(n403) );
  INVX1 U3758 ( .A(n403), .Y(n3990) );
  AND2X1 U3759 ( .A(mem[2]), .B(n5627), .Y(n385) );
  INVX1 U3760 ( .A(n385), .Y(n3991) );
  BUFX2 U3761 ( .A(n1482), .Y(n3992) );
  AND2X1 U3762 ( .A(n100), .B(n1786), .Y(n1785) );
  INVX1 U3763 ( .A(n1785), .Y(n3993) );
  AND2X1 U3764 ( .A(mem[1303]), .B(n5596), .Y(n1767) );
  INVX1 U3765 ( .A(n1767), .Y(n3994) );
  AND2X1 U3766 ( .A(mem[1286]), .B(n5596), .Y(n1750) );
  INVX1 U3767 ( .A(n1750), .Y(n3995) );
  AND2X1 U3768 ( .A(mem[1263]), .B(n5597), .Y(n1726) );
  INVX1 U3769 ( .A(n1726), .Y(n3996) );
  AND2X1 U3770 ( .A(mem[1246]), .B(n5597), .Y(n1709) );
  INVX1 U3771 ( .A(n1709), .Y(n3997) );
  AND2X1 U3772 ( .A(mem[1229]), .B(n5598), .Y(n1691) );
  INVX1 U3773 ( .A(n1691), .Y(n3998) );
  AND2X1 U3774 ( .A(mem[1219]), .B(n5598), .Y(n1681) );
  INVX1 U3775 ( .A(n1681), .Y(n3999) );
  AND2X1 U3776 ( .A(mem[1198]), .B(n5598), .Y(n1660) );
  INVX1 U3777 ( .A(n1660), .Y(n4000) );
  AND2X1 U3778 ( .A(mem[1179]), .B(n5599), .Y(n1640) );
  INVX1 U3779 ( .A(n1640), .Y(n4001) );
  AND2X1 U3780 ( .A(mem[1162]), .B(n5599), .Y(n1623) );
  INVX1 U3781 ( .A(n1623), .Y(n4002) );
  AND2X1 U3782 ( .A(mem[1143]), .B(n5600), .Y(n1603) );
  INVX1 U3783 ( .A(n1603), .Y(n4003) );
  AND2X1 U3784 ( .A(mem[1128]), .B(n5600), .Y(n1588) );
  INVX1 U3785 ( .A(n1588), .Y(n4004) );
  AND2X1 U3786 ( .A(mem[1114]), .B(n5600), .Y(n1574) );
  INVX1 U3787 ( .A(n1574), .Y(n4005) );
  AND2X1 U3788 ( .A(mem[1092]), .B(n5601), .Y(n1551) );
  INVX1 U3789 ( .A(n1551), .Y(n4006) );
  AND2X1 U3790 ( .A(mem[1079]), .B(n5601), .Y(n1538) );
  INVX1 U3791 ( .A(n1538), .Y(n4007) );
  AND2X1 U3792 ( .A(mem[1074]), .B(n5601), .Y(n1533) );
  INVX1 U3793 ( .A(n1533), .Y(n4008) );
  AND2X1 U3794 ( .A(mem[1059]), .B(n5602), .Y(n1517) );
  INVX1 U3795 ( .A(n1517), .Y(n4009) );
  AND2X1 U3796 ( .A(mem[1044]), .B(n5602), .Y(n1502) );
  INVX1 U3797 ( .A(n1502), .Y(n4010) );
  AND2X1 U3798 ( .A(mem[1030]), .B(n5602), .Y(n1488) );
  INVX1 U3799 ( .A(n1488), .Y(n4011) );
  AND2X1 U3800 ( .A(mem[1019]), .B(n5603), .Y(n1475) );
  INVX1 U3801 ( .A(n1475), .Y(n4012) );
  AND2X1 U3802 ( .A(mem[1004]), .B(n5603), .Y(n1460) );
  INVX1 U3803 ( .A(n1460), .Y(n4013) );
  AND2X1 U3804 ( .A(mem[990]), .B(n5603), .Y(n1446) );
  INVX1 U3805 ( .A(n1446), .Y(n4014) );
  AND2X1 U3806 ( .A(mem[971]), .B(n5604), .Y(n1426) );
  INVX1 U3807 ( .A(n1426), .Y(n4015) );
  AND2X1 U3808 ( .A(mem[954]), .B(n5604), .Y(n1409) );
  INVX1 U3809 ( .A(n1409), .Y(n4016) );
  AND2X1 U3810 ( .A(mem[945]), .B(n5604), .Y(n1400) );
  INVX1 U3811 ( .A(n1400), .Y(n4017) );
  AND2X1 U3812 ( .A(mem[931]), .B(n5605), .Y(n1385) );
  INVX1 U3813 ( .A(n1385), .Y(n4018) );
  AND2X1 U3814 ( .A(mem[914]), .B(n5605), .Y(n1368) );
  INVX1 U3815 ( .A(n1368), .Y(n4019) );
  AND2X1 U3816 ( .A(mem[905]), .B(n5605), .Y(n1359) );
  INVX1 U3817 ( .A(n1359), .Y(n4020) );
  AND2X1 U3818 ( .A(mem[886]), .B(n5606), .Y(n1339) );
  INVX1 U3819 ( .A(n1339), .Y(n4021) );
  AND2X1 U3820 ( .A(mem[865]), .B(n5606), .Y(n1318) );
  INVX1 U3821 ( .A(n1318), .Y(n4022) );
  AND2X1 U3822 ( .A(mem[861]), .B(n5606), .Y(n1314) );
  INVX1 U3823 ( .A(n1314), .Y(n4023) );
  AND2X1 U3824 ( .A(mem[847]), .B(n5607), .Y(n1299) );
  INVX1 U3825 ( .A(n1299), .Y(n4024) );
  AND2X1 U3826 ( .A(mem[830]), .B(n5607), .Y(n1282) );
  INVX1 U3827 ( .A(n1282), .Y(n4025) );
  AND2X1 U3828 ( .A(mem[821]), .B(n5607), .Y(n1273) );
  INVX1 U3829 ( .A(n1273), .Y(n4026) );
  AND2X1 U3830 ( .A(mem[811]), .B(n5608), .Y(n1262) );
  INVX1 U3831 ( .A(n1262), .Y(n4027) );
  AND2X1 U3832 ( .A(mem[794]), .B(n5608), .Y(n1245) );
  INVX1 U3833 ( .A(n1245), .Y(n4028) );
  AND2X1 U3834 ( .A(mem[771]), .B(n5609), .Y(n1221) );
  INVX1 U3835 ( .A(n1221), .Y(n4029) );
  AND2X1 U3836 ( .A(mem[754]), .B(n5609), .Y(n1204) );
  INVX1 U3837 ( .A(n1204), .Y(n4030) );
  AND2X1 U3838 ( .A(mem[737]), .B(n5610), .Y(n1186) );
  INVX1 U3839 ( .A(n1186), .Y(n4031) );
  AND2X1 U3840 ( .A(mem[727]), .B(n5610), .Y(n1176) );
  INVX1 U3841 ( .A(n1176), .Y(n4032) );
  AND2X1 U3842 ( .A(mem[706]), .B(n5610), .Y(n1155) );
  INVX1 U3843 ( .A(n1155), .Y(n4033) );
  AND2X1 U3844 ( .A(mem[687]), .B(n5611), .Y(n1134) );
  INVX1 U3845 ( .A(n1134), .Y(n4034) );
  AND2X1 U3846 ( .A(mem[670]), .B(n5611), .Y(n1117) );
  INVX1 U3847 ( .A(n1117), .Y(n4035) );
  AND2X1 U3848 ( .A(mem[651]), .B(n5612), .Y(n1097) );
  INVX1 U3849 ( .A(n1097), .Y(n4036) );
  AND2X1 U3850 ( .A(mem[636]), .B(n5612), .Y(n1082) );
  INVX1 U3851 ( .A(n1082), .Y(n4037) );
  AND2X1 U3852 ( .A(mem[622]), .B(n5612), .Y(n1068) );
  INVX1 U3853 ( .A(n1068), .Y(n4038) );
  AND2X1 U3854 ( .A(mem[600]), .B(n5613), .Y(n1045) );
  INVX1 U3855 ( .A(n1045), .Y(n4039) );
  AND2X1 U3856 ( .A(mem[587]), .B(n5613), .Y(n1032) );
  INVX1 U3857 ( .A(n1032), .Y(n4040) );
  AND2X1 U3858 ( .A(mem[582]), .B(n5613), .Y(n1027) );
  INVX1 U3859 ( .A(n1027), .Y(n4041) );
  AND2X1 U3860 ( .A(mem[567]), .B(n5614), .Y(n1011) );
  INVX1 U3861 ( .A(n1011), .Y(n4042) );
  AND2X1 U3862 ( .A(mem[552]), .B(n5614), .Y(n996) );
  INVX1 U3863 ( .A(n996), .Y(n4043) );
  AND2X1 U3864 ( .A(mem[538]), .B(n5614), .Y(n982) );
  INVX1 U3865 ( .A(n982), .Y(n4044) );
  AND2X1 U3866 ( .A(mem[527]), .B(n5615), .Y(n970) );
  INVX1 U3867 ( .A(n970), .Y(n4045) );
  AND2X1 U3868 ( .A(mem[512]), .B(n5615), .Y(n955) );
  INVX1 U3869 ( .A(n955), .Y(n4046) );
  AND2X1 U3870 ( .A(mem[498]), .B(n5615), .Y(n941) );
  INVX1 U3871 ( .A(n941), .Y(n4047) );
  AND2X1 U3872 ( .A(mem[479]), .B(n5616), .Y(n921) );
  INVX1 U3873 ( .A(n921), .Y(n4048) );
  AND2X1 U3874 ( .A(mem[462]), .B(n5616), .Y(n904) );
  INVX1 U3875 ( .A(n904), .Y(n4049) );
  AND2X1 U3876 ( .A(mem[453]), .B(n5616), .Y(n895) );
  INVX1 U3877 ( .A(n895), .Y(n4050) );
  AND2X1 U3878 ( .A(mem[439]), .B(n5617), .Y(n880) );
  INVX1 U3879 ( .A(n880), .Y(n4051) );
  AND2X1 U3880 ( .A(mem[422]), .B(n5617), .Y(n863) );
  INVX1 U3881 ( .A(n863), .Y(n4052) );
  AND2X1 U3882 ( .A(mem[413]), .B(n5617), .Y(n854) );
  INVX1 U3883 ( .A(n854), .Y(n4053) );
  AND2X1 U3884 ( .A(mem[394]), .B(n5618), .Y(n834) );
  INVX1 U3885 ( .A(n834), .Y(n4054) );
  AND2X1 U3886 ( .A(mem[373]), .B(n5618), .Y(n813) );
  INVX1 U3887 ( .A(n813), .Y(n4055) );
  AND2X1 U3888 ( .A(mem[369]), .B(n5618), .Y(n809) );
  INVX1 U3889 ( .A(n809), .Y(n4056) );
  AND2X1 U3890 ( .A(mem[355]), .B(n5619), .Y(n793) );
  INVX1 U3891 ( .A(n793), .Y(n4057) );
  AND2X1 U3892 ( .A(mem[338]), .B(n5619), .Y(n776) );
  INVX1 U3893 ( .A(n776), .Y(n4058) );
  AND2X1 U3894 ( .A(mem[329]), .B(n5619), .Y(n767) );
  INVX1 U3895 ( .A(n767), .Y(n4059) );
  AND2X1 U3896 ( .A(mem[323]), .B(n5620), .Y(n759) );
  INVX1 U3897 ( .A(n759), .Y(n4060) );
  AND2X1 U3898 ( .A(mem[308]), .B(n5620), .Y(n744) );
  INVX1 U3899 ( .A(n744), .Y(n4061) );
  AND2X1 U3900 ( .A(mem[294]), .B(n5620), .Y(n730) );
  INVX1 U3901 ( .A(n730), .Y(n4062) );
  AND2X1 U3902 ( .A(mem[272]), .B(n5621), .Y(n706) );
  INVX1 U3903 ( .A(n706), .Y(n4063) );
  AND2X1 U3904 ( .A(mem[259]), .B(n5621), .Y(n693) );
  INVX1 U3905 ( .A(n693), .Y(n4064) );
  AND2X1 U3906 ( .A(mem[254]), .B(n5621), .Y(n688) );
  INVX1 U3907 ( .A(n688), .Y(n4065) );
  AND2X1 U3908 ( .A(mem[239]), .B(n5622), .Y(n671) );
  INVX1 U3909 ( .A(n671), .Y(n4066) );
  AND2X1 U3910 ( .A(mem[224]), .B(n5622), .Y(n656) );
  INVX1 U3911 ( .A(n656), .Y(n4067) );
  AND2X1 U3912 ( .A(mem[210]), .B(n5622), .Y(n642) );
  INVX1 U3913 ( .A(n642), .Y(n4068) );
  AND2X1 U3914 ( .A(mem[199]), .B(n5623), .Y(n629) );
  INVX1 U3915 ( .A(n629), .Y(n4069) );
  AND2X1 U3916 ( .A(mem[184]), .B(n5623), .Y(n614) );
  INVX1 U3917 ( .A(n614), .Y(n4070) );
  AND2X1 U3918 ( .A(mem[170]), .B(n5623), .Y(n600) );
  INVX1 U3919 ( .A(n600), .Y(n4071) );
  AND2X1 U3920 ( .A(mem[151]), .B(n5624), .Y(n579) );
  INVX1 U3921 ( .A(n579), .Y(n4072) );
  AND2X1 U3922 ( .A(mem[134]), .B(n5624), .Y(n562) );
  INVX1 U3923 ( .A(n562), .Y(n4073) );
  AND2X1 U3924 ( .A(mem[125]), .B(n5624), .Y(n553) );
  INVX1 U3925 ( .A(n553), .Y(n4074) );
  AND2X1 U3926 ( .A(mem[111]), .B(n5625), .Y(n537) );
  INVX1 U3927 ( .A(n537), .Y(n4075) );
  AND2X1 U3928 ( .A(mem[94]), .B(n5625), .Y(n520) );
  INVX1 U3929 ( .A(n520), .Y(n4076) );
  AND2X1 U3930 ( .A(mem[85]), .B(n5625), .Y(n511) );
  INVX1 U3931 ( .A(n511), .Y(n4077) );
  AND2X1 U3932 ( .A(mem[66]), .B(n5626), .Y(n490) );
  INVX1 U3933 ( .A(n490), .Y(n4078) );
  AND2X1 U3934 ( .A(mem[45]), .B(n5626), .Y(n469) );
  INVX1 U3935 ( .A(n469), .Y(n4079) );
  AND2X1 U3936 ( .A(mem[41]), .B(n5626), .Y(n465) );
  INVX1 U3937 ( .A(n465), .Y(n4080) );
  AND2X1 U3938 ( .A(mem[27]), .B(n5627), .Y(n435) );
  INVX1 U3939 ( .A(n435), .Y(n4081) );
  AND2X1 U3940 ( .A(mem[10]), .B(n5627), .Y(n401) );
  INVX1 U3941 ( .A(n401), .Y(n4082) );
  AND2X1 U3942 ( .A(mem[1]), .B(n5627), .Y(n383) );
  INVX1 U3943 ( .A(n383), .Y(n4083) );
  INVX1 U3944 ( .A(n1778), .Y(n4084) );
  BUFX2 U3945 ( .A(n1145), .Y(n4085) );
  AND2X1 U3946 ( .A(mem[1304]), .B(n5596), .Y(n1768) );
  INVX1 U3947 ( .A(n1768), .Y(n4086) );
  AND2X1 U3948 ( .A(mem[1287]), .B(n5596), .Y(n1751) );
  INVX1 U3949 ( .A(n1751), .Y(n4087) );
  AND2X1 U3950 ( .A(mem[1262]), .B(n5597), .Y(n1725) );
  INVX1 U3951 ( .A(n1725), .Y(n4088) );
  AND2X1 U3952 ( .A(mem[1245]), .B(n5597), .Y(n1708) );
  INVX1 U3953 ( .A(n1708), .Y(n4089) );
  AND2X1 U3954 ( .A(mem[1220]), .B(n5598), .Y(n1682) );
  INVX1 U3955 ( .A(n1682), .Y(n4090) );
  AND2X1 U3956 ( .A(mem[1203]), .B(n5598), .Y(n1665) );
  INVX1 U3957 ( .A(n1665), .Y(n4091) );
  AND2X1 U3958 ( .A(mem[1188]), .B(n5599), .Y(n1649) );
  INVX1 U3959 ( .A(n1649), .Y(n4092) );
  AND2X1 U3960 ( .A(mem[1178]), .B(n5599), .Y(n1639) );
  INVX1 U3961 ( .A(n1639), .Y(n4093) );
  AND2X1 U3962 ( .A(mem[1157]), .B(n5599), .Y(n1618) );
  INVX1 U3963 ( .A(n1618), .Y(n4094) );
  AND2X1 U3964 ( .A(mem[1133]), .B(n5600), .Y(n1593) );
  INVX1 U3965 ( .A(n1593), .Y(n4095) );
  AND2X1 U3966 ( .A(mem[1120]), .B(n5600), .Y(n1580) );
  INVX1 U3967 ( .A(n1580), .Y(n4096) );
  AND2X1 U3968 ( .A(mem[1115]), .B(n5600), .Y(n1575) );
  INVX1 U3969 ( .A(n1575), .Y(n4097) );
  AND2X1 U3970 ( .A(mem[1102]), .B(n5601), .Y(n1561) );
  INVX1 U3971 ( .A(n1561), .Y(n4098) );
  AND2X1 U3972 ( .A(mem[1087]), .B(n5601), .Y(n1546) );
  INVX1 U3973 ( .A(n1546), .Y(n4099) );
  AND2X1 U3974 ( .A(mem[1073]), .B(n5601), .Y(n1532) );
  INVX1 U3975 ( .A(n1532), .Y(n4100) );
  AND2X1 U3976 ( .A(mem[1060]), .B(n5602), .Y(n1518) );
  INVX1 U3977 ( .A(n1518), .Y(n4101) );
  AND2X1 U3978 ( .A(mem[1045]), .B(n5602), .Y(n1503) );
  INVX1 U3979 ( .A(n1503), .Y(n4102) );
  AND2X1 U3980 ( .A(mem[1031]), .B(n5602), .Y(n1489) );
  INVX1 U3981 ( .A(n1489), .Y(n4103) );
  AND2X1 U3982 ( .A(mem[1018]), .B(n5603), .Y(n1474) );
  INVX1 U3983 ( .A(n1474), .Y(n4104) );
  AND2X1 U3984 ( .A(mem[1003]), .B(n5603), .Y(n1459) );
  INVX1 U3985 ( .A(n1459), .Y(n4105) );
  AND2X1 U3986 ( .A(mem[989]), .B(n5603), .Y(n1445) );
  INVX1 U3987 ( .A(n1445), .Y(n4106) );
  AND2X1 U3988 ( .A(mem[972]), .B(n5604), .Y(n1427) );
  INVX1 U3989 ( .A(n1427), .Y(n4107) );
  AND2X1 U3990 ( .A(mem[955]), .B(n5604), .Y(n1410) );
  INVX1 U3991 ( .A(n1410), .Y(n4108) );
  AND2X1 U3992 ( .A(mem[946]), .B(n5604), .Y(n1401) );
  INVX1 U3993 ( .A(n1401), .Y(n4109) );
  AND2X1 U3994 ( .A(mem[930]), .B(n5605), .Y(n1384) );
  INVX1 U3995 ( .A(n1384), .Y(n4110) );
  AND2X1 U3996 ( .A(mem[913]), .B(n5605), .Y(n1367) );
  INVX1 U3997 ( .A(n1367), .Y(n4111) );
  AND2X1 U3998 ( .A(mem[904]), .B(n5605), .Y(n1358) );
  INVX1 U3999 ( .A(n1358), .Y(n4112) );
  AND2X1 U4000 ( .A(mem[888]), .B(n5606), .Y(n1341) );
  INVX1 U4001 ( .A(n1341), .Y(n4113) );
  AND2X1 U4002 ( .A(mem[871]), .B(n5606), .Y(n1324) );
  INVX1 U4003 ( .A(n1324), .Y(n4114) );
  AND2X1 U4004 ( .A(mem[862]), .B(n5606), .Y(n1315) );
  INVX1 U4005 ( .A(n1315), .Y(n4115) );
  AND2X1 U4006 ( .A(mem[845]), .B(n5607), .Y(n1297) );
  INVX1 U4007 ( .A(n1297), .Y(n4116) );
  AND2X1 U4008 ( .A(mem[824]), .B(n5607), .Y(n1276) );
  INVX1 U4009 ( .A(n1276), .Y(n4117) );
  AND2X1 U4010 ( .A(mem[820]), .B(n5607), .Y(n1272) );
  INVX1 U4011 ( .A(n1272), .Y(n4118) );
  AND2X1 U4012 ( .A(mem[812]), .B(n5608), .Y(n1263) );
  INVX1 U4013 ( .A(n1263), .Y(n4119) );
  AND2X1 U4014 ( .A(mem[795]), .B(n5608), .Y(n1246) );
  INVX1 U4015 ( .A(n1246), .Y(n4120) );
  AND2X1 U4016 ( .A(mem[770]), .B(n5609), .Y(n1220) );
  INVX1 U4017 ( .A(n1220), .Y(n4121) );
  AND2X1 U4018 ( .A(mem[753]), .B(n5609), .Y(n1203) );
  INVX1 U4019 ( .A(n1203), .Y(n4122) );
  AND2X1 U4020 ( .A(mem[728]), .B(n5610), .Y(n1177) );
  INVX1 U4021 ( .A(n1177), .Y(n4123) );
  AND2X1 U4022 ( .A(mem[711]), .B(n5610), .Y(n1160) );
  INVX1 U4023 ( .A(n1160), .Y(n4124) );
  AND2X1 U4024 ( .A(mem[696]), .B(n5611), .Y(n1143) );
  INVX1 U4025 ( .A(n1143), .Y(n4125) );
  AND2X1 U4026 ( .A(mem[686]), .B(n5611), .Y(n1133) );
  INVX1 U4027 ( .A(n1133), .Y(n4126) );
  AND2X1 U4028 ( .A(mem[665]), .B(n5611), .Y(n1112) );
  INVX1 U4029 ( .A(n1112), .Y(n4127) );
  AND2X1 U4030 ( .A(mem[641]), .B(n5612), .Y(n1087) );
  INVX1 U4031 ( .A(n1087), .Y(n4128) );
  AND2X1 U4032 ( .A(mem[628]), .B(n5612), .Y(n1074) );
  INVX1 U4033 ( .A(n1074), .Y(n4129) );
  AND2X1 U4034 ( .A(mem[623]), .B(n5612), .Y(n1069) );
  INVX1 U4035 ( .A(n1069), .Y(n4130) );
  AND2X1 U4036 ( .A(mem[610]), .B(n5613), .Y(n1055) );
  INVX1 U4037 ( .A(n1055), .Y(n4131) );
  AND2X1 U4038 ( .A(mem[595]), .B(n5613), .Y(n1040) );
  INVX1 U4039 ( .A(n1040), .Y(n4132) );
  AND2X1 U4040 ( .A(mem[581]), .B(n5613), .Y(n1026) );
  INVX1 U4041 ( .A(n1026), .Y(n4133) );
  AND2X1 U4042 ( .A(mem[568]), .B(n5614), .Y(n1012) );
  INVX1 U4043 ( .A(n1012), .Y(n4134) );
  AND2X1 U4044 ( .A(mem[553]), .B(n5614), .Y(n997) );
  INVX1 U4045 ( .A(n997), .Y(n4135) );
  AND2X1 U4046 ( .A(mem[539]), .B(n5614), .Y(n983) );
  INVX1 U4047 ( .A(n983), .Y(n4136) );
  AND2X1 U4048 ( .A(mem[526]), .B(n5615), .Y(n969) );
  INVX1 U4049 ( .A(n969), .Y(n4137) );
  AND2X1 U4050 ( .A(mem[511]), .B(n5615), .Y(n954) );
  INVX1 U4051 ( .A(n954), .Y(n4138) );
  AND2X1 U4052 ( .A(mem[497]), .B(n5615), .Y(n940) );
  INVX1 U4053 ( .A(n940), .Y(n4139) );
  AND2X1 U4054 ( .A(mem[480]), .B(n5616), .Y(n922) );
  INVX1 U4055 ( .A(n922), .Y(n4140) );
  AND2X1 U4056 ( .A(mem[463]), .B(n5616), .Y(n905) );
  INVX1 U4057 ( .A(n905), .Y(n4141) );
  AND2X1 U4058 ( .A(mem[454]), .B(n5616), .Y(n896) );
  INVX1 U4059 ( .A(n896), .Y(n4142) );
  AND2X1 U4060 ( .A(mem[438]), .B(n5617), .Y(n879) );
  INVX1 U4061 ( .A(n879), .Y(n4143) );
  AND2X1 U4062 ( .A(mem[421]), .B(n5617), .Y(n862) );
  INVX1 U4063 ( .A(n862), .Y(n4144) );
  AND2X1 U4064 ( .A(mem[412]), .B(n5617), .Y(n853) );
  INVX1 U4065 ( .A(n853), .Y(n4145) );
  AND2X1 U4066 ( .A(mem[396]), .B(n5618), .Y(n836) );
  INVX1 U4067 ( .A(n836), .Y(n4146) );
  AND2X1 U4068 ( .A(mem[379]), .B(n5618), .Y(n819) );
  INVX1 U4069 ( .A(n819), .Y(n4147) );
  AND2X1 U4070 ( .A(mem[370]), .B(n5618), .Y(n810) );
  INVX1 U4071 ( .A(n810), .Y(n4148) );
  AND2X1 U4072 ( .A(mem[353]), .B(n5619), .Y(n791) );
  INVX1 U4073 ( .A(n791), .Y(n4149) );
  AND2X1 U4074 ( .A(mem[332]), .B(n5619), .Y(n770) );
  INVX1 U4075 ( .A(n770), .Y(n4150) );
  AND2X1 U4076 ( .A(mem[328]), .B(n5619), .Y(n766) );
  INVX1 U4077 ( .A(n766), .Y(n4151) );
  AND2X1 U4078 ( .A(mem[313]), .B(n5620), .Y(n749) );
  INVX1 U4079 ( .A(n749), .Y(n4152) );
  AND2X1 U4080 ( .A(mem[300]), .B(n5620), .Y(n736) );
  INVX1 U4081 ( .A(n736), .Y(n4153) );
  AND2X1 U4082 ( .A(mem[295]), .B(n5620), .Y(n731) );
  INVX1 U4083 ( .A(n731), .Y(n4154) );
  AND2X1 U4084 ( .A(mem[282]), .B(n5621), .Y(n716) );
  INVX1 U4085 ( .A(n716), .Y(n4155) );
  AND2X1 U4086 ( .A(mem[267]), .B(n5621), .Y(n701) );
  INVX1 U4087 ( .A(n701), .Y(n4156) );
  AND2X1 U4088 ( .A(mem[253]), .B(n5621), .Y(n687) );
  INVX1 U4089 ( .A(n687), .Y(n4157) );
  AND2X1 U4090 ( .A(mem[240]), .B(n5622), .Y(n672) );
  INVX1 U4091 ( .A(n672), .Y(n4158) );
  AND2X1 U4092 ( .A(mem[225]), .B(n5622), .Y(n657) );
  INVX1 U4093 ( .A(n657), .Y(n4159) );
  AND2X1 U4094 ( .A(mem[211]), .B(n5622), .Y(n643) );
  INVX1 U4095 ( .A(n643), .Y(n4160) );
  AND2X1 U4096 ( .A(mem[198]), .B(n5623), .Y(n628) );
  INVX1 U4097 ( .A(n628), .Y(n4161) );
  AND2X1 U4098 ( .A(mem[183]), .B(n5623), .Y(n613) );
  INVX1 U4099 ( .A(n613), .Y(n4162) );
  AND2X1 U4100 ( .A(mem[169]), .B(n5623), .Y(n599) );
  INVX1 U4101 ( .A(n599), .Y(n4163) );
  AND2X1 U4102 ( .A(mem[152]), .B(n5624), .Y(n580) );
  INVX1 U4103 ( .A(n580), .Y(n4164) );
  AND2X1 U4104 ( .A(mem[135]), .B(n5624), .Y(n563) );
  INVX1 U4105 ( .A(n563), .Y(n4165) );
  AND2X1 U4106 ( .A(mem[126]), .B(n5624), .Y(n554) );
  INVX1 U4107 ( .A(n554), .Y(n4166) );
  AND2X1 U4108 ( .A(mem[110]), .B(n5625), .Y(n536) );
  INVX1 U4109 ( .A(n536), .Y(n4167) );
  AND2X1 U4110 ( .A(mem[93]), .B(n5625), .Y(n519) );
  INVX1 U4111 ( .A(n519), .Y(n4168) );
  AND2X1 U4112 ( .A(mem[84]), .B(n5625), .Y(n510) );
  INVX1 U4113 ( .A(n510), .Y(n4169) );
  AND2X1 U4114 ( .A(mem[68]), .B(n5626), .Y(n492) );
  INVX1 U4115 ( .A(n492), .Y(n4170) );
  AND2X1 U4116 ( .A(mem[51]), .B(n5626), .Y(n475) );
  INVX1 U4117 ( .A(n475), .Y(n4171) );
  AND2X1 U4118 ( .A(mem[42]), .B(n5626), .Y(n466) );
  INVX1 U4119 ( .A(n466), .Y(n4172) );
  AND2X1 U4120 ( .A(mem[25]), .B(n5627), .Y(n431) );
  INVX1 U4121 ( .A(n431), .Y(n4173) );
  AND2X1 U4122 ( .A(mem[4]), .B(n5627), .Y(n389) );
  INVX1 U4123 ( .A(n389), .Y(n4174) );
  AND2X1 U4124 ( .A(mem[0]), .B(n5627), .Y(n381) );
  INVX1 U4125 ( .A(n381), .Y(n4175) );
  INVX1 U4126 ( .A(n1784), .Y(n4176) );
  INVX1 U4127 ( .A(n1832), .Y(n4177) );
  BUFX2 U4128 ( .A(n5721), .Y(empty_bar) );
  BUFX2 U4129 ( .A(n808), .Y(n4179) );
  INVX1 U4130 ( .A(n5500), .Y(n5513) );
  INVX1 U4131 ( .A(n5500), .Y(n5514) );
  INVX1 U4132 ( .A(n5500), .Y(n5515) );
  INVX1 U4133 ( .A(n5499), .Y(n5516) );
  INVX1 U4134 ( .A(n5499), .Y(n5517) );
  INVX1 U4135 ( .A(n5499), .Y(n5518) );
  INVX1 U4136 ( .A(n5498), .Y(n5519) );
  INVX1 U4137 ( .A(n5498), .Y(n5520) );
  INVX1 U4138 ( .A(n5498), .Y(n5521) );
  INVX1 U4139 ( .A(n5497), .Y(n5522) );
  INVX1 U4140 ( .A(n5497), .Y(n5523) );
  INVX1 U4141 ( .A(n5497), .Y(n5524) );
  INVX1 U4142 ( .A(n5496), .Y(n5525) );
  INVX1 U4143 ( .A(n5496), .Y(n5526) );
  INVX1 U4144 ( .A(n5496), .Y(n5527) );
  INVX1 U4145 ( .A(n5495), .Y(n5528) );
  INVX1 U4146 ( .A(n5495), .Y(n5529) );
  INVX1 U4147 ( .A(n5495), .Y(n5530) );
  INVX1 U4148 ( .A(n5502), .Y(n5531) );
  INVX1 U4149 ( .A(n5501), .Y(n5532) );
  INVX1 U4150 ( .A(n5503), .Y(n5533) );
  INVX1 U4151 ( .A(n5493), .Y(n5534) );
  INVX1 U4152 ( .A(n5500), .Y(n5535) );
  INVX1 U4153 ( .A(n5499), .Y(n5536) );
  INVX1 U4154 ( .A(n5492), .Y(n5537) );
  INVX1 U4155 ( .A(n5492), .Y(n5538) );
  INVX1 U4156 ( .A(n5494), .Y(n5539) );
  INVX1 U4157 ( .A(n5494), .Y(n5540) );
  INVX1 U4158 ( .A(n5494), .Y(n5541) );
  INVX1 U4159 ( .A(n5492), .Y(n5542) );
  INVX1 U4160 ( .A(n5494), .Y(n5543) );
  INVX1 U4161 ( .A(n5494), .Y(n5544) );
  INVX1 U4162 ( .A(n5494), .Y(n5545) );
  INVX1 U4163 ( .A(n5492), .Y(n5546) );
  INVX1 U4164 ( .A(n5494), .Y(n5547) );
  INVX1 U4165 ( .A(n5494), .Y(n5548) );
  INVX1 U4166 ( .A(n5493), .Y(n5549) );
  INVX1 U4167 ( .A(n5493), .Y(n5550) );
  INVX1 U4168 ( .A(n5493), .Y(n5551) );
  INVX1 U4169 ( .A(n5503), .Y(n5552) );
  INVX1 U4170 ( .A(n5502), .Y(n5553) );
  INVX1 U4171 ( .A(n5501), .Y(n5554) );
  INVX1 U4172 ( .A(n5492), .Y(n5555) );
  INVX1 U4173 ( .A(n5492), .Y(n5556) );
  INVX1 U4174 ( .A(n5492), .Y(n5557) );
  INVX1 U4175 ( .A(n5561), .Y(n5570) );
  INVX1 U4176 ( .A(n5561), .Y(n5571) );
  INVX1 U4177 ( .A(n5672), .Y(n5572) );
  INVX1 U4178 ( .A(n5672), .Y(n5573) );
  INVX1 U4179 ( .A(n5561), .Y(n5574) );
  INVX1 U4180 ( .A(n5561), .Y(n5575) );
  INVX1 U4181 ( .A(n5672), .Y(n5576) );
  INVX1 U4182 ( .A(n5561), .Y(n5577) );
  INVX1 U4183 ( .A(n5561), .Y(n5578) );
  INVX1 U4184 ( .A(n5672), .Y(n5579) );
  INVX1 U4185 ( .A(n5672), .Y(n5580) );
  INVX1 U4186 ( .A(n5561), .Y(n5581) );
  INVX1 U4187 ( .A(n5561), .Y(n5582) );
  INVX1 U4188 ( .A(n5561), .Y(n5583) );
  INVX1 U4189 ( .A(n5561), .Y(n5584) );
  INVX1 U4190 ( .A(n5561), .Y(n5585) );
  INVX1 U4191 ( .A(n5561), .Y(n5586) );
  INVX1 U4192 ( .A(n5561), .Y(n5587) );
  INVX1 U4193 ( .A(n5671), .Y(n5589) );
  INVX1 U4194 ( .A(n5671), .Y(n5590) );
  INVX1 U4195 ( .A(n5671), .Y(n5591) );
  INVX1 U4196 ( .A(n5671), .Y(n5592) );
  INVX1 U4197 ( .A(n5671), .Y(n5593) );
  INVX1 U4198 ( .A(n5671), .Y(n5594) );
  INVX1 U4199 ( .A(n5671), .Y(n5595) );
  INVX1 U4200 ( .A(n5503), .Y(n5505) );
  INVX1 U4201 ( .A(n5503), .Y(n5506) );
  INVX1 U4202 ( .A(n5502), .Y(n5507) );
  INVX1 U4203 ( .A(n5502), .Y(n5508) );
  INVX1 U4204 ( .A(n5502), .Y(n5509) );
  INVX1 U4205 ( .A(n5501), .Y(n5510) );
  INVX1 U4206 ( .A(n5501), .Y(n5511) );
  INVX1 U4207 ( .A(n5501), .Y(n5512) );
  INVX1 U4208 ( .A(n5503), .Y(n5504) );
  INVX1 U4209 ( .A(n5560), .Y(n5500) );
  INVX1 U4210 ( .A(n5560), .Y(n5499) );
  INVX1 U4211 ( .A(n5560), .Y(n5498) );
  INVX1 U4212 ( .A(n5559), .Y(n5497) );
  INVX1 U4213 ( .A(n5559), .Y(n5496) );
  INVX1 U4214 ( .A(n5559), .Y(n5495) );
  INVX1 U4215 ( .A(n12), .Y(n5494) );
  INVX1 U4216 ( .A(n5560), .Y(n5493) );
  INVX1 U4217 ( .A(n5672), .Y(n5562) );
  INVX1 U4218 ( .A(n5672), .Y(n5563) );
  INVX1 U4219 ( .A(n5561), .Y(n5564) );
  INVX1 U4220 ( .A(n5672), .Y(n5565) );
  INVX1 U4221 ( .A(n5561), .Y(n5566) );
  INVX1 U4222 ( .A(n5561), .Y(n5567) );
  INVX1 U4223 ( .A(n5672), .Y(n5568) );
  INVX1 U4224 ( .A(n5561), .Y(n5569) );
  INVX1 U4225 ( .A(n5492), .Y(n5558) );
  INVX1 U4226 ( .A(n12), .Y(n5492) );
  INVX1 U4227 ( .A(n5674), .Y(n5560) );
  INVX1 U4228 ( .A(n5674), .Y(n5559) );
  INVX1 U4229 ( .A(n12), .Y(n5503) );
  INVX1 U4230 ( .A(n12), .Y(n5502) );
  INVX1 U4231 ( .A(n12), .Y(n5501) );
  INVX1 U4232 ( .A(n462), .Y(n5627) );
  INVX1 U4233 ( .A(n5561), .Y(n5588) );
  INVX1 U4234 ( .A(n13), .Y(n5561) );
  INVX1 U4235 ( .A(n892), .Y(n5617) );
  INVX1 U4236 ( .A(n934), .Y(n5616) );
  INVX1 U4237 ( .A(n976), .Y(n5615) );
  INVX1 U4238 ( .A(n1018), .Y(n5614) );
  INVX1 U4239 ( .A(n1060), .Y(n5613) );
  INVX1 U4240 ( .A(n1102), .Y(n5612) );
  INVX1 U4241 ( .A(n1144), .Y(n5611) );
  INVX1 U4242 ( .A(n1187), .Y(n5610) );
  INVX1 U4243 ( .A(n1229), .Y(n5609) );
  INVX1 U4244 ( .A(n1271), .Y(n5608) );
  INVX1 U4245 ( .A(n1313), .Y(n5607) );
  INVX1 U4246 ( .A(n1355), .Y(n5606) );
  INVX1 U4247 ( .A(n1397), .Y(n5605) );
  INVX1 U4248 ( .A(n1439), .Y(n5604) );
  INVX1 U4249 ( .A(n1481), .Y(n5603) );
  INVX1 U4250 ( .A(n1524), .Y(n5602) );
  INVX1 U4251 ( .A(n1566), .Y(n5601) );
  INVX1 U4252 ( .A(n1608), .Y(n5600) );
  INVX1 U4253 ( .A(n1650), .Y(n5599) );
  INVX1 U4254 ( .A(n1692), .Y(n5598) );
  INVX1 U4255 ( .A(n1734), .Y(n5597) );
  INVX1 U4256 ( .A(n1776), .Y(n5596) );
  INVX1 U4257 ( .A(n506), .Y(n5626) );
  INVX1 U4258 ( .A(n592), .Y(n5624) );
  INVX1 U4259 ( .A(n678), .Y(n5622) );
  INVX1 U4260 ( .A(n764), .Y(n5620) );
  INVX1 U4261 ( .A(n549), .Y(n5625) );
  INVX1 U4262 ( .A(n635), .Y(n5623) );
  INVX1 U4263 ( .A(n721), .Y(n5621) );
  INVX1 U4264 ( .A(n807), .Y(n5619) );
  INVX1 U4265 ( .A(n850), .Y(n5618) );
  INVX1 U4266 ( .A(n5674), .Y(n5673) );
  INVX1 U4267 ( .A(n4181), .Y(n5630) );
  INVX1 U4268 ( .A(n4180), .Y(n5632) );
  INVX1 U4269 ( .A(n4182), .Y(n5629) );
  INVX1 U4270 ( .A(n4183), .Y(n5628) );
  INVX1 U4271 ( .A(n4184), .Y(n5657) );
  INVX1 U4272 ( .A(n4185), .Y(n5656) );
  INVX1 U4273 ( .A(n4186), .Y(n5655) );
  INVX1 U4274 ( .A(n4187), .Y(n5654) );
  INVX1 U4275 ( .A(n4188), .Y(n5653) );
  INVX1 U4276 ( .A(n4189), .Y(n5652) );
  INVX1 U4277 ( .A(n4190), .Y(n5651) );
  INVX1 U4278 ( .A(n4191), .Y(n5650) );
  INVX1 U4279 ( .A(n4192), .Y(n5649) );
  INVX1 U4280 ( .A(n4193), .Y(n5648) );
  INVX1 U4281 ( .A(n4194), .Y(n5647) );
  INVX1 U4282 ( .A(n4195), .Y(n5646) );
  INVX1 U4283 ( .A(n4196), .Y(n5645) );
  INVX1 U4284 ( .A(n4197), .Y(n5644) );
  INVX1 U4285 ( .A(n4198), .Y(n5643) );
  INVX1 U4286 ( .A(n4199), .Y(n5642) );
  INVX1 U4287 ( .A(n4200), .Y(n5641) );
  INVX1 U4288 ( .A(n4201), .Y(n5640) );
  INVX1 U4289 ( .A(n4202), .Y(n5639) );
  INVX1 U4290 ( .A(n4203), .Y(n5638) );
  INVX1 U4291 ( .A(n4204), .Y(n5637) );
  INVX1 U4292 ( .A(n4205), .Y(n5636) );
  INVX1 U4293 ( .A(n4206), .Y(n5635) );
  INVX1 U4294 ( .A(n4207), .Y(n5634) );
  INVX1 U4295 ( .A(n4208), .Y(n5633) );
  INVX1 U4296 ( .A(n4209), .Y(n5631) );
  INVX1 U4297 ( .A(n4210), .Y(n5668) );
  INVX1 U4298 ( .A(n4211), .Y(n5667) );
  INVX1 U4299 ( .A(n4212), .Y(n5666) );
  INVX1 U4300 ( .A(n4213), .Y(n5665) );
  INVX1 U4301 ( .A(n4214), .Y(n5664) );
  INVX1 U4302 ( .A(n4215), .Y(n5663) );
  INVX1 U4303 ( .A(n4216), .Y(n5662) );
  INVX1 U4304 ( .A(n4217), .Y(n5661) );
  INVX1 U4305 ( .A(n4218), .Y(n5660) );
  INVX1 U4306 ( .A(n4219), .Y(n5659) );
  INVX1 U4307 ( .A(n4220), .Y(n5658) );
  INVX1 U4308 ( .A(wr_ptr[2]), .Y(n5719) );
  INVX1 U4309 ( .A(wr_ptr[0]), .Y(n5716) );
  INVX1 U4310 ( .A(n1), .Y(n5675) );
  INVX1 U4311 ( .A(n5451), .Y(n96) );
  INVX1 U4312 ( .A(n2), .Y(n5676) );
  INVX1 U4313 ( .A(n5452), .Y(n95) );
  INVX1 U4314 ( .A(n3), .Y(n5677) );
  INVX1 U4315 ( .A(n5453), .Y(n94) );
  INVX1 U4316 ( .A(n4), .Y(n5678) );
  INVX1 U4317 ( .A(n5454), .Y(n93) );
  INVX1 U4318 ( .A(n5), .Y(n5679) );
  INVX1 U4319 ( .A(n5455), .Y(n92) );
  INVX1 U4320 ( .A(n6), .Y(n5680) );
  INVX1 U4321 ( .A(n5456), .Y(n91) );
  INVX1 U4322 ( .A(n7), .Y(n5681) );
  INVX1 U4323 ( .A(n5457), .Y(n90) );
  INVX1 U4324 ( .A(n8), .Y(n5682) );
  INVX1 U4325 ( .A(n5458), .Y(n89) );
  INVX1 U4326 ( .A(n9), .Y(n5683) );
  INVX1 U4327 ( .A(n5459), .Y(n88) );
  INVX1 U4328 ( .A(n10), .Y(n5684) );
  INVX1 U4329 ( .A(n5460), .Y(n87) );
  INVX1 U4330 ( .A(n11), .Y(n5685) );
  INVX1 U4331 ( .A(n5461), .Y(n86) );
  INVX1 U4332 ( .A(n17), .Y(n5686) );
  INVX1 U4333 ( .A(n5462), .Y(n85) );
  INVX1 U4334 ( .A(n46), .Y(n5711) );
  INVX1 U4335 ( .A(n5487), .Y(n60) );
  INVX1 U4336 ( .A(n47), .Y(n5712) );
  INVX1 U4337 ( .A(n5488), .Y(n59) );
  INVX1 U4338 ( .A(n48), .Y(n5713) );
  INVX1 U4339 ( .A(n5489), .Y(n58) );
  INVX1 U4340 ( .A(n49), .Y(n5714) );
  INVX1 U4341 ( .A(n5490), .Y(n57) );
  INVX1 U4342 ( .A(n50), .Y(n5715) );
  INVX1 U4343 ( .A(n5491), .Y(n56) );
  INVX1 U4344 ( .A(wr_ptr[1]), .Y(n5718) );
  INVX1 U4345 ( .A(wr_ptr[3]), .Y(n5720) );
  INVX1 U4346 ( .A(wr_ptr[4]), .Y(n5717) );
  INVX1 U4347 ( .A(n18), .Y(n5687) );
  INVX1 U4348 ( .A(n5463), .Y(n84) );
  INVX1 U4349 ( .A(n19), .Y(n5688) );
  INVX1 U4350 ( .A(n5464), .Y(n83) );
  INVX1 U4351 ( .A(n24), .Y(n5689) );
  INVX1 U4352 ( .A(n5465), .Y(n82) );
  INVX1 U4353 ( .A(n25), .Y(n5690) );
  INVX1 U4354 ( .A(n5466), .Y(n81) );
  INVX1 U4355 ( .A(n26), .Y(n5691) );
  INVX1 U4356 ( .A(n5467), .Y(n80) );
  INVX1 U4357 ( .A(n27), .Y(n5692) );
  INVX1 U4358 ( .A(n5468), .Y(n79) );
  INVX1 U4359 ( .A(n28), .Y(n5693) );
  INVX1 U4360 ( .A(n5469), .Y(n78) );
  INVX1 U4361 ( .A(n29), .Y(n5694) );
  INVX1 U4362 ( .A(n5470), .Y(n77) );
  INVX1 U4363 ( .A(n30), .Y(n5695) );
  INVX1 U4364 ( .A(n5471), .Y(n76) );
  INVX1 U4365 ( .A(n31), .Y(n5696) );
  INVX1 U4366 ( .A(n5472), .Y(n75) );
  INVX1 U4367 ( .A(n32), .Y(n5697) );
  INVX1 U4368 ( .A(n5473), .Y(n74) );
  INVX1 U4369 ( .A(n33), .Y(n5698) );
  INVX1 U4370 ( .A(n5474), .Y(n73) );
  INVX1 U4371 ( .A(n34), .Y(n5699) );
  INVX1 U4372 ( .A(n5475), .Y(n72) );
  INVX1 U4373 ( .A(n35), .Y(n5700) );
  INVX1 U4374 ( .A(n5476), .Y(n71) );
  INVX1 U4375 ( .A(n36), .Y(n5701) );
  INVX1 U4376 ( .A(n5477), .Y(n70) );
  INVX1 U4377 ( .A(n37), .Y(n5702) );
  INVX1 U4378 ( .A(n5478), .Y(n69) );
  INVX1 U4379 ( .A(n38), .Y(n5703) );
  INVX1 U4380 ( .A(n5479), .Y(n68) );
  INVX1 U4381 ( .A(n39), .Y(n5704) );
  INVX1 U4382 ( .A(n5480), .Y(n67) );
  INVX1 U4383 ( .A(n40), .Y(n5705) );
  INVX1 U4384 ( .A(n5481), .Y(n66) );
  INVX1 U4385 ( .A(n41), .Y(n5706) );
  INVX1 U4386 ( .A(n5482), .Y(n65) );
  INVX1 U4387 ( .A(n42), .Y(n5707) );
  INVX1 U4388 ( .A(n5483), .Y(n64) );
  INVX1 U4389 ( .A(n43), .Y(n5708) );
  INVX1 U4390 ( .A(n5484), .Y(n63) );
  INVX1 U4391 ( .A(n44), .Y(n5709) );
  INVX1 U4392 ( .A(n5485), .Y(n62) );
  INVX1 U4393 ( .A(n45), .Y(n5710) );
  INVX1 U4394 ( .A(n5486), .Y(n61) );
  INVX1 U4395 ( .A(n13), .Y(n5672) );
  INVX1 U4396 ( .A(n14), .Y(n5671) );
  INVX1 U4397 ( .A(n15), .Y(n5670) );
  INVX1 U4398 ( .A(n16), .Y(n5669) );
  INVX1 U4399 ( .A(n12), .Y(n5674) );
  INVX1 U4400 ( .A(sub_93_carry[5]), .Y(fillcount[5]) );
  AND2X1 U4401 ( .A(data_in[36]), .B(reset), .Y(n4180) );
  AND2X1 U4402 ( .A(data_in[38]), .B(reset), .Y(n4181) );
  AND2X1 U4403 ( .A(data_in[39]), .B(reset), .Y(n4182) );
  AND2X1 U4404 ( .A(data_in[40]), .B(reset), .Y(n4183) );
  AND2X1 U4405 ( .A(data_in[11]), .B(reset), .Y(n4184) );
  AND2X1 U4406 ( .A(data_in[12]), .B(reset), .Y(n4185) );
  AND2X1 U4407 ( .A(data_in[13]), .B(reset), .Y(n4186) );
  AND2X1 U4408 ( .A(data_in[14]), .B(reset), .Y(n4187) );
  AND2X1 U4409 ( .A(data_in[15]), .B(reset), .Y(n4188) );
  AND2X1 U4410 ( .A(data_in[16]), .B(reset), .Y(n4189) );
  AND2X1 U4411 ( .A(data_in[17]), .B(reset), .Y(n4190) );
  AND2X1 U4412 ( .A(data_in[18]), .B(reset), .Y(n4191) );
  AND2X1 U4413 ( .A(data_in[19]), .B(reset), .Y(n4192) );
  AND2X1 U4414 ( .A(data_in[20]), .B(reset), .Y(n4193) );
  AND2X1 U4415 ( .A(data_in[21]), .B(reset), .Y(n4194) );
  AND2X1 U4416 ( .A(data_in[22]), .B(reset), .Y(n4195) );
  AND2X1 U4417 ( .A(data_in[23]), .B(reset), .Y(n4196) );
  AND2X1 U4418 ( .A(data_in[24]), .B(reset), .Y(n4197) );
  AND2X1 U4419 ( .A(data_in[25]), .B(reset), .Y(n4198) );
  AND2X1 U4420 ( .A(data_in[26]), .B(reset), .Y(n4199) );
  AND2X1 U4421 ( .A(data_in[27]), .B(reset), .Y(n4200) );
  AND2X1 U4422 ( .A(data_in[28]), .B(reset), .Y(n4201) );
  AND2X1 U4423 ( .A(data_in[29]), .B(reset), .Y(n4202) );
  AND2X1 U4424 ( .A(data_in[30]), .B(reset), .Y(n4203) );
  AND2X1 U4425 ( .A(data_in[31]), .B(reset), .Y(n4204) );
  AND2X1 U4426 ( .A(data_in[32]), .B(reset), .Y(n4205) );
  AND2X1 U4427 ( .A(data_in[33]), .B(reset), .Y(n4206) );
  AND2X1 U4428 ( .A(data_in[34]), .B(reset), .Y(n4207) );
  AND2X1 U4429 ( .A(data_in[35]), .B(reset), .Y(n4208) );
  AND2X1 U4430 ( .A(data_in[37]), .B(reset), .Y(n4209) );
  AND2X1 U4431 ( .A(data_in[0]), .B(reset), .Y(n4210) );
  AND2X1 U4432 ( .A(data_in[1]), .B(reset), .Y(n4211) );
  AND2X1 U4433 ( .A(data_in[2]), .B(reset), .Y(n4212) );
  AND2X1 U4434 ( .A(data_in[3]), .B(reset), .Y(n4213) );
  AND2X1 U4435 ( .A(data_in[4]), .B(reset), .Y(n4214) );
  AND2X1 U4436 ( .A(data_in[5]), .B(reset), .Y(n4215) );
  AND2X1 U4437 ( .A(data_in[6]), .B(reset), .Y(n4216) );
  AND2X1 U4438 ( .A(data_in[7]), .B(reset), .Y(n4217) );
  AND2X1 U4439 ( .A(data_in[8]), .B(reset), .Y(n4218) );
  AND2X1 U4440 ( .A(data_in[9]), .B(reset), .Y(n4219) );
  AND2X1 U4441 ( .A(data_in[10]), .B(reset), .Y(n4220) );
  MUX2X1 U4442 ( .B(n4222), .A(n4223), .S(n5565), .Y(n4221) );
  MUX2X1 U4443 ( .B(n4225), .A(n4226), .S(n5576), .Y(n4224) );
  MUX2X1 U4444 ( .B(n4228), .A(n4229), .S(n5568), .Y(n4227) );
  MUX2X1 U4445 ( .B(n4231), .A(n4232), .S(n5563), .Y(n4230) );
  MUX2X1 U4446 ( .B(n4234), .A(n4235), .S(n15), .Y(n4233) );
  MUX2X1 U4447 ( .B(n4237), .A(n4238), .S(n5562), .Y(n4236) );
  MUX2X1 U4448 ( .B(n4240), .A(n4241), .S(n5562), .Y(n4239) );
  MUX2X1 U4449 ( .B(n4243), .A(n4244), .S(n5562), .Y(n4242) );
  MUX2X1 U4450 ( .B(n4246), .A(n4247), .S(n5562), .Y(n4245) );
  MUX2X1 U4451 ( .B(n4249), .A(n4250), .S(n15), .Y(n4248) );
  MUX2X1 U4452 ( .B(n4252), .A(n4253), .S(n5562), .Y(n4251) );
  MUX2X1 U4453 ( .B(n4255), .A(n4256), .S(n5562), .Y(n4254) );
  MUX2X1 U4454 ( .B(n4258), .A(n4259), .S(n5562), .Y(n4257) );
  MUX2X1 U4455 ( .B(n4261), .A(n4262), .S(n5562), .Y(n4260) );
  MUX2X1 U4456 ( .B(n4264), .A(n4265), .S(n15), .Y(n4263) );
  MUX2X1 U4457 ( .B(n4267), .A(n4268), .S(n5562), .Y(n4266) );
  MUX2X1 U4458 ( .B(n4270), .A(n4271), .S(n5562), .Y(n4269) );
  MUX2X1 U4459 ( .B(n4273), .A(n4274), .S(n5562), .Y(n4272) );
  MUX2X1 U4460 ( .B(n4276), .A(n4277), .S(n5562), .Y(n4275) );
  MUX2X1 U4461 ( .B(n4279), .A(n4280), .S(n15), .Y(n4278) );
  MUX2X1 U4462 ( .B(n4282), .A(n4283), .S(n5563), .Y(n4281) );
  MUX2X1 U4463 ( .B(n4285), .A(n4286), .S(n5563), .Y(n4284) );
  MUX2X1 U4464 ( .B(n4288), .A(n4289), .S(n5563), .Y(n4287) );
  MUX2X1 U4465 ( .B(n4291), .A(n4292), .S(n5563), .Y(n4290) );
  MUX2X1 U4466 ( .B(n4294), .A(n4295), .S(n15), .Y(n4293) );
  MUX2X1 U4467 ( .B(n4297), .A(n4298), .S(n5563), .Y(n4296) );
  MUX2X1 U4468 ( .B(n4300), .A(n4301), .S(n5563), .Y(n4299) );
  MUX2X1 U4469 ( .B(n4303), .A(n4304), .S(n5563), .Y(n4302) );
  MUX2X1 U4470 ( .B(n4306), .A(n4307), .S(n5563), .Y(n4305) );
  MUX2X1 U4471 ( .B(n4309), .A(n4310), .S(n15), .Y(n4308) );
  MUX2X1 U4472 ( .B(n4312), .A(n4313), .S(n5563), .Y(n4311) );
  MUX2X1 U4473 ( .B(n4315), .A(n4316), .S(n5563), .Y(n4314) );
  MUX2X1 U4474 ( .B(n4318), .A(n4319), .S(n5563), .Y(n4317) );
  MUX2X1 U4475 ( .B(n4321), .A(n4322), .S(n5563), .Y(n4320) );
  MUX2X1 U4476 ( .B(n4324), .A(n4325), .S(n15), .Y(n4323) );
  MUX2X1 U4477 ( .B(n4327), .A(n4328), .S(n5564), .Y(n4326) );
  MUX2X1 U4478 ( .B(n4330), .A(n4331), .S(n5564), .Y(n4329) );
  MUX2X1 U4479 ( .B(n4333), .A(n4334), .S(n5564), .Y(n4332) );
  MUX2X1 U4480 ( .B(n4336), .A(n4337), .S(n5564), .Y(n4335) );
  MUX2X1 U4481 ( .B(n4339), .A(n4340), .S(n15), .Y(n4338) );
  MUX2X1 U4482 ( .B(n4342), .A(n4343), .S(n5564), .Y(n4341) );
  MUX2X1 U4483 ( .B(n4345), .A(n4346), .S(n5564), .Y(n4344) );
  MUX2X1 U4484 ( .B(n4348), .A(n4349), .S(n5564), .Y(n4347) );
  MUX2X1 U4485 ( .B(n4351), .A(n4352), .S(n5564), .Y(n4350) );
  MUX2X1 U4486 ( .B(n4354), .A(n4355), .S(n15), .Y(n4353) );
  MUX2X1 U4487 ( .B(n4357), .A(n4358), .S(n5564), .Y(n4356) );
  MUX2X1 U4488 ( .B(n4360), .A(n4361), .S(n5564), .Y(n4359) );
  MUX2X1 U4489 ( .B(n4363), .A(n4364), .S(n5564), .Y(n4362) );
  MUX2X1 U4490 ( .B(n4366), .A(n4367), .S(n5564), .Y(n4365) );
  MUX2X1 U4491 ( .B(n4369), .A(n4370), .S(n15), .Y(n4368) );
  MUX2X1 U4492 ( .B(n4372), .A(n4373), .S(n5565), .Y(n4371) );
  MUX2X1 U4493 ( .B(n4375), .A(n4376), .S(n5565), .Y(n4374) );
  MUX2X1 U4494 ( .B(n4378), .A(n4379), .S(n5565), .Y(n4377) );
  MUX2X1 U4495 ( .B(n4381), .A(n4382), .S(n5565), .Y(n4380) );
  MUX2X1 U4496 ( .B(n4384), .A(n4385), .S(n15), .Y(n4383) );
  MUX2X1 U4497 ( .B(n4387), .A(n4388), .S(n5565), .Y(n4386) );
  MUX2X1 U4498 ( .B(n4390), .A(n4391), .S(n5565), .Y(n4389) );
  MUX2X1 U4499 ( .B(n4393), .A(n4394), .S(n5565), .Y(n4392) );
  MUX2X1 U4500 ( .B(n4396), .A(n4397), .S(n5565), .Y(n4395) );
  MUX2X1 U4501 ( .B(n4399), .A(n4400), .S(n15), .Y(n4398) );
  MUX2X1 U4502 ( .B(n4402), .A(n4403), .S(n5565), .Y(n4401) );
  MUX2X1 U4503 ( .B(n4405), .A(n4406), .S(n5565), .Y(n4404) );
  MUX2X1 U4504 ( .B(n4408), .A(n4409), .S(n5565), .Y(n4407) );
  MUX2X1 U4505 ( .B(n4411), .A(n4412), .S(n5565), .Y(n4410) );
  MUX2X1 U4506 ( .B(n4414), .A(n4415), .S(n15), .Y(n4413) );
  MUX2X1 U4507 ( .B(n4417), .A(n4418), .S(n5566), .Y(n4416) );
  MUX2X1 U4508 ( .B(n4420), .A(n4421), .S(n5566), .Y(n4419) );
  MUX2X1 U4509 ( .B(n4423), .A(n4424), .S(n5566), .Y(n4422) );
  MUX2X1 U4510 ( .B(n4426), .A(n4427), .S(n5566), .Y(n4425) );
  MUX2X1 U4511 ( .B(n4429), .A(n4430), .S(n15), .Y(n4428) );
  MUX2X1 U4512 ( .B(n4432), .A(n4433), .S(n5566), .Y(n4431) );
  MUX2X1 U4513 ( .B(n4435), .A(n4436), .S(n5566), .Y(n4434) );
  MUX2X1 U4514 ( .B(n4438), .A(n4439), .S(n5566), .Y(n4437) );
  MUX2X1 U4515 ( .B(n4441), .A(n4442), .S(n5566), .Y(n4440) );
  MUX2X1 U4516 ( .B(n4444), .A(n4445), .S(n15), .Y(n4443) );
  MUX2X1 U4517 ( .B(n4447), .A(n4448), .S(n5566), .Y(n4446) );
  MUX2X1 U4518 ( .B(n4450), .A(n4451), .S(n5566), .Y(n4449) );
  MUX2X1 U4519 ( .B(n4453), .A(n4454), .S(n5566), .Y(n4452) );
  MUX2X1 U4520 ( .B(n4456), .A(n4457), .S(n5566), .Y(n4455) );
  MUX2X1 U4521 ( .B(n4459), .A(n4460), .S(n15), .Y(n4458) );
  MUX2X1 U4522 ( .B(n4462), .A(n4463), .S(n5567), .Y(n4461) );
  MUX2X1 U4523 ( .B(n4465), .A(n4466), .S(n5567), .Y(n4464) );
  MUX2X1 U4524 ( .B(n4468), .A(n4469), .S(n5567), .Y(n4467) );
  MUX2X1 U4525 ( .B(n4471), .A(n4472), .S(n5567), .Y(n4470) );
  MUX2X1 U4526 ( .B(n4474), .A(n4475), .S(n15), .Y(n4473) );
  MUX2X1 U4527 ( .B(n4477), .A(n4478), .S(n5567), .Y(n4476) );
  MUX2X1 U4528 ( .B(n4480), .A(n4481), .S(n5567), .Y(n4479) );
  MUX2X1 U4529 ( .B(n4483), .A(n4484), .S(n5567), .Y(n4482) );
  MUX2X1 U4530 ( .B(n4486), .A(n4487), .S(n5567), .Y(n4485) );
  MUX2X1 U4531 ( .B(n4489), .A(n4490), .S(n15), .Y(n4488) );
  MUX2X1 U4532 ( .B(n4492), .A(n4493), .S(n5567), .Y(n4491) );
  MUX2X1 U4533 ( .B(n4495), .A(n4496), .S(n5567), .Y(n4494) );
  MUX2X1 U4534 ( .B(n4498), .A(n4499), .S(n5567), .Y(n4497) );
  MUX2X1 U4535 ( .B(n4501), .A(n4502), .S(n5567), .Y(n4500) );
  MUX2X1 U4536 ( .B(n4504), .A(n4505), .S(n15), .Y(n4503) );
  MUX2X1 U4537 ( .B(n4507), .A(n4508), .S(n5568), .Y(n4506) );
  MUX2X1 U4538 ( .B(n4510), .A(n4511), .S(n5568), .Y(n4509) );
  MUX2X1 U4539 ( .B(n4513), .A(n4514), .S(n5568), .Y(n4512) );
  MUX2X1 U4540 ( .B(n4516), .A(n4517), .S(n5568), .Y(n4515) );
  MUX2X1 U4541 ( .B(n4519), .A(n4520), .S(n15), .Y(n4518) );
  MUX2X1 U4542 ( .B(n4522), .A(n4523), .S(n5568), .Y(n4521) );
  MUX2X1 U4543 ( .B(n4525), .A(n4526), .S(n5568), .Y(n4524) );
  MUX2X1 U4544 ( .B(n4528), .A(n4529), .S(n5568), .Y(n4527) );
  MUX2X1 U4545 ( .B(n4531), .A(n4532), .S(n5568), .Y(n4530) );
  MUX2X1 U4546 ( .B(n4534), .A(n4535), .S(n15), .Y(n4533) );
  MUX2X1 U4547 ( .B(n4537), .A(n4538), .S(n5568), .Y(n4536) );
  MUX2X1 U4548 ( .B(n4540), .A(n4541), .S(n5568), .Y(n4539) );
  MUX2X1 U4549 ( .B(n4543), .A(n4544), .S(n5568), .Y(n4542) );
  MUX2X1 U4550 ( .B(n4546), .A(n4547), .S(n5568), .Y(n4545) );
  MUX2X1 U4551 ( .B(n4549), .A(n4550), .S(n15), .Y(n4548) );
  MUX2X1 U4552 ( .B(n4552), .A(n4553), .S(n5569), .Y(n4551) );
  MUX2X1 U4553 ( .B(n4555), .A(n4556), .S(n5569), .Y(n4554) );
  MUX2X1 U4554 ( .B(n4558), .A(n4559), .S(n5569), .Y(n4557) );
  MUX2X1 U4555 ( .B(n4561), .A(n4562), .S(n5569), .Y(n4560) );
  MUX2X1 U4556 ( .B(n4564), .A(n4565), .S(n15), .Y(n4563) );
  MUX2X1 U4557 ( .B(n4567), .A(n4568), .S(n5569), .Y(n4566) );
  MUX2X1 U4558 ( .B(n4570), .A(n4571), .S(n5569), .Y(n4569) );
  MUX2X1 U4559 ( .B(n4573), .A(n4574), .S(n5569), .Y(n4572) );
  MUX2X1 U4560 ( .B(n4576), .A(n4577), .S(n5569), .Y(n4575) );
  MUX2X1 U4561 ( .B(n4579), .A(n4580), .S(n15), .Y(n4578) );
  MUX2X1 U4562 ( .B(n4582), .A(n4583), .S(n5569), .Y(n4581) );
  MUX2X1 U4563 ( .B(n4585), .A(n4586), .S(n5569), .Y(n4584) );
  MUX2X1 U4564 ( .B(n4588), .A(n4589), .S(n5569), .Y(n4587) );
  MUX2X1 U4565 ( .B(n4591), .A(n4592), .S(n5569), .Y(n4590) );
  MUX2X1 U4566 ( .B(n4594), .A(n4595), .S(n15), .Y(n4593) );
  MUX2X1 U4567 ( .B(n4597), .A(n4598), .S(n5570), .Y(n4596) );
  MUX2X1 U4568 ( .B(n4600), .A(n4601), .S(n5570), .Y(n4599) );
  MUX2X1 U4569 ( .B(n4603), .A(n4604), .S(n5570), .Y(n4602) );
  MUX2X1 U4570 ( .B(n4606), .A(n4607), .S(n5570), .Y(n4605) );
  MUX2X1 U4571 ( .B(n4609), .A(n4610), .S(n15), .Y(n4608) );
  MUX2X1 U4572 ( .B(n4612), .A(n4613), .S(n5570), .Y(n4611) );
  MUX2X1 U4573 ( .B(n4615), .A(n4616), .S(n5570), .Y(n4614) );
  MUX2X1 U4574 ( .B(n4618), .A(n4619), .S(n5570), .Y(n4617) );
  MUX2X1 U4575 ( .B(n4621), .A(n4622), .S(n5570), .Y(n4620) );
  MUX2X1 U4576 ( .B(n4624), .A(n4625), .S(n15), .Y(n4623) );
  MUX2X1 U4577 ( .B(n4627), .A(n4628), .S(n5570), .Y(n4626) );
  MUX2X1 U4578 ( .B(n4630), .A(n4631), .S(n5570), .Y(n4629) );
  MUX2X1 U4579 ( .B(n4633), .A(n4634), .S(n5570), .Y(n4632) );
  MUX2X1 U4580 ( .B(n4636), .A(n4637), .S(n5570), .Y(n4635) );
  MUX2X1 U4581 ( .B(n4639), .A(n4640), .S(n15), .Y(n4638) );
  MUX2X1 U4582 ( .B(n4642), .A(n4643), .S(n5571), .Y(n4641) );
  MUX2X1 U4583 ( .B(n4645), .A(n4646), .S(n5571), .Y(n4644) );
  MUX2X1 U4584 ( .B(n4648), .A(n4649), .S(n5571), .Y(n4647) );
  MUX2X1 U4585 ( .B(n4651), .A(n4652), .S(n5571), .Y(n4650) );
  MUX2X1 U4586 ( .B(n4654), .A(n4655), .S(n15), .Y(n4653) );
  MUX2X1 U4587 ( .B(n4657), .A(n4658), .S(n5571), .Y(n4656) );
  MUX2X1 U4588 ( .B(n4660), .A(n4661), .S(n5571), .Y(n4659) );
  MUX2X1 U4589 ( .B(n4663), .A(n4664), .S(n5571), .Y(n4662) );
  MUX2X1 U4590 ( .B(n4666), .A(n4667), .S(n5571), .Y(n4665) );
  MUX2X1 U4591 ( .B(n4669), .A(n4670), .S(n15), .Y(n4668) );
  MUX2X1 U4592 ( .B(n4672), .A(n4673), .S(n5571), .Y(n4671) );
  MUX2X1 U4593 ( .B(n4675), .A(n4676), .S(n5571), .Y(n4674) );
  MUX2X1 U4594 ( .B(n4678), .A(n4679), .S(n5571), .Y(n4677) );
  MUX2X1 U4595 ( .B(n4681), .A(n4682), .S(n5571), .Y(n4680) );
  MUX2X1 U4596 ( .B(n4684), .A(n4685), .S(n15), .Y(n4683) );
  MUX2X1 U4597 ( .B(n4687), .A(n4688), .S(n5572), .Y(n4686) );
  MUX2X1 U4598 ( .B(n4690), .A(n4691), .S(n5572), .Y(n4689) );
  MUX2X1 U4599 ( .B(n4693), .A(n4694), .S(n5572), .Y(n4692) );
  MUX2X1 U4600 ( .B(n4696), .A(n4697), .S(n5572), .Y(n4695) );
  MUX2X1 U4601 ( .B(n4699), .A(n4700), .S(n15), .Y(n4698) );
  MUX2X1 U4602 ( .B(n4702), .A(n4703), .S(n5572), .Y(n4701) );
  MUX2X1 U4603 ( .B(n4705), .A(n4706), .S(n5572), .Y(n4704) );
  MUX2X1 U4604 ( .B(n4708), .A(n4709), .S(n5572), .Y(n4707) );
  MUX2X1 U4605 ( .B(n4711), .A(n4712), .S(n5572), .Y(n4710) );
  MUX2X1 U4606 ( .B(n4714), .A(n4715), .S(n15), .Y(n4713) );
  MUX2X1 U4607 ( .B(n4717), .A(n4718), .S(n5572), .Y(n4716) );
  MUX2X1 U4608 ( .B(n4720), .A(n4721), .S(n5572), .Y(n4719) );
  MUX2X1 U4609 ( .B(n4723), .A(n4724), .S(n5572), .Y(n4722) );
  MUX2X1 U4610 ( .B(n4726), .A(n4727), .S(n5572), .Y(n4725) );
  MUX2X1 U4611 ( .B(n4729), .A(n4730), .S(n15), .Y(n4728) );
  MUX2X1 U4612 ( .B(n4732), .A(n4733), .S(n5573), .Y(n4731) );
  MUX2X1 U4613 ( .B(n4735), .A(n4736), .S(n5573), .Y(n4734) );
  MUX2X1 U4614 ( .B(n4738), .A(n4739), .S(n5573), .Y(n4737) );
  MUX2X1 U4615 ( .B(n4741), .A(n4742), .S(n5573), .Y(n4740) );
  MUX2X1 U4616 ( .B(n4744), .A(n4745), .S(n15), .Y(n4743) );
  MUX2X1 U4617 ( .B(n4747), .A(n4748), .S(n5573), .Y(n4746) );
  MUX2X1 U4618 ( .B(n4750), .A(n4751), .S(n5573), .Y(n4749) );
  MUX2X1 U4619 ( .B(n4753), .A(n4754), .S(n5573), .Y(n4752) );
  MUX2X1 U4620 ( .B(n4756), .A(n4757), .S(n5573), .Y(n4755) );
  MUX2X1 U4621 ( .B(n4759), .A(n4760), .S(n15), .Y(n4758) );
  MUX2X1 U4622 ( .B(n4762), .A(n4763), .S(n5573), .Y(n4761) );
  MUX2X1 U4623 ( .B(n4765), .A(n4766), .S(n5573), .Y(n4764) );
  MUX2X1 U4624 ( .B(n4768), .A(n4769), .S(n5573), .Y(n4767) );
  MUX2X1 U4625 ( .B(n4771), .A(n4772), .S(n5573), .Y(n4770) );
  MUX2X1 U4626 ( .B(n4774), .A(n4775), .S(n15), .Y(n4773) );
  MUX2X1 U4627 ( .B(n4777), .A(n4778), .S(n5574), .Y(n4776) );
  MUX2X1 U4628 ( .B(n4780), .A(n4781), .S(n5574), .Y(n4779) );
  MUX2X1 U4629 ( .B(n4783), .A(n4784), .S(n5574), .Y(n4782) );
  MUX2X1 U4630 ( .B(n4786), .A(n4787), .S(n5574), .Y(n4785) );
  MUX2X1 U4631 ( .B(n4789), .A(n4790), .S(n15), .Y(n4788) );
  MUX2X1 U4632 ( .B(n4792), .A(n4793), .S(n5574), .Y(n4791) );
  MUX2X1 U4633 ( .B(n4795), .A(n4796), .S(n5574), .Y(n4794) );
  MUX2X1 U4634 ( .B(n4798), .A(n4799), .S(n5574), .Y(n4797) );
  MUX2X1 U4635 ( .B(n4801), .A(n4802), .S(n5574), .Y(n4800) );
  MUX2X1 U4636 ( .B(n4804), .A(n4805), .S(n15), .Y(n4803) );
  MUX2X1 U4637 ( .B(n4807), .A(n4808), .S(n5574), .Y(n4806) );
  MUX2X1 U4638 ( .B(n4810), .A(n4811), .S(n5574), .Y(n4809) );
  MUX2X1 U4639 ( .B(n4813), .A(n4814), .S(n5574), .Y(n4812) );
  MUX2X1 U4640 ( .B(n4816), .A(n4817), .S(n5574), .Y(n4815) );
  MUX2X1 U4641 ( .B(n4819), .A(n4820), .S(n15), .Y(n4818) );
  MUX2X1 U4642 ( .B(n4822), .A(n4823), .S(n5575), .Y(n4821) );
  MUX2X1 U4643 ( .B(n4825), .A(n4826), .S(n5575), .Y(n4824) );
  MUX2X1 U4644 ( .B(n4828), .A(n4829), .S(n5575), .Y(n4827) );
  MUX2X1 U4645 ( .B(n4831), .A(n4832), .S(n5575), .Y(n4830) );
  MUX2X1 U4646 ( .B(n4834), .A(n4835), .S(n15), .Y(n4833) );
  MUX2X1 U4647 ( .B(n4837), .A(n4838), .S(n5575), .Y(n4836) );
  MUX2X1 U4648 ( .B(n4840), .A(n4841), .S(n5575), .Y(n4839) );
  MUX2X1 U4649 ( .B(n4843), .A(n4844), .S(n5575), .Y(n4842) );
  MUX2X1 U4650 ( .B(n4846), .A(n4847), .S(n5575), .Y(n4845) );
  MUX2X1 U4651 ( .B(n4849), .A(n4850), .S(n15), .Y(n4848) );
  MUX2X1 U4652 ( .B(n4852), .A(n4853), .S(n5575), .Y(n4851) );
  MUX2X1 U4653 ( .B(n4855), .A(n4856), .S(n5575), .Y(n4854) );
  MUX2X1 U4654 ( .B(n4858), .A(n4859), .S(n5575), .Y(n4857) );
  MUX2X1 U4655 ( .B(n4861), .A(n4862), .S(n5575), .Y(n4860) );
  MUX2X1 U4656 ( .B(n4864), .A(n4865), .S(n15), .Y(n4863) );
  MUX2X1 U4657 ( .B(n4867), .A(n4868), .S(n5576), .Y(n4866) );
  MUX2X1 U4658 ( .B(n4870), .A(n4871), .S(n5576), .Y(n4869) );
  MUX2X1 U4659 ( .B(n4873), .A(n4874), .S(n5576), .Y(n4872) );
  MUX2X1 U4660 ( .B(n4876), .A(n4877), .S(n5576), .Y(n4875) );
  MUX2X1 U4661 ( .B(n4879), .A(n4880), .S(n15), .Y(n4878) );
  MUX2X1 U4662 ( .B(n4882), .A(n4883), .S(n5576), .Y(n4881) );
  MUX2X1 U4663 ( .B(n4885), .A(n4886), .S(n5576), .Y(n4884) );
  MUX2X1 U4664 ( .B(n4888), .A(n4889), .S(n5576), .Y(n4887) );
  MUX2X1 U4665 ( .B(n4891), .A(n4892), .S(n5576), .Y(n4890) );
  MUX2X1 U4666 ( .B(n4894), .A(n4895), .S(n15), .Y(n4893) );
  MUX2X1 U4667 ( .B(n4897), .A(n4898), .S(n5576), .Y(n4896) );
  MUX2X1 U4668 ( .B(n4900), .A(n4901), .S(n5576), .Y(n4899) );
  MUX2X1 U4669 ( .B(n4903), .A(n4904), .S(n5576), .Y(n4902) );
  MUX2X1 U4670 ( .B(n4906), .A(n4907), .S(n5576), .Y(n4905) );
  MUX2X1 U4671 ( .B(n4909), .A(n4910), .S(n15), .Y(n4908) );
  MUX2X1 U4672 ( .B(n4912), .A(n4913), .S(n5577), .Y(n4911) );
  MUX2X1 U4673 ( .B(n4915), .A(n4916), .S(n5577), .Y(n4914) );
  MUX2X1 U4674 ( .B(n4918), .A(n4919), .S(n5577), .Y(n4917) );
  MUX2X1 U4675 ( .B(n4921), .A(n4922), .S(n5577), .Y(n4920) );
  MUX2X1 U4676 ( .B(n4924), .A(n4925), .S(n15), .Y(n4923) );
  MUX2X1 U4677 ( .B(n4927), .A(n4928), .S(n5577), .Y(n4926) );
  MUX2X1 U4678 ( .B(n4930), .A(n4931), .S(n5577), .Y(n4929) );
  MUX2X1 U4679 ( .B(n4933), .A(n4934), .S(n5577), .Y(n4932) );
  MUX2X1 U4680 ( .B(n4936), .A(n4937), .S(n5577), .Y(n4935) );
  MUX2X1 U4681 ( .B(n4939), .A(n4940), .S(n15), .Y(n4938) );
  MUX2X1 U4682 ( .B(n4942), .A(n4943), .S(n5577), .Y(n4941) );
  MUX2X1 U4683 ( .B(n4945), .A(n4946), .S(n5577), .Y(n4944) );
  MUX2X1 U4684 ( .B(n4948), .A(n4949), .S(n5577), .Y(n4947) );
  MUX2X1 U4685 ( .B(n4951), .A(n4952), .S(n5577), .Y(n4950) );
  MUX2X1 U4686 ( .B(n4954), .A(n4955), .S(n15), .Y(n4953) );
  MUX2X1 U4687 ( .B(n4957), .A(n4958), .S(n5578), .Y(n4956) );
  MUX2X1 U4688 ( .B(n4960), .A(n4961), .S(n5578), .Y(n4959) );
  MUX2X1 U4689 ( .B(n4963), .A(n4964), .S(n5578), .Y(n4962) );
  MUX2X1 U4690 ( .B(n4966), .A(n4967), .S(n5578), .Y(n4965) );
  MUX2X1 U4691 ( .B(n4969), .A(n4970), .S(n15), .Y(n4968) );
  MUX2X1 U4692 ( .B(n4972), .A(n4973), .S(n5578), .Y(n4971) );
  MUX2X1 U4693 ( .B(n4975), .A(n4976), .S(n5578), .Y(n4974) );
  MUX2X1 U4694 ( .B(n4978), .A(n4979), .S(n5578), .Y(n4977) );
  MUX2X1 U4695 ( .B(n4981), .A(n4982), .S(n5578), .Y(n4980) );
  MUX2X1 U4696 ( .B(n4984), .A(n4985), .S(n15), .Y(n4983) );
  MUX2X1 U4697 ( .B(n4987), .A(n4988), .S(n5578), .Y(n4986) );
  MUX2X1 U4698 ( .B(n4990), .A(n4991), .S(n5578), .Y(n4989) );
  MUX2X1 U4699 ( .B(n4993), .A(n4994), .S(n5578), .Y(n4992) );
  MUX2X1 U4700 ( .B(n4996), .A(n4997), .S(n5578), .Y(n4995) );
  MUX2X1 U4701 ( .B(n4999), .A(n5000), .S(n15), .Y(n4998) );
  MUX2X1 U4702 ( .B(n5002), .A(n5003), .S(n5579), .Y(n5001) );
  MUX2X1 U4703 ( .B(n5005), .A(n5006), .S(n5579), .Y(n5004) );
  MUX2X1 U4704 ( .B(n5008), .A(n5009), .S(n5579), .Y(n5007) );
  MUX2X1 U4705 ( .B(n5011), .A(n5012), .S(n5579), .Y(n5010) );
  MUX2X1 U4706 ( .B(n5014), .A(n5015), .S(n15), .Y(n5013) );
  MUX2X1 U4707 ( .B(n5017), .A(n5018), .S(n5579), .Y(n5016) );
  MUX2X1 U4708 ( .B(n5020), .A(n5021), .S(n5579), .Y(n5019) );
  MUX2X1 U4709 ( .B(n5023), .A(n5024), .S(n5579), .Y(n5022) );
  MUX2X1 U4710 ( .B(n5026), .A(n5027), .S(n5579), .Y(n5025) );
  MUX2X1 U4711 ( .B(n5029), .A(n5030), .S(n15), .Y(n5028) );
  MUX2X1 U4712 ( .B(n5032), .A(n5033), .S(n5579), .Y(n5031) );
  MUX2X1 U4713 ( .B(n5035), .A(n5036), .S(n5579), .Y(n5034) );
  MUX2X1 U4714 ( .B(n5038), .A(n5039), .S(n5579), .Y(n5037) );
  MUX2X1 U4715 ( .B(n5041), .A(n5042), .S(n5579), .Y(n5040) );
  MUX2X1 U4716 ( .B(n5044), .A(n5045), .S(n15), .Y(n5043) );
  MUX2X1 U4717 ( .B(n5047), .A(n5048), .S(n5580), .Y(n5046) );
  MUX2X1 U4718 ( .B(n5050), .A(n5051), .S(n5580), .Y(n5049) );
  MUX2X1 U4719 ( .B(n5053), .A(n5054), .S(n5580), .Y(n5052) );
  MUX2X1 U4720 ( .B(n5056), .A(n5057), .S(n5580), .Y(n5055) );
  MUX2X1 U4721 ( .B(n5059), .A(n5060), .S(n15), .Y(n5058) );
  MUX2X1 U4722 ( .B(n5062), .A(n5063), .S(n5580), .Y(n5061) );
  MUX2X1 U4723 ( .B(n5065), .A(n5066), .S(n5580), .Y(n5064) );
  MUX2X1 U4724 ( .B(n5068), .A(n5069), .S(n5580), .Y(n5067) );
  MUX2X1 U4725 ( .B(n5071), .A(n5072), .S(n5580), .Y(n5070) );
  MUX2X1 U4726 ( .B(n5074), .A(n5075), .S(n15), .Y(n5073) );
  MUX2X1 U4727 ( .B(n5077), .A(n5078), .S(n5580), .Y(n5076) );
  MUX2X1 U4728 ( .B(n5080), .A(n5081), .S(n5580), .Y(n5079) );
  MUX2X1 U4729 ( .B(n5083), .A(n5084), .S(n5580), .Y(n5082) );
  MUX2X1 U4730 ( .B(n5086), .A(n5087), .S(n5580), .Y(n5085) );
  MUX2X1 U4731 ( .B(n5089), .A(n5090), .S(n15), .Y(n5088) );
  MUX2X1 U4732 ( .B(n5092), .A(n5093), .S(n5581), .Y(n5091) );
  MUX2X1 U4733 ( .B(n5095), .A(n5096), .S(n5581), .Y(n5094) );
  MUX2X1 U4734 ( .B(n5098), .A(n5099), .S(n5581), .Y(n5097) );
  MUX2X1 U4735 ( .B(n5101), .A(n5102), .S(n5581), .Y(n5100) );
  MUX2X1 U4736 ( .B(n5104), .A(n5105), .S(n15), .Y(n5103) );
  MUX2X1 U4737 ( .B(n5107), .A(n5108), .S(n5581), .Y(n5106) );
  MUX2X1 U4738 ( .B(n5110), .A(n5111), .S(n5581), .Y(n5109) );
  MUX2X1 U4739 ( .B(n5113), .A(n5114), .S(n5581), .Y(n5112) );
  MUX2X1 U4740 ( .B(n5116), .A(n5117), .S(n5581), .Y(n5115) );
  MUX2X1 U4741 ( .B(n5119), .A(n5120), .S(n15), .Y(n5118) );
  MUX2X1 U4742 ( .B(n5122), .A(n5123), .S(n5581), .Y(n5121) );
  MUX2X1 U4743 ( .B(n5125), .A(n5126), .S(n5581), .Y(n5124) );
  MUX2X1 U4744 ( .B(n5128), .A(n5129), .S(n5581), .Y(n5127) );
  MUX2X1 U4745 ( .B(n5131), .A(n5132), .S(n5581), .Y(n5130) );
  MUX2X1 U4746 ( .B(n5134), .A(n5135), .S(n15), .Y(n5133) );
  MUX2X1 U4747 ( .B(n5137), .A(n5138), .S(n5582), .Y(n5136) );
  MUX2X1 U4748 ( .B(n5140), .A(n5141), .S(n5582), .Y(n5139) );
  MUX2X1 U4749 ( .B(n5143), .A(n5144), .S(n5582), .Y(n5142) );
  MUX2X1 U4750 ( .B(n5146), .A(n5147), .S(n5582), .Y(n5145) );
  MUX2X1 U4751 ( .B(n5149), .A(n5150), .S(n15), .Y(n5148) );
  MUX2X1 U4752 ( .B(n5152), .A(n5153), .S(n5582), .Y(n5151) );
  MUX2X1 U4753 ( .B(n5155), .A(n5156), .S(n5582), .Y(n5154) );
  MUX2X1 U4754 ( .B(n5158), .A(n5159), .S(n5582), .Y(n5157) );
  MUX2X1 U4755 ( .B(n5161), .A(n5162), .S(n5582), .Y(n5160) );
  MUX2X1 U4756 ( .B(n5164), .A(n5165), .S(n15), .Y(n5163) );
  MUX2X1 U4757 ( .B(n5167), .A(n5168), .S(n5582), .Y(n5166) );
  MUX2X1 U4758 ( .B(n5170), .A(n5171), .S(n5582), .Y(n5169) );
  MUX2X1 U4759 ( .B(n5173), .A(n5174), .S(n5582), .Y(n5172) );
  MUX2X1 U4760 ( .B(n5176), .A(n5177), .S(n5582), .Y(n5175) );
  MUX2X1 U4761 ( .B(n5179), .A(n5180), .S(n15), .Y(n5178) );
  MUX2X1 U4762 ( .B(n5182), .A(n5183), .S(n5583), .Y(n5181) );
  MUX2X1 U4763 ( .B(n5185), .A(n5186), .S(n5583), .Y(n5184) );
  MUX2X1 U4764 ( .B(n5188), .A(n5189), .S(n5583), .Y(n5187) );
  MUX2X1 U4765 ( .B(n5191), .A(n5192), .S(n5583), .Y(n5190) );
  MUX2X1 U4766 ( .B(n5194), .A(n5195), .S(n15), .Y(n5193) );
  MUX2X1 U4767 ( .B(n5197), .A(n5198), .S(n5583), .Y(n5196) );
  MUX2X1 U4768 ( .B(n5200), .A(n5201), .S(n5583), .Y(n5199) );
  MUX2X1 U4769 ( .B(n5203), .A(n5204), .S(n5583), .Y(n5202) );
  MUX2X1 U4770 ( .B(n5206), .A(n5207), .S(n5583), .Y(n5205) );
  MUX2X1 U4771 ( .B(n5209), .A(n5210), .S(n15), .Y(n5208) );
  MUX2X1 U4772 ( .B(n5212), .A(n5213), .S(n5583), .Y(n5211) );
  MUX2X1 U4773 ( .B(n5215), .A(n5216), .S(n5583), .Y(n5214) );
  MUX2X1 U4774 ( .B(n5218), .A(n5219), .S(n5583), .Y(n5217) );
  MUX2X1 U4775 ( .B(n5221), .A(n5222), .S(n5583), .Y(n5220) );
  MUX2X1 U4776 ( .B(n5224), .A(n5225), .S(n15), .Y(n5223) );
  MUX2X1 U4777 ( .B(n5227), .A(n5228), .S(n5584), .Y(n5226) );
  MUX2X1 U4778 ( .B(n5230), .A(n5231), .S(n5584), .Y(n5229) );
  MUX2X1 U4779 ( .B(n5233), .A(n5234), .S(n5584), .Y(n5232) );
  MUX2X1 U4780 ( .B(n5236), .A(n5237), .S(n5584), .Y(n5235) );
  MUX2X1 U4781 ( .B(n5239), .A(n5240), .S(n15), .Y(n5238) );
  MUX2X1 U4782 ( .B(n5242), .A(n5243), .S(n5584), .Y(n5241) );
  MUX2X1 U4783 ( .B(n5245), .A(n5246), .S(n5584), .Y(n5244) );
  MUX2X1 U4784 ( .B(n5248), .A(n5249), .S(n5584), .Y(n5247) );
  MUX2X1 U4785 ( .B(n5251), .A(n5252), .S(n5584), .Y(n5250) );
  MUX2X1 U4786 ( .B(n5254), .A(n5255), .S(n15), .Y(n5253) );
  MUX2X1 U4787 ( .B(n5257), .A(n5258), .S(n5584), .Y(n5256) );
  MUX2X1 U4788 ( .B(n5260), .A(n5261), .S(n5584), .Y(n5259) );
  MUX2X1 U4789 ( .B(n5263), .A(n5264), .S(n5584), .Y(n5262) );
  MUX2X1 U4790 ( .B(n5266), .A(n5267), .S(n5584), .Y(n5265) );
  MUX2X1 U4791 ( .B(n5269), .A(n5270), .S(n15), .Y(n5268) );
  MUX2X1 U4792 ( .B(n5272), .A(n5273), .S(n5585), .Y(n5271) );
  MUX2X1 U4793 ( .B(n5275), .A(n5276), .S(n5585), .Y(n5274) );
  MUX2X1 U4794 ( .B(n5278), .A(n5279), .S(n5585), .Y(n5277) );
  MUX2X1 U4795 ( .B(n5281), .A(n5282), .S(n5585), .Y(n5280) );
  MUX2X1 U4796 ( .B(n5284), .A(n5285), .S(n15), .Y(n5283) );
  MUX2X1 U4797 ( .B(n5287), .A(n5288), .S(n5585), .Y(n5286) );
  MUX2X1 U4798 ( .B(n5290), .A(n5291), .S(n5585), .Y(n5289) );
  MUX2X1 U4799 ( .B(n5293), .A(n5294), .S(n5585), .Y(n5292) );
  MUX2X1 U4800 ( .B(n5296), .A(n5297), .S(n5585), .Y(n5295) );
  MUX2X1 U4801 ( .B(n5299), .A(n5300), .S(n15), .Y(n5298) );
  MUX2X1 U4802 ( .B(n5302), .A(n5303), .S(n5585), .Y(n5301) );
  MUX2X1 U4803 ( .B(n5305), .A(n5306), .S(n5585), .Y(n5304) );
  MUX2X1 U4804 ( .B(n5308), .A(n5309), .S(n5585), .Y(n5307) );
  MUX2X1 U4805 ( .B(n5311), .A(n5312), .S(n5585), .Y(n5310) );
  MUX2X1 U4806 ( .B(n5314), .A(n5315), .S(n15), .Y(n5313) );
  MUX2X1 U4807 ( .B(n5317), .A(n5318), .S(n5586), .Y(n5316) );
  MUX2X1 U4808 ( .B(n5320), .A(n5321), .S(n5586), .Y(n5319) );
  MUX2X1 U4809 ( .B(n5323), .A(n5324), .S(n5586), .Y(n5322) );
  MUX2X1 U4810 ( .B(n5326), .A(n5327), .S(n5586), .Y(n5325) );
  MUX2X1 U4811 ( .B(n5329), .A(n5330), .S(n15), .Y(n5328) );
  MUX2X1 U4812 ( .B(n5332), .A(n5333), .S(n5586), .Y(n5331) );
  MUX2X1 U4813 ( .B(n5335), .A(n5336), .S(n5586), .Y(n5334) );
  MUX2X1 U4814 ( .B(n5338), .A(n5339), .S(n5586), .Y(n5337) );
  MUX2X1 U4815 ( .B(n5341), .A(n5342), .S(n5586), .Y(n5340) );
  MUX2X1 U4816 ( .B(n5344), .A(n5345), .S(n15), .Y(n5343) );
  MUX2X1 U4817 ( .B(n5347), .A(n5348), .S(n5586), .Y(n5346) );
  MUX2X1 U4818 ( .B(n5350), .A(n5351), .S(n5586), .Y(n5349) );
  MUX2X1 U4819 ( .B(n5353), .A(n5354), .S(n5586), .Y(n5352) );
  MUX2X1 U4820 ( .B(n5356), .A(n5357), .S(n5586), .Y(n5355) );
  MUX2X1 U4821 ( .B(n5359), .A(n5360), .S(n15), .Y(n5358) );
  MUX2X1 U4822 ( .B(n5362), .A(n5363), .S(n5587), .Y(n5361) );
  MUX2X1 U4823 ( .B(n5365), .A(n5366), .S(n5587), .Y(n5364) );
  MUX2X1 U4824 ( .B(n5368), .A(n5369), .S(n5587), .Y(n5367) );
  MUX2X1 U4825 ( .B(n5371), .A(n5372), .S(n5587), .Y(n5370) );
  MUX2X1 U4826 ( .B(n5374), .A(n5375), .S(n15), .Y(n5373) );
  MUX2X1 U4827 ( .B(n5377), .A(n5378), .S(n5587), .Y(n5376) );
  MUX2X1 U4828 ( .B(n5380), .A(n5381), .S(n5587), .Y(n5379) );
  MUX2X1 U4829 ( .B(n5383), .A(n5384), .S(n5587), .Y(n5382) );
  MUX2X1 U4830 ( .B(n5386), .A(n5387), .S(n5587), .Y(n5385) );
  MUX2X1 U4831 ( .B(n5389), .A(n5390), .S(n15), .Y(n5388) );
  MUX2X1 U4832 ( .B(n5392), .A(n5393), .S(n5587), .Y(n5391) );
  MUX2X1 U4833 ( .B(n5395), .A(n5396), .S(n5587), .Y(n5394) );
  MUX2X1 U4834 ( .B(n5398), .A(n5399), .S(n5587), .Y(n5397) );
  MUX2X1 U4835 ( .B(n5401), .A(n5402), .S(n5587), .Y(n5400) );
  MUX2X1 U4836 ( .B(n5404), .A(n5405), .S(n15), .Y(n5403) );
  MUX2X1 U4837 ( .B(n5407), .A(n5408), .S(n5588), .Y(n5406) );
  MUX2X1 U4838 ( .B(n5410), .A(n5411), .S(n5588), .Y(n5409) );
  MUX2X1 U4839 ( .B(n5413), .A(n5414), .S(n5588), .Y(n5412) );
  MUX2X1 U4840 ( .B(n5416), .A(n5417), .S(n5588), .Y(n5415) );
  MUX2X1 U4841 ( .B(n5419), .A(n5420), .S(n15), .Y(n5418) );
  MUX2X1 U4842 ( .B(n5422), .A(n5423), .S(n5588), .Y(n5421) );
  MUX2X1 U4843 ( .B(n5425), .A(n5426), .S(n5588), .Y(n5424) );
  MUX2X1 U4844 ( .B(n5428), .A(n5429), .S(n5588), .Y(n5427) );
  MUX2X1 U4845 ( .B(n5431), .A(n5432), .S(n5588), .Y(n5430) );
  MUX2X1 U4846 ( .B(n5434), .A(n5435), .S(n15), .Y(n5433) );
  MUX2X1 U4847 ( .B(n5437), .A(n5438), .S(n5588), .Y(n5436) );
  MUX2X1 U4848 ( .B(n5440), .A(n5441), .S(n5588), .Y(n5439) );
  MUX2X1 U4849 ( .B(n5443), .A(n5444), .S(n5588), .Y(n5442) );
  MUX2X1 U4850 ( .B(n5446), .A(n5447), .S(n5588), .Y(n5445) );
  MUX2X1 U4851 ( .B(n5449), .A(n5450), .S(n15), .Y(n5448) );
  MUX2X1 U4852 ( .B(mem[1230]), .A(mem[1271]), .S(n5504), .Y(n4223) );
  MUX2X1 U4853 ( .B(mem[1148]), .A(mem[1189]), .S(n5504), .Y(n4222) );
  MUX2X1 U4854 ( .B(mem[1066]), .A(mem[1107]), .S(n5504), .Y(n4226) );
  MUX2X1 U4855 ( .B(mem[984]), .A(mem[1025]), .S(n5504), .Y(n4225) );
  MUX2X1 U4856 ( .B(n4224), .A(n4221), .S(n14), .Y(n4235) );
  MUX2X1 U4857 ( .B(mem[902]), .A(mem[943]), .S(n5504), .Y(n4229) );
  MUX2X1 U4858 ( .B(mem[820]), .A(mem[861]), .S(n5504), .Y(n4228) );
  MUX2X1 U4859 ( .B(mem[738]), .A(mem[779]), .S(n5504), .Y(n4232) );
  MUX2X1 U4860 ( .B(mem[656]), .A(mem[697]), .S(n5504), .Y(n4231) );
  MUX2X1 U4861 ( .B(n4230), .A(n4227), .S(n14), .Y(n4234) );
  MUX2X1 U4862 ( .B(mem[574]), .A(mem[615]), .S(n5505), .Y(n4238) );
  MUX2X1 U4863 ( .B(mem[492]), .A(mem[533]), .S(n5505), .Y(n4237) );
  MUX2X1 U4864 ( .B(mem[410]), .A(mem[451]), .S(n5505), .Y(n4241) );
  MUX2X1 U4865 ( .B(mem[328]), .A(mem[369]), .S(n5505), .Y(n4240) );
  MUX2X1 U4866 ( .B(n4239), .A(n4236), .S(n14), .Y(n4250) );
  MUX2X1 U4867 ( .B(mem[246]), .A(mem[287]), .S(n5505), .Y(n4244) );
  MUX2X1 U4868 ( .B(mem[164]), .A(mem[205]), .S(n5505), .Y(n4243) );
  MUX2X1 U4869 ( .B(mem[82]), .A(mem[123]), .S(n5505), .Y(n4247) );
  MUX2X1 U4870 ( .B(mem[0]), .A(mem[41]), .S(n5505), .Y(n4246) );
  MUX2X1 U4871 ( .B(n4245), .A(n4242), .S(n14), .Y(n4249) );
  MUX2X1 U4872 ( .B(n4248), .A(n4233), .S(n16), .Y(n5451) );
  MUX2X1 U4873 ( .B(mem[1231]), .A(mem[1272]), .S(n5505), .Y(n4253) );
  MUX2X1 U4874 ( .B(mem[1149]), .A(mem[1190]), .S(n5505), .Y(n4252) );
  MUX2X1 U4875 ( .B(mem[1067]), .A(mem[1108]), .S(n5505), .Y(n4256) );
  MUX2X1 U4876 ( .B(mem[985]), .A(mem[1026]), .S(n5505), .Y(n4255) );
  MUX2X1 U4877 ( .B(n4254), .A(n4251), .S(n14), .Y(n4265) );
  MUX2X1 U4878 ( .B(mem[903]), .A(mem[944]), .S(n5506), .Y(n4259) );
  MUX2X1 U4879 ( .B(mem[821]), .A(mem[862]), .S(n5506), .Y(n4258) );
  MUX2X1 U4880 ( .B(mem[739]), .A(mem[780]), .S(n5506), .Y(n4262) );
  MUX2X1 U4881 ( .B(mem[657]), .A(mem[698]), .S(n5506), .Y(n4261) );
  MUX2X1 U4882 ( .B(n4260), .A(n4257), .S(n14), .Y(n4264) );
  MUX2X1 U4883 ( .B(mem[575]), .A(mem[616]), .S(n5506), .Y(n4268) );
  MUX2X1 U4884 ( .B(mem[493]), .A(mem[534]), .S(n5506), .Y(n4267) );
  MUX2X1 U4885 ( .B(mem[411]), .A(mem[452]), .S(n5506), .Y(n4271) );
  MUX2X1 U4886 ( .B(mem[329]), .A(mem[370]), .S(n5506), .Y(n4270) );
  MUX2X1 U4887 ( .B(n4269), .A(n4266), .S(n14), .Y(n4280) );
  MUX2X1 U4888 ( .B(mem[247]), .A(mem[288]), .S(n5506), .Y(n4274) );
  MUX2X1 U4889 ( .B(mem[165]), .A(mem[206]), .S(n5506), .Y(n4273) );
  MUX2X1 U4890 ( .B(mem[83]), .A(mem[124]), .S(n5506), .Y(n4277) );
  MUX2X1 U4891 ( .B(mem[1]), .A(mem[42]), .S(n5506), .Y(n4276) );
  MUX2X1 U4892 ( .B(n4275), .A(n4272), .S(n14), .Y(n4279) );
  MUX2X1 U4893 ( .B(n4278), .A(n4263), .S(n16), .Y(n5452) );
  MUX2X1 U4894 ( .B(mem[1232]), .A(mem[1273]), .S(n5507), .Y(n4283) );
  MUX2X1 U4895 ( .B(mem[1150]), .A(mem[1191]), .S(n5507), .Y(n4282) );
  MUX2X1 U4896 ( .B(mem[1068]), .A(mem[1109]), .S(n5507), .Y(n4286) );
  MUX2X1 U4897 ( .B(mem[986]), .A(mem[1027]), .S(n5507), .Y(n4285) );
  MUX2X1 U4898 ( .B(n4284), .A(n4281), .S(n5589), .Y(n4295) );
  MUX2X1 U4899 ( .B(mem[904]), .A(mem[945]), .S(n5507), .Y(n4289) );
  MUX2X1 U4900 ( .B(mem[822]), .A(mem[863]), .S(n5507), .Y(n4288) );
  MUX2X1 U4901 ( .B(mem[740]), .A(mem[781]), .S(n5507), .Y(n4292) );
  MUX2X1 U4902 ( .B(mem[658]), .A(mem[699]), .S(n5507), .Y(n4291) );
  MUX2X1 U4903 ( .B(n4290), .A(n4287), .S(n5589), .Y(n4294) );
  MUX2X1 U4904 ( .B(mem[576]), .A(mem[617]), .S(n5507), .Y(n4298) );
  MUX2X1 U4905 ( .B(mem[494]), .A(mem[535]), .S(n5507), .Y(n4297) );
  MUX2X1 U4906 ( .B(mem[412]), .A(mem[453]), .S(n5507), .Y(n4301) );
  MUX2X1 U4907 ( .B(mem[330]), .A(mem[371]), .S(n5507), .Y(n4300) );
  MUX2X1 U4908 ( .B(n4299), .A(n4296), .S(n5589), .Y(n4310) );
  MUX2X1 U4909 ( .B(mem[248]), .A(mem[289]), .S(n5508), .Y(n4304) );
  MUX2X1 U4910 ( .B(mem[166]), .A(mem[207]), .S(n5508), .Y(n4303) );
  MUX2X1 U4911 ( .B(mem[84]), .A(mem[125]), .S(n5508), .Y(n4307) );
  MUX2X1 U4912 ( .B(mem[2]), .A(mem[43]), .S(n5508), .Y(n4306) );
  MUX2X1 U4913 ( .B(n4305), .A(n4302), .S(n5589), .Y(n4309) );
  MUX2X1 U4914 ( .B(n4308), .A(n4293), .S(n16), .Y(n5453) );
  MUX2X1 U4915 ( .B(mem[1233]), .A(mem[1274]), .S(n5508), .Y(n4313) );
  MUX2X1 U4916 ( .B(mem[1151]), .A(mem[1192]), .S(n5508), .Y(n4312) );
  MUX2X1 U4917 ( .B(mem[1069]), .A(mem[1110]), .S(n5508), .Y(n4316) );
  MUX2X1 U4918 ( .B(mem[987]), .A(mem[1028]), .S(n5508), .Y(n4315) );
  MUX2X1 U4919 ( .B(n4314), .A(n4311), .S(n5589), .Y(n4325) );
  MUX2X1 U4920 ( .B(mem[905]), .A(mem[946]), .S(n5508), .Y(n4319) );
  MUX2X1 U4921 ( .B(mem[823]), .A(mem[864]), .S(n5508), .Y(n4318) );
  MUX2X1 U4922 ( .B(mem[741]), .A(mem[782]), .S(n5508), .Y(n4322) );
  MUX2X1 U4923 ( .B(mem[659]), .A(mem[700]), .S(n5508), .Y(n4321) );
  MUX2X1 U4924 ( .B(n4320), .A(n4317), .S(n5589), .Y(n4324) );
  MUX2X1 U4925 ( .B(mem[577]), .A(mem[618]), .S(n5509), .Y(n4328) );
  MUX2X1 U4926 ( .B(mem[495]), .A(mem[536]), .S(n5509), .Y(n4327) );
  MUX2X1 U4927 ( .B(mem[413]), .A(mem[454]), .S(n5509), .Y(n4331) );
  MUX2X1 U4928 ( .B(mem[331]), .A(mem[372]), .S(n5509), .Y(n4330) );
  MUX2X1 U4929 ( .B(n4329), .A(n4326), .S(n5589), .Y(n4340) );
  MUX2X1 U4930 ( .B(mem[249]), .A(mem[290]), .S(n5509), .Y(n4334) );
  MUX2X1 U4931 ( .B(mem[167]), .A(mem[208]), .S(n5509), .Y(n4333) );
  MUX2X1 U4932 ( .B(mem[85]), .A(mem[126]), .S(n5509), .Y(n4337) );
  MUX2X1 U4933 ( .B(mem[3]), .A(mem[44]), .S(n5509), .Y(n4336) );
  MUX2X1 U4934 ( .B(n4335), .A(n4332), .S(n5589), .Y(n4339) );
  MUX2X1 U4935 ( .B(n4338), .A(n4323), .S(n16), .Y(n5454) );
  MUX2X1 U4936 ( .B(mem[1234]), .A(mem[1275]), .S(n5509), .Y(n4343) );
  MUX2X1 U4937 ( .B(mem[1152]), .A(mem[1193]), .S(n5509), .Y(n4342) );
  MUX2X1 U4938 ( .B(mem[1070]), .A(mem[1111]), .S(n5509), .Y(n4346) );
  MUX2X1 U4939 ( .B(mem[988]), .A(mem[1029]), .S(n5509), .Y(n4345) );
  MUX2X1 U4940 ( .B(n4344), .A(n4341), .S(n5589), .Y(n4355) );
  MUX2X1 U4941 ( .B(mem[906]), .A(mem[947]), .S(n5510), .Y(n4349) );
  MUX2X1 U4942 ( .B(mem[824]), .A(mem[865]), .S(n5510), .Y(n4348) );
  MUX2X1 U4943 ( .B(mem[742]), .A(mem[783]), .S(n5510), .Y(n4352) );
  MUX2X1 U4944 ( .B(mem[660]), .A(mem[701]), .S(n5510), .Y(n4351) );
  MUX2X1 U4945 ( .B(n4350), .A(n4347), .S(n5589), .Y(n4354) );
  MUX2X1 U4946 ( .B(mem[578]), .A(mem[619]), .S(n5510), .Y(n4358) );
  MUX2X1 U4947 ( .B(mem[496]), .A(mem[537]), .S(n5510), .Y(n4357) );
  MUX2X1 U4948 ( .B(mem[414]), .A(mem[455]), .S(n5510), .Y(n4361) );
  MUX2X1 U4949 ( .B(mem[332]), .A(mem[373]), .S(n5510), .Y(n4360) );
  MUX2X1 U4950 ( .B(n4359), .A(n4356), .S(n5589), .Y(n4370) );
  MUX2X1 U4951 ( .B(mem[250]), .A(mem[291]), .S(n5510), .Y(n4364) );
  MUX2X1 U4952 ( .B(mem[168]), .A(mem[209]), .S(n5510), .Y(n4363) );
  MUX2X1 U4953 ( .B(mem[86]), .A(mem[127]), .S(n5510), .Y(n4367) );
  MUX2X1 U4954 ( .B(mem[4]), .A(mem[45]), .S(n5510), .Y(n4366) );
  MUX2X1 U4955 ( .B(n4365), .A(n4362), .S(n5589), .Y(n4369) );
  MUX2X1 U4956 ( .B(n4368), .A(n4353), .S(n16), .Y(n5455) );
  MUX2X1 U4957 ( .B(mem[1235]), .A(mem[1276]), .S(n5511), .Y(n4373) );
  MUX2X1 U4958 ( .B(mem[1153]), .A(mem[1194]), .S(n5511), .Y(n4372) );
  MUX2X1 U4959 ( .B(mem[1071]), .A(mem[1112]), .S(n5511), .Y(n4376) );
  MUX2X1 U4960 ( .B(mem[989]), .A(mem[1030]), .S(n5511), .Y(n4375) );
  MUX2X1 U4961 ( .B(n4374), .A(n4371), .S(n5590), .Y(n4385) );
  MUX2X1 U4962 ( .B(mem[907]), .A(mem[948]), .S(n5511), .Y(n4379) );
  MUX2X1 U4963 ( .B(mem[825]), .A(mem[866]), .S(n5511), .Y(n4378) );
  MUX2X1 U4964 ( .B(mem[743]), .A(mem[784]), .S(n5511), .Y(n4382) );
  MUX2X1 U4965 ( .B(mem[661]), .A(mem[702]), .S(n5511), .Y(n4381) );
  MUX2X1 U4966 ( .B(n4380), .A(n4377), .S(n5590), .Y(n4384) );
  MUX2X1 U4967 ( .B(mem[579]), .A(mem[620]), .S(n5511), .Y(n4388) );
  MUX2X1 U4968 ( .B(mem[497]), .A(mem[538]), .S(n5511), .Y(n4387) );
  MUX2X1 U4969 ( .B(mem[415]), .A(mem[456]), .S(n5511), .Y(n4391) );
  MUX2X1 U4970 ( .B(mem[333]), .A(mem[374]), .S(n5511), .Y(n4390) );
  MUX2X1 U4971 ( .B(n4389), .A(n4386), .S(n5590), .Y(n4400) );
  MUX2X1 U4972 ( .B(mem[251]), .A(mem[292]), .S(n5512), .Y(n4394) );
  MUX2X1 U4973 ( .B(mem[169]), .A(mem[210]), .S(n5512), .Y(n4393) );
  MUX2X1 U4974 ( .B(mem[87]), .A(mem[128]), .S(n5512), .Y(n4397) );
  MUX2X1 U4975 ( .B(mem[5]), .A(mem[46]), .S(n5512), .Y(n4396) );
  MUX2X1 U4976 ( .B(n4395), .A(n4392), .S(n5590), .Y(n4399) );
  MUX2X1 U4977 ( .B(n4398), .A(n4383), .S(n16), .Y(n5456) );
  MUX2X1 U4978 ( .B(mem[1236]), .A(mem[1277]), .S(n5512), .Y(n4403) );
  MUX2X1 U4979 ( .B(mem[1154]), .A(mem[1195]), .S(n5512), .Y(n4402) );
  MUX2X1 U4980 ( .B(mem[1072]), .A(mem[1113]), .S(n5512), .Y(n4406) );
  MUX2X1 U4981 ( .B(mem[990]), .A(mem[1031]), .S(n5512), .Y(n4405) );
  MUX2X1 U4982 ( .B(n4404), .A(n4401), .S(n5590), .Y(n4415) );
  MUX2X1 U4983 ( .B(mem[908]), .A(mem[949]), .S(n5512), .Y(n4409) );
  MUX2X1 U4984 ( .B(mem[826]), .A(mem[867]), .S(n5512), .Y(n4408) );
  MUX2X1 U4985 ( .B(mem[744]), .A(mem[785]), .S(n5512), .Y(n4412) );
  MUX2X1 U4986 ( .B(mem[662]), .A(mem[703]), .S(n5512), .Y(n4411) );
  MUX2X1 U4987 ( .B(n4410), .A(n4407), .S(n5590), .Y(n4414) );
  MUX2X1 U4988 ( .B(mem[580]), .A(mem[621]), .S(n5513), .Y(n4418) );
  MUX2X1 U4989 ( .B(mem[498]), .A(mem[539]), .S(n5513), .Y(n4417) );
  MUX2X1 U4990 ( .B(mem[416]), .A(mem[457]), .S(n5513), .Y(n4421) );
  MUX2X1 U4991 ( .B(mem[334]), .A(mem[375]), .S(n5513), .Y(n4420) );
  MUX2X1 U4992 ( .B(n4419), .A(n4416), .S(n5590), .Y(n4430) );
  MUX2X1 U4993 ( .B(mem[252]), .A(mem[293]), .S(n5513), .Y(n4424) );
  MUX2X1 U4994 ( .B(mem[170]), .A(mem[211]), .S(n5513), .Y(n4423) );
  MUX2X1 U4995 ( .B(mem[88]), .A(mem[129]), .S(n5513), .Y(n4427) );
  MUX2X1 U4996 ( .B(mem[6]), .A(mem[47]), .S(n5513), .Y(n4426) );
  MUX2X1 U4997 ( .B(n4425), .A(n4422), .S(n5590), .Y(n4429) );
  MUX2X1 U4998 ( .B(n4428), .A(n4413), .S(n16), .Y(n5457) );
  MUX2X1 U4999 ( .B(mem[1237]), .A(mem[1278]), .S(n5513), .Y(n4433) );
  MUX2X1 U5000 ( .B(mem[1155]), .A(mem[1196]), .S(n5513), .Y(n4432) );
  MUX2X1 U5001 ( .B(mem[1073]), .A(mem[1114]), .S(n5513), .Y(n4436) );
  MUX2X1 U5002 ( .B(mem[991]), .A(mem[1032]), .S(n5513), .Y(n4435) );
  MUX2X1 U5003 ( .B(n4434), .A(n4431), .S(n5590), .Y(n4445) );
  MUX2X1 U5004 ( .B(mem[909]), .A(mem[950]), .S(n5514), .Y(n4439) );
  MUX2X1 U5005 ( .B(mem[827]), .A(mem[868]), .S(n5514), .Y(n4438) );
  MUX2X1 U5006 ( .B(mem[745]), .A(mem[786]), .S(n5514), .Y(n4442) );
  MUX2X1 U5007 ( .B(mem[663]), .A(mem[704]), .S(n5514), .Y(n4441) );
  MUX2X1 U5008 ( .B(n4440), .A(n4437), .S(n5590), .Y(n4444) );
  MUX2X1 U5009 ( .B(mem[581]), .A(mem[622]), .S(n5514), .Y(n4448) );
  MUX2X1 U5010 ( .B(mem[499]), .A(mem[540]), .S(n5514), .Y(n4447) );
  MUX2X1 U5011 ( .B(mem[417]), .A(mem[458]), .S(n5514), .Y(n4451) );
  MUX2X1 U5012 ( .B(mem[335]), .A(mem[376]), .S(n5514), .Y(n4450) );
  MUX2X1 U5013 ( .B(n4449), .A(n4446), .S(n5590), .Y(n4460) );
  MUX2X1 U5014 ( .B(mem[253]), .A(mem[294]), .S(n5514), .Y(n4454) );
  MUX2X1 U5015 ( .B(mem[171]), .A(mem[212]), .S(n5514), .Y(n4453) );
  MUX2X1 U5016 ( .B(mem[89]), .A(mem[130]), .S(n5514), .Y(n4457) );
  MUX2X1 U5017 ( .B(mem[7]), .A(mem[48]), .S(n5514), .Y(n4456) );
  MUX2X1 U5018 ( .B(n4455), .A(n4452), .S(n5590), .Y(n4459) );
  MUX2X1 U5019 ( .B(n4458), .A(n4443), .S(n16), .Y(n5458) );
  MUX2X1 U5020 ( .B(mem[1238]), .A(mem[1279]), .S(n5515), .Y(n4463) );
  MUX2X1 U5021 ( .B(mem[1156]), .A(mem[1197]), .S(n5515), .Y(n4462) );
  MUX2X1 U5022 ( .B(mem[1074]), .A(mem[1115]), .S(n5515), .Y(n4466) );
  MUX2X1 U5023 ( .B(mem[992]), .A(mem[1033]), .S(n5515), .Y(n4465) );
  MUX2X1 U5024 ( .B(n4464), .A(n4461), .S(n5591), .Y(n4475) );
  MUX2X1 U5025 ( .B(mem[910]), .A(mem[951]), .S(n5515), .Y(n4469) );
  MUX2X1 U5026 ( .B(mem[828]), .A(mem[869]), .S(n5515), .Y(n4468) );
  MUX2X1 U5027 ( .B(mem[746]), .A(mem[787]), .S(n5515), .Y(n4472) );
  MUX2X1 U5028 ( .B(mem[664]), .A(mem[705]), .S(n5515), .Y(n4471) );
  MUX2X1 U5029 ( .B(n4470), .A(n4467), .S(n5591), .Y(n4474) );
  MUX2X1 U5030 ( .B(mem[582]), .A(mem[623]), .S(n5515), .Y(n4478) );
  MUX2X1 U5031 ( .B(mem[500]), .A(mem[541]), .S(n5515), .Y(n4477) );
  MUX2X1 U5032 ( .B(mem[418]), .A(mem[459]), .S(n5515), .Y(n4481) );
  MUX2X1 U5033 ( .B(mem[336]), .A(mem[377]), .S(n5515), .Y(n4480) );
  MUX2X1 U5034 ( .B(n4479), .A(n4476), .S(n5591), .Y(n4490) );
  MUX2X1 U5035 ( .B(mem[254]), .A(mem[295]), .S(n5516), .Y(n4484) );
  MUX2X1 U5036 ( .B(mem[172]), .A(mem[213]), .S(n5516), .Y(n4483) );
  MUX2X1 U5037 ( .B(mem[90]), .A(mem[131]), .S(n5516), .Y(n4487) );
  MUX2X1 U5038 ( .B(mem[8]), .A(mem[49]), .S(n5516), .Y(n4486) );
  MUX2X1 U5039 ( .B(n4485), .A(n4482), .S(n5591), .Y(n4489) );
  MUX2X1 U5040 ( .B(n4488), .A(n4473), .S(n16), .Y(n5459) );
  MUX2X1 U5041 ( .B(mem[1239]), .A(mem[1280]), .S(n5516), .Y(n4493) );
  MUX2X1 U5042 ( .B(mem[1157]), .A(mem[1198]), .S(n5516), .Y(n4492) );
  MUX2X1 U5043 ( .B(mem[1075]), .A(mem[1116]), .S(n5516), .Y(n4496) );
  MUX2X1 U5044 ( .B(mem[993]), .A(mem[1034]), .S(n5516), .Y(n4495) );
  MUX2X1 U5045 ( .B(n4494), .A(n4491), .S(n5591), .Y(n4505) );
  MUX2X1 U5046 ( .B(mem[911]), .A(mem[952]), .S(n5516), .Y(n4499) );
  MUX2X1 U5047 ( .B(mem[829]), .A(mem[870]), .S(n5516), .Y(n4498) );
  MUX2X1 U5048 ( .B(mem[747]), .A(mem[788]), .S(n5516), .Y(n4502) );
  MUX2X1 U5049 ( .B(mem[665]), .A(mem[706]), .S(n5516), .Y(n4501) );
  MUX2X1 U5050 ( .B(n4500), .A(n4497), .S(n5591), .Y(n4504) );
  MUX2X1 U5051 ( .B(mem[583]), .A(mem[624]), .S(n5517), .Y(n4508) );
  MUX2X1 U5052 ( .B(mem[501]), .A(mem[542]), .S(n5517), .Y(n4507) );
  MUX2X1 U5053 ( .B(mem[419]), .A(mem[460]), .S(n5517), .Y(n4511) );
  MUX2X1 U5054 ( .B(mem[337]), .A(mem[378]), .S(n5517), .Y(n4510) );
  MUX2X1 U5055 ( .B(n4509), .A(n4506), .S(n5591), .Y(n4520) );
  MUX2X1 U5056 ( .B(mem[255]), .A(mem[296]), .S(n5517), .Y(n4514) );
  MUX2X1 U5057 ( .B(mem[173]), .A(mem[214]), .S(n5517), .Y(n4513) );
  MUX2X1 U5058 ( .B(mem[91]), .A(mem[132]), .S(n5517), .Y(n4517) );
  MUX2X1 U5059 ( .B(mem[9]), .A(mem[50]), .S(n5517), .Y(n4516) );
  MUX2X1 U5060 ( .B(n4515), .A(n4512), .S(n5591), .Y(n4519) );
  MUX2X1 U5061 ( .B(n4518), .A(n4503), .S(n16), .Y(n5460) );
  MUX2X1 U5062 ( .B(mem[1240]), .A(mem[1281]), .S(n5517), .Y(n4523) );
  MUX2X1 U5063 ( .B(mem[1158]), .A(mem[1199]), .S(n5517), .Y(n4522) );
  MUX2X1 U5064 ( .B(mem[1076]), .A(mem[1117]), .S(n5517), .Y(n4526) );
  MUX2X1 U5065 ( .B(mem[994]), .A(mem[1035]), .S(n5517), .Y(n4525) );
  MUX2X1 U5066 ( .B(n4524), .A(n4521), .S(n5591), .Y(n4535) );
  MUX2X1 U5067 ( .B(mem[912]), .A(mem[953]), .S(n5518), .Y(n4529) );
  MUX2X1 U5068 ( .B(mem[830]), .A(mem[871]), .S(n5518), .Y(n4528) );
  MUX2X1 U5069 ( .B(mem[748]), .A(mem[789]), .S(n5518), .Y(n4532) );
  MUX2X1 U5070 ( .B(mem[666]), .A(mem[707]), .S(n5518), .Y(n4531) );
  MUX2X1 U5071 ( .B(n4530), .A(n4527), .S(n5591), .Y(n4534) );
  MUX2X1 U5072 ( .B(mem[584]), .A(mem[625]), .S(n5518), .Y(n4538) );
  MUX2X1 U5073 ( .B(mem[502]), .A(mem[543]), .S(n5518), .Y(n4537) );
  MUX2X1 U5074 ( .B(mem[420]), .A(mem[461]), .S(n5518), .Y(n4541) );
  MUX2X1 U5075 ( .B(mem[338]), .A(mem[379]), .S(n5518), .Y(n4540) );
  MUX2X1 U5076 ( .B(n4539), .A(n4536), .S(n5591), .Y(n4550) );
  MUX2X1 U5077 ( .B(mem[256]), .A(mem[297]), .S(n5518), .Y(n4544) );
  MUX2X1 U5078 ( .B(mem[174]), .A(mem[215]), .S(n5518), .Y(n4543) );
  MUX2X1 U5079 ( .B(mem[92]), .A(mem[133]), .S(n5518), .Y(n4547) );
  MUX2X1 U5080 ( .B(mem[10]), .A(mem[51]), .S(n5518), .Y(n4546) );
  MUX2X1 U5081 ( .B(n4545), .A(n4542), .S(n5591), .Y(n4549) );
  MUX2X1 U5082 ( .B(n4548), .A(n4533), .S(n16), .Y(n5461) );
  MUX2X1 U5083 ( .B(mem[1241]), .A(mem[1282]), .S(n5519), .Y(n4553) );
  MUX2X1 U5084 ( .B(mem[1159]), .A(mem[1200]), .S(n5519), .Y(n4552) );
  MUX2X1 U5085 ( .B(mem[1077]), .A(mem[1118]), .S(n5519), .Y(n4556) );
  MUX2X1 U5086 ( .B(mem[995]), .A(mem[1036]), .S(n5519), .Y(n4555) );
  MUX2X1 U5087 ( .B(n4554), .A(n4551), .S(n5592), .Y(n4565) );
  MUX2X1 U5088 ( .B(mem[913]), .A(mem[954]), .S(n5519), .Y(n4559) );
  MUX2X1 U5089 ( .B(mem[831]), .A(mem[872]), .S(n5519), .Y(n4558) );
  MUX2X1 U5090 ( .B(mem[749]), .A(mem[790]), .S(n5519), .Y(n4562) );
  MUX2X1 U5091 ( .B(mem[667]), .A(mem[708]), .S(n5519), .Y(n4561) );
  MUX2X1 U5092 ( .B(n4560), .A(n4557), .S(n5592), .Y(n4564) );
  MUX2X1 U5093 ( .B(mem[585]), .A(mem[626]), .S(n5519), .Y(n4568) );
  MUX2X1 U5094 ( .B(mem[503]), .A(mem[544]), .S(n5519), .Y(n4567) );
  MUX2X1 U5095 ( .B(mem[421]), .A(mem[462]), .S(n5519), .Y(n4571) );
  MUX2X1 U5096 ( .B(mem[339]), .A(mem[380]), .S(n5519), .Y(n4570) );
  MUX2X1 U5097 ( .B(n4569), .A(n4566), .S(n5592), .Y(n4580) );
  MUX2X1 U5098 ( .B(mem[257]), .A(mem[298]), .S(n5520), .Y(n4574) );
  MUX2X1 U5099 ( .B(mem[175]), .A(mem[216]), .S(n5520), .Y(n4573) );
  MUX2X1 U5100 ( .B(mem[93]), .A(mem[134]), .S(n5520), .Y(n4577) );
  MUX2X1 U5101 ( .B(mem[11]), .A(mem[52]), .S(n5520), .Y(n4576) );
  MUX2X1 U5102 ( .B(n4575), .A(n4572), .S(n5592), .Y(n4579) );
  MUX2X1 U5103 ( .B(n4578), .A(n4563), .S(n16), .Y(n5462) );
  MUX2X1 U5104 ( .B(mem[1242]), .A(mem[1283]), .S(n5520), .Y(n4583) );
  MUX2X1 U5105 ( .B(mem[1160]), .A(mem[1201]), .S(n5520), .Y(n4582) );
  MUX2X1 U5106 ( .B(mem[1078]), .A(mem[1119]), .S(n5520), .Y(n4586) );
  MUX2X1 U5107 ( .B(mem[996]), .A(mem[1037]), .S(n5520), .Y(n4585) );
  MUX2X1 U5108 ( .B(n4584), .A(n4581), .S(n5592), .Y(n4595) );
  MUX2X1 U5109 ( .B(mem[914]), .A(mem[955]), .S(n5520), .Y(n4589) );
  MUX2X1 U5110 ( .B(mem[832]), .A(mem[873]), .S(n5520), .Y(n4588) );
  MUX2X1 U5111 ( .B(mem[750]), .A(mem[791]), .S(n5520), .Y(n4592) );
  MUX2X1 U5112 ( .B(mem[668]), .A(mem[709]), .S(n5520), .Y(n4591) );
  MUX2X1 U5113 ( .B(n4590), .A(n4587), .S(n5592), .Y(n4594) );
  MUX2X1 U5114 ( .B(mem[586]), .A(mem[627]), .S(n5521), .Y(n4598) );
  MUX2X1 U5115 ( .B(mem[504]), .A(mem[545]), .S(n5521), .Y(n4597) );
  MUX2X1 U5116 ( .B(mem[422]), .A(mem[463]), .S(n5521), .Y(n4601) );
  MUX2X1 U5117 ( .B(mem[340]), .A(mem[381]), .S(n5521), .Y(n4600) );
  MUX2X1 U5118 ( .B(n4599), .A(n4596), .S(n5592), .Y(n4610) );
  MUX2X1 U5119 ( .B(mem[258]), .A(mem[299]), .S(n5521), .Y(n4604) );
  MUX2X1 U5120 ( .B(mem[176]), .A(mem[217]), .S(n5521), .Y(n4603) );
  MUX2X1 U5121 ( .B(mem[94]), .A(mem[135]), .S(n5521), .Y(n4607) );
  MUX2X1 U5122 ( .B(mem[12]), .A(mem[53]), .S(n5521), .Y(n4606) );
  MUX2X1 U5123 ( .B(n4605), .A(n4602), .S(n5592), .Y(n4609) );
  MUX2X1 U5124 ( .B(n4608), .A(n4593), .S(n16), .Y(n5463) );
  MUX2X1 U5125 ( .B(mem[1243]), .A(mem[1284]), .S(n5521), .Y(n4613) );
  MUX2X1 U5126 ( .B(mem[1161]), .A(mem[1202]), .S(n5521), .Y(n4612) );
  MUX2X1 U5127 ( .B(mem[1079]), .A(mem[1120]), .S(n5521), .Y(n4616) );
  MUX2X1 U5128 ( .B(mem[997]), .A(mem[1038]), .S(n5521), .Y(n4615) );
  MUX2X1 U5129 ( .B(n4614), .A(n4611), .S(n5592), .Y(n4625) );
  MUX2X1 U5130 ( .B(mem[915]), .A(mem[956]), .S(n5522), .Y(n4619) );
  MUX2X1 U5131 ( .B(mem[833]), .A(mem[874]), .S(n5522), .Y(n4618) );
  MUX2X1 U5132 ( .B(mem[751]), .A(mem[792]), .S(n5522), .Y(n4622) );
  MUX2X1 U5133 ( .B(mem[669]), .A(mem[710]), .S(n5522), .Y(n4621) );
  MUX2X1 U5134 ( .B(n4620), .A(n4617), .S(n5592), .Y(n4624) );
  MUX2X1 U5135 ( .B(mem[587]), .A(mem[628]), .S(n5522), .Y(n4628) );
  MUX2X1 U5136 ( .B(mem[505]), .A(mem[546]), .S(n5522), .Y(n4627) );
  MUX2X1 U5137 ( .B(mem[423]), .A(mem[464]), .S(n5522), .Y(n4631) );
  MUX2X1 U5138 ( .B(mem[341]), .A(mem[382]), .S(n5522), .Y(n4630) );
  MUX2X1 U5139 ( .B(n4629), .A(n4626), .S(n5592), .Y(n4640) );
  MUX2X1 U5140 ( .B(mem[259]), .A(mem[300]), .S(n5522), .Y(n4634) );
  MUX2X1 U5141 ( .B(mem[177]), .A(mem[218]), .S(n5522), .Y(n4633) );
  MUX2X1 U5142 ( .B(mem[95]), .A(mem[136]), .S(n5522), .Y(n4637) );
  MUX2X1 U5143 ( .B(mem[13]), .A(mem[54]), .S(n5522), .Y(n4636) );
  MUX2X1 U5144 ( .B(n4635), .A(n4632), .S(n5592), .Y(n4639) );
  MUX2X1 U5145 ( .B(n4638), .A(n4623), .S(n16), .Y(n5464) );
  MUX2X1 U5146 ( .B(mem[1244]), .A(mem[1285]), .S(n5523), .Y(n4643) );
  MUX2X1 U5147 ( .B(mem[1162]), .A(mem[1203]), .S(n5523), .Y(n4642) );
  MUX2X1 U5148 ( .B(mem[1080]), .A(mem[1121]), .S(n5523), .Y(n4646) );
  MUX2X1 U5149 ( .B(mem[998]), .A(mem[1039]), .S(n5523), .Y(n4645) );
  MUX2X1 U5150 ( .B(n4644), .A(n4641), .S(n5593), .Y(n4655) );
  MUX2X1 U5151 ( .B(mem[916]), .A(mem[957]), .S(n5523), .Y(n4649) );
  MUX2X1 U5152 ( .B(mem[834]), .A(mem[875]), .S(n5523), .Y(n4648) );
  MUX2X1 U5153 ( .B(mem[752]), .A(mem[793]), .S(n5523), .Y(n4652) );
  MUX2X1 U5154 ( .B(mem[670]), .A(mem[711]), .S(n5523), .Y(n4651) );
  MUX2X1 U5155 ( .B(n4650), .A(n4647), .S(n5593), .Y(n4654) );
  MUX2X1 U5156 ( .B(mem[588]), .A(mem[629]), .S(n5523), .Y(n4658) );
  MUX2X1 U5157 ( .B(mem[506]), .A(mem[547]), .S(n5523), .Y(n4657) );
  MUX2X1 U5158 ( .B(mem[424]), .A(mem[465]), .S(n5523), .Y(n4661) );
  MUX2X1 U5159 ( .B(mem[342]), .A(mem[383]), .S(n5523), .Y(n4660) );
  MUX2X1 U5160 ( .B(n4659), .A(n4656), .S(n5593), .Y(n4670) );
  MUX2X1 U5161 ( .B(mem[260]), .A(mem[301]), .S(n5524), .Y(n4664) );
  MUX2X1 U5162 ( .B(mem[178]), .A(mem[219]), .S(n5524), .Y(n4663) );
  MUX2X1 U5163 ( .B(mem[96]), .A(mem[137]), .S(n5524), .Y(n4667) );
  MUX2X1 U5164 ( .B(mem[14]), .A(mem[55]), .S(n5524), .Y(n4666) );
  MUX2X1 U5165 ( .B(n4665), .A(n4662), .S(n5593), .Y(n4669) );
  MUX2X1 U5166 ( .B(n4668), .A(n4653), .S(n16), .Y(n5465) );
  MUX2X1 U5167 ( .B(mem[1245]), .A(mem[1286]), .S(n5524), .Y(n4673) );
  MUX2X1 U5168 ( .B(mem[1163]), .A(mem[1204]), .S(n5524), .Y(n4672) );
  MUX2X1 U5169 ( .B(mem[1081]), .A(mem[1122]), .S(n5524), .Y(n4676) );
  MUX2X1 U5170 ( .B(mem[999]), .A(mem[1040]), .S(n5524), .Y(n4675) );
  MUX2X1 U5171 ( .B(n4674), .A(n4671), .S(n5593), .Y(n4685) );
  MUX2X1 U5172 ( .B(mem[917]), .A(mem[958]), .S(n5524), .Y(n4679) );
  MUX2X1 U5173 ( .B(mem[835]), .A(mem[876]), .S(n5524), .Y(n4678) );
  MUX2X1 U5174 ( .B(mem[753]), .A(mem[794]), .S(n5524), .Y(n4682) );
  MUX2X1 U5175 ( .B(mem[671]), .A(mem[712]), .S(n5524), .Y(n4681) );
  MUX2X1 U5176 ( .B(n4680), .A(n4677), .S(n5593), .Y(n4684) );
  MUX2X1 U5177 ( .B(mem[589]), .A(mem[630]), .S(n5525), .Y(n4688) );
  MUX2X1 U5178 ( .B(mem[507]), .A(mem[548]), .S(n5525), .Y(n4687) );
  MUX2X1 U5179 ( .B(mem[425]), .A(mem[466]), .S(n5525), .Y(n4691) );
  MUX2X1 U5180 ( .B(mem[343]), .A(mem[384]), .S(n5525), .Y(n4690) );
  MUX2X1 U5181 ( .B(n4689), .A(n4686), .S(n5593), .Y(n4700) );
  MUX2X1 U5182 ( .B(mem[261]), .A(mem[302]), .S(n5525), .Y(n4694) );
  MUX2X1 U5183 ( .B(mem[179]), .A(mem[220]), .S(n5525), .Y(n4693) );
  MUX2X1 U5184 ( .B(mem[97]), .A(mem[138]), .S(n5525), .Y(n4697) );
  MUX2X1 U5185 ( .B(mem[15]), .A(mem[56]), .S(n5525), .Y(n4696) );
  MUX2X1 U5186 ( .B(n4695), .A(n4692), .S(n5593), .Y(n4699) );
  MUX2X1 U5187 ( .B(n4698), .A(n4683), .S(n16), .Y(n5466) );
  MUX2X1 U5188 ( .B(mem[1246]), .A(mem[1287]), .S(n5525), .Y(n4703) );
  MUX2X1 U5189 ( .B(mem[1164]), .A(mem[1205]), .S(n5525), .Y(n4702) );
  MUX2X1 U5190 ( .B(mem[1082]), .A(mem[1123]), .S(n5525), .Y(n4706) );
  MUX2X1 U5191 ( .B(mem[1000]), .A(mem[1041]), .S(n5525), .Y(n4705) );
  MUX2X1 U5192 ( .B(n4704), .A(n4701), .S(n5593), .Y(n4715) );
  MUX2X1 U5193 ( .B(mem[918]), .A(mem[959]), .S(n5526), .Y(n4709) );
  MUX2X1 U5194 ( .B(mem[836]), .A(mem[877]), .S(n5526), .Y(n4708) );
  MUX2X1 U5195 ( .B(mem[754]), .A(mem[795]), .S(n5526), .Y(n4712) );
  MUX2X1 U5196 ( .B(mem[672]), .A(mem[713]), .S(n5526), .Y(n4711) );
  MUX2X1 U5197 ( .B(n4710), .A(n4707), .S(n5593), .Y(n4714) );
  MUX2X1 U5198 ( .B(mem[590]), .A(mem[631]), .S(n5526), .Y(n4718) );
  MUX2X1 U5199 ( .B(mem[508]), .A(mem[549]), .S(n5526), .Y(n4717) );
  MUX2X1 U5200 ( .B(mem[426]), .A(mem[467]), .S(n5526), .Y(n4721) );
  MUX2X1 U5201 ( .B(mem[344]), .A(mem[385]), .S(n5526), .Y(n4720) );
  MUX2X1 U5202 ( .B(n4719), .A(n4716), .S(n5593), .Y(n4730) );
  MUX2X1 U5203 ( .B(mem[262]), .A(mem[303]), .S(n5526), .Y(n4724) );
  MUX2X1 U5204 ( .B(mem[180]), .A(mem[221]), .S(n5526), .Y(n4723) );
  MUX2X1 U5205 ( .B(mem[98]), .A(mem[139]), .S(n5526), .Y(n4727) );
  MUX2X1 U5206 ( .B(mem[16]), .A(mem[57]), .S(n5526), .Y(n4726) );
  MUX2X1 U5207 ( .B(n4725), .A(n4722), .S(n5593), .Y(n4729) );
  MUX2X1 U5208 ( .B(n4728), .A(n4713), .S(n16), .Y(n5467) );
  MUX2X1 U5209 ( .B(mem[1247]), .A(mem[1288]), .S(n5527), .Y(n4733) );
  MUX2X1 U5210 ( .B(mem[1165]), .A(mem[1206]), .S(n5527), .Y(n4732) );
  MUX2X1 U5211 ( .B(mem[1083]), .A(mem[1124]), .S(n5527), .Y(n4736) );
  MUX2X1 U5212 ( .B(mem[1001]), .A(mem[1042]), .S(n5527), .Y(n4735) );
  MUX2X1 U5213 ( .B(n4734), .A(n4731), .S(n5594), .Y(n4745) );
  MUX2X1 U5214 ( .B(mem[919]), .A(mem[960]), .S(n5527), .Y(n4739) );
  MUX2X1 U5215 ( .B(mem[837]), .A(mem[878]), .S(n5527), .Y(n4738) );
  MUX2X1 U5216 ( .B(mem[755]), .A(mem[796]), .S(n5527), .Y(n4742) );
  MUX2X1 U5217 ( .B(mem[673]), .A(mem[714]), .S(n5527), .Y(n4741) );
  MUX2X1 U5218 ( .B(n4740), .A(n4737), .S(n5594), .Y(n4744) );
  MUX2X1 U5219 ( .B(mem[591]), .A(mem[632]), .S(n5527), .Y(n4748) );
  MUX2X1 U5220 ( .B(mem[509]), .A(mem[550]), .S(n5527), .Y(n4747) );
  MUX2X1 U5221 ( .B(mem[427]), .A(mem[468]), .S(n5527), .Y(n4751) );
  MUX2X1 U5222 ( .B(mem[345]), .A(mem[386]), .S(n5527), .Y(n4750) );
  MUX2X1 U5223 ( .B(n4749), .A(n4746), .S(n5594), .Y(n4760) );
  MUX2X1 U5224 ( .B(mem[263]), .A(mem[304]), .S(n5528), .Y(n4754) );
  MUX2X1 U5225 ( .B(mem[181]), .A(mem[222]), .S(n5528), .Y(n4753) );
  MUX2X1 U5226 ( .B(mem[99]), .A(mem[140]), .S(n5528), .Y(n4757) );
  MUX2X1 U5227 ( .B(mem[17]), .A(mem[58]), .S(n5528), .Y(n4756) );
  MUX2X1 U5228 ( .B(n4755), .A(n4752), .S(n5594), .Y(n4759) );
  MUX2X1 U5229 ( .B(n4758), .A(n4743), .S(n16), .Y(n5468) );
  MUX2X1 U5230 ( .B(mem[1248]), .A(mem[1289]), .S(n5528), .Y(n4763) );
  MUX2X1 U5231 ( .B(mem[1166]), .A(mem[1207]), .S(n5528), .Y(n4762) );
  MUX2X1 U5232 ( .B(mem[1084]), .A(mem[1125]), .S(n5528), .Y(n4766) );
  MUX2X1 U5233 ( .B(mem[1002]), .A(mem[1043]), .S(n5528), .Y(n4765) );
  MUX2X1 U5234 ( .B(n4764), .A(n4761), .S(n5594), .Y(n4775) );
  MUX2X1 U5235 ( .B(mem[920]), .A(mem[961]), .S(n5528), .Y(n4769) );
  MUX2X1 U5236 ( .B(mem[838]), .A(mem[879]), .S(n5528), .Y(n4768) );
  MUX2X1 U5237 ( .B(mem[756]), .A(mem[797]), .S(n5528), .Y(n4772) );
  MUX2X1 U5238 ( .B(mem[674]), .A(mem[715]), .S(n5528), .Y(n4771) );
  MUX2X1 U5239 ( .B(n4770), .A(n4767), .S(n5594), .Y(n4774) );
  MUX2X1 U5240 ( .B(mem[592]), .A(mem[633]), .S(n5529), .Y(n4778) );
  MUX2X1 U5241 ( .B(mem[510]), .A(mem[551]), .S(n5529), .Y(n4777) );
  MUX2X1 U5242 ( .B(mem[428]), .A(mem[469]), .S(n5529), .Y(n4781) );
  MUX2X1 U5243 ( .B(mem[346]), .A(mem[387]), .S(n5529), .Y(n4780) );
  MUX2X1 U5244 ( .B(n4779), .A(n4776), .S(n5594), .Y(n4790) );
  MUX2X1 U5245 ( .B(mem[264]), .A(mem[305]), .S(n5529), .Y(n4784) );
  MUX2X1 U5246 ( .B(mem[182]), .A(mem[223]), .S(n5529), .Y(n4783) );
  MUX2X1 U5247 ( .B(mem[100]), .A(mem[141]), .S(n5529), .Y(n4787) );
  MUX2X1 U5248 ( .B(mem[18]), .A(mem[59]), .S(n5529), .Y(n4786) );
  MUX2X1 U5249 ( .B(n4785), .A(n4782), .S(n5594), .Y(n4789) );
  MUX2X1 U5250 ( .B(n4788), .A(n4773), .S(n16), .Y(n5469) );
  MUX2X1 U5251 ( .B(mem[1249]), .A(mem[1290]), .S(n5529), .Y(n4793) );
  MUX2X1 U5252 ( .B(mem[1167]), .A(mem[1208]), .S(n5529), .Y(n4792) );
  MUX2X1 U5253 ( .B(mem[1085]), .A(mem[1126]), .S(n5529), .Y(n4796) );
  MUX2X1 U5254 ( .B(mem[1003]), .A(mem[1044]), .S(n5529), .Y(n4795) );
  MUX2X1 U5255 ( .B(n4794), .A(n4791), .S(n5594), .Y(n4805) );
  MUX2X1 U5256 ( .B(mem[921]), .A(mem[962]), .S(n5530), .Y(n4799) );
  MUX2X1 U5257 ( .B(mem[839]), .A(mem[880]), .S(n5530), .Y(n4798) );
  MUX2X1 U5258 ( .B(mem[757]), .A(mem[798]), .S(n5530), .Y(n4802) );
  MUX2X1 U5259 ( .B(mem[675]), .A(mem[716]), .S(n5530), .Y(n4801) );
  MUX2X1 U5260 ( .B(n4800), .A(n4797), .S(n5594), .Y(n4804) );
  MUX2X1 U5261 ( .B(mem[593]), .A(mem[634]), .S(n5530), .Y(n4808) );
  MUX2X1 U5262 ( .B(mem[511]), .A(mem[552]), .S(n5530), .Y(n4807) );
  MUX2X1 U5263 ( .B(mem[429]), .A(mem[470]), .S(n5530), .Y(n4811) );
  MUX2X1 U5264 ( .B(mem[347]), .A(mem[388]), .S(n5530), .Y(n4810) );
  MUX2X1 U5265 ( .B(n4809), .A(n4806), .S(n5594), .Y(n4820) );
  MUX2X1 U5266 ( .B(mem[265]), .A(mem[306]), .S(n5530), .Y(n4814) );
  MUX2X1 U5267 ( .B(mem[183]), .A(mem[224]), .S(n5530), .Y(n4813) );
  MUX2X1 U5268 ( .B(mem[101]), .A(mem[142]), .S(n5530), .Y(n4817) );
  MUX2X1 U5269 ( .B(mem[19]), .A(mem[60]), .S(n5530), .Y(n4816) );
  MUX2X1 U5270 ( .B(n4815), .A(n4812), .S(n5594), .Y(n4819) );
  MUX2X1 U5271 ( .B(n4818), .A(n4803), .S(n16), .Y(n5470) );
  MUX2X1 U5272 ( .B(mem[1250]), .A(mem[1291]), .S(n5531), .Y(n4823) );
  MUX2X1 U5273 ( .B(mem[1168]), .A(mem[1209]), .S(n5531), .Y(n4822) );
  MUX2X1 U5274 ( .B(mem[1086]), .A(mem[1127]), .S(n5531), .Y(n4826) );
  MUX2X1 U5275 ( .B(mem[1004]), .A(mem[1045]), .S(n5531), .Y(n4825) );
  MUX2X1 U5276 ( .B(n4824), .A(n4821), .S(n5595), .Y(n4835) );
  MUX2X1 U5277 ( .B(mem[922]), .A(mem[963]), .S(n5531), .Y(n4829) );
  MUX2X1 U5278 ( .B(mem[840]), .A(mem[881]), .S(n5531), .Y(n4828) );
  MUX2X1 U5279 ( .B(mem[758]), .A(mem[799]), .S(n5531), .Y(n4832) );
  MUX2X1 U5280 ( .B(mem[676]), .A(mem[717]), .S(n5531), .Y(n4831) );
  MUX2X1 U5281 ( .B(n4830), .A(n4827), .S(n5595), .Y(n4834) );
  MUX2X1 U5282 ( .B(mem[594]), .A(mem[635]), .S(n5531), .Y(n4838) );
  MUX2X1 U5283 ( .B(mem[512]), .A(mem[553]), .S(n5531), .Y(n4837) );
  MUX2X1 U5284 ( .B(mem[430]), .A(mem[471]), .S(n5531), .Y(n4841) );
  MUX2X1 U5285 ( .B(mem[348]), .A(mem[389]), .S(n5531), .Y(n4840) );
  MUX2X1 U5286 ( .B(n4839), .A(n4836), .S(n5595), .Y(n4850) );
  MUX2X1 U5287 ( .B(mem[266]), .A(mem[307]), .S(n5532), .Y(n4844) );
  MUX2X1 U5288 ( .B(mem[184]), .A(mem[225]), .S(n5532), .Y(n4843) );
  MUX2X1 U5289 ( .B(mem[102]), .A(mem[143]), .S(n5532), .Y(n4847) );
  MUX2X1 U5290 ( .B(mem[20]), .A(mem[61]), .S(n5532), .Y(n4846) );
  MUX2X1 U5291 ( .B(n4845), .A(n4842), .S(n5595), .Y(n4849) );
  MUX2X1 U5292 ( .B(n4848), .A(n4833), .S(n16), .Y(n5471) );
  MUX2X1 U5293 ( .B(mem[1251]), .A(mem[1292]), .S(n5532), .Y(n4853) );
  MUX2X1 U5294 ( .B(mem[1169]), .A(mem[1210]), .S(n5532), .Y(n4852) );
  MUX2X1 U5295 ( .B(mem[1087]), .A(mem[1128]), .S(n5532), .Y(n4856) );
  MUX2X1 U5296 ( .B(mem[1005]), .A(mem[1046]), .S(n5532), .Y(n4855) );
  MUX2X1 U5297 ( .B(n4854), .A(n4851), .S(n5595), .Y(n4865) );
  MUX2X1 U5298 ( .B(mem[923]), .A(mem[964]), .S(n5532), .Y(n4859) );
  MUX2X1 U5299 ( .B(mem[841]), .A(mem[882]), .S(n5532), .Y(n4858) );
  MUX2X1 U5300 ( .B(mem[759]), .A(mem[800]), .S(n5532), .Y(n4862) );
  MUX2X1 U5301 ( .B(mem[677]), .A(mem[718]), .S(n5532), .Y(n4861) );
  MUX2X1 U5302 ( .B(n4860), .A(n4857), .S(n5595), .Y(n4864) );
  MUX2X1 U5303 ( .B(mem[595]), .A(mem[636]), .S(n5533), .Y(n4868) );
  MUX2X1 U5304 ( .B(mem[513]), .A(mem[554]), .S(n5533), .Y(n4867) );
  MUX2X1 U5305 ( .B(mem[431]), .A(mem[472]), .S(n5533), .Y(n4871) );
  MUX2X1 U5306 ( .B(mem[349]), .A(mem[390]), .S(n5533), .Y(n4870) );
  MUX2X1 U5307 ( .B(n4869), .A(n4866), .S(n5595), .Y(n4880) );
  MUX2X1 U5308 ( .B(mem[267]), .A(mem[308]), .S(n5533), .Y(n4874) );
  MUX2X1 U5309 ( .B(mem[185]), .A(mem[226]), .S(n5533), .Y(n4873) );
  MUX2X1 U5310 ( .B(mem[103]), .A(mem[144]), .S(n5533), .Y(n4877) );
  MUX2X1 U5311 ( .B(mem[21]), .A(mem[62]), .S(n5533), .Y(n4876) );
  MUX2X1 U5312 ( .B(n4875), .A(n4872), .S(n5595), .Y(n4879) );
  MUX2X1 U5313 ( .B(n4878), .A(n4863), .S(n16), .Y(n5472) );
  MUX2X1 U5314 ( .B(mem[1252]), .A(mem[1293]), .S(n5533), .Y(n4883) );
  MUX2X1 U5315 ( .B(mem[1170]), .A(mem[1211]), .S(n5533), .Y(n4882) );
  MUX2X1 U5316 ( .B(mem[1088]), .A(mem[1129]), .S(n5533), .Y(n4886) );
  MUX2X1 U5317 ( .B(mem[1006]), .A(mem[1047]), .S(n5533), .Y(n4885) );
  MUX2X1 U5318 ( .B(n4884), .A(n4881), .S(n5595), .Y(n4895) );
  MUX2X1 U5319 ( .B(mem[924]), .A(mem[965]), .S(n5534), .Y(n4889) );
  MUX2X1 U5320 ( .B(mem[842]), .A(mem[883]), .S(n5534), .Y(n4888) );
  MUX2X1 U5321 ( .B(mem[760]), .A(mem[801]), .S(n5534), .Y(n4892) );
  MUX2X1 U5322 ( .B(mem[678]), .A(mem[719]), .S(n5534), .Y(n4891) );
  MUX2X1 U5323 ( .B(n4890), .A(n4887), .S(n5595), .Y(n4894) );
  MUX2X1 U5324 ( .B(mem[596]), .A(mem[637]), .S(n5534), .Y(n4898) );
  MUX2X1 U5325 ( .B(mem[514]), .A(mem[555]), .S(n5534), .Y(n4897) );
  MUX2X1 U5326 ( .B(mem[432]), .A(mem[473]), .S(n5534), .Y(n4901) );
  MUX2X1 U5327 ( .B(mem[350]), .A(mem[391]), .S(n5534), .Y(n4900) );
  MUX2X1 U5328 ( .B(n4899), .A(n4896), .S(n5595), .Y(n4910) );
  MUX2X1 U5329 ( .B(mem[268]), .A(mem[309]), .S(n5534), .Y(n4904) );
  MUX2X1 U5330 ( .B(mem[186]), .A(mem[227]), .S(n5534), .Y(n4903) );
  MUX2X1 U5331 ( .B(mem[104]), .A(mem[145]), .S(n5534), .Y(n4907) );
  MUX2X1 U5332 ( .B(mem[22]), .A(mem[63]), .S(n5534), .Y(n4906) );
  MUX2X1 U5333 ( .B(n4905), .A(n4902), .S(n5595), .Y(n4909) );
  MUX2X1 U5334 ( .B(n4908), .A(n4893), .S(n16), .Y(n5473) );
  MUX2X1 U5335 ( .B(mem[1253]), .A(mem[1294]), .S(n5535), .Y(n4913) );
  MUX2X1 U5336 ( .B(mem[1171]), .A(mem[1212]), .S(n5535), .Y(n4912) );
  MUX2X1 U5337 ( .B(mem[1089]), .A(mem[1130]), .S(n5535), .Y(n4916) );
  MUX2X1 U5338 ( .B(mem[1007]), .A(mem[1048]), .S(n5535), .Y(n4915) );
  MUX2X1 U5339 ( .B(n4914), .A(n4911), .S(n14), .Y(n4925) );
  MUX2X1 U5340 ( .B(mem[925]), .A(mem[966]), .S(n5535), .Y(n4919) );
  MUX2X1 U5341 ( .B(mem[843]), .A(mem[884]), .S(n5535), .Y(n4918) );
  MUX2X1 U5342 ( .B(mem[761]), .A(mem[802]), .S(n5535), .Y(n4922) );
  MUX2X1 U5343 ( .B(mem[679]), .A(mem[720]), .S(n5535), .Y(n4921) );
  MUX2X1 U5344 ( .B(n4920), .A(n4917), .S(n14), .Y(n4924) );
  MUX2X1 U5345 ( .B(mem[597]), .A(mem[638]), .S(n5535), .Y(n4928) );
  MUX2X1 U5346 ( .B(mem[515]), .A(mem[556]), .S(n5535), .Y(n4927) );
  MUX2X1 U5347 ( .B(mem[433]), .A(mem[474]), .S(n5535), .Y(n4931) );
  MUX2X1 U5348 ( .B(mem[351]), .A(mem[392]), .S(n5535), .Y(n4930) );
  MUX2X1 U5349 ( .B(n4929), .A(n4926), .S(n14), .Y(n4940) );
  MUX2X1 U5350 ( .B(mem[269]), .A(mem[310]), .S(n5536), .Y(n4934) );
  MUX2X1 U5351 ( .B(mem[187]), .A(mem[228]), .S(n5536), .Y(n4933) );
  MUX2X1 U5352 ( .B(mem[105]), .A(mem[146]), .S(n5536), .Y(n4937) );
  MUX2X1 U5353 ( .B(mem[23]), .A(mem[64]), .S(n5536), .Y(n4936) );
  MUX2X1 U5354 ( .B(n4935), .A(n4932), .S(n14), .Y(n4939) );
  MUX2X1 U5355 ( .B(n4938), .A(n4923), .S(n16), .Y(n5474) );
  MUX2X1 U5356 ( .B(mem[1254]), .A(mem[1295]), .S(n5536), .Y(n4943) );
  MUX2X1 U5357 ( .B(mem[1172]), .A(mem[1213]), .S(n5536), .Y(n4942) );
  MUX2X1 U5358 ( .B(mem[1090]), .A(mem[1131]), .S(n5536), .Y(n4946) );
  MUX2X1 U5359 ( .B(mem[1008]), .A(mem[1049]), .S(n5536), .Y(n4945) );
  MUX2X1 U5360 ( .B(n4944), .A(n4941), .S(n14), .Y(n4955) );
  MUX2X1 U5361 ( .B(mem[926]), .A(mem[967]), .S(n5536), .Y(n4949) );
  MUX2X1 U5362 ( .B(mem[844]), .A(mem[885]), .S(n5536), .Y(n4948) );
  MUX2X1 U5363 ( .B(mem[762]), .A(mem[803]), .S(n5536), .Y(n4952) );
  MUX2X1 U5364 ( .B(mem[680]), .A(mem[721]), .S(n5536), .Y(n4951) );
  MUX2X1 U5365 ( .B(n4950), .A(n4947), .S(n14), .Y(n4954) );
  MUX2X1 U5366 ( .B(mem[598]), .A(mem[639]), .S(n5537), .Y(n4958) );
  MUX2X1 U5367 ( .B(mem[516]), .A(mem[557]), .S(n5537), .Y(n4957) );
  MUX2X1 U5368 ( .B(mem[434]), .A(mem[475]), .S(n5537), .Y(n4961) );
  MUX2X1 U5369 ( .B(mem[352]), .A(mem[393]), .S(n5537), .Y(n4960) );
  MUX2X1 U5370 ( .B(n4959), .A(n4956), .S(n14), .Y(n4970) );
  MUX2X1 U5371 ( .B(mem[270]), .A(mem[311]), .S(n5537), .Y(n4964) );
  MUX2X1 U5372 ( .B(mem[188]), .A(mem[229]), .S(n5537), .Y(n4963) );
  MUX2X1 U5373 ( .B(mem[106]), .A(mem[147]), .S(n5537), .Y(n4967) );
  MUX2X1 U5374 ( .B(mem[24]), .A(mem[65]), .S(n5537), .Y(n4966) );
  MUX2X1 U5375 ( .B(n4965), .A(n4962), .S(n14), .Y(n4969) );
  MUX2X1 U5376 ( .B(n4968), .A(n4953), .S(n16), .Y(n5475) );
  MUX2X1 U5377 ( .B(mem[1255]), .A(mem[1296]), .S(n5537), .Y(n4973) );
  MUX2X1 U5378 ( .B(mem[1173]), .A(mem[1214]), .S(n5537), .Y(n4972) );
  MUX2X1 U5379 ( .B(mem[1091]), .A(mem[1132]), .S(n5537), .Y(n4976) );
  MUX2X1 U5380 ( .B(mem[1009]), .A(mem[1050]), .S(n5537), .Y(n4975) );
  MUX2X1 U5381 ( .B(n4974), .A(n4971), .S(n14), .Y(n4985) );
  MUX2X1 U5382 ( .B(mem[927]), .A(mem[968]), .S(n5538), .Y(n4979) );
  MUX2X1 U5383 ( .B(mem[845]), .A(mem[886]), .S(n5538), .Y(n4978) );
  MUX2X1 U5384 ( .B(mem[763]), .A(mem[804]), .S(n5538), .Y(n4982) );
  MUX2X1 U5385 ( .B(mem[681]), .A(mem[722]), .S(n5538), .Y(n4981) );
  MUX2X1 U5386 ( .B(n4980), .A(n4977), .S(n14), .Y(n4984) );
  MUX2X1 U5387 ( .B(mem[599]), .A(mem[640]), .S(n5538), .Y(n4988) );
  MUX2X1 U5388 ( .B(mem[517]), .A(mem[558]), .S(n5538), .Y(n4987) );
  MUX2X1 U5389 ( .B(mem[435]), .A(mem[476]), .S(n5538), .Y(n4991) );
  MUX2X1 U5390 ( .B(mem[353]), .A(mem[394]), .S(n5538), .Y(n4990) );
  MUX2X1 U5391 ( .B(n4989), .A(n4986), .S(n14), .Y(n5000) );
  MUX2X1 U5392 ( .B(mem[271]), .A(mem[312]), .S(n5538), .Y(n4994) );
  MUX2X1 U5393 ( .B(mem[189]), .A(mem[230]), .S(n5538), .Y(n4993) );
  MUX2X1 U5394 ( .B(mem[107]), .A(mem[148]), .S(n5538), .Y(n4997) );
  MUX2X1 U5395 ( .B(mem[25]), .A(mem[66]), .S(n5538), .Y(n4996) );
  MUX2X1 U5396 ( .B(n4995), .A(n4992), .S(n14), .Y(n4999) );
  MUX2X1 U5397 ( .B(n4998), .A(n4983), .S(n16), .Y(n5476) );
  MUX2X1 U5398 ( .B(mem[1256]), .A(mem[1297]), .S(n5539), .Y(n5003) );
  MUX2X1 U5399 ( .B(mem[1174]), .A(mem[1215]), .S(n5539), .Y(n5002) );
  MUX2X1 U5400 ( .B(mem[1092]), .A(mem[1133]), .S(n5539), .Y(n5006) );
  MUX2X1 U5401 ( .B(mem[1010]), .A(mem[1051]), .S(n5539), .Y(n5005) );
  MUX2X1 U5402 ( .B(n5004), .A(n5001), .S(n14), .Y(n5015) );
  MUX2X1 U5403 ( .B(mem[928]), .A(mem[969]), .S(n5539), .Y(n5009) );
  MUX2X1 U5404 ( .B(mem[846]), .A(mem[887]), .S(n5539), .Y(n5008) );
  MUX2X1 U5405 ( .B(mem[764]), .A(mem[805]), .S(n5539), .Y(n5012) );
  MUX2X1 U5406 ( .B(mem[682]), .A(mem[723]), .S(n5539), .Y(n5011) );
  MUX2X1 U5407 ( .B(n5010), .A(n5007), .S(n14), .Y(n5014) );
  MUX2X1 U5408 ( .B(mem[600]), .A(mem[641]), .S(n5539), .Y(n5018) );
  MUX2X1 U5409 ( .B(mem[518]), .A(mem[559]), .S(n5539), .Y(n5017) );
  MUX2X1 U5410 ( .B(mem[436]), .A(mem[477]), .S(n5539), .Y(n5021) );
  MUX2X1 U5411 ( .B(mem[354]), .A(mem[395]), .S(n5539), .Y(n5020) );
  MUX2X1 U5412 ( .B(n5019), .A(n5016), .S(n14), .Y(n5030) );
  MUX2X1 U5413 ( .B(mem[272]), .A(mem[313]), .S(n5540), .Y(n5024) );
  MUX2X1 U5414 ( .B(mem[190]), .A(mem[231]), .S(n5540), .Y(n5023) );
  MUX2X1 U5415 ( .B(mem[108]), .A(mem[149]), .S(n5540), .Y(n5027) );
  MUX2X1 U5416 ( .B(mem[26]), .A(mem[67]), .S(n5540), .Y(n5026) );
  MUX2X1 U5417 ( .B(n5025), .A(n5022), .S(n14), .Y(n5029) );
  MUX2X1 U5418 ( .B(n5028), .A(n5013), .S(n16), .Y(n5477) );
  MUX2X1 U5419 ( .B(mem[1257]), .A(mem[1298]), .S(n5540), .Y(n5033) );
  MUX2X1 U5420 ( .B(mem[1175]), .A(mem[1216]), .S(n5540), .Y(n5032) );
  MUX2X1 U5421 ( .B(mem[1093]), .A(mem[1134]), .S(n5540), .Y(n5036) );
  MUX2X1 U5422 ( .B(mem[1011]), .A(mem[1052]), .S(n5540), .Y(n5035) );
  MUX2X1 U5423 ( .B(n5034), .A(n5031), .S(n14), .Y(n5045) );
  MUX2X1 U5424 ( .B(mem[929]), .A(mem[970]), .S(n5540), .Y(n5039) );
  MUX2X1 U5425 ( .B(mem[847]), .A(mem[888]), .S(n5540), .Y(n5038) );
  MUX2X1 U5426 ( .B(mem[765]), .A(mem[806]), .S(n5540), .Y(n5042) );
  MUX2X1 U5427 ( .B(mem[683]), .A(mem[724]), .S(n5540), .Y(n5041) );
  MUX2X1 U5428 ( .B(n5040), .A(n5037), .S(n14), .Y(n5044) );
  MUX2X1 U5429 ( .B(mem[601]), .A(mem[642]), .S(n5541), .Y(n5048) );
  MUX2X1 U5430 ( .B(mem[519]), .A(mem[560]), .S(n5541), .Y(n5047) );
  MUX2X1 U5431 ( .B(mem[437]), .A(mem[478]), .S(n5541), .Y(n5051) );
  MUX2X1 U5432 ( .B(mem[355]), .A(mem[396]), .S(n5541), .Y(n5050) );
  MUX2X1 U5433 ( .B(n5049), .A(n5046), .S(n14), .Y(n5060) );
  MUX2X1 U5434 ( .B(mem[273]), .A(mem[314]), .S(n5541), .Y(n5054) );
  MUX2X1 U5435 ( .B(mem[191]), .A(mem[232]), .S(n5541), .Y(n5053) );
  MUX2X1 U5436 ( .B(mem[109]), .A(mem[150]), .S(n5541), .Y(n5057) );
  MUX2X1 U5437 ( .B(mem[27]), .A(mem[68]), .S(n5541), .Y(n5056) );
  MUX2X1 U5438 ( .B(n5055), .A(n5052), .S(n14), .Y(n5059) );
  MUX2X1 U5439 ( .B(n5058), .A(n5043), .S(n16), .Y(n5478) );
  MUX2X1 U5440 ( .B(mem[1258]), .A(mem[1299]), .S(n5541), .Y(n5063) );
  MUX2X1 U5441 ( .B(mem[1176]), .A(mem[1217]), .S(n5541), .Y(n5062) );
  MUX2X1 U5442 ( .B(mem[1094]), .A(mem[1135]), .S(n5541), .Y(n5066) );
  MUX2X1 U5443 ( .B(mem[1012]), .A(mem[1053]), .S(n5541), .Y(n5065) );
  MUX2X1 U5444 ( .B(n5064), .A(n5061), .S(n14), .Y(n5075) );
  MUX2X1 U5445 ( .B(mem[930]), .A(mem[971]), .S(n5542), .Y(n5069) );
  MUX2X1 U5446 ( .B(mem[848]), .A(mem[889]), .S(n5542), .Y(n5068) );
  MUX2X1 U5447 ( .B(mem[766]), .A(mem[807]), .S(n5542), .Y(n5072) );
  MUX2X1 U5448 ( .B(mem[684]), .A(mem[725]), .S(n5542), .Y(n5071) );
  MUX2X1 U5449 ( .B(n5070), .A(n5067), .S(n14), .Y(n5074) );
  MUX2X1 U5450 ( .B(mem[602]), .A(mem[643]), .S(n5542), .Y(n5078) );
  MUX2X1 U5451 ( .B(mem[520]), .A(mem[561]), .S(n5542), .Y(n5077) );
  MUX2X1 U5452 ( .B(mem[438]), .A(mem[479]), .S(n5542), .Y(n5081) );
  MUX2X1 U5453 ( .B(mem[356]), .A(mem[397]), .S(n5542), .Y(n5080) );
  MUX2X1 U5454 ( .B(n5079), .A(n5076), .S(n14), .Y(n5090) );
  MUX2X1 U5455 ( .B(mem[274]), .A(mem[315]), .S(n5542), .Y(n5084) );
  MUX2X1 U5456 ( .B(mem[192]), .A(mem[233]), .S(n5542), .Y(n5083) );
  MUX2X1 U5457 ( .B(mem[110]), .A(mem[151]), .S(n5542), .Y(n5087) );
  MUX2X1 U5458 ( .B(mem[28]), .A(mem[69]), .S(n5542), .Y(n5086) );
  MUX2X1 U5459 ( .B(n5085), .A(n5082), .S(n14), .Y(n5089) );
  MUX2X1 U5460 ( .B(n5088), .A(n5073), .S(n16), .Y(n5479) );
  MUX2X1 U5461 ( .B(mem[1259]), .A(mem[1300]), .S(n5543), .Y(n5093) );
  MUX2X1 U5462 ( .B(mem[1177]), .A(mem[1218]), .S(n5543), .Y(n5092) );
  MUX2X1 U5463 ( .B(mem[1095]), .A(mem[1136]), .S(n5543), .Y(n5096) );
  MUX2X1 U5464 ( .B(mem[1013]), .A(mem[1054]), .S(n5543), .Y(n5095) );
  MUX2X1 U5465 ( .B(n5094), .A(n5091), .S(n14), .Y(n5105) );
  MUX2X1 U5466 ( .B(mem[931]), .A(mem[972]), .S(n5543), .Y(n5099) );
  MUX2X1 U5467 ( .B(mem[849]), .A(mem[890]), .S(n5543), .Y(n5098) );
  MUX2X1 U5468 ( .B(mem[767]), .A(mem[808]), .S(n5543), .Y(n5102) );
  MUX2X1 U5469 ( .B(mem[685]), .A(mem[726]), .S(n5543), .Y(n5101) );
  MUX2X1 U5470 ( .B(n5100), .A(n5097), .S(n14), .Y(n5104) );
  MUX2X1 U5471 ( .B(mem[603]), .A(mem[644]), .S(n5543), .Y(n5108) );
  MUX2X1 U5472 ( .B(mem[521]), .A(mem[562]), .S(n5543), .Y(n5107) );
  MUX2X1 U5473 ( .B(mem[439]), .A(mem[480]), .S(n5543), .Y(n5111) );
  MUX2X1 U5474 ( .B(mem[357]), .A(mem[398]), .S(n5543), .Y(n5110) );
  MUX2X1 U5475 ( .B(n5109), .A(n5106), .S(n14), .Y(n5120) );
  MUX2X1 U5476 ( .B(mem[275]), .A(mem[316]), .S(n5544), .Y(n5114) );
  MUX2X1 U5477 ( .B(mem[193]), .A(mem[234]), .S(n5544), .Y(n5113) );
  MUX2X1 U5478 ( .B(mem[111]), .A(mem[152]), .S(n5544), .Y(n5117) );
  MUX2X1 U5479 ( .B(mem[29]), .A(mem[70]), .S(n5544), .Y(n5116) );
  MUX2X1 U5480 ( .B(n5115), .A(n5112), .S(n14), .Y(n5119) );
  MUX2X1 U5481 ( .B(n5118), .A(n5103), .S(n16), .Y(n5480) );
  MUX2X1 U5482 ( .B(mem[1260]), .A(mem[1301]), .S(n5544), .Y(n5123) );
  MUX2X1 U5483 ( .B(mem[1178]), .A(mem[1219]), .S(n5544), .Y(n5122) );
  MUX2X1 U5484 ( .B(mem[1096]), .A(mem[1137]), .S(n5544), .Y(n5126) );
  MUX2X1 U5485 ( .B(mem[1014]), .A(mem[1055]), .S(n5544), .Y(n5125) );
  MUX2X1 U5486 ( .B(n5124), .A(n5121), .S(n14), .Y(n5135) );
  MUX2X1 U5487 ( .B(mem[932]), .A(mem[973]), .S(n5544), .Y(n5129) );
  MUX2X1 U5488 ( .B(mem[850]), .A(mem[891]), .S(n5544), .Y(n5128) );
  MUX2X1 U5489 ( .B(mem[768]), .A(mem[809]), .S(n5544), .Y(n5132) );
  MUX2X1 U5490 ( .B(mem[686]), .A(mem[727]), .S(n5544), .Y(n5131) );
  MUX2X1 U5491 ( .B(n5130), .A(n5127), .S(n14), .Y(n5134) );
  MUX2X1 U5492 ( .B(mem[604]), .A(mem[645]), .S(n5545), .Y(n5138) );
  MUX2X1 U5493 ( .B(mem[522]), .A(mem[563]), .S(n5545), .Y(n5137) );
  MUX2X1 U5494 ( .B(mem[440]), .A(mem[481]), .S(n5545), .Y(n5141) );
  MUX2X1 U5495 ( .B(mem[358]), .A(mem[399]), .S(n5545), .Y(n5140) );
  MUX2X1 U5496 ( .B(n5139), .A(n5136), .S(n14), .Y(n5150) );
  MUX2X1 U5497 ( .B(mem[276]), .A(mem[317]), .S(n5545), .Y(n5144) );
  MUX2X1 U5498 ( .B(mem[194]), .A(mem[235]), .S(n5545), .Y(n5143) );
  MUX2X1 U5499 ( .B(mem[112]), .A(mem[153]), .S(n5545), .Y(n5147) );
  MUX2X1 U5500 ( .B(mem[30]), .A(mem[71]), .S(n5545), .Y(n5146) );
  MUX2X1 U5501 ( .B(n5145), .A(n5142), .S(n14), .Y(n5149) );
  MUX2X1 U5502 ( .B(n5148), .A(n5133), .S(n16), .Y(n5481) );
  MUX2X1 U5503 ( .B(mem[1261]), .A(mem[1302]), .S(n5545), .Y(n5153) );
  MUX2X1 U5504 ( .B(mem[1179]), .A(mem[1220]), .S(n5545), .Y(n5152) );
  MUX2X1 U5505 ( .B(mem[1097]), .A(mem[1138]), .S(n5545), .Y(n5156) );
  MUX2X1 U5506 ( .B(mem[1015]), .A(mem[1056]), .S(n5545), .Y(n5155) );
  MUX2X1 U5507 ( .B(n5154), .A(n5151), .S(n14), .Y(n5165) );
  MUX2X1 U5508 ( .B(mem[933]), .A(mem[974]), .S(n5546), .Y(n5159) );
  MUX2X1 U5509 ( .B(mem[851]), .A(mem[892]), .S(n5546), .Y(n5158) );
  MUX2X1 U5510 ( .B(mem[769]), .A(mem[810]), .S(n5546), .Y(n5162) );
  MUX2X1 U5511 ( .B(mem[687]), .A(mem[728]), .S(n5546), .Y(n5161) );
  MUX2X1 U5512 ( .B(n5160), .A(n5157), .S(n14), .Y(n5164) );
  MUX2X1 U5513 ( .B(mem[605]), .A(mem[646]), .S(n5546), .Y(n5168) );
  MUX2X1 U5514 ( .B(mem[523]), .A(mem[564]), .S(n5546), .Y(n5167) );
  MUX2X1 U5515 ( .B(mem[441]), .A(mem[482]), .S(n5546), .Y(n5171) );
  MUX2X1 U5516 ( .B(mem[359]), .A(mem[400]), .S(n5546), .Y(n5170) );
  MUX2X1 U5517 ( .B(n5169), .A(n5166), .S(n14), .Y(n5180) );
  MUX2X1 U5518 ( .B(mem[277]), .A(mem[318]), .S(n5546), .Y(n5174) );
  MUX2X1 U5519 ( .B(mem[195]), .A(mem[236]), .S(n5546), .Y(n5173) );
  MUX2X1 U5520 ( .B(mem[113]), .A(mem[154]), .S(n5546), .Y(n5177) );
  MUX2X1 U5521 ( .B(mem[31]), .A(mem[72]), .S(n5546), .Y(n5176) );
  MUX2X1 U5522 ( .B(n5175), .A(n5172), .S(n14), .Y(n5179) );
  MUX2X1 U5523 ( .B(n5178), .A(n5163), .S(n16), .Y(n5482) );
  MUX2X1 U5524 ( .B(mem[1262]), .A(mem[1303]), .S(n5547), .Y(n5183) );
  MUX2X1 U5525 ( .B(mem[1180]), .A(mem[1221]), .S(n5547), .Y(n5182) );
  MUX2X1 U5526 ( .B(mem[1098]), .A(mem[1139]), .S(n5547), .Y(n5186) );
  MUX2X1 U5527 ( .B(mem[1016]), .A(mem[1057]), .S(n5547), .Y(n5185) );
  MUX2X1 U5528 ( .B(n5184), .A(n5181), .S(n14), .Y(n5195) );
  MUX2X1 U5529 ( .B(mem[934]), .A(mem[975]), .S(n5547), .Y(n5189) );
  MUX2X1 U5530 ( .B(mem[852]), .A(mem[893]), .S(n5547), .Y(n5188) );
  MUX2X1 U5531 ( .B(mem[770]), .A(mem[811]), .S(n5547), .Y(n5192) );
  MUX2X1 U5532 ( .B(mem[688]), .A(mem[729]), .S(n5547), .Y(n5191) );
  MUX2X1 U5533 ( .B(n5190), .A(n5187), .S(n14), .Y(n5194) );
  MUX2X1 U5534 ( .B(mem[606]), .A(mem[647]), .S(n5547), .Y(n5198) );
  MUX2X1 U5535 ( .B(mem[524]), .A(mem[565]), .S(n5547), .Y(n5197) );
  MUX2X1 U5536 ( .B(mem[442]), .A(mem[483]), .S(n5547), .Y(n5201) );
  MUX2X1 U5537 ( .B(mem[360]), .A(mem[401]), .S(n5547), .Y(n5200) );
  MUX2X1 U5538 ( .B(n5199), .A(n5196), .S(n14), .Y(n5210) );
  MUX2X1 U5539 ( .B(mem[278]), .A(mem[319]), .S(n5548), .Y(n5204) );
  MUX2X1 U5540 ( .B(mem[196]), .A(mem[237]), .S(n5548), .Y(n5203) );
  MUX2X1 U5541 ( .B(mem[114]), .A(mem[155]), .S(n5548), .Y(n5207) );
  MUX2X1 U5542 ( .B(mem[32]), .A(mem[73]), .S(n5548), .Y(n5206) );
  MUX2X1 U5543 ( .B(n5205), .A(n5202), .S(n14), .Y(n5209) );
  MUX2X1 U5544 ( .B(n5208), .A(n5193), .S(n16), .Y(n5483) );
  MUX2X1 U5545 ( .B(mem[1263]), .A(mem[1304]), .S(n5548), .Y(n5213) );
  MUX2X1 U5546 ( .B(mem[1181]), .A(mem[1222]), .S(n5548), .Y(n5212) );
  MUX2X1 U5547 ( .B(mem[1099]), .A(mem[1140]), .S(n5548), .Y(n5216) );
  MUX2X1 U5548 ( .B(mem[1017]), .A(mem[1058]), .S(n5548), .Y(n5215) );
  MUX2X1 U5549 ( .B(n5214), .A(n5211), .S(n14), .Y(n5225) );
  MUX2X1 U5550 ( .B(mem[935]), .A(mem[976]), .S(n5548), .Y(n5219) );
  MUX2X1 U5551 ( .B(mem[853]), .A(mem[894]), .S(n5548), .Y(n5218) );
  MUX2X1 U5552 ( .B(mem[771]), .A(mem[812]), .S(n5548), .Y(n5222) );
  MUX2X1 U5553 ( .B(mem[689]), .A(mem[730]), .S(n5548), .Y(n5221) );
  MUX2X1 U5554 ( .B(n5220), .A(n5217), .S(n14), .Y(n5224) );
  MUX2X1 U5555 ( .B(mem[607]), .A(mem[648]), .S(n5549), .Y(n5228) );
  MUX2X1 U5556 ( .B(mem[525]), .A(mem[566]), .S(n5549), .Y(n5227) );
  MUX2X1 U5557 ( .B(mem[443]), .A(mem[484]), .S(n5549), .Y(n5231) );
  MUX2X1 U5558 ( .B(mem[361]), .A(mem[402]), .S(n5549), .Y(n5230) );
  MUX2X1 U5559 ( .B(n5229), .A(n5226), .S(n14), .Y(n5240) );
  MUX2X1 U5560 ( .B(mem[279]), .A(mem[320]), .S(n5549), .Y(n5234) );
  MUX2X1 U5561 ( .B(mem[197]), .A(mem[238]), .S(n5549), .Y(n5233) );
  MUX2X1 U5562 ( .B(mem[115]), .A(mem[156]), .S(n5549), .Y(n5237) );
  MUX2X1 U5563 ( .B(mem[33]), .A(mem[74]), .S(n5549), .Y(n5236) );
  MUX2X1 U5564 ( .B(n5235), .A(n5232), .S(n14), .Y(n5239) );
  MUX2X1 U5565 ( .B(n5238), .A(n5223), .S(n16), .Y(n5484) );
  MUX2X1 U5566 ( .B(mem[1264]), .A(mem[1305]), .S(n5549), .Y(n5243) );
  MUX2X1 U5567 ( .B(mem[1182]), .A(mem[1223]), .S(n5549), .Y(n5242) );
  MUX2X1 U5568 ( .B(mem[1100]), .A(mem[1141]), .S(n5549), .Y(n5246) );
  MUX2X1 U5569 ( .B(mem[1018]), .A(mem[1059]), .S(n5549), .Y(n5245) );
  MUX2X1 U5570 ( .B(n5244), .A(n5241), .S(n14), .Y(n5255) );
  MUX2X1 U5571 ( .B(mem[936]), .A(mem[977]), .S(n5550), .Y(n5249) );
  MUX2X1 U5572 ( .B(mem[854]), .A(mem[895]), .S(n5550), .Y(n5248) );
  MUX2X1 U5573 ( .B(mem[772]), .A(mem[813]), .S(n5550), .Y(n5252) );
  MUX2X1 U5574 ( .B(mem[690]), .A(mem[731]), .S(n5550), .Y(n5251) );
  MUX2X1 U5575 ( .B(n5250), .A(n5247), .S(n14), .Y(n5254) );
  MUX2X1 U5576 ( .B(mem[608]), .A(mem[649]), .S(n5550), .Y(n5258) );
  MUX2X1 U5577 ( .B(mem[526]), .A(mem[567]), .S(n5550), .Y(n5257) );
  MUX2X1 U5578 ( .B(mem[444]), .A(mem[485]), .S(n5550), .Y(n5261) );
  MUX2X1 U5579 ( .B(mem[362]), .A(mem[403]), .S(n5550), .Y(n5260) );
  MUX2X1 U5580 ( .B(n5259), .A(n5256), .S(n14), .Y(n5270) );
  MUX2X1 U5581 ( .B(mem[280]), .A(mem[321]), .S(n5550), .Y(n5264) );
  MUX2X1 U5582 ( .B(mem[198]), .A(mem[239]), .S(n5550), .Y(n5263) );
  MUX2X1 U5583 ( .B(mem[116]), .A(mem[157]), .S(n5550), .Y(n5267) );
  MUX2X1 U5584 ( .B(mem[34]), .A(mem[75]), .S(n5550), .Y(n5266) );
  MUX2X1 U5585 ( .B(n5265), .A(n5262), .S(n14), .Y(n5269) );
  MUX2X1 U5586 ( .B(n5268), .A(n5253), .S(n16), .Y(n5485) );
  MUX2X1 U5587 ( .B(mem[1265]), .A(mem[1306]), .S(n5551), .Y(n5273) );
  MUX2X1 U5588 ( .B(mem[1183]), .A(mem[1224]), .S(n5551), .Y(n5272) );
  MUX2X1 U5589 ( .B(mem[1101]), .A(mem[1142]), .S(n5551), .Y(n5276) );
  MUX2X1 U5590 ( .B(mem[1019]), .A(mem[1060]), .S(n5551), .Y(n5275) );
  MUX2X1 U5591 ( .B(n5274), .A(n5271), .S(n14), .Y(n5285) );
  MUX2X1 U5592 ( .B(mem[937]), .A(mem[978]), .S(n5551), .Y(n5279) );
  MUX2X1 U5593 ( .B(mem[855]), .A(mem[896]), .S(n5551), .Y(n5278) );
  MUX2X1 U5594 ( .B(mem[773]), .A(mem[814]), .S(n5551), .Y(n5282) );
  MUX2X1 U5595 ( .B(mem[691]), .A(mem[732]), .S(n5551), .Y(n5281) );
  MUX2X1 U5596 ( .B(n5280), .A(n5277), .S(n14), .Y(n5284) );
  MUX2X1 U5597 ( .B(mem[609]), .A(mem[650]), .S(n5551), .Y(n5288) );
  MUX2X1 U5598 ( .B(mem[527]), .A(mem[568]), .S(n5551), .Y(n5287) );
  MUX2X1 U5599 ( .B(mem[445]), .A(mem[486]), .S(n5551), .Y(n5291) );
  MUX2X1 U5600 ( .B(mem[363]), .A(mem[404]), .S(n5551), .Y(n5290) );
  MUX2X1 U5601 ( .B(n5289), .A(n5286), .S(n14), .Y(n5300) );
  MUX2X1 U5602 ( .B(mem[281]), .A(mem[322]), .S(n5552), .Y(n5294) );
  MUX2X1 U5603 ( .B(mem[199]), .A(mem[240]), .S(n5552), .Y(n5293) );
  MUX2X1 U5604 ( .B(mem[117]), .A(mem[158]), .S(n5552), .Y(n5297) );
  MUX2X1 U5605 ( .B(mem[35]), .A(mem[76]), .S(n5552), .Y(n5296) );
  MUX2X1 U5606 ( .B(n5295), .A(n5292), .S(n14), .Y(n5299) );
  MUX2X1 U5607 ( .B(n5298), .A(n5283), .S(n16), .Y(n5486) );
  MUX2X1 U5608 ( .B(mem[1266]), .A(mem[1307]), .S(n5552), .Y(n5303) );
  MUX2X1 U5609 ( .B(mem[1184]), .A(mem[1225]), .S(n5552), .Y(n5302) );
  MUX2X1 U5610 ( .B(mem[1102]), .A(mem[1143]), .S(n5552), .Y(n5306) );
  MUX2X1 U5611 ( .B(mem[1020]), .A(mem[1061]), .S(n5552), .Y(n5305) );
  MUX2X1 U5612 ( .B(n5304), .A(n5301), .S(n14), .Y(n5315) );
  MUX2X1 U5613 ( .B(mem[938]), .A(mem[979]), .S(n5552), .Y(n5309) );
  MUX2X1 U5614 ( .B(mem[856]), .A(mem[897]), .S(n5552), .Y(n5308) );
  MUX2X1 U5615 ( .B(mem[774]), .A(mem[815]), .S(n5552), .Y(n5312) );
  MUX2X1 U5616 ( .B(mem[692]), .A(mem[733]), .S(n5552), .Y(n5311) );
  MUX2X1 U5617 ( .B(n5310), .A(n5307), .S(n14), .Y(n5314) );
  MUX2X1 U5618 ( .B(mem[610]), .A(mem[651]), .S(n5553), .Y(n5318) );
  MUX2X1 U5619 ( .B(mem[528]), .A(mem[569]), .S(n5553), .Y(n5317) );
  MUX2X1 U5620 ( .B(mem[446]), .A(mem[487]), .S(n5553), .Y(n5321) );
  MUX2X1 U5621 ( .B(mem[364]), .A(mem[405]), .S(n5553), .Y(n5320) );
  MUX2X1 U5622 ( .B(n5319), .A(n5316), .S(n14), .Y(n5330) );
  MUX2X1 U5623 ( .B(mem[282]), .A(mem[323]), .S(n5553), .Y(n5324) );
  MUX2X1 U5624 ( .B(mem[200]), .A(mem[241]), .S(n5553), .Y(n5323) );
  MUX2X1 U5625 ( .B(mem[118]), .A(mem[159]), .S(n5553), .Y(n5327) );
  MUX2X1 U5626 ( .B(mem[36]), .A(mem[77]), .S(n5553), .Y(n5326) );
  MUX2X1 U5627 ( .B(n5325), .A(n5322), .S(n14), .Y(n5329) );
  MUX2X1 U5628 ( .B(n5328), .A(n5313), .S(n16), .Y(n5487) );
  MUX2X1 U5629 ( .B(mem[1267]), .A(mem[1308]), .S(n5553), .Y(n5333) );
  MUX2X1 U5630 ( .B(mem[1185]), .A(mem[1226]), .S(n5553), .Y(n5332) );
  MUX2X1 U5631 ( .B(mem[1103]), .A(mem[1144]), .S(n5553), .Y(n5336) );
  MUX2X1 U5632 ( .B(mem[1021]), .A(mem[1062]), .S(n5553), .Y(n5335) );
  MUX2X1 U5633 ( .B(n5334), .A(n5331), .S(n14), .Y(n5345) );
  MUX2X1 U5634 ( .B(mem[939]), .A(mem[980]), .S(n5554), .Y(n5339) );
  MUX2X1 U5635 ( .B(mem[857]), .A(mem[898]), .S(n5554), .Y(n5338) );
  MUX2X1 U5636 ( .B(mem[775]), .A(mem[816]), .S(n5554), .Y(n5342) );
  MUX2X1 U5637 ( .B(mem[693]), .A(mem[734]), .S(n5554), .Y(n5341) );
  MUX2X1 U5638 ( .B(n5340), .A(n5337), .S(n14), .Y(n5344) );
  MUX2X1 U5639 ( .B(mem[611]), .A(mem[652]), .S(n5554), .Y(n5348) );
  MUX2X1 U5640 ( .B(mem[529]), .A(mem[570]), .S(n5554), .Y(n5347) );
  MUX2X1 U5641 ( .B(mem[447]), .A(mem[488]), .S(n5554), .Y(n5351) );
  MUX2X1 U5642 ( .B(mem[365]), .A(mem[406]), .S(n5554), .Y(n5350) );
  MUX2X1 U5643 ( .B(n5349), .A(n5346), .S(n14), .Y(n5360) );
  MUX2X1 U5644 ( .B(mem[283]), .A(mem[324]), .S(n5554), .Y(n5354) );
  MUX2X1 U5645 ( .B(mem[201]), .A(mem[242]), .S(n5554), .Y(n5353) );
  MUX2X1 U5646 ( .B(mem[119]), .A(mem[160]), .S(n5554), .Y(n5357) );
  MUX2X1 U5647 ( .B(mem[37]), .A(mem[78]), .S(n5554), .Y(n5356) );
  MUX2X1 U5648 ( .B(n5355), .A(n5352), .S(n14), .Y(n5359) );
  MUX2X1 U5649 ( .B(n5358), .A(n5343), .S(n16), .Y(n5488) );
  MUX2X1 U5650 ( .B(mem[1268]), .A(mem[1309]), .S(n5555), .Y(n5363) );
  MUX2X1 U5651 ( .B(mem[1186]), .A(mem[1227]), .S(n5555), .Y(n5362) );
  MUX2X1 U5652 ( .B(mem[1104]), .A(mem[1145]), .S(n5555), .Y(n5366) );
  MUX2X1 U5653 ( .B(mem[1022]), .A(mem[1063]), .S(n5555), .Y(n5365) );
  MUX2X1 U5654 ( .B(n5364), .A(n5361), .S(n14), .Y(n5375) );
  MUX2X1 U5655 ( .B(mem[940]), .A(mem[981]), .S(n5555), .Y(n5369) );
  MUX2X1 U5656 ( .B(mem[858]), .A(mem[899]), .S(n5555), .Y(n5368) );
  MUX2X1 U5657 ( .B(mem[776]), .A(mem[817]), .S(n5555), .Y(n5372) );
  MUX2X1 U5658 ( .B(mem[694]), .A(mem[735]), .S(n5555), .Y(n5371) );
  MUX2X1 U5659 ( .B(n5370), .A(n5367), .S(n14), .Y(n5374) );
  MUX2X1 U5660 ( .B(mem[612]), .A(mem[653]), .S(n5555), .Y(n5378) );
  MUX2X1 U5661 ( .B(mem[530]), .A(mem[571]), .S(n5555), .Y(n5377) );
  MUX2X1 U5662 ( .B(mem[448]), .A(mem[489]), .S(n5555), .Y(n5381) );
  MUX2X1 U5663 ( .B(mem[366]), .A(mem[407]), .S(n5555), .Y(n5380) );
  MUX2X1 U5664 ( .B(n5379), .A(n5376), .S(n14), .Y(n5390) );
  MUX2X1 U5665 ( .B(mem[284]), .A(mem[325]), .S(n5556), .Y(n5384) );
  MUX2X1 U5666 ( .B(mem[202]), .A(mem[243]), .S(n5556), .Y(n5383) );
  MUX2X1 U5667 ( .B(mem[120]), .A(mem[161]), .S(n5556), .Y(n5387) );
  MUX2X1 U5668 ( .B(mem[38]), .A(mem[79]), .S(n5556), .Y(n5386) );
  MUX2X1 U5669 ( .B(n5385), .A(n5382), .S(n14), .Y(n5389) );
  MUX2X1 U5670 ( .B(n5388), .A(n5373), .S(n16), .Y(n5489) );
  MUX2X1 U5671 ( .B(mem[1269]), .A(mem[1310]), .S(n5556), .Y(n5393) );
  MUX2X1 U5672 ( .B(mem[1187]), .A(mem[1228]), .S(n5556), .Y(n5392) );
  MUX2X1 U5673 ( .B(mem[1105]), .A(mem[1146]), .S(n5556), .Y(n5396) );
  MUX2X1 U5674 ( .B(mem[1023]), .A(mem[1064]), .S(n5556), .Y(n5395) );
  MUX2X1 U5675 ( .B(n5394), .A(n5391), .S(n14), .Y(n5405) );
  MUX2X1 U5676 ( .B(mem[941]), .A(mem[982]), .S(n5556), .Y(n5399) );
  MUX2X1 U5677 ( .B(mem[859]), .A(mem[900]), .S(n5556), .Y(n5398) );
  MUX2X1 U5678 ( .B(mem[777]), .A(mem[818]), .S(n5556), .Y(n5402) );
  MUX2X1 U5679 ( .B(mem[695]), .A(mem[736]), .S(n5556), .Y(n5401) );
  MUX2X1 U5680 ( .B(n5400), .A(n5397), .S(n14), .Y(n5404) );
  MUX2X1 U5681 ( .B(mem[613]), .A(mem[654]), .S(n5557), .Y(n5408) );
  MUX2X1 U5682 ( .B(mem[531]), .A(mem[572]), .S(n5557), .Y(n5407) );
  MUX2X1 U5683 ( .B(mem[449]), .A(mem[490]), .S(n5557), .Y(n5411) );
  MUX2X1 U5684 ( .B(mem[367]), .A(mem[408]), .S(n5557), .Y(n5410) );
  MUX2X1 U5685 ( .B(n5409), .A(n5406), .S(n14), .Y(n5420) );
  MUX2X1 U5686 ( .B(mem[285]), .A(mem[326]), .S(n5557), .Y(n5414) );
  MUX2X1 U5687 ( .B(mem[203]), .A(mem[244]), .S(n5557), .Y(n5413) );
  MUX2X1 U5688 ( .B(mem[121]), .A(mem[162]), .S(n5557), .Y(n5417) );
  MUX2X1 U5689 ( .B(mem[39]), .A(mem[80]), .S(n5557), .Y(n5416) );
  MUX2X1 U5690 ( .B(n5415), .A(n5412), .S(n14), .Y(n5419) );
  MUX2X1 U5691 ( .B(n5418), .A(n5403), .S(n16), .Y(n5490) );
  MUX2X1 U5692 ( .B(mem[1270]), .A(mem[1311]), .S(n5557), .Y(n5423) );
  MUX2X1 U5693 ( .B(mem[1188]), .A(mem[1229]), .S(n5557), .Y(n5422) );
  MUX2X1 U5694 ( .B(mem[1106]), .A(mem[1147]), .S(n5557), .Y(n5426) );
  MUX2X1 U5695 ( .B(mem[1024]), .A(mem[1065]), .S(n5557), .Y(n5425) );
  MUX2X1 U5696 ( .B(n5424), .A(n5421), .S(n14), .Y(n5435) );
  MUX2X1 U5697 ( .B(mem[942]), .A(mem[983]), .S(n5558), .Y(n5429) );
  MUX2X1 U5698 ( .B(mem[860]), .A(mem[901]), .S(n5558), .Y(n5428) );
  MUX2X1 U5699 ( .B(mem[778]), .A(mem[819]), .S(n5558), .Y(n5432) );
  MUX2X1 U5700 ( .B(mem[696]), .A(mem[737]), .S(n5558), .Y(n5431) );
  MUX2X1 U5701 ( .B(n5430), .A(n5427), .S(n14), .Y(n5434) );
  MUX2X1 U5702 ( .B(mem[614]), .A(mem[655]), .S(n5558), .Y(n5438) );
  MUX2X1 U5703 ( .B(mem[532]), .A(mem[573]), .S(n5558), .Y(n5437) );
  MUX2X1 U5704 ( .B(mem[450]), .A(mem[491]), .S(n5558), .Y(n5441) );
  MUX2X1 U5705 ( .B(mem[368]), .A(mem[409]), .S(n5558), .Y(n5440) );
  MUX2X1 U5706 ( .B(n5439), .A(n5436), .S(n14), .Y(n5450) );
  MUX2X1 U5707 ( .B(mem[286]), .A(mem[327]), .S(n5558), .Y(n5444) );
  MUX2X1 U5708 ( .B(mem[204]), .A(mem[245]), .S(n5558), .Y(n5443) );
  MUX2X1 U5709 ( .B(mem[122]), .A(mem[163]), .S(n5558), .Y(n5447) );
  MUX2X1 U5710 ( .B(mem[40]), .A(mem[81]), .S(n5558), .Y(n5446) );
  MUX2X1 U5711 ( .B(n5445), .A(n5442), .S(n14), .Y(n5449) );
  MUX2X1 U5712 ( .B(n5448), .A(n5433), .S(n16), .Y(n5491) );
  OR2X1 U5713 ( .A(n5674), .B(wr_ptr[0]), .Y(sub_93_carry[1]) );
  XNOR2X1 U5714 ( .A(wr_ptr[0]), .B(n5674), .Y(fillcount[0]) );
  XOR2X1 U5715 ( .A(add_51_carry[4]), .B(wr_ptr[4]), .Y(n23) );
  XOR2X1 U5716 ( .A(add_57_carry[4]), .B(n16), .Y(n101) );
endmodule


module ddr3_init_engine_DW01_inc_0 ( A, SUM );
  input [18:0] A;
  output [18:0] SUM;

  wire   [18:2] carry;

  HAX1 U1_1_17 ( .A(A[17]), .B(carry[17]), .YC(carry[18]), .YS(SUM[17]) );
  HAX1 U1_1_16 ( .A(A[16]), .B(carry[16]), .YC(carry[17]), .YS(SUM[16]) );
  HAX1 U1_1_15 ( .A(A[15]), .B(carry[15]), .YC(carry[16]), .YS(SUM[15]) );
  HAX1 U1_1_14 ( .A(A[14]), .B(carry[14]), .YC(carry[15]), .YS(SUM[14]) );
  HAX1 U1_1_13 ( .A(A[13]), .B(carry[13]), .YC(carry[14]), .YS(SUM[13]) );
  HAX1 U1_1_12 ( .A(A[12]), .B(carry[12]), .YC(carry[13]), .YS(SUM[12]) );
  HAX1 U1_1_11 ( .A(A[11]), .B(carry[11]), .YC(carry[12]), .YS(SUM[11]) );
  HAX1 U1_1_10 ( .A(A[10]), .B(carry[10]), .YC(carry[11]), .YS(SUM[10]) );
  HAX1 U1_1_9 ( .A(A[9]), .B(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  HAX1 U1_1_8 ( .A(A[8]), .B(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  HAX1 U1_1_7 ( .A(A[7]), .B(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  HAX1 U1_1_6 ( .A(A[6]), .B(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  HAX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry[2]), .YS(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[18]), .B(A[18]), .Y(SUM[18]) );
endmodule


module ddr3_init_engine ( ready, csbar, rasbar, casbar, webar, ba, a, odt, 
        ts_con, cke, clk, resetbar, init, ck, Port15 );
  output [2:0] ba;
  output [13:0] a;
  input clk, resetbar, init, ck;
  output ready, csbar, rasbar, casbar, webar, odt, ts_con, cke;
  inout Port15;
  wire   flag, RESET, INIT, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n244, n252, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n245;
  wire   [18:0] counter;
  assign csbar = 1'b0;
  assign ba[2] = 1'b0;
  assign a[13] = 1'b0;
  assign a[12] = 1'b0;
  assign a[11] = 1'b0;
  assign a[9] = 1'b0;
  assign a[7] = 1'b0;
  assign a[6] = 1'b0;
  assign a[5] = 1'b0;
  assign a[3] = 1'b0;
  assign a[2] = 1'b0;
  assign a[1] = 1'b0;
  assign a[0] = 1'b0;
  assign odt = 1'b0;
  assign ts_con = 1'b0;

  DFFPOSX1 RESET_reg ( .D(resetbar), .CLK(clk), .Q(RESET) );
  DFFPOSX1 INIT_reg ( .D(init), .CLK(clk), .Q(INIT) );
  DFFPOSX1 flag_reg ( .D(n173), .CLK(clk), .Q(flag) );
  DFFPOSX1 counter_reg_0_ ( .D(n172), .CLK(clk), .Q(counter[0]) );
  DFFPOSX1 counter_reg_1_ ( .D(n171), .CLK(clk), .Q(counter[1]) );
  DFFPOSX1 counter_reg_2_ ( .D(n170), .CLK(clk), .Q(counter[2]) );
  DFFPOSX1 counter_reg_3_ ( .D(n169), .CLK(clk), .Q(counter[3]) );
  DFFPOSX1 counter_reg_4_ ( .D(n168), .CLK(clk), .Q(counter[4]) );
  DFFPOSX1 counter_reg_5_ ( .D(n167), .CLK(clk), .Q(counter[5]) );
  DFFPOSX1 counter_reg_6_ ( .D(n166), .CLK(clk), .Q(counter[6]) );
  DFFPOSX1 counter_reg_7_ ( .D(n165), .CLK(clk), .Q(counter[7]) );
  DFFPOSX1 counter_reg_8_ ( .D(n164), .CLK(clk), .Q(counter[8]) );
  DFFPOSX1 counter_reg_9_ ( .D(n163), .CLK(clk), .Q(counter[9]) );
  DFFPOSX1 counter_reg_10_ ( .D(n162), .CLK(clk), .Q(counter[10]) );
  DFFPOSX1 counter_reg_11_ ( .D(n161), .CLK(clk), .Q(counter[11]) );
  DFFPOSX1 counter_reg_12_ ( .D(n160), .CLK(clk), .Q(counter[12]) );
  DFFPOSX1 counter_reg_13_ ( .D(n159), .CLK(clk), .Q(counter[13]) );
  DFFPOSX1 counter_reg_14_ ( .D(n158), .CLK(clk), .Q(counter[14]) );
  DFFPOSX1 counter_reg_15_ ( .D(n157), .CLK(clk), .Q(counter[15]) );
  DFFPOSX1 counter_reg_16_ ( .D(n156), .CLK(clk), .Q(counter[16]) );
  DFFPOSX1 counter_reg_17_ ( .D(n155), .CLK(clk), .Q(counter[17]) );
  DFFPOSX1 counter_reg_18_ ( .D(n154), .CLK(clk), .Q(counter[18]) );
  DFFPOSX1 ready_reg ( .D(n153), .CLK(clk), .Q(ready) );
  DFFPOSX1 casbar_reg ( .D(n150), .CLK(clk), .Q(casbar) );
  DFFPOSX1 webar_reg ( .D(n4), .CLK(clk), .Q(webar) );
  DFFPOSX1 rasbar_reg ( .D(n5), .CLK(clk), .Q(rasbar) );
  DFFPOSX1 cke_reg ( .D(n149), .CLK(clk), .Q(cke) );
  DFFPOSX1 a_reg_10_ ( .D(n148), .CLK(clk), .Q(a[10]) );
  DFFPOSX1 a_reg_8_ ( .D(n6), .CLK(clk), .Q(a[8]) );
  DFFPOSX1 a_reg_4_ ( .D(n3), .CLK(clk), .Q(a[4]) );
  DFFPOSX1 ba_reg_1_ ( .D(n145), .CLK(clk), .Q(ba[1]) );
  DFFPOSX1 ba_reg_0_ ( .D(n7), .CLK(clk), .Q(ba[0]) );
  NAND3X1 U59 ( .A(n55), .B(n218), .C(n57), .Y(n54) );
  OAI21X1 U61 ( .A(n213), .B(n58), .C(n181), .Y(n145) );
  OAI21X1 U63 ( .A(n208), .B(n61), .C(n218), .Y(n58) );
  NAND3X1 U64 ( .A(n36), .B(n43), .C(n40), .Y(n146) );
  NAND3X1 U66 ( .A(n57), .B(n219), .C(n66), .Y(n62) );
  NAND3X1 U69 ( .A(n57), .B(n219), .C(n68), .Y(n63) );
  OAI21X1 U70 ( .A(n213), .B(n69), .C(n202), .Y(n148) );
  OAI21X1 U72 ( .A(n222), .B(n68), .C(n217), .Y(n69) );
  AOI21X1 U73 ( .A(n72), .B(n222), .C(n219), .Y(n71) );
  OAI21X1 U74 ( .A(n73), .B(n213), .C(n175), .Y(n149) );
  NAND3X1 U76 ( .A(n72), .B(n224), .C(n225), .Y(n75) );
  OAI21X1 U77 ( .A(n46), .B(n45), .C(n9), .Y(n150) );
  NAND3X1 U80 ( .A(n207), .B(n77), .C(n57), .Y(n81) );
  NAND3X1 U83 ( .A(n207), .B(n44), .C(n57), .Y(n83) );
  OAI21X1 U85 ( .A(n188), .B(n213), .C(n187), .Y(n153) );
  AOI21X1 U87 ( .A(n72), .B(n223), .C(n216), .Y(n85) );
  OAI21X1 U88 ( .A(n173), .B(n245), .C(n210), .Y(n154) );
  OAI21X1 U90 ( .A(n173), .B(n243), .C(n201), .Y(n155) );
  OAI21X1 U92 ( .A(n173), .B(n242), .C(n196), .Y(n156) );
  OAI21X1 U94 ( .A(n173), .B(n241), .C(n190), .Y(n157) );
  OAI21X1 U96 ( .A(n173), .B(n240), .C(n185), .Y(n158) );
  OAI21X1 U98 ( .A(n173), .B(n239), .C(n180), .Y(n159) );
  OAI21X1 U100 ( .A(n173), .B(n238), .C(n174), .Y(n160) );
  OAI21X1 U102 ( .A(n173), .B(n237), .C(n51), .Y(n161) );
  OAI21X1 U104 ( .A(n173), .B(n236), .C(n50), .Y(n162) );
  OAI21X1 U106 ( .A(n173), .B(n235), .C(n209), .Y(n163) );
  OAI21X1 U108 ( .A(n173), .B(n234), .C(n200), .Y(n164) );
  OAI21X1 U110 ( .A(n173), .B(n232), .C(n195), .Y(n165) );
  OAI21X1 U112 ( .A(n173), .B(n231), .C(n189), .Y(n166) );
  OAI21X1 U114 ( .A(n173), .B(n230), .C(n184), .Y(n167) );
  OAI21X1 U116 ( .A(n173), .B(n229), .C(n49), .Y(n168) );
  OAI21X1 U118 ( .A(n173), .B(n227), .C(n48), .Y(n169) );
  OAI21X1 U120 ( .A(n173), .B(n226), .C(n47), .Y(n170) );
  OAI21X1 U122 ( .A(n173), .B(n224), .C(n179), .Y(n171) );
  OAI21X1 U124 ( .A(n173), .B(n221), .C(n52), .Y(n172) );
  OAI21X1 U126 ( .A(n216), .B(n204), .C(n213), .Y(n173) );
  NAND3X1 U130 ( .A(n42), .B(n46), .C(n39), .Y(n108) );
  NAND3X1 U133 ( .A(n111), .B(n112), .C(n38), .Y(n110) );
  NOR3X1 U136 ( .A(n116), .B(n223), .C(n117), .Y(n115) );
  NOR3X1 U137 ( .A(n182), .B(n186), .C(n206), .Y(n117) );
  AOI22X1 U138 ( .A(n121), .B(n122), .C(counter[3]), .D(n233), .Y(n119) );
  NOR3X1 U139 ( .A(counter[11]), .B(counter[8]), .C(counter[3]), .Y(n122) );
  NOR3X1 U140 ( .A(n235), .B(counter[10]), .C(n232), .Y(n121) );
  NAND3X1 U142 ( .A(counter[11]), .B(n124), .C(n178), .Y(n123) );
  NOR3X1 U144 ( .A(n211), .B(n226), .C(n198), .Y(n116) );
  AOI22X1 U146 ( .A(counter[1]), .B(n37), .C(n124), .D(n111), .Y(n114) );
  NOR3X1 U147 ( .A(n226), .B(n234), .C(n206), .Y(n124) );
  NAND3X1 U148 ( .A(n224), .B(n229), .C(counter[6]), .Y(n120) );
  NAND3X1 U149 ( .A(n197), .B(n192), .C(n131), .Y(n129) );
  NAND3X1 U150 ( .A(n111), .B(counter[4]), .C(n133), .Y(n76) );
  NOR3X1 U151 ( .A(n226), .B(counter[8]), .C(counter[6]), .Y(n133) );
  NOR3X1 U152 ( .A(n236), .B(counter[11]), .C(n205), .Y(n111) );
  NAND3X1 U153 ( .A(counter[7]), .B(counter[5]), .C(n134), .Y(n126) );
  AOI21X1 U155 ( .A(n72), .B(n208), .C(n219), .Y(n56) );
  NAND3X1 U157 ( .A(n228), .B(n226), .C(counter[4]), .Y(n130) );
  AOI21X1 U158 ( .A(n72), .B(n68), .C(n194), .Y(n65) );
  OAI21X1 U160 ( .A(n66), .B(n61), .C(n72), .Y(n135) );
  NOR3X1 U161 ( .A(counter[2]), .B(counter[4]), .C(n224), .Y(n112) );
  NAND3X1 U162 ( .A(counter[5]), .B(counter[3]), .C(n136), .Y(n128) );
  NOR3X1 U163 ( .A(n212), .B(counter[4]), .C(n224), .Y(n66) );
  NOR3X1 U164 ( .A(n212), .B(counter[1]), .C(n229), .Y(n68) );
  NAND3X1 U165 ( .A(counter[6]), .B(counter[2]), .C(n138), .Y(n132) );
  NOR3X1 U166 ( .A(n191), .B(counter[5]), .C(counter[3]), .Y(n138) );
  NAND3X1 U167 ( .A(counter[8]), .B(counter[10]), .C(n139), .Y(n137) );
  NOR3X1 U168 ( .A(counter[11]), .B(counter[9]), .C(counter[7]), .Y(n139) );
  NOR3X1 U169 ( .A(n41), .B(counter[12]), .C(counter[0]), .Y(n141) );
  NAND3X1 U170 ( .A(n242), .B(n243), .C(n239), .Y(n142) );
  NOR3X1 U171 ( .A(n203), .B(n245), .C(n213), .Y(n140) );
  ddr3_init_engine_DW01_inc_0 add_80 ( .A(counter), .SUM({n28, n27, n26, n25, 
        n24, n23, n22, n21, n20, n19, n18, n17, n16, n15, n14, n13, n12, n11, 
        n10}) );
  OR2X1 U18 ( .A(n229), .B(n212), .Y(n131) );
  AND2X1 U19 ( .A(n2), .B(n115), .Y(n84) );
  AND2X1 U20 ( .A(n173), .B(n204), .Y(n88) );
  OR2X1 U21 ( .A(n192), .B(counter[1]), .Y(n60) );
  AND2X1 U22 ( .A(n72), .B(n8), .Y(n78) );
  AND2X1 U23 ( .A(a[10]), .B(n183), .Y(n70) );
  AND2X1 U24 ( .A(n176), .B(RESET), .Y(n73) );
  AND2X1 U25 ( .A(ready), .B(n188), .Y(n86) );
  AND2X1 U26 ( .A(n45), .B(RESET), .Y(n252) );
  OR2X1 U27 ( .A(n44), .B(n222), .Y(n77) );
  BUFX2 U28 ( .A(n110), .Y(n1) );
  BUFX2 U29 ( .A(n114), .Y(n2) );
  BUFX2 U30 ( .A(n146), .Y(n3) );
  AND2X1 U31 ( .A(n33), .B(n29), .Y(n152) );
  INVX1 U32 ( .A(n152), .Y(n4) );
  AND2X1 U33 ( .A(n34), .B(n30), .Y(n151) );
  INVX1 U34 ( .A(n151), .Y(n5) );
  AND2X1 U35 ( .A(n43), .B(n32), .Y(n147) );
  INVX1 U36 ( .A(n147), .Y(n6) );
  AND2X1 U37 ( .A(n35), .B(n31), .Y(n144) );
  INVX1 U38 ( .A(n144), .Y(n7) );
  BUFX2 U39 ( .A(n108), .Y(n8) );
  AND2X1 U40 ( .A(casbar), .B(n45), .Y(n79) );
  INVX1 U41 ( .A(n79), .Y(n9) );
  BUFX2 U42 ( .A(n83), .Y(n29) );
  BUFX2 U43 ( .A(n81), .Y(n30) );
  BUFX2 U44 ( .A(n54), .Y(n31) );
  AND2X1 U45 ( .A(a[8]), .B(n193), .Y(n67) );
  INVX1 U46 ( .A(n67), .Y(n32) );
  AND2X1 U47 ( .A(webar), .B(n252), .Y(n82) );
  INVX1 U48 ( .A(n82), .Y(n33) );
  AND2X1 U49 ( .A(rasbar), .B(n252), .Y(n80) );
  INVX1 U50 ( .A(n80), .Y(n34) );
  AND2X1 U51 ( .A(ba[0]), .B(n199), .Y(n53) );
  INVX1 U52 ( .A(n53), .Y(n35) );
  BUFX2 U53 ( .A(n62), .Y(n36) );
  BUFX2 U54 ( .A(n129), .Y(n37) );
  OR2X1 U55 ( .A(n231), .B(n234), .Y(n113) );
  INVX1 U56 ( .A(n113), .Y(n38) );
  OR2X1 U57 ( .A(n61), .B(n68), .Y(n109) );
  INVX1 U58 ( .A(n109), .Y(n39) );
  AND2X1 U60 ( .A(a[4]), .B(n193), .Y(n64) );
  INVX1 U62 ( .A(n64), .Y(n40) );
  BUFX2 U65 ( .A(n142), .Y(n41) );
  OR2X1 U67 ( .A(n66), .B(n208), .Y(n55) );
  INVX1 U68 ( .A(n55), .Y(n42) );
  BUFX2 U71 ( .A(n63), .Y(n43) );
  INVX1 U75 ( .A(n84), .Y(n44) );
  INVX1 U78 ( .A(n78), .Y(n45) );
  INVX1 U79 ( .A(n77), .Y(n46) );
  AND2X1 U81 ( .A(n12), .B(n214), .Y(n104) );
  INVX1 U82 ( .A(n104), .Y(n47) );
  AND2X1 U84 ( .A(n13), .B(n214), .Y(n103) );
  INVX1 U86 ( .A(n103), .Y(n48) );
  AND2X1 U89 ( .A(n14), .B(n214), .Y(n102) );
  INVX1 U91 ( .A(n102), .Y(n49) );
  AND2X1 U93 ( .A(n20), .B(n215), .Y(n96) );
  INVX1 U95 ( .A(n96), .Y(n50) );
  AND2X1 U97 ( .A(n21), .B(n215), .Y(n95) );
  INVX1 U99 ( .A(n95), .Y(n51) );
  AND2X1 U101 ( .A(n10), .B(n214), .Y(n106) );
  INVX1 U103 ( .A(n106), .Y(n52) );
  AND2X1 U105 ( .A(n22), .B(n215), .Y(n94) );
  INVX1 U107 ( .A(n94), .Y(n174) );
  AND2X1 U109 ( .A(cke), .B(n73), .Y(n74) );
  INVX1 U111 ( .A(n74), .Y(n175) );
  BUFX2 U113 ( .A(n75), .Y(n176) );
  BUFX2 U115 ( .A(n123), .Y(n177) );
  OR2X1 U117 ( .A(counter[10]), .B(n205), .Y(n125) );
  INVX1 U119 ( .A(n125), .Y(n178) );
  AND2X1 U121 ( .A(n11), .B(n214), .Y(n105) );
  INVX1 U123 ( .A(n105), .Y(n179) );
  AND2X1 U125 ( .A(n23), .B(n215), .Y(n93) );
  INVX1 U127 ( .A(n93), .Y(n180) );
  AND2X1 U128 ( .A(ba[1]), .B(n199), .Y(n59) );
  INVX1 U129 ( .A(n59), .Y(n181) );
  AND2X1 U131 ( .A(n226), .B(n230), .Y(n118) );
  INVX1 U132 ( .A(n118), .Y(n182) );
  BUFX2 U134 ( .A(n71), .Y(n183) );
  AND2X1 U135 ( .A(n15), .B(n214), .Y(n101) );
  INVX1 U141 ( .A(n101), .Y(n184) );
  AND2X1 U143 ( .A(n24), .B(n215), .Y(n92) );
  INVX1 U145 ( .A(n92), .Y(n185) );
  BUFX2 U154 ( .A(n119), .Y(n186) );
  INVX1 U156 ( .A(n86), .Y(n187) );
  BUFX2 U159 ( .A(n85), .Y(n188) );
  AND2X1 U172 ( .A(n16), .B(n214), .Y(n100) );
  INVX1 U173 ( .A(n100), .Y(n189) );
  AND2X1 U174 ( .A(n25), .B(n215), .Y(n91) );
  INVX1 U175 ( .A(n91), .Y(n190) );
  BUFX2 U176 ( .A(n137), .Y(n191) );
  BUFX2 U177 ( .A(n130), .Y(n192) );
  BUFX2 U178 ( .A(n65), .Y(n193) );
  AND2X1 U179 ( .A(n135), .B(RESET), .Y(n244) );
  INVX1 U180 ( .A(n244), .Y(n194) );
  AND2X1 U181 ( .A(n17), .B(n214), .Y(n99) );
  INVX1 U182 ( .A(n99), .Y(n195) );
  AND2X1 U183 ( .A(n26), .B(n215), .Y(n90) );
  INVX1 U184 ( .A(n90), .Y(n196) );
  BUFX2 U185 ( .A(n76), .Y(n197) );
  BUFX2 U186 ( .A(n128), .Y(n198) );
  BUFX2 U187 ( .A(n56), .Y(n199) );
  AND2X1 U188 ( .A(n18), .B(n214), .Y(n98) );
  INVX1 U189 ( .A(n98), .Y(n200) );
  AND2X1 U190 ( .A(n27), .B(n215), .Y(n89) );
  INVX1 U191 ( .A(n89), .Y(n201) );
  INVX1 U192 ( .A(n70), .Y(n202) );
  AND2X1 U193 ( .A(counter[15]), .B(counter[14]), .Y(n143) );
  INVX1 U194 ( .A(n143), .Y(n203) );
  AND2X1 U195 ( .A(INIT), .B(n220), .Y(n107) );
  INVX1 U196 ( .A(n107), .Y(n204) );
  BUFX2 U197 ( .A(n126), .Y(n205) );
  BUFX2 U198 ( .A(n120), .Y(n206) );
  INVX1 U199 ( .A(n252), .Y(n207) );
  INVX1 U200 ( .A(n60), .Y(n208) );
  AND2X1 U201 ( .A(n19), .B(n214), .Y(n97) );
  INVX1 U202 ( .A(n97), .Y(n209) );
  AND2X1 U203 ( .A(n28), .B(n215), .Y(n87) );
  INVX1 U204 ( .A(n87), .Y(n210) );
  AND2X1 U205 ( .A(n224), .B(n229), .Y(n127) );
  INVX1 U206 ( .A(n127), .Y(n211) );
  BUFX2 U207 ( .A(n132), .Y(n212) );
  AND2X1 U208 ( .A(flag), .B(RESET), .Y(n57) );
  INVX1 U209 ( .A(n57), .Y(n213) );
  BUFX2 U210 ( .A(n88), .Y(n214) );
  BUFX2 U211 ( .A(n88), .Y(n215) );
  INVX1 U212 ( .A(n199), .Y(n218) );
  INVX1 U213 ( .A(n193), .Y(n219) );
  AND2X1 U214 ( .A(n228), .B(n112), .Y(n61) );
  INVX1 U215 ( .A(n191), .Y(n233) );
  INVX1 U216 ( .A(n198), .Y(n228) );
  INVX1 U217 ( .A(n1), .Y(n222) );
  INVX1 U218 ( .A(n197), .Y(n225) );
  AND2X1 U219 ( .A(n231), .B(n233), .Y(n136) );
  AND2X1 U220 ( .A(n235), .B(n227), .Y(n134) );
  INVX1 U221 ( .A(flag), .Y(n220) );
  AND2X1 U222 ( .A(n140), .B(n141), .Y(n72) );
  INVX1 U223 ( .A(counter[1]), .Y(n224) );
  INVX1 U224 ( .A(counter[14]), .Y(n240) );
  INVX1 U225 ( .A(counter[15]), .Y(n241) );
  INVX1 U226 ( .A(counter[12]), .Y(n238) );
  INVX1 U227 ( .A(counter[11]), .Y(n237) );
  INVX1 U228 ( .A(counter[0]), .Y(n221) );
  INVX1 U229 ( .A(counter[2]), .Y(n226) );
  INVX1 U230 ( .A(n183), .Y(n217) );
  INVX1 U231 ( .A(counter[4]), .Y(n229) );
  INVX1 U232 ( .A(counter[8]), .Y(n234) );
  INVX1 U233 ( .A(counter[3]), .Y(n227) );
  INVX1 U234 ( .A(counter[6]), .Y(n231) );
  INVX1 U235 ( .A(counter[10]), .Y(n236) );
  INVX1 U236 ( .A(counter[5]), .Y(n230) );
  INVX1 U237 ( .A(n177), .Y(n223) );
  INVX1 U238 ( .A(counter[7]), .Y(n232) );
  INVX1 U239 ( .A(counter[9]), .Y(n235) );
  INVX1 U240 ( .A(RESET), .Y(n216) );
  INVX1 U241 ( .A(counter[18]), .Y(n245) );
  INVX1 U242 ( .A(counter[13]), .Y(n239) );
  INVX1 U243 ( .A(counter[17]), .Y(n243) );
  INVX1 U244 ( .A(counter[16]), .Y(n242) );
endmodule


module SSTL18DDR3DIFF ( PAD, PADN, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD,  PADN;
  wire   n1, n2, n3, n5;

  TBUFX2 b2 ( .A(A), .EN(TS), .Y(PADN) );
  TBUFX2 b1 ( .A(n5), .EN(TS), .Y(PAD) );
  NAND3X1 U2 ( .A(PAD), .B(n2), .C(RI), .Y(n1) );
  BUFX2 U1 ( .A(n1), .Y(n3) );
  INVX1 U3 ( .A(n3), .Y(Z) );
  INVX1 U4 ( .A(A), .Y(n5) );
  INVX1 U5 ( .A(PADN), .Y(n2) );
endmodule


module SSTL18DDR3_45 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_44 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_43 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_42 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_41 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_40 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_39 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_38 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_37 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_36 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_35 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_34 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_33 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_32 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_31 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_30 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_29 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_28 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_27 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_26 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_25 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_24 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_23 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_22 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_21 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_20 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_19 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_18 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_17 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_16 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_15 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_14 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_13 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_12 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_11 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_10 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_9 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_8 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_7 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_6 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_5 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_4 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_3 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_2 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_1 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_0 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3INTERFACE ( ck_pad, ckbar_pad, cke_pad, csbar_pad, rasbar_pad, 
        casbar_pad, webar_pad, ba_pad, a_pad, dm_pad, odt_pad, resetbar_pad, 
        dq_o, dqs_o, dqsbar_o, dq_pad, dqs_pad, dqsbar_pad, ri_i, ts_i, ck_i, 
        cke_i, csbar_i, rasbar_i, casbar_i, webar_i, ba_i, a_i, dq_i, dqs_i, 
        dqsbar_i, dm_i, odt_i, resetbar_i );
  output [2:0] ba_pad;
  output [13:0] a_pad;
  output [1:0] dm_pad;
  output [15:0] dq_o;
  output [1:0] dqs_o;
  output [1:0] dqsbar_o;
  inout [15:0] dq_pad;
  inout [1:0] dqs_pad;
  inout [1:0] dqsbar_pad;
  input [2:0] ba_i;
  input [13:0] a_i;
  input [15:0] dq_i;
  input [1:0] dqs_i;
  input [1:0] dqsbar_i;
  input [1:0] dm_i;
  input ri_i, ts_i, ck_i, cke_i, csbar_i, rasbar_i, casbar_i, webar_i, odt_i,
         resetbar_i;
  output ck_pad, ckbar_pad, cke_pad, csbar_pad, rasbar_pad, casbar_pad,
         webar_pad, odt_pad, resetbar_pad;


  SSTL18DDR3DIFF ck_sstl ( .PAD(ck_pad), .PADN(ckbar_pad), .Z(), .A(ck_i), 
        .RI(1'b0), .TS(1'b1) );
  SSTL18DDR3_45 cke_sstl ( .PAD(cke_pad), .Z(), .A(cke_i), .RI(1'b0), .TS(1'b1) );
  SSTL18DDR3_44 casbar_sstl ( .PAD(casbar_pad), .Z(), .A(casbar_i), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_43 rasbar_sstl ( .PAD(rasbar_pad), .Z(), .A(rasbar_i), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_42 csbar_sstl ( .PAD(csbar_pad), .Z(), .A(csbar_i), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_41 webar_sstl ( .PAD(webar_pad), .Z(), .A(webar_i), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_40 odt_sstl ( .PAD(odt_pad), .Z(), .A(odt_i), .RI(1'b0), .TS(1'b1) );
  SSTL18DDR3_39 resetbar_sstl ( .PAD(resetbar_pad), .Z(), .A(resetbar_i), .RI(
        1'b0), .TS(1'b1) );
  SSTL18DDR3_38 BA_0__sstl_ba ( .PAD(ba_pad[0]), .Z(), .A(ba_i[0]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_37 BA_1__sstl_ba ( .PAD(ba_pad[1]), .Z(), .A(ba_i[1]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_36 BA_2__sstl_ba ( .PAD(ba_pad[2]), .Z(), .A(ba_i[2]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_35 A_0__sstl_a ( .PAD(a_pad[0]), .Z(), .A(a_i[0]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_34 A_1__sstl_a ( .PAD(a_pad[1]), .Z(), .A(a_i[1]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_33 A_2__sstl_a ( .PAD(a_pad[2]), .Z(), .A(a_i[2]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_32 A_3__sstl_a ( .PAD(a_pad[3]), .Z(), .A(a_i[3]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_31 A_4__sstl_a ( .PAD(a_pad[4]), .Z(), .A(a_i[4]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_30 A_5__sstl_a ( .PAD(a_pad[5]), .Z(), .A(a_i[5]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_29 A_6__sstl_a ( .PAD(a_pad[6]), .Z(), .A(a_i[6]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_28 A_7__sstl_a ( .PAD(a_pad[7]), .Z(), .A(a_i[7]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_27 A_8__sstl_a ( .PAD(a_pad[8]), .Z(), .A(a_i[8]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_26 A_9__sstl_a ( .PAD(a_pad[9]), .Z(), .A(a_i[9]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_25 A_10__sstl_a ( .PAD(a_pad[10]), .Z(), .A(a_i[10]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_24 A_11__sstl_a ( .PAD(a_pad[11]), .Z(), .A(a_i[11]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_23 A_12__sstl_a ( .PAD(a_pad[12]), .Z(), .A(a_i[12]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_22 A_13__sstl_a ( .PAD(a_pad[13]), .Z(), .A(a_i[13]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_21 DQ_0__sstl_dq ( .PAD(dq_pad[0]), .Z(dq_o[0]), .A(dq_i[0]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_20 DQ_1__sstl_dq ( .PAD(dq_pad[1]), .Z(dq_o[1]), .A(dq_i[1]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_19 DQ_2__sstl_dq ( .PAD(dq_pad[2]), .Z(dq_o[2]), .A(dq_i[2]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_18 DQ_3__sstl_dq ( .PAD(dq_pad[3]), .Z(dq_o[3]), .A(dq_i[3]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_17 DQ_4__sstl_dq ( .PAD(dq_pad[4]), .Z(dq_o[4]), .A(dq_i[4]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_16 DQ_5__sstl_dq ( .PAD(dq_pad[5]), .Z(dq_o[5]), .A(dq_i[5]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_15 DQ_6__sstl_dq ( .PAD(dq_pad[6]), .Z(dq_o[6]), .A(dq_i[6]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_14 DQ_7__sstl_dq ( .PAD(dq_pad[7]), .Z(dq_o[7]), .A(dq_i[7]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_13 DQ_8__sstl_dq ( .PAD(dq_pad[8]), .Z(dq_o[8]), .A(dq_i[8]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_12 DQ_9__sstl_dq ( .PAD(dq_pad[9]), .Z(dq_o[9]), .A(dq_i[9]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_11 DQ_10__sstl_dq ( .PAD(dq_pad[10]), .Z(dq_o[10]), .A(dq_i[10]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_10 DQ_11__sstl_dq ( .PAD(dq_pad[11]), .Z(dq_o[11]), .A(dq_i[11]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_9 DQ_12__sstl_dq ( .PAD(dq_pad[12]), .Z(dq_o[12]), .A(dq_i[12]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_8 DQ_13__sstl_dq ( .PAD(dq_pad[13]), .Z(dq_o[13]), .A(dq_i[13]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_7 DQ_14__sstl_dq ( .PAD(dq_pad[14]), .Z(dq_o[14]), .A(dq_i[14]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_6 DQ_15__sstl_dq ( .PAD(dq_pad[15]), .Z(dq_o[15]), .A(dq_i[15]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_5 DQS_0__sstl_dqs ( .PAD(dqs_pad[0]), .Z(dqs_o[0]), .A(dqs_i[0]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_4 DQS_1__sstl_dqs ( .PAD(dqs_pad[1]), .Z(dqs_o[1]), .A(dqs_i[1]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_3 DQSBAR_0__sstl_dqsbar ( .PAD(dqsbar_pad[0]), .Z(dqsbar_o[0]), 
        .A(dqsbar_i[0]), .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_2 DQSBAR_1__sstl_dqsbar ( .PAD(dqsbar_pad[1]), .Z(dqsbar_o[1]), 
        .A(dqsbar_i[1]), .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_1 DM_0__sstl_dm ( .PAD(dm_pad[0]), .Z(), .A(dm_i[0]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_0 DM_1__sstl_dm ( .PAD(dm_pad[1]), .Z(), .A(dm_i[1]), .RI(1'b0), 
        .TS(1'b1) );
endmodule


module ddr3_controller ( dout, raddr, fillcount, notfull, ready, ck_pad, 
        ckbar_pad, cke_pad, csbar_pad, rasbar_pad, casbar_pad, webar_pad, 
        ba_pad, a_pad, dm_pad, odt_pad, notempty, resetbar_pad, dq_pad, 
        dqs_pad, dqsbar_pad, clk, resetbar, read, cmd, din, addr, initddr );
  output [15:0] dout;
  output [24:0] raddr;
  output [5:0] fillcount;
  output [2:0] ba_pad;
  output [13:0] a_pad;
  output [1:0] dm_pad;
  inout [15:0] dq_pad;
  inout [1:0] dqs_pad;
  inout [1:0] dqsbar_pad;
  input [2:0] cmd;
  input [15:0] din;
  input [24:0] addr;
  input clk, resetbar, read, initddr;
  output notfull, ready, ck_pad, ckbar_pad, cke_pad, csbar_pad, rasbar_pad,
         casbar_pad, webar_pad, odt_pad, notempty, resetbar_pad;
  wire   ck_i, n6, init_rasbar, init_casbar, init_webar, init_cke, rasbar_i,
         casbar_i, webar_i, n3, n4, n7, SYNOPSYS_UNCONNECTED_1,
         SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3,
         SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5,
         SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7,
         SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9,
         SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11,
         SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13,
         SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15,
         SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17,
         SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19,
         SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21,
         SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23,
         SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25,
         SYNOPSYS_UNCONNECTED_26, SYNOPSYS_UNCONNECTED_27,
         SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29,
         SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31,
         SYNOPSYS_UNCONNECTED_32, SYNOPSYS_UNCONNECTED_33,
         SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35,
         SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37,
         SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39,
         SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41,
         SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_43,
         SYNOPSYS_UNCONNECTED_44, SYNOPSYS_UNCONNECTED_45,
         SYNOPSYS_UNCONNECTED_46, SYNOPSYS_UNCONNECTED_47,
         SYNOPSYS_UNCONNECTED_48, SYNOPSYS_UNCONNECTED_49,
         SYNOPSYS_UNCONNECTED_50, SYNOPSYS_UNCONNECTED_51,
         SYNOPSYS_UNCONNECTED_52, SYNOPSYS_UNCONNECTED_53,
         SYNOPSYS_UNCONNECTED_54, SYNOPSYS_UNCONNECTED_55,
         SYNOPSYS_UNCONNECTED_56, SYNOPSYS_UNCONNECTED_57,
         SYNOPSYS_UNCONNECTED_58, SYNOPSYS_UNCONNECTED_59,
         SYNOPSYS_UNCONNECTED_60, SYNOPSYS_UNCONNECTED_61,
         SYNOPSYS_UNCONNECTED_62, SYNOPSYS_UNCONNECTED_63,
         SYNOPSYS_UNCONNECTED_64, SYNOPSYS_UNCONNECTED_65,
         SYNOPSYS_UNCONNECTED_66, SYNOPSYS_UNCONNECTED_67,
         SYNOPSYS_UNCONNECTED_68, SYNOPSYS_UNCONNECTED_69,
         SYNOPSYS_UNCONNECTED_70, SYNOPSYS_UNCONNECTED_71,
         SYNOPSYS_UNCONNECTED_72, SYNOPSYS_UNCONNECTED_73,
         SYNOPSYS_UNCONNECTED_74, SYNOPSYS_UNCONNECTED_75,
         SYNOPSYS_UNCONNECTED_76, SYNOPSYS_UNCONNECTED_77,
         SYNOPSYS_UNCONNECTED_78, SYNOPSYS_UNCONNECTED_79,
         SYNOPSYS_UNCONNECTED_80, SYNOPSYS_UNCONNECTED_81,
         SYNOPSYS_UNCONNECTED_82, SYNOPSYS_UNCONNECTED_83,
         SYNOPSYS_UNCONNECTED_84, SYNOPSYS_UNCONNECTED_85,
         SYNOPSYS_UNCONNECTED_86, SYNOPSYS_UNCONNECTED_87,
         SYNOPSYS_UNCONNECTED_88, SYNOPSYS_UNCONNECTED_89,
         SYNOPSYS_UNCONNECTED_90, SYNOPSYS_UNCONNECTED_91,
         SYNOPSYS_UNCONNECTED_92, SYNOPSYS_UNCONNECTED_93,
         SYNOPSYS_UNCONNECTED_94, SYNOPSYS_UNCONNECTED_95,
         SYNOPSYS_UNCONNECTED_96, SYNOPSYS_UNCONNECTED_97,
         SYNOPSYS_UNCONNECTED_98, SYNOPSYS_UNCONNECTED_99,
         SYNOPSYS_UNCONNECTED_100, SYNOPSYS_UNCONNECTED_101,
         SYNOPSYS_UNCONNECTED_102, SYNOPSYS_UNCONNECTED_103,
         SYNOPSYS_UNCONNECTED_104, SYNOPSYS_UNCONNECTED_105,
         SYNOPSYS_UNCONNECTED_106, SYNOPSYS_UNCONNECTED_107,
         SYNOPSYS_UNCONNECTED_108, SYNOPSYS_UNCONNECTED_109,
         SYNOPSYS_UNCONNECTED_110, SYNOPSYS_UNCONNECTED_111,
         SYNOPSYS_UNCONNECTED_112, SYNOPSYS_UNCONNECTED_113,
         SYNOPSYS_UNCONNECTED_114, SYNOPSYS_UNCONNECTED_115,
         SYNOPSYS_UNCONNECTED_116, SYNOPSYS_UNCONNECTED_117,
         SYNOPSYS_UNCONNECTED_118;
  wire   [32:0] CMD_data_in;
  wire   [40:0] RETURN_data_in;
  wire   [1:0] init_ba;
  wire   [10:4] init_a;
  wire   [10:4] a_i;
  wire   [1:0] ba_i;
  wire   [15:0] dq_i;
  wire   [1:0] dqs_i;
  wire   [1:0] dqsbar_i;
  wire   [1:0] dm_i;

  DFFPOSX1 ck_i_reg ( .D(n3), .CLK(clk), .Q(ck_i) );
  FIFO_DEPTH_P25_WIDTH16 FIFO_IN ( .clk(clk), .reset(resetbar), .data_in(din), 
        .put(1'b0), .get(1'b0), .data_out(dout), .empty_bar(notempty), 
        .full_bar(notfull), .fillcount(fillcount) );
  FIFO_DEPTH_P25_WIDTH33 FIFO_CMD ( .clk(clk), .reset(resetbar), .data_in({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .put(1'b0), 
        .get(1'b0), .data_out({SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, 
        SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, 
        SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, 
        SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10, 
        SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12, 
        SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14, 
        SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16, 
        SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18, 
        SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20, 
        SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22, 
        SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24, 
        SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26, 
        SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28, 
        SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30, 
        SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32, 
        SYNOPSYS_UNCONNECTED_33}), .empty_bar(), .full_bar(), .fillcount({
        SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35, 
        SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37, 
        SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39}) );
  FIFO_DEPTH_P25_WIDTH41 FIFO_RETURN ( .clk(clk), .reset(resetbar), .data_in({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .put(1'b0), .get(1'b0), .data_out({
        SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41, 
        SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_43, 
        SYNOPSYS_UNCONNECTED_44, SYNOPSYS_UNCONNECTED_45, 
        SYNOPSYS_UNCONNECTED_46, SYNOPSYS_UNCONNECTED_47, 
        SYNOPSYS_UNCONNECTED_48, SYNOPSYS_UNCONNECTED_49, 
        SYNOPSYS_UNCONNECTED_50, SYNOPSYS_UNCONNECTED_51, 
        SYNOPSYS_UNCONNECTED_52, SYNOPSYS_UNCONNECTED_53, 
        SYNOPSYS_UNCONNECTED_54, SYNOPSYS_UNCONNECTED_55, 
        SYNOPSYS_UNCONNECTED_56, SYNOPSYS_UNCONNECTED_57, 
        SYNOPSYS_UNCONNECTED_58, SYNOPSYS_UNCONNECTED_59, 
        SYNOPSYS_UNCONNECTED_60, SYNOPSYS_UNCONNECTED_61, 
        SYNOPSYS_UNCONNECTED_62, SYNOPSYS_UNCONNECTED_63, 
        SYNOPSYS_UNCONNECTED_64, SYNOPSYS_UNCONNECTED_65, 
        SYNOPSYS_UNCONNECTED_66, SYNOPSYS_UNCONNECTED_67, 
        SYNOPSYS_UNCONNECTED_68, SYNOPSYS_UNCONNECTED_69, 
        SYNOPSYS_UNCONNECTED_70, SYNOPSYS_UNCONNECTED_71, 
        SYNOPSYS_UNCONNECTED_72, SYNOPSYS_UNCONNECTED_73, 
        SYNOPSYS_UNCONNECTED_74, SYNOPSYS_UNCONNECTED_75, 
        SYNOPSYS_UNCONNECTED_76, SYNOPSYS_UNCONNECTED_77, 
        SYNOPSYS_UNCONNECTED_78, SYNOPSYS_UNCONNECTED_79, 
        SYNOPSYS_UNCONNECTED_80}), .empty_bar(), .full_bar(), .fillcount({
        SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82, 
        SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84, 
        SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86}) );
  ddr3_init_engine XINIT ( .ready(ready), .csbar(), .rasbar(init_rasbar), 
        .casbar(init_casbar), .webar(init_webar), .ba({SYNOPSYS_UNCONNECTED_87, 
        init_ba}), .a({SYNOPSYS_UNCONNECTED_88, SYNOPSYS_UNCONNECTED_89, 
        SYNOPSYS_UNCONNECTED_90, init_a[10], SYNOPSYS_UNCONNECTED_91, 
        init_a[8], SYNOPSYS_UNCONNECTED_92, SYNOPSYS_UNCONNECTED_93, 
        SYNOPSYS_UNCONNECTED_94, init_a[4], SYNOPSYS_UNCONNECTED_95, 
        SYNOPSYS_UNCONNECTED_96, SYNOPSYS_UNCONNECTED_97, 
        SYNOPSYS_UNCONNECTED_98}), .odt(), .ts_con(), .cke(init_cke), .clk(clk), .resetbar(resetbar), .init(initddr), .ck(1'b0), .Port15() );
  SSTL18DDR3INTERFACE XSSTL ( .ck_pad(ck_pad), .ckbar_pad(ckbar_pad), 
        .cke_pad(cke_pad), .csbar_pad(csbar_pad), .rasbar_pad(rasbar_pad), 
        .casbar_pad(casbar_pad), .webar_pad(webar_pad), .ba_pad(ba_pad), 
        .a_pad(a_pad), .dm_pad(dm_pad), .odt_pad(odt_pad), .resetbar_pad(
        resetbar_pad), .dq_o({SYNOPSYS_UNCONNECTED_99, 
        SYNOPSYS_UNCONNECTED_100, SYNOPSYS_UNCONNECTED_101, 
        SYNOPSYS_UNCONNECTED_102, SYNOPSYS_UNCONNECTED_103, 
        SYNOPSYS_UNCONNECTED_104, SYNOPSYS_UNCONNECTED_105, 
        SYNOPSYS_UNCONNECTED_106, SYNOPSYS_UNCONNECTED_107, 
        SYNOPSYS_UNCONNECTED_108, SYNOPSYS_UNCONNECTED_109, 
        SYNOPSYS_UNCONNECTED_110, SYNOPSYS_UNCONNECTED_111, 
        SYNOPSYS_UNCONNECTED_112, SYNOPSYS_UNCONNECTED_113, 
        SYNOPSYS_UNCONNECTED_114}), .dqs_o({SYNOPSYS_UNCONNECTED_115, 
        SYNOPSYS_UNCONNECTED_116}), .dqsbar_o({SYNOPSYS_UNCONNECTED_117, 
        SYNOPSYS_UNCONNECTED_118}), .dq_pad(dq_pad), .dqs_pad(dqs_pad), 
        .dqsbar_pad(dqsbar_pad), .ri_i(1'b0), .ts_i(1'b0), .ck_i(ck_i), 
        .cke_i(init_cke), .csbar_i(1'b0), .rasbar_i(rasbar_i), .casbar_i(
        casbar_i), .webar_i(webar_i), .ba_i({1'b0, ba_i}), .a_i({1'b0, 1'b0, 
        1'b0, a_i[10], 1'b0, a_i[8], 1'b0, 1'b0, 1'b0, a_i[4], 1'b0, 1'b0, 
        1'b0, 1'b0}), .dq_i({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .dqs_i({1'b0, 1'b0}), 
        .dqsbar_i({1'b0, 1'b0}), .dm_i({1'b0, 1'b0}), .odt_i(1'b0), 
        .resetbar_i(1'b0) );
  OR2X1 U27 ( .A(ck_i), .B(n4), .Y(n6) );
  INVX1 U28 ( .A(n6), .Y(n3) );
  INVX1 U29 ( .A(ready), .Y(n7) );
  AND2X1 U30 ( .A(init_casbar), .B(n7), .Y(casbar_i) );
  AND2X1 U31 ( .A(init_rasbar), .B(n7), .Y(rasbar_i) );
  AND2X1 U32 ( .A(init_webar), .B(n7), .Y(webar_i) );
  AND2X1 U33 ( .A(init_ba[0]), .B(n7), .Y(ba_i[0]) );
  AND2X1 U34 ( .A(init_ba[1]), .B(n7), .Y(ba_i[1]) );
  AND2X1 U35 ( .A(init_a[4]), .B(n7), .Y(a_i[4]) );
  AND2X1 U36 ( .A(init_a[8]), .B(n7), .Y(a_i[8]) );
  AND2X1 U37 ( .A(init_a[10]), .B(n7), .Y(a_i[10]) );
  INVX1 U38 ( .A(resetbar), .Y(n4) );
endmodule

