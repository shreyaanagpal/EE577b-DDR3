
module FIFO_2clk ( rclk, wclk, reset, we, re, data_in, empty_bar, full_bar, 
        data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input rclk, wclk, reset, we, re;
  output empty_bar, full_bar;
  wire   n14, n15, n16, n17, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, rd_ptr_bin_ss_1_,
         rd_ptr_bin_4_, n19, n20, n21, n22, n23, n24, n25, n26, n36, n37, n38,
         n39, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n108, n109, n110, n111, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1399, n1400, n1401, n1402, n1403,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749;
  wire   [3:0] wr_ptr_gray;
  wire   [3:0] wr_ptr_gray_ss;
  wire   [3:0] wr_ptr_gray_s;
  wire   [3:0] rd_ptr_gray;
  wire   [3:0] rd_ptr_gray_ss;
  wire   [3:0] rd_ptr_gray_s;
  wire   [4:0] wr_ptr_bin;
  wire   [4:1] full_check;
  wire   [511:0] fifo;
  wire   [4:2] add_169_carry;
  wire   [4:2] add_148_carry;
  wire   [4:1] sub_125_carry;

  DFFSR rd_ptr_gray_s_reg_0_ ( .D(n1967), .CLK(wclk), .R(n3643), .S(1'b1), .Q(
        rd_ptr_gray_s[0]) );
  DFFSR rd_ptr_gray_ss_reg_0_ ( .D(n1980), .CLK(wclk), .R(n3643), .S(1'b1), 
        .Q(rd_ptr_gray_ss[0]) );
  DFFSR rd_ptr_gray_s_reg_1_ ( .D(n1966), .CLK(wclk), .R(n3642), .S(1'b1), .Q(
        rd_ptr_gray_s[1]) );
  DFFSR rd_ptr_gray_ss_reg_1_ ( .D(n1979), .CLK(wclk), .R(n3642), .S(1'b1), 
        .Q(rd_ptr_gray_ss[1]) );
  DFFSR rd_ptr_gray_s_reg_2_ ( .D(n1965), .CLK(wclk), .R(n3642), .S(1'b1), .Q(
        rd_ptr_gray_s[2]) );
  DFFSR rd_ptr_gray_ss_reg_2_ ( .D(n1978), .CLK(wclk), .R(n3642), .S(1'b1), 
        .Q(rd_ptr_gray_ss[2]) );
  DFFSR rd_ptr_gray_s_reg_3_ ( .D(n1968), .CLK(wclk), .R(n3642), .S(1'b1), .Q(
        rd_ptr_gray_s[3]) );
  DFFSR rd_ptr_gray_ss_reg_3_ ( .D(n1977), .CLK(wclk), .R(n3642), .S(1'b1), 
        .Q(rd_ptr_gray_ss[3]) );
  DFFSR wr_ptr_bin_reg_4_ ( .D(n1922), .CLK(wclk), .R(n3642), .S(1'b1), .Q(
        wr_ptr_bin[4]) );
  DFFSR wr_ptr_bin_reg_0_ ( .D(n1921), .CLK(wclk), .R(n3641), .S(1'b1), .Q(
        wr_ptr_bin[0]) );
  DFFSR wr_ptr_bin_reg_1_ ( .D(n1920), .CLK(wclk), .R(n3641), .S(1'b1), .Q(
        wr_ptr_bin[1]) );
  DFFSR wr_ptr_gray_reg_0_ ( .D(n23), .CLK(wclk), .R(n3641), .S(1'b1), .Q(
        wr_ptr_gray[0]) );
  DFFSR wr_ptr_gray_s_reg_0_ ( .D(n1976), .CLK(rclk), .R(n3641), .S(1'b1), .Q(
        wr_ptr_gray_s[0]) );
  DFFSR wr_ptr_bin_reg_2_ ( .D(n1919), .CLK(wclk), .R(n3641), .S(1'b1), .Q(
        wr_ptr_bin[2]) );
  DFFSR wr_ptr_gray_reg_1_ ( .D(n1981), .CLK(wclk), .R(n3641), .S(1'b1), .Q(
        wr_ptr_gray[1]) );
  DFFSR wr_ptr_gray_s_reg_1_ ( .D(n1974), .CLK(rclk), .R(n3641), .S(1'b1), .Q(
        wr_ptr_gray_s[1]) );
  DFFSR wr_ptr_bin_reg_3_ ( .D(n1918), .CLK(wclk), .R(n3641), .S(1'b1), .Q(
        wr_ptr_bin[3]) );
  DFFSR wr_ptr_gray_reg_2_ ( .D(n25), .CLK(wclk), .R(n3641), .S(1'b1), .Q(
        wr_ptr_gray[2]) );
  DFFSR wr_ptr_gray_s_reg_2_ ( .D(n1972), .CLK(rclk), .R(n3641), .S(1'b1), .Q(
        wr_ptr_gray_s[2]) );
  DFFSR wr_ptr_gray_reg_3_ ( .D(n26), .CLK(wclk), .R(n3640), .S(1'b1), .Q(
        wr_ptr_gray[3]) );
  DFFSR wr_ptr_gray_s_reg_3_ ( .D(n1970), .CLK(rclk), .R(n3640), .S(1'b1), .Q(
        wr_ptr_gray_s[3]) );
  DFFSR fifo_reg_0__31_ ( .D(n1406), .CLK(wclk), .R(n3640), .S(1'b1), .Q(
        fifo[511]) );
  DFFSR fifo_reg_0__30_ ( .D(n1407), .CLK(wclk), .R(n3640), .S(1'b1), .Q(
        fifo[510]) );
  DFFSR fifo_reg_0__29_ ( .D(n1408), .CLK(wclk), .R(n3640), .S(1'b1), .Q(
        fifo[509]) );
  DFFSR fifo_reg_0__28_ ( .D(n1409), .CLK(wclk), .R(n3640), .S(1'b1), .Q(
        fifo[508]) );
  DFFSR fifo_reg_0__27_ ( .D(n1410), .CLK(wclk), .R(n3640), .S(1'b1), .Q(
        fifo[507]) );
  DFFSR fifo_reg_0__26_ ( .D(n1411), .CLK(wclk), .R(n3640), .S(1'b1), .Q(
        fifo[506]) );
  DFFSR fifo_reg_0__25_ ( .D(n1412), .CLK(wclk), .R(n3640), .S(1'b1), .Q(
        fifo[505]) );
  DFFSR fifo_reg_0__24_ ( .D(n1413), .CLK(wclk), .R(n3640), .S(1'b1), .Q(
        fifo[504]) );
  DFFSR fifo_reg_0__23_ ( .D(n1414), .CLK(wclk), .R(n3639), .S(1'b1), .Q(
        fifo[503]) );
  DFFSR fifo_reg_0__22_ ( .D(n1415), .CLK(wclk), .R(n3639), .S(1'b1), .Q(
        fifo[502]) );
  DFFSR fifo_reg_0__21_ ( .D(n1416), .CLK(wclk), .R(n3639), .S(1'b1), .Q(
        fifo[501]) );
  DFFSR fifo_reg_0__20_ ( .D(n1417), .CLK(wclk), .R(n3639), .S(1'b1), .Q(
        fifo[500]) );
  DFFSR fifo_reg_0__19_ ( .D(n1418), .CLK(wclk), .R(n3639), .S(1'b1), .Q(
        fifo[499]) );
  DFFSR fifo_reg_0__18_ ( .D(n1419), .CLK(wclk), .R(n3639), .S(1'b1), .Q(
        fifo[498]) );
  DFFSR fifo_reg_0__17_ ( .D(n1420), .CLK(wclk), .R(n3639), .S(1'b1), .Q(
        fifo[497]) );
  DFFSR fifo_reg_0__16_ ( .D(n1421), .CLK(wclk), .R(n3639), .S(1'b1), .Q(
        fifo[496]) );
  DFFSR fifo_reg_0__15_ ( .D(n1422), .CLK(wclk), .R(n3639), .S(1'b1), .Q(
        fifo[495]) );
  DFFSR fifo_reg_0__14_ ( .D(n1423), .CLK(wclk), .R(n3639), .S(1'b1), .Q(
        fifo[494]) );
  DFFSR fifo_reg_0__13_ ( .D(n1424), .CLK(wclk), .R(n3639), .S(1'b1), .Q(
        fifo[493]) );
  DFFSR fifo_reg_0__12_ ( .D(n1425), .CLK(wclk), .R(n3639), .S(1'b1), .Q(
        fifo[492]) );
  DFFSR fifo_reg_0__11_ ( .D(n1426), .CLK(wclk), .R(n3638), .S(1'b1), .Q(
        fifo[491]) );
  DFFSR fifo_reg_0__10_ ( .D(n1427), .CLK(wclk), .R(n3638), .S(1'b1), .Q(
        fifo[490]) );
  DFFSR fifo_reg_0__9_ ( .D(n1428), .CLK(wclk), .R(n3638), .S(1'b1), .Q(
        fifo[489]) );
  DFFSR fifo_reg_0__8_ ( .D(n1429), .CLK(wclk), .R(n3638), .S(1'b1), .Q(
        fifo[488]) );
  DFFSR fifo_reg_0__7_ ( .D(n1430), .CLK(wclk), .R(n3638), .S(1'b1), .Q(
        fifo[487]) );
  DFFSR fifo_reg_0__6_ ( .D(n1431), .CLK(wclk), .R(n3638), .S(1'b1), .Q(
        fifo[486]) );
  DFFSR fifo_reg_0__5_ ( .D(n1432), .CLK(wclk), .R(n3638), .S(1'b1), .Q(
        fifo[485]) );
  DFFSR fifo_reg_0__4_ ( .D(n1433), .CLK(wclk), .R(n3638), .S(1'b1), .Q(
        fifo[484]) );
  DFFSR fifo_reg_0__3_ ( .D(n1434), .CLK(wclk), .R(n3638), .S(1'b1), .Q(
        fifo[483]) );
  DFFSR fifo_reg_0__2_ ( .D(n1435), .CLK(wclk), .R(n3638), .S(1'b1), .Q(
        fifo[482]) );
  DFFSR fifo_reg_0__1_ ( .D(n1436), .CLK(wclk), .R(n3638), .S(1'b1), .Q(
        fifo[481]) );
  DFFSR fifo_reg_0__0_ ( .D(n1437), .CLK(wclk), .R(n3638), .S(1'b1), .Q(
        fifo[480]) );
  DFFSR fifo_reg_2__31_ ( .D(n1470), .CLK(wclk), .R(n3637), .S(1'b1), .Q(
        fifo[447]) );
  DFFSR fifo_reg_2__30_ ( .D(n1471), .CLK(wclk), .R(n3637), .S(1'b1), .Q(
        fifo[446]) );
  DFFSR fifo_reg_2__29_ ( .D(n1472), .CLK(wclk), .R(n3637), .S(1'b1), .Q(
        fifo[445]) );
  DFFSR fifo_reg_2__28_ ( .D(n1473), .CLK(wclk), .R(n3637), .S(1'b1), .Q(
        fifo[444]) );
  DFFSR fifo_reg_2__27_ ( .D(n1474), .CLK(wclk), .R(n3637), .S(1'b1), .Q(
        fifo[443]) );
  DFFSR fifo_reg_2__26_ ( .D(n1475), .CLK(wclk), .R(n3637), .S(1'b1), .Q(
        fifo[442]) );
  DFFSR fifo_reg_2__25_ ( .D(n1476), .CLK(wclk), .R(n3637), .S(1'b1), .Q(
        fifo[441]) );
  DFFSR fifo_reg_2__24_ ( .D(n1477), .CLK(wclk), .R(n3637), .S(1'b1), .Q(
        fifo[440]) );
  DFFSR fifo_reg_2__23_ ( .D(n1478), .CLK(wclk), .R(n3637), .S(1'b1), .Q(
        fifo[439]) );
  DFFSR fifo_reg_2__22_ ( .D(n1479), .CLK(wclk), .R(n3637), .S(1'b1), .Q(
        fifo[438]) );
  DFFSR fifo_reg_2__21_ ( .D(n1480), .CLK(wclk), .R(n3637), .S(1'b1), .Q(
        fifo[437]) );
  DFFSR fifo_reg_2__20_ ( .D(n1481), .CLK(wclk), .R(n3637), .S(1'b1), .Q(
        fifo[436]) );
  DFFSR fifo_reg_2__19_ ( .D(n1482), .CLK(wclk), .R(n3636), .S(1'b1), .Q(
        fifo[435]) );
  DFFSR fifo_reg_2__18_ ( .D(n1483), .CLK(wclk), .R(n3636), .S(1'b1), .Q(
        fifo[434]) );
  DFFSR fifo_reg_2__17_ ( .D(n1484), .CLK(wclk), .R(n3636), .S(1'b1), .Q(
        fifo[433]) );
  DFFSR fifo_reg_2__16_ ( .D(n1485), .CLK(wclk), .R(n3636), .S(1'b1), .Q(
        fifo[432]) );
  DFFSR fifo_reg_2__15_ ( .D(n1486), .CLK(wclk), .R(n3636), .S(1'b1), .Q(
        fifo[431]) );
  DFFSR fifo_reg_2__14_ ( .D(n1487), .CLK(wclk), .R(n3636), .S(1'b1), .Q(
        fifo[430]) );
  DFFSR fifo_reg_2__13_ ( .D(n1488), .CLK(wclk), .R(n3636), .S(1'b1), .Q(
        fifo[429]) );
  DFFSR fifo_reg_2__12_ ( .D(n1489), .CLK(wclk), .R(n3636), .S(1'b1), .Q(
        fifo[428]) );
  DFFSR fifo_reg_2__11_ ( .D(n1490), .CLK(wclk), .R(n3636), .S(1'b1), .Q(
        fifo[427]) );
  DFFSR fifo_reg_2__10_ ( .D(n1491), .CLK(wclk), .R(n3636), .S(1'b1), .Q(
        fifo[426]) );
  DFFSR fifo_reg_2__9_ ( .D(n1492), .CLK(wclk), .R(n3636), .S(1'b1), .Q(
        fifo[425]) );
  DFFSR fifo_reg_2__8_ ( .D(n1493), .CLK(wclk), .R(n3636), .S(1'b1), .Q(
        fifo[424]) );
  DFFSR fifo_reg_2__7_ ( .D(n1494), .CLK(wclk), .R(n3635), .S(1'b1), .Q(
        fifo[423]) );
  DFFSR fifo_reg_2__6_ ( .D(n1495), .CLK(wclk), .R(n3635), .S(1'b1), .Q(
        fifo[422]) );
  DFFSR fifo_reg_2__5_ ( .D(n1496), .CLK(wclk), .R(n3635), .S(1'b1), .Q(
        fifo[421]) );
  DFFSR fifo_reg_2__4_ ( .D(n1497), .CLK(wclk), .R(n3635), .S(1'b1), .Q(
        fifo[420]) );
  DFFSR fifo_reg_2__3_ ( .D(n1498), .CLK(wclk), .R(n3635), .S(1'b1), .Q(
        fifo[419]) );
  DFFSR fifo_reg_2__2_ ( .D(n1499), .CLK(wclk), .R(n3635), .S(1'b1), .Q(
        fifo[418]) );
  DFFSR fifo_reg_2__1_ ( .D(n1500), .CLK(wclk), .R(n3635), .S(1'b1), .Q(
        fifo[417]) );
  DFFSR fifo_reg_2__0_ ( .D(n1501), .CLK(wclk), .R(n3635), .S(1'b1), .Q(
        fifo[416]) );
  DFFSR fifo_reg_4__31_ ( .D(n1534), .CLK(wclk), .R(n3635), .S(1'b1), .Q(
        fifo[383]) );
  DFFSR fifo_reg_4__30_ ( .D(n1535), .CLK(wclk), .R(n3635), .S(1'b1), .Q(
        fifo[382]) );
  DFFSR fifo_reg_4__29_ ( .D(n1536), .CLK(wclk), .R(n3635), .S(1'b1), .Q(
        fifo[381]) );
  DFFSR fifo_reg_4__28_ ( .D(n1537), .CLK(wclk), .R(n3635), .S(1'b1), .Q(
        fifo[380]) );
  DFFSR fifo_reg_4__27_ ( .D(n1538), .CLK(wclk), .R(n3634), .S(1'b1), .Q(
        fifo[379]) );
  DFFSR fifo_reg_4__26_ ( .D(n1539), .CLK(wclk), .R(n3634), .S(1'b1), .Q(
        fifo[378]) );
  DFFSR fifo_reg_4__25_ ( .D(n1540), .CLK(wclk), .R(n3634), .S(1'b1), .Q(
        fifo[377]) );
  DFFSR fifo_reg_4__24_ ( .D(n1541), .CLK(wclk), .R(n3634), .S(1'b1), .Q(
        fifo[376]) );
  DFFSR fifo_reg_4__23_ ( .D(n1542), .CLK(wclk), .R(n3634), .S(1'b1), .Q(
        fifo[375]) );
  DFFSR fifo_reg_4__22_ ( .D(n1543), .CLK(wclk), .R(n3634), .S(1'b1), .Q(
        fifo[374]) );
  DFFSR fifo_reg_4__21_ ( .D(n1544), .CLK(wclk), .R(n3634), .S(1'b1), .Q(
        fifo[373]) );
  DFFSR fifo_reg_4__20_ ( .D(n1545), .CLK(wclk), .R(n3634), .S(1'b1), .Q(
        fifo[372]) );
  DFFSR fifo_reg_4__19_ ( .D(n1546), .CLK(wclk), .R(n3634), .S(1'b1), .Q(
        fifo[371]) );
  DFFSR fifo_reg_4__18_ ( .D(n1547), .CLK(wclk), .R(n3634), .S(1'b1), .Q(
        fifo[370]) );
  DFFSR fifo_reg_4__17_ ( .D(n1548), .CLK(wclk), .R(n3634), .S(1'b1), .Q(
        fifo[369]) );
  DFFSR fifo_reg_4__16_ ( .D(n1549), .CLK(wclk), .R(n3634), .S(1'b1), .Q(
        fifo[368]) );
  DFFSR fifo_reg_4__15_ ( .D(n1550), .CLK(wclk), .R(n3633), .S(1'b1), .Q(
        fifo[367]) );
  DFFSR fifo_reg_4__14_ ( .D(n1551), .CLK(wclk), .R(n3633), .S(1'b1), .Q(
        fifo[366]) );
  DFFSR fifo_reg_4__13_ ( .D(n1552), .CLK(wclk), .R(n3633), .S(1'b1), .Q(
        fifo[365]) );
  DFFSR fifo_reg_4__12_ ( .D(n1553), .CLK(wclk), .R(n3633), .S(1'b1), .Q(
        fifo[364]) );
  DFFSR fifo_reg_4__11_ ( .D(n1554), .CLK(wclk), .R(n3633), .S(1'b1), .Q(
        fifo[363]) );
  DFFSR fifo_reg_4__10_ ( .D(n1555), .CLK(wclk), .R(n3633), .S(1'b1), .Q(
        fifo[362]) );
  DFFSR fifo_reg_4__9_ ( .D(n1556), .CLK(wclk), .R(n3633), .S(1'b1), .Q(
        fifo[361]) );
  DFFSR fifo_reg_4__8_ ( .D(n1557), .CLK(wclk), .R(n3633), .S(1'b1), .Q(
        fifo[360]) );
  DFFSR fifo_reg_4__7_ ( .D(n1558), .CLK(wclk), .R(n3633), .S(1'b1), .Q(
        fifo[359]) );
  DFFSR fifo_reg_4__6_ ( .D(n1559), .CLK(wclk), .R(n3633), .S(1'b1), .Q(
        fifo[358]) );
  DFFSR fifo_reg_4__5_ ( .D(n1560), .CLK(wclk), .R(n3633), .S(1'b1), .Q(
        fifo[357]) );
  DFFSR fifo_reg_4__4_ ( .D(n1561), .CLK(wclk), .R(n3633), .S(1'b1), .Q(
        fifo[356]) );
  DFFSR fifo_reg_4__3_ ( .D(n1562), .CLK(wclk), .R(n3632), .S(1'b1), .Q(
        fifo[355]) );
  DFFSR fifo_reg_4__2_ ( .D(n1563), .CLK(wclk), .R(n3632), .S(1'b1), .Q(
        fifo[354]) );
  DFFSR fifo_reg_4__1_ ( .D(n1564), .CLK(wclk), .R(n3632), .S(1'b1), .Q(
        fifo[353]) );
  DFFSR fifo_reg_4__0_ ( .D(n1565), .CLK(wclk), .R(n3632), .S(1'b1), .Q(
        fifo[352]) );
  DFFSR fifo_reg_6__31_ ( .D(n1598), .CLK(wclk), .R(n3632), .S(1'b1), .Q(
        fifo[319]) );
  DFFSR fifo_reg_6__30_ ( .D(n1599), .CLK(wclk), .R(n3632), .S(1'b1), .Q(
        fifo[318]) );
  DFFSR fifo_reg_6__29_ ( .D(n1600), .CLK(wclk), .R(n3632), .S(1'b1), .Q(
        fifo[317]) );
  DFFSR fifo_reg_6__28_ ( .D(n1601), .CLK(wclk), .R(n3632), .S(1'b1), .Q(
        fifo[316]) );
  DFFSR fifo_reg_6__27_ ( .D(n1602), .CLK(wclk), .R(n3632), .S(1'b1), .Q(
        fifo[315]) );
  DFFSR fifo_reg_6__26_ ( .D(n1603), .CLK(wclk), .R(n3632), .S(1'b1), .Q(
        fifo[314]) );
  DFFSR fifo_reg_6__25_ ( .D(n1604), .CLK(wclk), .R(n3632), .S(1'b1), .Q(
        fifo[313]) );
  DFFSR fifo_reg_6__24_ ( .D(n1605), .CLK(wclk), .R(n3632), .S(1'b1), .Q(
        fifo[312]) );
  DFFSR fifo_reg_6__23_ ( .D(n1606), .CLK(wclk), .R(n3631), .S(1'b1), .Q(
        fifo[311]) );
  DFFSR fifo_reg_6__22_ ( .D(n1607), .CLK(wclk), .R(n3631), .S(1'b1), .Q(
        fifo[310]) );
  DFFSR fifo_reg_6__21_ ( .D(n1608), .CLK(wclk), .R(n3631), .S(1'b1), .Q(
        fifo[309]) );
  DFFSR fifo_reg_6__20_ ( .D(n1609), .CLK(wclk), .R(n3631), .S(1'b1), .Q(
        fifo[308]) );
  DFFSR fifo_reg_6__19_ ( .D(n1610), .CLK(wclk), .R(n3631), .S(1'b1), .Q(
        fifo[307]) );
  DFFSR fifo_reg_6__18_ ( .D(n1611), .CLK(wclk), .R(n3631), .S(1'b1), .Q(
        fifo[306]) );
  DFFSR fifo_reg_6__17_ ( .D(n1612), .CLK(wclk), .R(n3631), .S(1'b1), .Q(
        fifo[305]) );
  DFFSR fifo_reg_6__16_ ( .D(n1613), .CLK(wclk), .R(n3631), .S(1'b1), .Q(
        fifo[304]) );
  DFFSR fifo_reg_6__15_ ( .D(n1614), .CLK(wclk), .R(n3631), .S(1'b1), .Q(
        fifo[303]) );
  DFFSR fifo_reg_6__14_ ( .D(n1615), .CLK(wclk), .R(n3631), .S(1'b1), .Q(
        fifo[302]) );
  DFFSR fifo_reg_6__13_ ( .D(n1616), .CLK(wclk), .R(n3631), .S(1'b1), .Q(
        fifo[301]) );
  DFFSR fifo_reg_6__12_ ( .D(n1617), .CLK(wclk), .R(n3631), .S(1'b1), .Q(
        fifo[300]) );
  DFFSR fifo_reg_6__11_ ( .D(n1618), .CLK(wclk), .R(n3630), .S(1'b1), .Q(
        fifo[299]) );
  DFFSR fifo_reg_6__10_ ( .D(n1619), .CLK(wclk), .R(n3630), .S(1'b1), .Q(
        fifo[298]) );
  DFFSR fifo_reg_6__9_ ( .D(n1620), .CLK(wclk), .R(n3630), .S(1'b1), .Q(
        fifo[297]) );
  DFFSR fifo_reg_6__8_ ( .D(n1621), .CLK(wclk), .R(n3630), .S(1'b1), .Q(
        fifo[296]) );
  DFFSR fifo_reg_6__7_ ( .D(n1622), .CLK(wclk), .R(n3630), .S(1'b1), .Q(
        fifo[295]) );
  DFFSR fifo_reg_6__6_ ( .D(n1623), .CLK(wclk), .R(n3630), .S(1'b1), .Q(
        fifo[294]) );
  DFFSR fifo_reg_6__5_ ( .D(n1624), .CLK(wclk), .R(n3630), .S(1'b1), .Q(
        fifo[293]) );
  DFFSR fifo_reg_6__4_ ( .D(n1625), .CLK(wclk), .R(n3630), .S(1'b1), .Q(
        fifo[292]) );
  DFFSR fifo_reg_6__3_ ( .D(n1626), .CLK(wclk), .R(n3630), .S(1'b1), .Q(
        fifo[291]) );
  DFFSR fifo_reg_6__2_ ( .D(n1627), .CLK(wclk), .R(n3630), .S(1'b1), .Q(
        fifo[290]) );
  DFFSR fifo_reg_6__1_ ( .D(n1628), .CLK(wclk), .R(n3630), .S(1'b1), .Q(
        fifo[289]) );
  DFFSR fifo_reg_6__0_ ( .D(n1629), .CLK(wclk), .R(n3630), .S(1'b1), .Q(
        fifo[288]) );
  DFFSR fifo_reg_1__31_ ( .D(n1438), .CLK(wclk), .R(n3629), .S(1'b1), .Q(
        fifo[479]) );
  DFFSR fifo_reg_1__30_ ( .D(n1439), .CLK(wclk), .R(n3629), .S(1'b1), .Q(
        fifo[478]) );
  DFFSR fifo_reg_1__29_ ( .D(n1440), .CLK(wclk), .R(n3629), .S(1'b1), .Q(
        fifo[477]) );
  DFFSR fifo_reg_1__28_ ( .D(n1441), .CLK(wclk), .R(n3629), .S(1'b1), .Q(
        fifo[476]) );
  DFFSR fifo_reg_1__27_ ( .D(n1442), .CLK(wclk), .R(n3629), .S(1'b1), .Q(
        fifo[475]) );
  DFFSR fifo_reg_1__26_ ( .D(n1443), .CLK(wclk), .R(n3629), .S(1'b1), .Q(
        fifo[474]) );
  DFFSR fifo_reg_1__25_ ( .D(n1444), .CLK(wclk), .R(n3629), .S(1'b1), .Q(
        fifo[473]) );
  DFFSR fifo_reg_1__24_ ( .D(n1445), .CLK(wclk), .R(n3629), .S(1'b1), .Q(
        fifo[472]) );
  DFFSR fifo_reg_1__23_ ( .D(n1446), .CLK(wclk), .R(n3629), .S(1'b1), .Q(
        fifo[471]) );
  DFFSR fifo_reg_1__22_ ( .D(n1447), .CLK(wclk), .R(n3629), .S(1'b1), .Q(
        fifo[470]) );
  DFFSR fifo_reg_1__21_ ( .D(n1448), .CLK(wclk), .R(n3629), .S(1'b1), .Q(
        fifo[469]) );
  DFFSR fifo_reg_1__20_ ( .D(n1449), .CLK(wclk), .R(n3629), .S(1'b1), .Q(
        fifo[468]) );
  DFFSR fifo_reg_1__19_ ( .D(n1450), .CLK(wclk), .R(n3628), .S(1'b1), .Q(
        fifo[467]) );
  DFFSR fifo_reg_1__18_ ( .D(n1451), .CLK(wclk), .R(n3628), .S(1'b1), .Q(
        fifo[466]) );
  DFFSR fifo_reg_1__17_ ( .D(n1452), .CLK(wclk), .R(n3628), .S(1'b1), .Q(
        fifo[465]) );
  DFFSR fifo_reg_1__16_ ( .D(n1453), .CLK(wclk), .R(n3628), .S(1'b1), .Q(
        fifo[464]) );
  DFFSR fifo_reg_1__15_ ( .D(n1454), .CLK(wclk), .R(n3628), .S(1'b1), .Q(
        fifo[463]) );
  DFFSR fifo_reg_1__14_ ( .D(n1455), .CLK(wclk), .R(n3628), .S(1'b1), .Q(
        fifo[462]) );
  DFFSR fifo_reg_1__13_ ( .D(n1456), .CLK(wclk), .R(n3628), .S(1'b1), .Q(
        fifo[461]) );
  DFFSR fifo_reg_1__12_ ( .D(n1457), .CLK(wclk), .R(n3628), .S(1'b1), .Q(
        fifo[460]) );
  DFFSR fifo_reg_1__11_ ( .D(n1458), .CLK(wclk), .R(n3628), .S(1'b1), .Q(
        fifo[459]) );
  DFFSR fifo_reg_1__10_ ( .D(n1459), .CLK(wclk), .R(n3628), .S(1'b1), .Q(
        fifo[458]) );
  DFFSR fifo_reg_1__9_ ( .D(n1460), .CLK(wclk), .R(n3628), .S(1'b1), .Q(
        fifo[457]) );
  DFFSR fifo_reg_1__8_ ( .D(n1461), .CLK(wclk), .R(n3628), .S(1'b1), .Q(
        fifo[456]) );
  DFFSR fifo_reg_1__7_ ( .D(n1462), .CLK(wclk), .R(n3627), .S(1'b1), .Q(
        fifo[455]) );
  DFFSR fifo_reg_1__6_ ( .D(n1463), .CLK(wclk), .R(n3627), .S(1'b1), .Q(
        fifo[454]) );
  DFFSR fifo_reg_1__5_ ( .D(n1464), .CLK(wclk), .R(n3627), .S(1'b1), .Q(
        fifo[453]) );
  DFFSR fifo_reg_1__4_ ( .D(n1465), .CLK(wclk), .R(n3627), .S(1'b1), .Q(
        fifo[452]) );
  DFFSR fifo_reg_1__3_ ( .D(n1466), .CLK(wclk), .R(n3627), .S(1'b1), .Q(
        fifo[451]) );
  DFFSR fifo_reg_1__2_ ( .D(n1467), .CLK(wclk), .R(n3627), .S(1'b1), .Q(
        fifo[450]) );
  DFFSR fifo_reg_1__1_ ( .D(n1468), .CLK(wclk), .R(n3627), .S(1'b1), .Q(
        fifo[449]) );
  DFFSR fifo_reg_1__0_ ( .D(n1469), .CLK(wclk), .R(n3627), .S(1'b1), .Q(
        fifo[448]) );
  DFFSR fifo_reg_3__31_ ( .D(n1502), .CLK(wclk), .R(n3627), .S(1'b1), .Q(
        fifo[415]) );
  DFFSR fifo_reg_3__30_ ( .D(n1503), .CLK(wclk), .R(n3627), .S(1'b1), .Q(
        fifo[414]) );
  DFFSR fifo_reg_3__29_ ( .D(n1504), .CLK(wclk), .R(n3627), .S(1'b1), .Q(
        fifo[413]) );
  DFFSR fifo_reg_3__28_ ( .D(n1505), .CLK(wclk), .R(n3627), .S(1'b1), .Q(
        fifo[412]) );
  DFFSR fifo_reg_3__27_ ( .D(n1506), .CLK(wclk), .R(n3626), .S(1'b1), .Q(
        fifo[411]) );
  DFFSR fifo_reg_3__26_ ( .D(n1507), .CLK(wclk), .R(n3626), .S(1'b1), .Q(
        fifo[410]) );
  DFFSR fifo_reg_3__25_ ( .D(n1508), .CLK(wclk), .R(n3626), .S(1'b1), .Q(
        fifo[409]) );
  DFFSR fifo_reg_3__24_ ( .D(n1509), .CLK(wclk), .R(n3626), .S(1'b1), .Q(
        fifo[408]) );
  DFFSR fifo_reg_3__23_ ( .D(n1510), .CLK(wclk), .R(n3626), .S(1'b1), .Q(
        fifo[407]) );
  DFFSR fifo_reg_3__22_ ( .D(n1511), .CLK(wclk), .R(n3626), .S(1'b1), .Q(
        fifo[406]) );
  DFFSR fifo_reg_3__21_ ( .D(n1512), .CLK(wclk), .R(n3626), .S(1'b1), .Q(
        fifo[405]) );
  DFFSR fifo_reg_3__20_ ( .D(n1513), .CLK(wclk), .R(n3626), .S(1'b1), .Q(
        fifo[404]) );
  DFFSR fifo_reg_3__19_ ( .D(n1514), .CLK(wclk), .R(n3626), .S(1'b1), .Q(
        fifo[403]) );
  DFFSR fifo_reg_3__18_ ( .D(n1515), .CLK(wclk), .R(n3626), .S(1'b1), .Q(
        fifo[402]) );
  DFFSR fifo_reg_3__17_ ( .D(n1516), .CLK(wclk), .R(n3626), .S(1'b1), .Q(
        fifo[401]) );
  DFFSR fifo_reg_3__16_ ( .D(n1517), .CLK(wclk), .R(n3626), .S(1'b1), .Q(
        fifo[400]) );
  DFFSR fifo_reg_3__15_ ( .D(n1518), .CLK(wclk), .R(n3625), .S(1'b1), .Q(
        fifo[399]) );
  DFFSR fifo_reg_3__14_ ( .D(n1519), .CLK(wclk), .R(n3625), .S(1'b1), .Q(
        fifo[398]) );
  DFFSR fifo_reg_3__13_ ( .D(n1520), .CLK(wclk), .R(n3625), .S(1'b1), .Q(
        fifo[397]) );
  DFFSR fifo_reg_3__12_ ( .D(n1521), .CLK(wclk), .R(n3625), .S(1'b1), .Q(
        fifo[396]) );
  DFFSR fifo_reg_3__11_ ( .D(n1522), .CLK(wclk), .R(n3625), .S(1'b1), .Q(
        fifo[395]) );
  DFFSR fifo_reg_3__10_ ( .D(n1523), .CLK(wclk), .R(n3625), .S(1'b1), .Q(
        fifo[394]) );
  DFFSR fifo_reg_3__9_ ( .D(n1524), .CLK(wclk), .R(n3625), .S(1'b1), .Q(
        fifo[393]) );
  DFFSR fifo_reg_3__8_ ( .D(n1525), .CLK(wclk), .R(n3625), .S(1'b1), .Q(
        fifo[392]) );
  DFFSR fifo_reg_3__7_ ( .D(n1526), .CLK(wclk), .R(n3625), .S(1'b1), .Q(
        fifo[391]) );
  DFFSR fifo_reg_3__6_ ( .D(n1527), .CLK(wclk), .R(n3625), .S(1'b1), .Q(
        fifo[390]) );
  DFFSR fifo_reg_3__5_ ( .D(n1528), .CLK(wclk), .R(n3625), .S(1'b1), .Q(
        fifo[389]) );
  DFFSR fifo_reg_3__4_ ( .D(n1529), .CLK(wclk), .R(n3625), .S(1'b1), .Q(
        fifo[388]) );
  DFFSR fifo_reg_3__3_ ( .D(n1530), .CLK(wclk), .R(n3624), .S(1'b1), .Q(
        fifo[387]) );
  DFFSR fifo_reg_3__2_ ( .D(n1531), .CLK(wclk), .R(n3624), .S(1'b1), .Q(
        fifo[386]) );
  DFFSR fifo_reg_3__1_ ( .D(n1532), .CLK(wclk), .R(n3624), .S(1'b1), .Q(
        fifo[385]) );
  DFFSR fifo_reg_3__0_ ( .D(n1533), .CLK(wclk), .R(n3624), .S(1'b1), .Q(
        fifo[384]) );
  DFFSR fifo_reg_5__31_ ( .D(n1566), .CLK(wclk), .R(n3624), .S(1'b1), .Q(
        fifo[351]) );
  DFFSR fifo_reg_5__30_ ( .D(n1567), .CLK(wclk), .R(n3624), .S(1'b1), .Q(
        fifo[350]) );
  DFFSR fifo_reg_5__29_ ( .D(n1568), .CLK(wclk), .R(n3624), .S(1'b1), .Q(
        fifo[349]) );
  DFFSR fifo_reg_5__28_ ( .D(n1569), .CLK(wclk), .R(n3624), .S(1'b1), .Q(
        fifo[348]) );
  DFFSR fifo_reg_5__27_ ( .D(n1570), .CLK(wclk), .R(n3624), .S(1'b1), .Q(
        fifo[347]) );
  DFFSR fifo_reg_5__26_ ( .D(n1571), .CLK(wclk), .R(n3624), .S(1'b1), .Q(
        fifo[346]) );
  DFFSR fifo_reg_5__25_ ( .D(n1572), .CLK(wclk), .R(n3624), .S(1'b1), .Q(
        fifo[345]) );
  DFFSR fifo_reg_5__24_ ( .D(n1573), .CLK(wclk), .R(n3624), .S(1'b1), .Q(
        fifo[344]) );
  DFFSR fifo_reg_5__23_ ( .D(n1574), .CLK(wclk), .R(n3623), .S(1'b1), .Q(
        fifo[343]) );
  DFFSR fifo_reg_5__22_ ( .D(n1575), .CLK(wclk), .R(n3623), .S(1'b1), .Q(
        fifo[342]) );
  DFFSR fifo_reg_5__21_ ( .D(n1576), .CLK(wclk), .R(n3623), .S(1'b1), .Q(
        fifo[341]) );
  DFFSR fifo_reg_5__20_ ( .D(n1577), .CLK(wclk), .R(n3623), .S(1'b1), .Q(
        fifo[340]) );
  DFFSR fifo_reg_5__19_ ( .D(n1578), .CLK(wclk), .R(n3623), .S(1'b1), .Q(
        fifo[339]) );
  DFFSR fifo_reg_5__18_ ( .D(n1579), .CLK(wclk), .R(n3623), .S(1'b1), .Q(
        fifo[338]) );
  DFFSR fifo_reg_5__17_ ( .D(n1580), .CLK(wclk), .R(n3623), .S(1'b1), .Q(
        fifo[337]) );
  DFFSR fifo_reg_5__16_ ( .D(n1581), .CLK(wclk), .R(n3623), .S(1'b1), .Q(
        fifo[336]) );
  DFFSR fifo_reg_5__15_ ( .D(n1582), .CLK(wclk), .R(n3623), .S(1'b1), .Q(
        fifo[335]) );
  DFFSR fifo_reg_5__14_ ( .D(n1583), .CLK(wclk), .R(n3623), .S(1'b1), .Q(
        fifo[334]) );
  DFFSR fifo_reg_5__13_ ( .D(n1584), .CLK(wclk), .R(n3623), .S(1'b1), .Q(
        fifo[333]) );
  DFFSR fifo_reg_5__12_ ( .D(n1585), .CLK(wclk), .R(n3623), .S(1'b1), .Q(
        fifo[332]) );
  DFFSR fifo_reg_5__11_ ( .D(n1586), .CLK(wclk), .R(n3622), .S(1'b1), .Q(
        fifo[331]) );
  DFFSR fifo_reg_5__10_ ( .D(n1587), .CLK(wclk), .R(n3622), .S(1'b1), .Q(
        fifo[330]) );
  DFFSR fifo_reg_5__9_ ( .D(n1588), .CLK(wclk), .R(n3622), .S(1'b1), .Q(
        fifo[329]) );
  DFFSR fifo_reg_5__8_ ( .D(n1589), .CLK(wclk), .R(n3622), .S(1'b1), .Q(
        fifo[328]) );
  DFFSR fifo_reg_5__7_ ( .D(n1590), .CLK(wclk), .R(n3622), .S(1'b1), .Q(
        fifo[327]) );
  DFFSR fifo_reg_5__6_ ( .D(n1591), .CLK(wclk), .R(n3622), .S(1'b1), .Q(
        fifo[326]) );
  DFFSR fifo_reg_5__5_ ( .D(n1592), .CLK(wclk), .R(n3622), .S(1'b1), .Q(
        fifo[325]) );
  DFFSR fifo_reg_5__4_ ( .D(n1593), .CLK(wclk), .R(n3622), .S(1'b1), .Q(
        fifo[324]) );
  DFFSR fifo_reg_5__3_ ( .D(n1594), .CLK(wclk), .R(n3622), .S(1'b1), .Q(
        fifo[323]) );
  DFFSR fifo_reg_5__2_ ( .D(n1595), .CLK(wclk), .R(n3622), .S(1'b1), .Q(
        fifo[322]) );
  DFFSR fifo_reg_5__1_ ( .D(n1596), .CLK(wclk), .R(n3622), .S(1'b1), .Q(
        fifo[321]) );
  DFFSR fifo_reg_5__0_ ( .D(n1597), .CLK(wclk), .R(n3622), .S(1'b1), .Q(
        fifo[320]) );
  DFFSR fifo_reg_7__31_ ( .D(n1630), .CLK(wclk), .R(n3621), .S(1'b1), .Q(
        fifo[287]) );
  DFFSR fifo_reg_7__30_ ( .D(n1631), .CLK(wclk), .R(n3621), .S(1'b1), .Q(
        fifo[286]) );
  DFFSR fifo_reg_7__29_ ( .D(n1632), .CLK(wclk), .R(n3621), .S(1'b1), .Q(
        fifo[285]) );
  DFFSR fifo_reg_7__28_ ( .D(n1633), .CLK(wclk), .R(n3621), .S(1'b1), .Q(
        fifo[284]) );
  DFFSR fifo_reg_7__27_ ( .D(n1634), .CLK(wclk), .R(n3621), .S(1'b1), .Q(
        fifo[283]) );
  DFFSR fifo_reg_7__26_ ( .D(n1635), .CLK(wclk), .R(n3621), .S(1'b1), .Q(
        fifo[282]) );
  DFFSR fifo_reg_7__25_ ( .D(n1636), .CLK(wclk), .R(n3621), .S(1'b1), .Q(
        fifo[281]) );
  DFFSR fifo_reg_7__24_ ( .D(n1637), .CLK(wclk), .R(n3621), .S(1'b1), .Q(
        fifo[280]) );
  DFFSR fifo_reg_7__23_ ( .D(n1638), .CLK(wclk), .R(n3621), .S(1'b1), .Q(
        fifo[279]) );
  DFFSR fifo_reg_7__22_ ( .D(n1639), .CLK(wclk), .R(n3621), .S(1'b1), .Q(
        fifo[278]) );
  DFFSR fifo_reg_7__21_ ( .D(n1640), .CLK(wclk), .R(n3621), .S(1'b1), .Q(
        fifo[277]) );
  DFFSR fifo_reg_7__20_ ( .D(n1641), .CLK(wclk), .R(n3621), .S(1'b1), .Q(
        fifo[276]) );
  DFFSR fifo_reg_7__19_ ( .D(n1642), .CLK(wclk), .R(n3620), .S(1'b1), .Q(
        fifo[275]) );
  DFFSR fifo_reg_7__18_ ( .D(n1643), .CLK(wclk), .R(n3620), .S(1'b1), .Q(
        fifo[274]) );
  DFFSR fifo_reg_7__17_ ( .D(n1644), .CLK(wclk), .R(n3620), .S(1'b1), .Q(
        fifo[273]) );
  DFFSR fifo_reg_7__16_ ( .D(n1645), .CLK(wclk), .R(n3620), .S(1'b1), .Q(
        fifo[272]) );
  DFFSR fifo_reg_7__15_ ( .D(n1646), .CLK(wclk), .R(n3620), .S(1'b1), .Q(
        fifo[271]) );
  DFFSR fifo_reg_7__14_ ( .D(n1647), .CLK(wclk), .R(n3620), .S(1'b1), .Q(
        fifo[270]) );
  DFFSR fifo_reg_7__13_ ( .D(n1648), .CLK(wclk), .R(n3620), .S(1'b1), .Q(
        fifo[269]) );
  DFFSR fifo_reg_7__12_ ( .D(n1649), .CLK(wclk), .R(n3620), .S(1'b1), .Q(
        fifo[268]) );
  DFFSR fifo_reg_7__11_ ( .D(n1650), .CLK(wclk), .R(n3620), .S(1'b1), .Q(
        fifo[267]) );
  DFFSR fifo_reg_7__10_ ( .D(n1651), .CLK(wclk), .R(n3620), .S(1'b1), .Q(
        fifo[266]) );
  DFFSR fifo_reg_7__9_ ( .D(n1652), .CLK(wclk), .R(n3620), .S(1'b1), .Q(
        fifo[265]) );
  DFFSR fifo_reg_7__8_ ( .D(n1653), .CLK(wclk), .R(n3620), .S(1'b1), .Q(
        fifo[264]) );
  DFFSR fifo_reg_7__7_ ( .D(n1654), .CLK(wclk), .R(n3619), .S(1'b1), .Q(
        fifo[263]) );
  DFFSR fifo_reg_7__6_ ( .D(n1655), .CLK(wclk), .R(n3619), .S(1'b1), .Q(
        fifo[262]) );
  DFFSR fifo_reg_7__5_ ( .D(n1656), .CLK(wclk), .R(n3619), .S(1'b1), .Q(
        fifo[261]) );
  DFFSR fifo_reg_7__4_ ( .D(n1657), .CLK(wclk), .R(n3619), .S(1'b1), .Q(
        fifo[260]) );
  DFFSR fifo_reg_7__3_ ( .D(n1658), .CLK(wclk), .R(n3619), .S(1'b1), .Q(
        fifo[259]) );
  DFFSR fifo_reg_7__2_ ( .D(n1659), .CLK(wclk), .R(n3619), .S(1'b1), .Q(
        fifo[258]) );
  DFFSR fifo_reg_7__1_ ( .D(n1660), .CLK(wclk), .R(n3619), .S(1'b1), .Q(
        fifo[257]) );
  DFFSR fifo_reg_7__0_ ( .D(n1661), .CLK(wclk), .R(n3619), .S(1'b1), .Q(
        fifo[256]) );
  DFFSR fifo_reg_8__31_ ( .D(n1662), .CLK(wclk), .R(n3619), .S(1'b1), .Q(
        fifo[255]) );
  DFFSR fifo_reg_8__30_ ( .D(n1663), .CLK(wclk), .R(n3619), .S(1'b1), .Q(
        fifo[254]) );
  DFFSR fifo_reg_8__29_ ( .D(n1664), .CLK(wclk), .R(n3619), .S(1'b1), .Q(
        fifo[253]) );
  DFFSR fifo_reg_8__28_ ( .D(n1665), .CLK(wclk), .R(n3619), .S(1'b1), .Q(
        fifo[252]) );
  DFFSR fifo_reg_8__27_ ( .D(n1666), .CLK(wclk), .R(n3618), .S(1'b1), .Q(
        fifo[251]) );
  DFFSR fifo_reg_8__26_ ( .D(n1667), .CLK(wclk), .R(n3618), .S(1'b1), .Q(
        fifo[250]) );
  DFFSR fifo_reg_8__25_ ( .D(n1668), .CLK(wclk), .R(n3618), .S(1'b1), .Q(
        fifo[249]) );
  DFFSR fifo_reg_8__24_ ( .D(n1669), .CLK(wclk), .R(n3618), .S(1'b1), .Q(
        fifo[248]) );
  DFFSR fifo_reg_8__23_ ( .D(n1670), .CLK(wclk), .R(n3618), .S(1'b1), .Q(
        fifo[247]) );
  DFFSR fifo_reg_8__22_ ( .D(n1671), .CLK(wclk), .R(n3618), .S(1'b1), .Q(
        fifo[246]) );
  DFFSR fifo_reg_8__21_ ( .D(n1672), .CLK(wclk), .R(n3618), .S(1'b1), .Q(
        fifo[245]) );
  DFFSR fifo_reg_8__20_ ( .D(n1673), .CLK(wclk), .R(n3618), .S(1'b1), .Q(
        fifo[244]) );
  DFFSR fifo_reg_8__19_ ( .D(n1674), .CLK(wclk), .R(n3618), .S(1'b1), .Q(
        fifo[243]) );
  DFFSR fifo_reg_8__18_ ( .D(n1675), .CLK(wclk), .R(n3618), .S(1'b1), .Q(
        fifo[242]) );
  DFFSR fifo_reg_8__17_ ( .D(n1676), .CLK(wclk), .R(n3618), .S(1'b1), .Q(
        fifo[241]) );
  DFFSR fifo_reg_8__16_ ( .D(n1677), .CLK(wclk), .R(n3618), .S(1'b1), .Q(
        fifo[240]) );
  DFFSR fifo_reg_8__15_ ( .D(n1678), .CLK(wclk), .R(n3617), .S(1'b1), .Q(
        fifo[239]) );
  DFFSR fifo_reg_8__14_ ( .D(n1679), .CLK(wclk), .R(n3617), .S(1'b1), .Q(
        fifo[238]) );
  DFFSR fifo_reg_8__13_ ( .D(n1680), .CLK(wclk), .R(n3617), .S(1'b1), .Q(
        fifo[237]) );
  DFFSR fifo_reg_8__12_ ( .D(n1681), .CLK(wclk), .R(n3617), .S(1'b1), .Q(
        fifo[236]) );
  DFFSR fifo_reg_8__11_ ( .D(n1682), .CLK(wclk), .R(n3617), .S(1'b1), .Q(
        fifo[235]) );
  DFFSR fifo_reg_8__10_ ( .D(n1683), .CLK(wclk), .R(n3617), .S(1'b1), .Q(
        fifo[234]) );
  DFFSR fifo_reg_8__9_ ( .D(n1684), .CLK(wclk), .R(n3617), .S(1'b1), .Q(
        fifo[233]) );
  DFFSR fifo_reg_8__8_ ( .D(n1685), .CLK(wclk), .R(n3617), .S(1'b1), .Q(
        fifo[232]) );
  DFFSR fifo_reg_8__7_ ( .D(n1686), .CLK(wclk), .R(n3617), .S(1'b1), .Q(
        fifo[231]) );
  DFFSR fifo_reg_8__6_ ( .D(n1687), .CLK(wclk), .R(n3617), .S(1'b1), .Q(
        fifo[230]) );
  DFFSR fifo_reg_8__5_ ( .D(n1688), .CLK(wclk), .R(n3617), .S(1'b1), .Q(
        fifo[229]) );
  DFFSR fifo_reg_8__4_ ( .D(n1689), .CLK(wclk), .R(n3617), .S(1'b1), .Q(
        fifo[228]) );
  DFFSR fifo_reg_8__3_ ( .D(n1690), .CLK(wclk), .R(n3616), .S(1'b1), .Q(
        fifo[227]) );
  DFFSR fifo_reg_8__2_ ( .D(n1691), .CLK(wclk), .R(n3616), .S(1'b1), .Q(
        fifo[226]) );
  DFFSR fifo_reg_8__1_ ( .D(n1692), .CLK(wclk), .R(n3616), .S(1'b1), .Q(
        fifo[225]) );
  DFFSR fifo_reg_8__0_ ( .D(n1693), .CLK(wclk), .R(n3616), .S(1'b1), .Q(
        fifo[224]) );
  DFFSR fifo_reg_10__31_ ( .D(n1726), .CLK(wclk), .R(n3616), .S(1'b1), .Q(
        fifo[191]) );
  DFFSR fifo_reg_10__30_ ( .D(n1727), .CLK(wclk), .R(n3616), .S(1'b1), .Q(
        fifo[190]) );
  DFFSR fifo_reg_10__29_ ( .D(n1728), .CLK(wclk), .R(n3616), .S(1'b1), .Q(
        fifo[189]) );
  DFFSR fifo_reg_10__28_ ( .D(n1729), .CLK(wclk), .R(n3616), .S(1'b1), .Q(
        fifo[188]) );
  DFFSR fifo_reg_10__27_ ( .D(n1730), .CLK(wclk), .R(n3616), .S(1'b1), .Q(
        fifo[187]) );
  DFFSR fifo_reg_10__26_ ( .D(n1731), .CLK(wclk), .R(n3616), .S(1'b1), .Q(
        fifo[186]) );
  DFFSR fifo_reg_10__25_ ( .D(n1732), .CLK(wclk), .R(n3616), .S(1'b1), .Q(
        fifo[185]) );
  DFFSR fifo_reg_10__24_ ( .D(n1733), .CLK(wclk), .R(n3616), .S(1'b1), .Q(
        fifo[184]) );
  DFFSR fifo_reg_10__23_ ( .D(n1734), .CLK(wclk), .R(n3615), .S(1'b1), .Q(
        fifo[183]) );
  DFFSR fifo_reg_10__22_ ( .D(n1735), .CLK(wclk), .R(n3615), .S(1'b1), .Q(
        fifo[182]) );
  DFFSR fifo_reg_10__21_ ( .D(n1736), .CLK(wclk), .R(n3615), .S(1'b1), .Q(
        fifo[181]) );
  DFFSR fifo_reg_10__20_ ( .D(n1737), .CLK(wclk), .R(n3615), .S(1'b1), .Q(
        fifo[180]) );
  DFFSR fifo_reg_10__19_ ( .D(n1738), .CLK(wclk), .R(n3615), .S(1'b1), .Q(
        fifo[179]) );
  DFFSR fifo_reg_10__18_ ( .D(n1739), .CLK(wclk), .R(n3615), .S(1'b1), .Q(
        fifo[178]) );
  DFFSR fifo_reg_10__17_ ( .D(n1740), .CLK(wclk), .R(n3615), .S(1'b1), .Q(
        fifo[177]) );
  DFFSR fifo_reg_10__16_ ( .D(n1741), .CLK(wclk), .R(n3615), .S(1'b1), .Q(
        fifo[176]) );
  DFFSR fifo_reg_10__15_ ( .D(n1742), .CLK(wclk), .R(n3615), .S(1'b1), .Q(
        fifo[175]) );
  DFFSR fifo_reg_10__14_ ( .D(n1743), .CLK(wclk), .R(n3615), .S(1'b1), .Q(
        fifo[174]) );
  DFFSR fifo_reg_10__13_ ( .D(n1744), .CLK(wclk), .R(n3615), .S(1'b1), .Q(
        fifo[173]) );
  DFFSR fifo_reg_10__12_ ( .D(n1745), .CLK(wclk), .R(n3615), .S(1'b1), .Q(
        fifo[172]) );
  DFFSR fifo_reg_10__11_ ( .D(n1746), .CLK(wclk), .R(n3614), .S(1'b1), .Q(
        fifo[171]) );
  DFFSR fifo_reg_10__10_ ( .D(n1747), .CLK(wclk), .R(n3614), .S(1'b1), .Q(
        fifo[170]) );
  DFFSR fifo_reg_10__9_ ( .D(n1748), .CLK(wclk), .R(n3614), .S(1'b1), .Q(
        fifo[169]) );
  DFFSR fifo_reg_10__8_ ( .D(n1749), .CLK(wclk), .R(n3614), .S(1'b1), .Q(
        fifo[168]) );
  DFFSR fifo_reg_10__7_ ( .D(n1750), .CLK(wclk), .R(n3614), .S(1'b1), .Q(
        fifo[167]) );
  DFFSR fifo_reg_10__6_ ( .D(n1751), .CLK(wclk), .R(n3614), .S(1'b1), .Q(
        fifo[166]) );
  DFFSR fifo_reg_10__5_ ( .D(n1752), .CLK(wclk), .R(n3614), .S(1'b1), .Q(
        fifo[165]) );
  DFFSR fifo_reg_10__4_ ( .D(n1753), .CLK(wclk), .R(n3614), .S(1'b1), .Q(
        fifo[164]) );
  DFFSR fifo_reg_10__3_ ( .D(n1754), .CLK(wclk), .R(n3614), .S(1'b1), .Q(
        fifo[163]) );
  DFFSR fifo_reg_10__2_ ( .D(n1755), .CLK(wclk), .R(n3614), .S(1'b1), .Q(
        fifo[162]) );
  DFFSR fifo_reg_10__1_ ( .D(n1756), .CLK(wclk), .R(n3614), .S(1'b1), .Q(
        fifo[161]) );
  DFFSR fifo_reg_10__0_ ( .D(n1757), .CLK(wclk), .R(n3614), .S(1'b1), .Q(
        fifo[160]) );
  DFFSR fifo_reg_12__31_ ( .D(n1790), .CLK(wclk), .R(n3613), .S(1'b1), .Q(
        fifo[127]) );
  DFFSR fifo_reg_12__30_ ( .D(n1791), .CLK(wclk), .R(n3613), .S(1'b1), .Q(
        fifo[126]) );
  DFFSR fifo_reg_12__29_ ( .D(n1792), .CLK(wclk), .R(n3613), .S(1'b1), .Q(
        fifo[125]) );
  DFFSR fifo_reg_12__28_ ( .D(n1793), .CLK(wclk), .R(n3613), .S(1'b1), .Q(
        fifo[124]) );
  DFFSR fifo_reg_12__27_ ( .D(n1794), .CLK(wclk), .R(n3613), .S(1'b1), .Q(
        fifo[123]) );
  DFFSR fifo_reg_12__26_ ( .D(n1795), .CLK(wclk), .R(n3613), .S(1'b1), .Q(
        fifo[122]) );
  DFFSR fifo_reg_12__25_ ( .D(n1796), .CLK(wclk), .R(n3613), .S(1'b1), .Q(
        fifo[121]) );
  DFFSR fifo_reg_12__24_ ( .D(n1797), .CLK(wclk), .R(n3613), .S(1'b1), .Q(
        fifo[120]) );
  DFFSR fifo_reg_12__23_ ( .D(n1798), .CLK(wclk), .R(n3613), .S(1'b1), .Q(
        fifo[119]) );
  DFFSR fifo_reg_12__22_ ( .D(n1799), .CLK(wclk), .R(n3613), .S(1'b1), .Q(
        fifo[118]) );
  DFFSR fifo_reg_12__21_ ( .D(n1800), .CLK(wclk), .R(n3613), .S(1'b1), .Q(
        fifo[117]) );
  DFFSR fifo_reg_12__20_ ( .D(n1801), .CLK(wclk), .R(n3613), .S(1'b1), .Q(
        fifo[116]) );
  DFFSR fifo_reg_12__19_ ( .D(n1802), .CLK(wclk), .R(n3612), .S(1'b1), .Q(
        fifo[115]) );
  DFFSR fifo_reg_12__18_ ( .D(n1803), .CLK(wclk), .R(n3612), .S(1'b1), .Q(
        fifo[114]) );
  DFFSR fifo_reg_12__17_ ( .D(n1804), .CLK(wclk), .R(n3612), .S(1'b1), .Q(
        fifo[113]) );
  DFFSR fifo_reg_12__16_ ( .D(n1805), .CLK(wclk), .R(n3612), .S(1'b1), .Q(
        fifo[112]) );
  DFFSR fifo_reg_12__15_ ( .D(n1806), .CLK(wclk), .R(n3612), .S(1'b1), .Q(
        fifo[111]) );
  DFFSR fifo_reg_12__14_ ( .D(n1807), .CLK(wclk), .R(n3612), .S(1'b1), .Q(
        fifo[110]) );
  DFFSR fifo_reg_12__13_ ( .D(n1808), .CLK(wclk), .R(n3612), .S(1'b1), .Q(
        fifo[109]) );
  DFFSR fifo_reg_12__12_ ( .D(n1809), .CLK(wclk), .R(n3612), .S(1'b1), .Q(
        fifo[108]) );
  DFFSR fifo_reg_12__11_ ( .D(n1810), .CLK(wclk), .R(n3612), .S(1'b1), .Q(
        fifo[107]) );
  DFFSR fifo_reg_12__10_ ( .D(n1811), .CLK(wclk), .R(n3612), .S(1'b1), .Q(
        fifo[106]) );
  DFFSR fifo_reg_12__9_ ( .D(n1812), .CLK(wclk), .R(n3612), .S(1'b1), .Q(
        fifo[105]) );
  DFFSR fifo_reg_12__8_ ( .D(n1813), .CLK(wclk), .R(n3612), .S(1'b1), .Q(
        fifo[104]) );
  DFFSR fifo_reg_12__7_ ( .D(n1814), .CLK(wclk), .R(n3611), .S(1'b1), .Q(
        fifo[103]) );
  DFFSR fifo_reg_12__6_ ( .D(n1815), .CLK(wclk), .R(n3611), .S(1'b1), .Q(
        fifo[102]) );
  DFFSR fifo_reg_12__5_ ( .D(n1816), .CLK(wclk), .R(n3611), .S(1'b1), .Q(
        fifo[101]) );
  DFFSR fifo_reg_12__4_ ( .D(n1817), .CLK(wclk), .R(n3611), .S(1'b1), .Q(
        fifo[100]) );
  DFFSR fifo_reg_12__3_ ( .D(n1818), .CLK(wclk), .R(n3611), .S(1'b1), .Q(
        fifo[99]) );
  DFFSR fifo_reg_12__2_ ( .D(n1819), .CLK(wclk), .R(n3611), .S(1'b1), .Q(
        fifo[98]) );
  DFFSR fifo_reg_12__1_ ( .D(n1820), .CLK(wclk), .R(n3611), .S(1'b1), .Q(
        fifo[97]) );
  DFFSR fifo_reg_12__0_ ( .D(n1821), .CLK(wclk), .R(n3611), .S(1'b1), .Q(
        fifo[96]) );
  DFFSR fifo_reg_14__31_ ( .D(n1854), .CLK(wclk), .R(n3611), .S(1'b1), .Q(
        fifo[63]) );
  DFFSR fifo_reg_14__30_ ( .D(n1855), .CLK(wclk), .R(n3611), .S(1'b1), .Q(
        fifo[62]) );
  DFFSR fifo_reg_14__29_ ( .D(n1856), .CLK(wclk), .R(n3611), .S(1'b1), .Q(
        fifo[61]) );
  DFFSR fifo_reg_14__28_ ( .D(n1857), .CLK(wclk), .R(n3611), .S(1'b1), .Q(
        fifo[60]) );
  DFFSR fifo_reg_14__27_ ( .D(n1858), .CLK(wclk), .R(n3610), .S(1'b1), .Q(
        fifo[59]) );
  DFFSR fifo_reg_14__26_ ( .D(n1859), .CLK(wclk), .R(n3610), .S(1'b1), .Q(
        fifo[58]) );
  DFFSR fifo_reg_14__25_ ( .D(n1860), .CLK(wclk), .R(n3610), .S(1'b1), .Q(
        fifo[57]) );
  DFFSR fifo_reg_14__24_ ( .D(n1861), .CLK(wclk), .R(n3610), .S(1'b1), .Q(
        fifo[56]) );
  DFFSR fifo_reg_14__23_ ( .D(n1862), .CLK(wclk), .R(n3610), .S(1'b1), .Q(
        fifo[55]) );
  DFFSR fifo_reg_14__22_ ( .D(n1863), .CLK(wclk), .R(n3610), .S(1'b1), .Q(
        fifo[54]) );
  DFFSR fifo_reg_14__21_ ( .D(n1864), .CLK(wclk), .R(n3610), .S(1'b1), .Q(
        fifo[53]) );
  DFFSR fifo_reg_14__20_ ( .D(n1865), .CLK(wclk), .R(n3610), .S(1'b1), .Q(
        fifo[52]) );
  DFFSR fifo_reg_14__19_ ( .D(n1866), .CLK(wclk), .R(n3610), .S(1'b1), .Q(
        fifo[51]) );
  DFFSR fifo_reg_14__18_ ( .D(n1867), .CLK(wclk), .R(n3610), .S(1'b1), .Q(
        fifo[50]) );
  DFFSR fifo_reg_14__17_ ( .D(n1868), .CLK(wclk), .R(n3610), .S(1'b1), .Q(
        fifo[49]) );
  DFFSR fifo_reg_14__16_ ( .D(n1869), .CLK(wclk), .R(n3610), .S(1'b1), .Q(
        fifo[48]) );
  DFFSR fifo_reg_14__15_ ( .D(n1870), .CLK(wclk), .R(n3609), .S(1'b1), .Q(
        fifo[47]) );
  DFFSR fifo_reg_14__14_ ( .D(n1871), .CLK(wclk), .R(n3609), .S(1'b1), .Q(
        fifo[46]) );
  DFFSR fifo_reg_14__13_ ( .D(n1872), .CLK(wclk), .R(n3609), .S(1'b1), .Q(
        fifo[45]) );
  DFFSR fifo_reg_14__12_ ( .D(n1873), .CLK(wclk), .R(n3609), .S(1'b1), .Q(
        fifo[44]) );
  DFFSR fifo_reg_14__11_ ( .D(n1874), .CLK(wclk), .R(n3609), .S(1'b1), .Q(
        fifo[43]) );
  DFFSR fifo_reg_14__10_ ( .D(n1875), .CLK(wclk), .R(n3609), .S(1'b1), .Q(
        fifo[42]) );
  DFFSR fifo_reg_14__9_ ( .D(n1876), .CLK(wclk), .R(n3609), .S(1'b1), .Q(
        fifo[41]) );
  DFFSR fifo_reg_14__8_ ( .D(n1877), .CLK(wclk), .R(n3609), .S(1'b1), .Q(
        fifo[40]) );
  DFFSR fifo_reg_14__7_ ( .D(n1878), .CLK(wclk), .R(n3609), .S(1'b1), .Q(
        fifo[39]) );
  DFFSR fifo_reg_14__6_ ( .D(n1879), .CLK(wclk), .R(n3609), .S(1'b1), .Q(
        fifo[38]) );
  DFFSR fifo_reg_14__5_ ( .D(n1880), .CLK(wclk), .R(n3609), .S(1'b1), .Q(
        fifo[37]) );
  DFFSR fifo_reg_14__4_ ( .D(n1881), .CLK(wclk), .R(n3609), .S(1'b1), .Q(
        fifo[36]) );
  DFFSR fifo_reg_14__3_ ( .D(n1882), .CLK(wclk), .R(n3608), .S(1'b1), .Q(
        fifo[35]) );
  DFFSR fifo_reg_14__2_ ( .D(n1883), .CLK(wclk), .R(n3608), .S(1'b1), .Q(
        fifo[34]) );
  DFFSR fifo_reg_14__1_ ( .D(n1884), .CLK(wclk), .R(n3608), .S(1'b1), .Q(
        fifo[33]) );
  DFFSR fifo_reg_14__0_ ( .D(n1885), .CLK(wclk), .R(n3608), .S(1'b1), .Q(
        fifo[32]) );
  DFFSR fifo_reg_9__31_ ( .D(n1694), .CLK(wclk), .R(n3608), .S(1'b1), .Q(
        fifo[223]) );
  DFFSR fifo_reg_9__30_ ( .D(n1695), .CLK(wclk), .R(n3608), .S(1'b1), .Q(
        fifo[222]) );
  DFFSR fifo_reg_9__29_ ( .D(n1696), .CLK(wclk), .R(n3608), .S(1'b1), .Q(
        fifo[221]) );
  DFFSR fifo_reg_9__28_ ( .D(n1697), .CLK(wclk), .R(n3608), .S(1'b1), .Q(
        fifo[220]) );
  DFFSR fifo_reg_9__27_ ( .D(n1698), .CLK(wclk), .R(n3608), .S(1'b1), .Q(
        fifo[219]) );
  DFFSR fifo_reg_9__26_ ( .D(n1699), .CLK(wclk), .R(n3608), .S(1'b1), .Q(
        fifo[218]) );
  DFFSR fifo_reg_9__25_ ( .D(n1700), .CLK(wclk), .R(n3608), .S(1'b1), .Q(
        fifo[217]) );
  DFFSR fifo_reg_9__24_ ( .D(n1701), .CLK(wclk), .R(n3608), .S(1'b1), .Q(
        fifo[216]) );
  DFFSR fifo_reg_9__23_ ( .D(n1702), .CLK(wclk), .R(n3607), .S(1'b1), .Q(
        fifo[215]) );
  DFFSR fifo_reg_9__22_ ( .D(n1703), .CLK(wclk), .R(n3607), .S(1'b1), .Q(
        fifo[214]) );
  DFFSR fifo_reg_9__21_ ( .D(n1704), .CLK(wclk), .R(n3607), .S(1'b1), .Q(
        fifo[213]) );
  DFFSR fifo_reg_9__20_ ( .D(n1705), .CLK(wclk), .R(n3607), .S(1'b1), .Q(
        fifo[212]) );
  DFFSR fifo_reg_9__19_ ( .D(n1706), .CLK(wclk), .R(n3607), .S(1'b1), .Q(
        fifo[211]) );
  DFFSR fifo_reg_9__18_ ( .D(n1707), .CLK(wclk), .R(n3607), .S(1'b1), .Q(
        fifo[210]) );
  DFFSR fifo_reg_9__17_ ( .D(n1708), .CLK(wclk), .R(n3607), .S(1'b1), .Q(
        fifo[209]) );
  DFFSR fifo_reg_9__16_ ( .D(n1709), .CLK(wclk), .R(n3607), .S(1'b1), .Q(
        fifo[208]) );
  DFFSR fifo_reg_9__15_ ( .D(n1710), .CLK(wclk), .R(n3607), .S(1'b1), .Q(
        fifo[207]) );
  DFFSR fifo_reg_9__14_ ( .D(n1711), .CLK(wclk), .R(n3607), .S(1'b1), .Q(
        fifo[206]) );
  DFFSR fifo_reg_9__13_ ( .D(n1712), .CLK(wclk), .R(n3607), .S(1'b1), .Q(
        fifo[205]) );
  DFFSR fifo_reg_9__12_ ( .D(n1713), .CLK(wclk), .R(n3607), .S(1'b1), .Q(
        fifo[204]) );
  DFFSR fifo_reg_9__11_ ( .D(n1714), .CLK(wclk), .R(n3606), .S(1'b1), .Q(
        fifo[203]) );
  DFFSR fifo_reg_9__10_ ( .D(n1715), .CLK(wclk), .R(n3606), .S(1'b1), .Q(
        fifo[202]) );
  DFFSR fifo_reg_9__9_ ( .D(n1716), .CLK(wclk), .R(n3606), .S(1'b1), .Q(
        fifo[201]) );
  DFFSR fifo_reg_9__8_ ( .D(n1717), .CLK(wclk), .R(n3606), .S(1'b1), .Q(
        fifo[200]) );
  DFFSR fifo_reg_9__7_ ( .D(n1718), .CLK(wclk), .R(n3606), .S(1'b1), .Q(
        fifo[199]) );
  DFFSR fifo_reg_9__6_ ( .D(n1719), .CLK(wclk), .R(n3606), .S(1'b1), .Q(
        fifo[198]) );
  DFFSR fifo_reg_9__5_ ( .D(n1720), .CLK(wclk), .R(n3606), .S(1'b1), .Q(
        fifo[197]) );
  DFFSR fifo_reg_9__4_ ( .D(n1721), .CLK(wclk), .R(n3606), .S(1'b1), .Q(
        fifo[196]) );
  DFFSR fifo_reg_9__3_ ( .D(n1722), .CLK(wclk), .R(n3606), .S(1'b1), .Q(
        fifo[195]) );
  DFFSR fifo_reg_9__2_ ( .D(n1723), .CLK(wclk), .R(n3606), .S(1'b1), .Q(
        fifo[194]) );
  DFFSR fifo_reg_9__1_ ( .D(n1724), .CLK(wclk), .R(n3606), .S(1'b1), .Q(
        fifo[193]) );
  DFFSR fifo_reg_9__0_ ( .D(n1725), .CLK(wclk), .R(n3606), .S(1'b1), .Q(
        fifo[192]) );
  DFFSR fifo_reg_11__31_ ( .D(n1758), .CLK(wclk), .R(n3605), .S(1'b1), .Q(
        fifo[159]) );
  DFFSR fifo_reg_11__30_ ( .D(n1759), .CLK(wclk), .R(n3605), .S(1'b1), .Q(
        fifo[158]) );
  DFFSR fifo_reg_11__29_ ( .D(n1760), .CLK(wclk), .R(n3605), .S(1'b1), .Q(
        fifo[157]) );
  DFFSR fifo_reg_11__28_ ( .D(n1761), .CLK(wclk), .R(n3605), .S(1'b1), .Q(
        fifo[156]) );
  DFFSR fifo_reg_11__27_ ( .D(n1762), .CLK(wclk), .R(n3605), .S(1'b1), .Q(
        fifo[155]) );
  DFFSR fifo_reg_11__26_ ( .D(n1763), .CLK(wclk), .R(n3605), .S(1'b1), .Q(
        fifo[154]) );
  DFFSR fifo_reg_11__25_ ( .D(n1764), .CLK(wclk), .R(n3605), .S(1'b1), .Q(
        fifo[153]) );
  DFFSR fifo_reg_11__24_ ( .D(n1765), .CLK(wclk), .R(n3605), .S(1'b1), .Q(
        fifo[152]) );
  DFFSR fifo_reg_11__23_ ( .D(n1766), .CLK(wclk), .R(n3605), .S(1'b1), .Q(
        fifo[151]) );
  DFFSR fifo_reg_11__22_ ( .D(n1767), .CLK(wclk), .R(n3605), .S(1'b1), .Q(
        fifo[150]) );
  DFFSR fifo_reg_11__21_ ( .D(n1768), .CLK(wclk), .R(n3605), .S(1'b1), .Q(
        fifo[149]) );
  DFFSR fifo_reg_11__20_ ( .D(n1769), .CLK(wclk), .R(n3605), .S(1'b1), .Q(
        fifo[148]) );
  DFFSR fifo_reg_11__19_ ( .D(n1770), .CLK(wclk), .R(n3604), .S(1'b1), .Q(
        fifo[147]) );
  DFFSR fifo_reg_11__18_ ( .D(n1771), .CLK(wclk), .R(n3604), .S(1'b1), .Q(
        fifo[146]) );
  DFFSR fifo_reg_11__17_ ( .D(n1772), .CLK(wclk), .R(n3604), .S(1'b1), .Q(
        fifo[145]) );
  DFFSR fifo_reg_11__16_ ( .D(n1773), .CLK(wclk), .R(n3604), .S(1'b1), .Q(
        fifo[144]) );
  DFFSR fifo_reg_11__15_ ( .D(n1774), .CLK(wclk), .R(n3604), .S(1'b1), .Q(
        fifo[143]) );
  DFFSR fifo_reg_11__14_ ( .D(n1775), .CLK(wclk), .R(n3604), .S(1'b1), .Q(
        fifo[142]) );
  DFFSR fifo_reg_11__13_ ( .D(n1776), .CLK(wclk), .R(n3604), .S(1'b1), .Q(
        fifo[141]) );
  DFFSR fifo_reg_11__12_ ( .D(n1777), .CLK(wclk), .R(n3604), .S(1'b1), .Q(
        fifo[140]) );
  DFFSR fifo_reg_11__11_ ( .D(n1778), .CLK(wclk), .R(n3604), .S(1'b1), .Q(
        fifo[139]) );
  DFFSR fifo_reg_11__10_ ( .D(n1779), .CLK(wclk), .R(n3604), .S(1'b1), .Q(
        fifo[138]) );
  DFFSR fifo_reg_11__9_ ( .D(n1780), .CLK(wclk), .R(n3604), .S(1'b1), .Q(
        fifo[137]) );
  DFFSR fifo_reg_11__8_ ( .D(n1781), .CLK(wclk), .R(n3604), .S(1'b1), .Q(
        fifo[136]) );
  DFFSR fifo_reg_11__7_ ( .D(n1782), .CLK(wclk), .R(n3603), .S(1'b1), .Q(
        fifo[135]) );
  DFFSR fifo_reg_11__6_ ( .D(n1783), .CLK(wclk), .R(n3603), .S(1'b1), .Q(
        fifo[134]) );
  DFFSR fifo_reg_11__5_ ( .D(n1784), .CLK(wclk), .R(n3603), .S(1'b1), .Q(
        fifo[133]) );
  DFFSR fifo_reg_11__4_ ( .D(n1785), .CLK(wclk), .R(n3603), .S(1'b1), .Q(
        fifo[132]) );
  DFFSR fifo_reg_11__3_ ( .D(n1786), .CLK(wclk), .R(n3603), .S(1'b1), .Q(
        fifo[131]) );
  DFFSR fifo_reg_11__2_ ( .D(n1787), .CLK(wclk), .R(n3603), .S(1'b1), .Q(
        fifo[130]) );
  DFFSR fifo_reg_11__1_ ( .D(n1788), .CLK(wclk), .R(n3603), .S(1'b1), .Q(
        fifo[129]) );
  DFFSR fifo_reg_11__0_ ( .D(n1789), .CLK(wclk), .R(n3603), .S(1'b1), .Q(
        fifo[128]) );
  DFFSR fifo_reg_13__31_ ( .D(n1822), .CLK(wclk), .R(n3603), .S(1'b1), .Q(
        fifo[95]) );
  DFFSR fifo_reg_13__30_ ( .D(n1823), .CLK(wclk), .R(n3603), .S(1'b1), .Q(
        fifo[94]) );
  DFFSR fifo_reg_13__29_ ( .D(n1824), .CLK(wclk), .R(n3603), .S(1'b1), .Q(
        fifo[93]) );
  DFFSR fifo_reg_13__28_ ( .D(n1825), .CLK(wclk), .R(n3603), .S(1'b1), .Q(
        fifo[92]) );
  DFFSR fifo_reg_13__27_ ( .D(n1826), .CLK(wclk), .R(n3602), .S(1'b1), .Q(
        fifo[91]) );
  DFFSR fifo_reg_13__26_ ( .D(n1827), .CLK(wclk), .R(n3602), .S(1'b1), .Q(
        fifo[90]) );
  DFFSR fifo_reg_13__25_ ( .D(n1828), .CLK(wclk), .R(n3602), .S(1'b1), .Q(
        fifo[89]) );
  DFFSR fifo_reg_13__24_ ( .D(n1829), .CLK(wclk), .R(n3602), .S(1'b1), .Q(
        fifo[88]) );
  DFFSR fifo_reg_13__23_ ( .D(n1830), .CLK(wclk), .R(n3602), .S(1'b1), .Q(
        fifo[87]) );
  DFFSR fifo_reg_13__22_ ( .D(n1831), .CLK(wclk), .R(n3602), .S(1'b1), .Q(
        fifo[86]) );
  DFFSR fifo_reg_13__21_ ( .D(n1832), .CLK(wclk), .R(n3602), .S(1'b1), .Q(
        fifo[85]) );
  DFFSR fifo_reg_13__20_ ( .D(n1833), .CLK(wclk), .R(n3602), .S(1'b1), .Q(
        fifo[84]) );
  DFFSR fifo_reg_13__19_ ( .D(n1834), .CLK(wclk), .R(n3602), .S(1'b1), .Q(
        fifo[83]) );
  DFFSR fifo_reg_13__18_ ( .D(n1835), .CLK(wclk), .R(n3602), .S(1'b1), .Q(
        fifo[82]) );
  DFFSR fifo_reg_13__17_ ( .D(n1836), .CLK(wclk), .R(n3602), .S(1'b1), .Q(
        fifo[81]) );
  DFFSR fifo_reg_13__16_ ( .D(n1837), .CLK(wclk), .R(n3602), .S(1'b1), .Q(
        fifo[80]) );
  DFFSR fifo_reg_13__15_ ( .D(n1838), .CLK(wclk), .R(n3601), .S(1'b1), .Q(
        fifo[79]) );
  DFFSR fifo_reg_13__14_ ( .D(n1839), .CLK(wclk), .R(n3601), .S(1'b1), .Q(
        fifo[78]) );
  DFFSR fifo_reg_13__13_ ( .D(n1840), .CLK(wclk), .R(n3601), .S(1'b1), .Q(
        fifo[77]) );
  DFFSR fifo_reg_13__12_ ( .D(n1841), .CLK(wclk), .R(n3601), .S(1'b1), .Q(
        fifo[76]) );
  DFFSR fifo_reg_13__11_ ( .D(n1842), .CLK(wclk), .R(n3601), .S(1'b1), .Q(
        fifo[75]) );
  DFFSR fifo_reg_13__10_ ( .D(n1843), .CLK(wclk), .R(n3601), .S(1'b1), .Q(
        fifo[74]) );
  DFFSR fifo_reg_13__9_ ( .D(n1844), .CLK(wclk), .R(n3601), .S(1'b1), .Q(
        fifo[73]) );
  DFFSR fifo_reg_13__8_ ( .D(n1845), .CLK(wclk), .R(n3601), .S(1'b1), .Q(
        fifo[72]) );
  DFFSR fifo_reg_13__7_ ( .D(n1846), .CLK(wclk), .R(n3601), .S(1'b1), .Q(
        fifo[71]) );
  DFFSR fifo_reg_13__6_ ( .D(n1847), .CLK(wclk), .R(n3601), .S(1'b1), .Q(
        fifo[70]) );
  DFFSR fifo_reg_13__5_ ( .D(n1848), .CLK(wclk), .R(n3601), .S(1'b1), .Q(
        fifo[69]) );
  DFFSR fifo_reg_13__4_ ( .D(n1849), .CLK(wclk), .R(n3601), .S(1'b1), .Q(
        fifo[68]) );
  DFFSR fifo_reg_13__3_ ( .D(n1850), .CLK(wclk), .R(n3600), .S(1'b1), .Q(
        fifo[67]) );
  DFFSR fifo_reg_13__2_ ( .D(n1851), .CLK(wclk), .R(n3600), .S(1'b1), .Q(
        fifo[66]) );
  DFFSR fifo_reg_13__1_ ( .D(n1852), .CLK(wclk), .R(n3600), .S(1'b1), .Q(
        fifo[65]) );
  DFFSR fifo_reg_13__0_ ( .D(n1853), .CLK(wclk), .R(n3600), .S(1'b1), .Q(
        fifo[64]) );
  DFFSR fifo_reg_15__31_ ( .D(n1886), .CLK(wclk), .R(n3600), .S(1'b1), .Q(
        fifo[31]) );
  DFFSR fifo_reg_15__30_ ( .D(n1887), .CLK(wclk), .R(n3600), .S(1'b1), .Q(
        fifo[30]) );
  DFFSR fifo_reg_15__29_ ( .D(n1888), .CLK(wclk), .R(n3600), .S(1'b1), .Q(
        fifo[29]) );
  DFFSR fifo_reg_15__28_ ( .D(n1889), .CLK(wclk), .R(n3600), .S(1'b1), .Q(
        fifo[28]) );
  DFFSR fifo_reg_15__27_ ( .D(n1890), .CLK(wclk), .R(n3600), .S(1'b1), .Q(
        fifo[27]) );
  DFFSR fifo_reg_15__26_ ( .D(n1891), .CLK(wclk), .R(n3600), .S(1'b1), .Q(
        fifo[26]) );
  DFFSR fifo_reg_15__25_ ( .D(n1892), .CLK(wclk), .R(n3600), .S(1'b1), .Q(
        fifo[25]) );
  DFFSR fifo_reg_15__24_ ( .D(n1893), .CLK(wclk), .R(n3600), .S(1'b1), .Q(
        fifo[24]) );
  DFFSR fifo_reg_15__23_ ( .D(n1894), .CLK(wclk), .R(n3599), .S(1'b1), .Q(
        fifo[23]) );
  DFFSR fifo_reg_15__22_ ( .D(n1895), .CLK(wclk), .R(n3599), .S(1'b1), .Q(
        fifo[22]) );
  DFFSR fifo_reg_15__21_ ( .D(n1896), .CLK(wclk), .R(n3599), .S(1'b1), .Q(
        fifo[21]) );
  DFFSR fifo_reg_15__20_ ( .D(n1897), .CLK(wclk), .R(n3599), .S(1'b1), .Q(
        fifo[20]) );
  DFFSR fifo_reg_15__19_ ( .D(n1898), .CLK(wclk), .R(n3599), .S(1'b1), .Q(
        fifo[19]) );
  DFFSR fifo_reg_15__18_ ( .D(n1899), .CLK(wclk), .R(n3599), .S(1'b1), .Q(
        fifo[18]) );
  DFFSR fifo_reg_15__17_ ( .D(n1900), .CLK(wclk), .R(n3599), .S(1'b1), .Q(
        fifo[17]) );
  DFFSR fifo_reg_15__16_ ( .D(n1901), .CLK(wclk), .R(n3599), .S(1'b1), .Q(
        fifo[16]) );
  DFFSR fifo_reg_15__15_ ( .D(n1902), .CLK(wclk), .R(n3599), .S(1'b1), .Q(
        fifo[15]) );
  DFFSR fifo_reg_15__14_ ( .D(n1903), .CLK(wclk), .R(n3599), .S(1'b1), .Q(
        fifo[14]) );
  DFFSR fifo_reg_15__13_ ( .D(n1904), .CLK(wclk), .R(n3599), .S(1'b1), .Q(
        fifo[13]) );
  DFFSR fifo_reg_15__12_ ( .D(n1905), .CLK(wclk), .R(n3599), .S(1'b1), .Q(
        fifo[12]) );
  DFFSR fifo_reg_15__11_ ( .D(n1906), .CLK(wclk), .R(n3598), .S(1'b1), .Q(
        fifo[11]) );
  DFFSR fifo_reg_15__10_ ( .D(n1907), .CLK(wclk), .R(n3598), .S(1'b1), .Q(
        fifo[10]) );
  DFFSR fifo_reg_15__9_ ( .D(n1908), .CLK(wclk), .R(n3598), .S(1'b1), .Q(
        fifo[9]) );
  DFFSR fifo_reg_15__8_ ( .D(n1909), .CLK(wclk), .R(n3598), .S(1'b1), .Q(
        fifo[8]) );
  DFFSR fifo_reg_15__7_ ( .D(n1910), .CLK(wclk), .R(n3598), .S(1'b1), .Q(
        fifo[7]) );
  DFFSR fifo_reg_15__6_ ( .D(n1911), .CLK(wclk), .R(n3598), .S(1'b1), .Q(
        fifo[6]) );
  DFFSR fifo_reg_15__5_ ( .D(n1912), .CLK(wclk), .R(n3598), .S(1'b1), .Q(
        fifo[5]) );
  DFFSR fifo_reg_15__4_ ( .D(n1913), .CLK(wclk), .R(n3598), .S(1'b1), .Q(
        fifo[4]) );
  DFFSR fifo_reg_15__3_ ( .D(n1914), .CLK(wclk), .R(n3598), .S(1'b1), .Q(
        fifo[3]) );
  DFFSR fifo_reg_15__2_ ( .D(n1915), .CLK(wclk), .R(n3598), .S(1'b1), .Q(
        fifo[2]) );
  DFFSR fifo_reg_15__1_ ( .D(n1916), .CLK(wclk), .R(n3598), .S(1'b1), .Q(
        fifo[1]) );
  DFFSR fifo_reg_15__0_ ( .D(n1917), .CLK(wclk), .R(n3598), .S(1'b1), .Q(
        fifo[0]) );
  FAX1 U673 ( .A(n3108), .B(n2854), .C(n2634), .YC(), .YS(rd_ptr_bin_ss_1_) );
  OAI21X1 U675 ( .A(n3672), .B(n3712), .C(n2290), .Y(n1406) );
  OAI21X1 U677 ( .A(n3672), .B(n3713), .C(n2058), .Y(n1407) );
  OAI21X1 U679 ( .A(n3672), .B(n3714), .C(n2176), .Y(n1408) );
  OAI21X1 U681 ( .A(n3672), .B(n3715), .C(n2203), .Y(n1409) );
  OAI21X1 U683 ( .A(n3672), .B(n3716), .C(n2151), .Y(n1410) );
  OAI21X1 U685 ( .A(n3672), .B(n3717), .C(n2379), .Y(n1411) );
  OAI21X1 U687 ( .A(n3672), .B(n3718), .C(n2413), .Y(n1412) );
  OAI21X1 U689 ( .A(n3672), .B(n3719), .C(n2445), .Y(n1413) );
  OAI21X1 U691 ( .A(n3672), .B(n3720), .C(n2347), .Y(n1414) );
  OAI21X1 U693 ( .A(n3672), .B(n3721), .C(n2316), .Y(n1415) );
  OAI21X1 U695 ( .A(n3672), .B(n3722), .C(n2057), .Y(n1416) );
  OAI21X1 U697 ( .A(n3672), .B(n3723), .C(n2859), .Y(n1417) );
  OAI21X1 U699 ( .A(n3672), .B(n3724), .C(n2056), .Y(n1418) );
  OAI21X1 U701 ( .A(n3672), .B(n3725), .C(n2542), .Y(n1419) );
  OAI21X1 U703 ( .A(n3672), .B(n3726), .C(n2055), .Y(n1420) );
  OAI21X1 U705 ( .A(n3672), .B(n3727), .C(n2348), .Y(n1421) );
  OAI21X1 U707 ( .A(n3672), .B(n3728), .C(n2054), .Y(n1422) );
  OAI21X1 U709 ( .A(n3672), .B(n3729), .C(n2317), .Y(n1423) );
  OAI21X1 U711 ( .A(n3672), .B(n3730), .C(n2053), .Y(n1424) );
  OAI21X1 U713 ( .A(n3672), .B(n3731), .C(n2052), .Y(n1425) );
  OAI21X1 U715 ( .A(n3672), .B(n3732), .C(n2860), .Y(n1426) );
  OAI21X1 U717 ( .A(n3672), .B(n3733), .C(n2051), .Y(n1427) );
  OAI21X1 U719 ( .A(n3672), .B(n3734), .C(n2128), .Y(n1428) );
  OAI21X1 U721 ( .A(n3672), .B(n3735), .C(n2050), .Y(n1429) );
  OAI21X1 U723 ( .A(n3672), .B(n3736), .C(n2106), .Y(n1430) );
  OAI21X1 U725 ( .A(n3672), .B(n3737), .C(n2177), .Y(n1431) );
  OAI21X1 U727 ( .A(n3672), .B(n3738), .C(n2204), .Y(n1432) );
  OAI21X1 U729 ( .A(n3672), .B(n3739), .C(n2152), .Y(n1433) );
  OAI21X1 U731 ( .A(n3672), .B(n3740), .C(n2049), .Y(n1434) );
  OAI21X1 U733 ( .A(n3672), .B(n3741), .C(n2048), .Y(n1435) );
  OAI21X1 U735 ( .A(n3672), .B(n3742), .C(n2129), .Y(n1436) );
  OAI21X1 U737 ( .A(n3672), .B(n3743), .C(n2107), .Y(n1437) );
  OAI21X1 U740 ( .A(n3712), .B(n3671), .C(n2322), .Y(n1438) );
  OAI21X1 U742 ( .A(n3713), .B(n3671), .C(n2047), .Y(n1439) );
  OAI21X1 U744 ( .A(n3714), .B(n3671), .C(n2136), .Y(n1440) );
  OAI21X1 U746 ( .A(n3715), .B(n3671), .C(n2115), .Y(n1441) );
  OAI21X1 U748 ( .A(n3716), .B(n3671), .C(n2266), .Y(n1442) );
  OAI21X1 U750 ( .A(n3717), .B(n3671), .C(n2046), .Y(n1443) );
  OAI21X1 U752 ( .A(n3718), .B(n3671), .C(n2292), .Y(n1444) );
  OAI21X1 U754 ( .A(n3719), .B(n3671), .C(n2323), .Y(n1445) );
  OAI21X1 U756 ( .A(n3720), .B(n3671), .C(n2385), .Y(n1446) );
  OAI21X1 U758 ( .A(n3721), .B(n3671), .C(n2419), .Y(n1447) );
  OAI21X1 U760 ( .A(n3722), .B(n3671), .C(n2549), .Y(n1448) );
  OAI21X1 U762 ( .A(n3723), .B(n3671), .C(n2637), .Y(n1449) );
  OAI21X1 U764 ( .A(n3724), .B(n3671), .C(n2452), .Y(n1450) );
  OAI21X1 U766 ( .A(n3725), .B(n3671), .C(n2354), .Y(n1451) );
  OAI21X1 U768 ( .A(n3726), .B(n3671), .C(n2045), .Y(n1452) );
  OAI21X1 U770 ( .A(n3727), .B(n3671), .C(n2386), .Y(n1453) );
  OAI21X1 U772 ( .A(n3728), .B(n3671), .C(n2184), .Y(n1454) );
  OAI21X1 U774 ( .A(n3729), .B(n3671), .C(n2420), .Y(n1455) );
  OAI21X1 U776 ( .A(n3730), .B(n3671), .C(n2550), .Y(n1456) );
  OAI21X1 U778 ( .A(n3731), .B(n3671), .C(n2159), .Y(n1457) );
  OAI21X1 U780 ( .A(n3732), .B(n3671), .C(n2638), .Y(n1458) );
  OAI21X1 U782 ( .A(n3733), .B(n3671), .C(n2453), .Y(n1459) );
  OAI21X1 U784 ( .A(n3734), .B(n3671), .C(n2240), .Y(n1460) );
  OAI21X1 U786 ( .A(n3735), .B(n3671), .C(n2044), .Y(n1461) );
  OAI21X1 U788 ( .A(n3736), .B(n3671), .C(n2210), .Y(n1462) );
  OAI21X1 U790 ( .A(n3737), .B(n3671), .C(n2137), .Y(n1463) );
  OAI21X1 U792 ( .A(n3738), .B(n3671), .C(n2116), .Y(n1464) );
  OAI21X1 U794 ( .A(n3739), .B(n3671), .C(n2267), .Y(n1465) );
  OAI21X1 U796 ( .A(n3740), .B(n3671), .C(n2185), .Y(n1466) );
  OAI21X1 U798 ( .A(n3741), .B(n3671), .C(n2160), .Y(n1467) );
  OAI21X1 U800 ( .A(n3742), .B(n3671), .C(n2241), .Y(n1468) );
  OAI21X1 U802 ( .A(n3743), .B(n3671), .C(n2211), .Y(n1469) );
  OAI21X1 U805 ( .A(n3712), .B(n3670), .C(n2414), .Y(n1470) );
  OAI21X1 U807 ( .A(n3713), .B(n3670), .C(n2043), .Y(n1471) );
  OAI21X1 U809 ( .A(n3714), .B(n3670), .C(n2153), .Y(n1472) );
  OAI21X1 U811 ( .A(n3715), .B(n3670), .C(n2234), .Y(n1473) );
  OAI21X1 U813 ( .A(n3716), .B(n3670), .C(n2178), .Y(n1474) );
  OAI21X1 U815 ( .A(n3717), .B(n3670), .C(n2205), .Y(n1475) );
  OAI21X1 U817 ( .A(n3718), .B(n3670), .C(n2349), .Y(n1476) );
  OAI21X1 U819 ( .A(n3719), .B(n3670), .C(n2415), .Y(n1477) );
  OAI21X1 U821 ( .A(n3720), .B(n3670), .C(n2543), .Y(n1478) );
  OAI21X1 U823 ( .A(n3721), .B(n3670), .C(n2446), .Y(n1479) );
  OAI21X1 U825 ( .A(n3722), .B(n3670), .C(n2318), .Y(n1480) );
  OAI21X1 U827 ( .A(n3723), .B(n3670), .C(n2042), .Y(n1481) );
  OAI21X1 U829 ( .A(n3724), .B(n3670), .C(n2861), .Y(n1482) );
  OAI21X1 U831 ( .A(n3725), .B(n3670), .C(n2380), .Y(n1483) );
  OAI21X1 U833 ( .A(n3726), .B(n3670), .C(n2041), .Y(n1484) );
  OAI21X1 U835 ( .A(n3727), .B(n3670), .C(n2544), .Y(n1485) );
  OAI21X1 U837 ( .A(n3728), .B(n3670), .C(n2040), .Y(n1486) );
  OAI21X1 U839 ( .A(n3729), .B(n3670), .C(n2447), .Y(n1487) );
  OAI21X1 U841 ( .A(n3730), .B(n3670), .C(n2319), .Y(n1488) );
  OAI21X1 U843 ( .A(n3731), .B(n3670), .C(n2039), .Y(n1489) );
  OAI21X1 U845 ( .A(n3732), .B(n3670), .C(n2038), .Y(n1490) );
  OAI21X1 U847 ( .A(n3733), .B(n3670), .C(n2862), .Y(n1491) );
  OAI21X1 U849 ( .A(n3734), .B(n3670), .C(n2108), .Y(n1492) );
  OAI21X1 U851 ( .A(n3735), .B(n3670), .C(n2037), .Y(n1493) );
  OAI21X1 U853 ( .A(n3736), .B(n3670), .C(n2130), .Y(n1494) );
  OAI21X1 U855 ( .A(n3737), .B(n3670), .C(n2154), .Y(n1495) );
  OAI21X1 U857 ( .A(n3738), .B(n3670), .C(n2235), .Y(n1496) );
  OAI21X1 U859 ( .A(n3739), .B(n3670), .C(n2179), .Y(n1497) );
  OAI21X1 U861 ( .A(n3740), .B(n3670), .C(n2036), .Y(n1498) );
  OAI21X1 U863 ( .A(n3741), .B(n3670), .C(n2035), .Y(n1499) );
  OAI21X1 U865 ( .A(n3742), .B(n3670), .C(n2109), .Y(n1500) );
  OAI21X1 U867 ( .A(n3743), .B(n3670), .C(n2131), .Y(n1501) );
  OAI21X1 U870 ( .A(n3712), .B(n3669), .C(n2034), .Y(n1502) );
  OAI21X1 U872 ( .A(n3713), .B(n3669), .C(n2551), .Y(n1503) );
  OAI21X1 U874 ( .A(n3714), .B(n3669), .C(n2387), .Y(n1504) );
  OAI21X1 U876 ( .A(n3715), .B(n3669), .C(n2138), .Y(n1505) );
  OAI21X1 U878 ( .A(n3716), .B(n3669), .C(n2293), .Y(n1506) );
  OAI21X1 U880 ( .A(n3717), .B(n3669), .C(n2033), .Y(n1507) );
  OAI21X1 U882 ( .A(n3718), .B(n3669), .C(n2032), .Y(n1508) );
  OAI21X1 U884 ( .A(n3719), .B(n3669), .C(n2031), .Y(n1509) );
  OAI21X1 U886 ( .A(n3720), .B(n3669), .C(n2324), .Y(n1510) );
  OAI21X1 U888 ( .A(n3721), .B(n3669), .C(n2355), .Y(n1511) );
  OAI21X1 U890 ( .A(n3722), .B(n3669), .C(n2421), .Y(n1512) );
  OAI21X1 U892 ( .A(n3723), .B(n3669), .C(n2454), .Y(n1513) );
  OAI21X1 U894 ( .A(n3724), .B(n3669), .C(n2639), .Y(n1514) );
  OAI21X1 U896 ( .A(n3725), .B(n3669), .C(n2268), .Y(n1515) );
  OAI21X1 U898 ( .A(n3726), .B(n3669), .C(n2552), .Y(n1516) );
  OAI21X1 U900 ( .A(n3727), .B(n3669), .C(n2325), .Y(n1517) );
  OAI21X1 U902 ( .A(n3728), .B(n3669), .C(n2161), .Y(n1518) );
  OAI21X1 U904 ( .A(n3729), .B(n3669), .C(n2356), .Y(n1519) );
  OAI21X1 U906 ( .A(n3730), .B(n3669), .C(n2422), .Y(n1520) );
  OAI21X1 U908 ( .A(n3731), .B(n3669), .C(n2186), .Y(n1521) );
  OAI21X1 U910 ( .A(n3732), .B(n3669), .C(n2455), .Y(n1522) );
  OAI21X1 U912 ( .A(n3733), .B(n3669), .C(n2640), .Y(n1523) );
  OAI21X1 U914 ( .A(n3734), .B(n3669), .C(n2212), .Y(n1524) );
  OAI21X1 U916 ( .A(n3735), .B(n3669), .C(n2553), .Y(n1525) );
  OAI21X1 U918 ( .A(n3736), .B(n3669), .C(n2242), .Y(n1526) );
  OAI21X1 U920 ( .A(n3737), .B(n3669), .C(n2388), .Y(n1527) );
  OAI21X1 U922 ( .A(n3738), .B(n3669), .C(n2139), .Y(n1528) );
  OAI21X1 U924 ( .A(n3739), .B(n3669), .C(n2294), .Y(n1529) );
  OAI21X1 U926 ( .A(n3740), .B(n3669), .C(n2162), .Y(n1530) );
  OAI21X1 U928 ( .A(n3741), .B(n3669), .C(n2187), .Y(n1531) );
  OAI21X1 U930 ( .A(n3742), .B(n3669), .C(n2213), .Y(n1532) );
  OAI21X1 U932 ( .A(n3743), .B(n3669), .C(n2243), .Y(n1533) );
  OAI21X1 U935 ( .A(n3712), .B(n3668), .C(n2381), .Y(n1534) );
  OAI21X1 U937 ( .A(n3713), .B(n3668), .C(n2863), .Y(n1535) );
  OAI21X1 U939 ( .A(n3714), .B(n3668), .C(n2030), .Y(n1536) );
  OAI21X1 U941 ( .A(n3715), .B(n3668), .C(n2029), .Y(n1537) );
  OAI21X1 U943 ( .A(n3716), .B(n3668), .C(n2110), .Y(n1538) );
  OAI21X1 U945 ( .A(n3717), .B(n3668), .C(n2264), .Y(n1539) );
  OAI21X1 U947 ( .A(n3718), .B(n3668), .C(n2320), .Y(n1540) );
  OAI21X1 U949 ( .A(n3719), .B(n3668), .C(n2382), .Y(n1541) );
  OAI21X1 U951 ( .A(n3720), .B(n3668), .C(n2448), .Y(n1542) );
  OAI21X1 U953 ( .A(n3721), .B(n3668), .C(n2545), .Y(n1543) );
  OAI21X1 U955 ( .A(n3722), .B(n3668), .C(n2350), .Y(n1544) );
  OAI21X1 U957 ( .A(n3723), .B(n3668), .C(n2028), .Y(n1545) );
  OAI21X1 U959 ( .A(n3724), .B(n3668), .C(n2132), .Y(n1546) );
  OAI21X1 U961 ( .A(n3725), .B(n3668), .C(n2416), .Y(n1547) );
  OAI21X1 U963 ( .A(n3726), .B(n3668), .C(n2864), .Y(n1548) );
  OAI21X1 U965 ( .A(n3727), .B(n3668), .C(n2449), .Y(n1549) );
  OAI21X1 U967 ( .A(n3728), .B(n3668), .C(n2236), .Y(n1550) );
  OAI21X1 U969 ( .A(n3729), .B(n3668), .C(n2546), .Y(n1551) );
  OAI21X1 U971 ( .A(n3730), .B(n3668), .C(n2351), .Y(n1552) );
  OAI21X1 U973 ( .A(n3731), .B(n3668), .C(n2206), .Y(n1553) );
  OAI21X1 U975 ( .A(n3732), .B(n3668), .C(n2027), .Y(n1554) );
  OAI21X1 U977 ( .A(n3733), .B(n3668), .C(n2133), .Y(n1555) );
  OAI21X1 U979 ( .A(n3734), .B(n3668), .C(n2180), .Y(n1556) );
  OAI21X1 U981 ( .A(n3735), .B(n3668), .C(n2865), .Y(n1557) );
  OAI21X1 U983 ( .A(n3736), .B(n3668), .C(n2155), .Y(n1558) );
  OAI21X1 U985 ( .A(n3737), .B(n3668), .C(n2026), .Y(n1559) );
  OAI21X1 U987 ( .A(n3738), .B(n3668), .C(n2025), .Y(n1560) );
  OAI21X1 U989 ( .A(n3739), .B(n3668), .C(n2111), .Y(n1561) );
  OAI21X1 U991 ( .A(n3740), .B(n3668), .C(n2237), .Y(n1562) );
  OAI21X1 U993 ( .A(n3741), .B(n3668), .C(n2207), .Y(n1563) );
  OAI21X1 U995 ( .A(n3742), .B(n3668), .C(n2181), .Y(n1564) );
  OAI21X1 U997 ( .A(n3743), .B(n3668), .C(n2156), .Y(n1565) );
  OAI21X1 U1000 ( .A(n3712), .B(n3667), .C(n2244), .Y(n1566) );
  OAI21X1 U1002 ( .A(n3713), .B(n3667), .C(n2641), .Y(n1567) );
  OAI21X1 U1004 ( .A(n3714), .B(n3667), .C(n2423), .Y(n1568) );
  OAI21X1 U1006 ( .A(n3715), .B(n3667), .C(n2456), .Y(n1569) );
  OAI21X1 U1008 ( .A(n3716), .B(n3667), .C(n2214), .Y(n1570) );
  OAI21X1 U1010 ( .A(n3717), .B(n3667), .C(n2024), .Y(n1571) );
  OAI21X1 U1012 ( .A(n3718), .B(n3667), .C(n2023), .Y(n1572) );
  OAI21X1 U1014 ( .A(n3719), .B(n3667), .C(n2245), .Y(n1573) );
  OAI21X1 U1016 ( .A(n3720), .B(n3667), .C(n2022), .Y(n1574) );
  OAI21X1 U1018 ( .A(n3721), .B(n3667), .C(n2021), .Y(n1575) );
  OAI21X1 U1020 ( .A(n3722), .B(n3667), .C(n2020), .Y(n1576) );
  OAI21X1 U1022 ( .A(n3723), .B(n3667), .C(n2389), .Y(n1577) );
  OAI21X1 U1024 ( .A(n3724), .B(n3667), .C(n2554), .Y(n1578) );
  OAI21X1 U1026 ( .A(n3725), .B(n3667), .C(n2019), .Y(n1579) );
  OAI21X1 U1028 ( .A(n3726), .B(n3667), .C(n2642), .Y(n1580) );
  OAI21X1 U1030 ( .A(n3727), .B(n3667), .C(n2018), .Y(n1581) );
  OAI21X1 U1032 ( .A(n3728), .B(n3667), .C(n2357), .Y(n1582) );
  OAI21X1 U1034 ( .A(n3729), .B(n3667), .C(n2017), .Y(n1583) );
  OAI21X1 U1036 ( .A(n3730), .B(n3667), .C(n2016), .Y(n1584) );
  OAI21X1 U1038 ( .A(n3731), .B(n3667), .C(n2326), .Y(n1585) );
  OAI21X1 U1040 ( .A(n3732), .B(n3667), .C(n2390), .Y(n1586) );
  OAI21X1 U1042 ( .A(n3733), .B(n3667), .C(n2555), .Y(n1587) );
  OAI21X1 U1044 ( .A(n3734), .B(n3667), .C(n2295), .Y(n1588) );
  OAI21X1 U1046 ( .A(n3735), .B(n3667), .C(n2643), .Y(n1589) );
  OAI21X1 U1048 ( .A(n3736), .B(n3667), .C(n2269), .Y(n1590) );
  OAI21X1 U1050 ( .A(n3737), .B(n3667), .C(n2424), .Y(n1591) );
  OAI21X1 U1052 ( .A(n3738), .B(n3667), .C(n2457), .Y(n1592) );
  OAI21X1 U1054 ( .A(n3739), .B(n3667), .C(n2215), .Y(n1593) );
  OAI21X1 U1056 ( .A(n3740), .B(n3667), .C(n2358), .Y(n1594) );
  OAI21X1 U1058 ( .A(n3741), .B(n3667), .C(n2327), .Y(n1595) );
  OAI21X1 U1060 ( .A(n3742), .B(n3667), .C(n2296), .Y(n1596) );
  OAI21X1 U1062 ( .A(n3743), .B(n3667), .C(n2270), .Y(n1597) );
  OAI21X1 U1065 ( .A(n3712), .B(n3666), .C(n2352), .Y(n1598) );
  OAI21X1 U1067 ( .A(n3713), .B(n3666), .C(n2112), .Y(n1599) );
  OAI21X1 U1069 ( .A(n3714), .B(n3666), .C(n2866), .Y(n1600) );
  OAI21X1 U1071 ( .A(n3715), .B(n3666), .C(n2015), .Y(n1601) );
  OAI21X1 U1073 ( .A(n3716), .B(n3666), .C(n2134), .Y(n1602) );
  OAI21X1 U1075 ( .A(n3717), .B(n3666), .C(n2291), .Y(n1603) );
  OAI21X1 U1077 ( .A(n3718), .B(n3666), .C(n2265), .Y(n1604) );
  OAI21X1 U1079 ( .A(n3719), .B(n3666), .C(n2353), .Y(n1605) );
  OAI21X1 U1081 ( .A(n3720), .B(n3666), .C(n2417), .Y(n1606) );
  OAI21X1 U1083 ( .A(n3721), .B(n3666), .C(n2383), .Y(n1607) );
  OAI21X1 U1085 ( .A(n3722), .B(n3666), .C(n2450), .Y(n1608) );
  OAI21X1 U1087 ( .A(n3723), .B(n3666), .C(n2547), .Y(n1609) );
  OAI21X1 U1089 ( .A(n3724), .B(n3666), .C(n2014), .Y(n1610) );
  OAI21X1 U1091 ( .A(n3725), .B(n3666), .C(n2321), .Y(n1611) );
  OAI21X1 U1093 ( .A(n3726), .B(n3666), .C(n2113), .Y(n1612) );
  OAI21X1 U1095 ( .A(n3727), .B(n3666), .C(n2418), .Y(n1613) );
  OAI21X1 U1097 ( .A(n3728), .B(n3666), .C(n2208), .Y(n1614) );
  OAI21X1 U1099 ( .A(n3729), .B(n3666), .C(n2384), .Y(n1615) );
  OAI21X1 U1101 ( .A(n3730), .B(n3666), .C(n2451), .Y(n1616) );
  OAI21X1 U1103 ( .A(n3731), .B(n3666), .C(n2238), .Y(n1617) );
  OAI21X1 U1105 ( .A(n3732), .B(n3666), .C(n2548), .Y(n1618) );
  OAI21X1 U1107 ( .A(n3733), .B(n3666), .C(n2013), .Y(n1619) );
  OAI21X1 U1109 ( .A(n3734), .B(n3666), .C(n2157), .Y(n1620) );
  OAI21X1 U1111 ( .A(n3735), .B(n3666), .C(n2114), .Y(n1621) );
  OAI21X1 U1113 ( .A(n3736), .B(n3666), .C(n2182), .Y(n1622) );
  OAI21X1 U1115 ( .A(n3737), .B(n3666), .C(n2867), .Y(n1623) );
  OAI21X1 U1117 ( .A(n3738), .B(n3666), .C(n2012), .Y(n1624) );
  OAI21X1 U1119 ( .A(n3739), .B(n3666), .C(n2135), .Y(n1625) );
  OAI21X1 U1121 ( .A(n3740), .B(n3666), .C(n2209), .Y(n1626) );
  OAI21X1 U1123 ( .A(n3741), .B(n3666), .C(n2239), .Y(n1627) );
  OAI21X1 U1125 ( .A(n3742), .B(n3666), .C(n2158), .Y(n1628) );
  OAI21X1 U1127 ( .A(n3743), .B(n3666), .C(n2183), .Y(n1629) );
  OAI21X1 U1130 ( .A(n3712), .B(n3665), .C(n2216), .Y(n1630) );
  OAI21X1 U1132 ( .A(n3713), .B(n3665), .C(n2458), .Y(n1631) );
  OAI21X1 U1134 ( .A(n3714), .B(n3665), .C(n2644), .Y(n1632) );
  OAI21X1 U1136 ( .A(n3715), .B(n3665), .C(n2556), .Y(n1633) );
  OAI21X1 U1138 ( .A(n3716), .B(n3665), .C(n2246), .Y(n1634) );
  OAI21X1 U1140 ( .A(n3717), .B(n3665), .C(n2011), .Y(n1635) );
  OAI21X1 U1142 ( .A(n3718), .B(n3665), .C(n2010), .Y(n1636) );
  OAI21X1 U1144 ( .A(n3719), .B(n3665), .C(n2217), .Y(n1637) );
  OAI21X1 U1146 ( .A(n3720), .B(n3665), .C(n2009), .Y(n1638) );
  OAI21X1 U1148 ( .A(n3721), .B(n3665), .C(n2008), .Y(n1639) );
  OAI21X1 U1150 ( .A(n3722), .B(n3665), .C(n2391), .Y(n1640) );
  OAI21X1 U1152 ( .A(n3723), .B(n3665), .C(n2425), .Y(n1641) );
  OAI21X1 U1154 ( .A(n3724), .B(n3665), .C(n2188), .Y(n1642) );
  OAI21X1 U1156 ( .A(n3725), .B(n3665), .C(n2007), .Y(n1643) );
  OAI21X1 U1158 ( .A(n3726), .B(n3665), .C(n2459), .Y(n1644) );
  OAI21X1 U1160 ( .A(n3727), .B(n3665), .C(n2006), .Y(n1645) );
  OAI21X1 U1162 ( .A(n3728), .B(n3665), .C(n2328), .Y(n1646) );
  OAI21X1 U1164 ( .A(n3729), .B(n3665), .C(n2005), .Y(n1647) );
  OAI21X1 U1166 ( .A(n3730), .B(n3665), .C(n2392), .Y(n1648) );
  OAI21X1 U1168 ( .A(n3731), .B(n3665), .C(n2359), .Y(n1649) );
  OAI21X1 U1170 ( .A(n3732), .B(n3665), .C(n2426), .Y(n1650) );
  OAI21X1 U1172 ( .A(n3733), .B(n3665), .C(n2189), .Y(n1651) );
  OAI21X1 U1174 ( .A(n3734), .B(n3665), .C(n2271), .Y(n1652) );
  OAI21X1 U1176 ( .A(n3735), .B(n3665), .C(n2460), .Y(n1653) );
  OAI21X1 U1178 ( .A(n3736), .B(n3665), .C(n2297), .Y(n1654) );
  OAI21X1 U1180 ( .A(n3737), .B(n3665), .C(n2645), .Y(n1655) );
  OAI21X1 U1182 ( .A(n3738), .B(n3665), .C(n2557), .Y(n1656) );
  OAI21X1 U1184 ( .A(n3739), .B(n3665), .C(n2247), .Y(n1657) );
  OAI21X1 U1186 ( .A(n3740), .B(n3665), .C(n2329), .Y(n1658) );
  OAI21X1 U1188 ( .A(n3741), .B(n3665), .C(n2360), .Y(n1659) );
  OAI21X1 U1190 ( .A(n3742), .B(n3665), .C(n2272), .Y(n1660) );
  OAI21X1 U1192 ( .A(n3743), .B(n3665), .C(n2298), .Y(n1661) );
  OAI21X1 U1195 ( .A(n3712), .B(n3664), .C(n2190), .Y(n1662) );
  OAI21X1 U1197 ( .A(n3713), .B(n3664), .C(n2393), .Y(n1663) );
  OAI21X1 U1199 ( .A(n3714), .B(n3664), .C(n2558), .Y(n1664) );
  OAI21X1 U1201 ( .A(n3715), .B(n3664), .C(n2868), .Y(n1665) );
  OAI21X1 U1203 ( .A(n3716), .B(n3664), .C(n2646), .Y(n1666) );
  OAI21X1 U1205 ( .A(n3717), .B(n3664), .C(n2191), .Y(n1667) );
  OAI21X1 U1207 ( .A(n3718), .B(n3664), .C(n2004), .Y(n1668) );
  OAI21X1 U1209 ( .A(n3719), .B(n3664), .C(n2003), .Y(n1669) );
  OAI21X1 U1211 ( .A(n3720), .B(n3664), .C(n2218), .Y(n1670) );
  OAI21X1 U1213 ( .A(n3721), .B(n3664), .C(n2002), .Y(n1671) );
  OAI21X1 U1215 ( .A(n3722), .B(n3664), .C(n2117), .Y(n1672) );
  OAI21X1 U1217 ( .A(n3723), .B(n3664), .C(n2163), .Y(n1673) );
  OAI21X1 U1219 ( .A(n3724), .B(n3664), .C(n2427), .Y(n1674) );
  OAI21X1 U1221 ( .A(n3725), .B(n3664), .C(n2248), .Y(n1675) );
  OAI21X1 U1223 ( .A(n3726), .B(n3664), .C(n2394), .Y(n1676) );
  OAI21X1 U1225 ( .A(n3727), .B(n3664), .C(n2219), .Y(n1677) );
  OAI21X1 U1227 ( .A(n3728), .B(n3664), .C(n2299), .Y(n1678) );
  OAI21X1 U1229 ( .A(n3729), .B(n3664), .C(n2001), .Y(n1679) );
  OAI21X1 U1231 ( .A(n3730), .B(n3664), .C(n2118), .Y(n1680) );
  OAI21X1 U1233 ( .A(n3731), .B(n3664), .C(n2273), .Y(n1681) );
  OAI21X1 U1235 ( .A(n3732), .B(n3664), .C(n2164), .Y(n1682) );
  OAI21X1 U1237 ( .A(n3733), .B(n3664), .C(n2428), .Y(n1683) );
  OAI21X1 U1239 ( .A(n3734), .B(n3664), .C(n2361), .Y(n1684) );
  OAI21X1 U1241 ( .A(n3735), .B(n3664), .C(n2395), .Y(n1685) );
  OAI21X1 U1243 ( .A(n3736), .B(n3664), .C(n2330), .Y(n1686) );
  OAI21X1 U1245 ( .A(n3737), .B(n3664), .C(n2559), .Y(n1687) );
  OAI21X1 U1247 ( .A(n3738), .B(n3664), .C(n2869), .Y(n1688) );
  OAI21X1 U1249 ( .A(n3739), .B(n3664), .C(n2647), .Y(n1689) );
  OAI21X1 U1251 ( .A(n3740), .B(n3664), .C(n2300), .Y(n1690) );
  OAI21X1 U1253 ( .A(n3741), .B(n3664), .C(n2274), .Y(n1691) );
  OAI21X1 U1255 ( .A(n3742), .B(n3664), .C(n2362), .Y(n1692) );
  OAI21X1 U1257 ( .A(n3743), .B(n3664), .C(n2331), .Y(n1693) );
  OAI21X1 U1260 ( .A(n3712), .B(n3663), .C(n2145), .Y(n1694) );
  OAI21X1 U1262 ( .A(n3713), .B(n3663), .C(n2369), .Y(n1695) );
  OAI21X1 U1264 ( .A(n3714), .B(n3663), .C(n2281), .Y(n1696) );
  OAI21X1 U1266 ( .A(n3715), .B(n3663), .C(n2436), .Y(n1697) );
  OAI21X1 U1268 ( .A(n3716), .B(n3663), .C(n2338), .Y(n1698) );
  OAI21X1 U1270 ( .A(n3717), .B(n3663), .C(n2000), .Y(n1699) );
  OAI21X1 U1272 ( .A(n3718), .B(n3663), .C(n2146), .Y(n1700) );
  OAI21X1 U1274 ( .A(n3719), .B(n3663), .C(n1999), .Y(n1701) );
  OAI21X1 U1276 ( .A(n3720), .B(n3663), .C(n2122), .Y(n1702) );
  OAI21X1 U1278 ( .A(n3721), .B(n3663), .C(n2256), .Y(n1703) );
  OAI21X1 U1280 ( .A(n3722), .B(n3663), .C(n2169), .Y(n1704) );
  OAI21X1 U1282 ( .A(n3723), .B(n3663), .C(n2307), .Y(n1705) );
  OAI21X1 U1284 ( .A(n3724), .B(n3663), .C(n2226), .Y(n1706) );
  OAI21X1 U1286 ( .A(n3725), .B(n3663), .C(n2196), .Y(n1707) );
  OAI21X1 U1288 ( .A(n3726), .B(n3663), .C(n2370), .Y(n1708) );
  OAI21X1 U1290 ( .A(n3727), .B(n3663), .C(n2123), .Y(n1709) );
  OAI21X1 U1292 ( .A(n3728), .B(n3663), .C(n2563), .Y(n1710) );
  OAI21X1 U1294 ( .A(n3729), .B(n3663), .C(n2257), .Y(n1711) );
  OAI21X1 U1296 ( .A(n3730), .B(n3663), .C(n2170), .Y(n1712) );
  OAI21X1 U1298 ( .A(n3731), .B(n3663), .C(n2402), .Y(n1713) );
  OAI21X1 U1300 ( .A(n3732), .B(n3663), .C(n2308), .Y(n1714) );
  OAI21X1 U1302 ( .A(n3733), .B(n3663), .C(n2227), .Y(n1715) );
  OAI21X1 U1304 ( .A(n3734), .B(n3663), .C(n2876), .Y(n1716) );
  OAI21X1 U1306 ( .A(n3735), .B(n3663), .C(n2371), .Y(n1717) );
  OAI21X1 U1308 ( .A(n3736), .B(n3663), .C(n2466), .Y(n1718) );
  OAI21X1 U1310 ( .A(n3737), .B(n3663), .C(n2282), .Y(n1719) );
  OAI21X1 U1312 ( .A(n3738), .B(n3663), .C(n2437), .Y(n1720) );
  OAI21X1 U1314 ( .A(n3739), .B(n3663), .C(n2339), .Y(n1721) );
  OAI21X1 U1316 ( .A(n3740), .B(n3663), .C(n2564), .Y(n1722) );
  OAI21X1 U1318 ( .A(n3741), .B(n3663), .C(n2403), .Y(n1723) );
  OAI21X1 U1320 ( .A(n3742), .B(n3663), .C(n2877), .Y(n1724) );
  OAI21X1 U1322 ( .A(n3743), .B(n3663), .C(n2467), .Y(n1725) );
  OAI21X1 U1326 ( .A(n3712), .B(n3662), .C(n2165), .Y(n1726) );
  OAI21X1 U1328 ( .A(n3713), .B(n3662), .C(n2429), .Y(n1727) );
  OAI21X1 U1330 ( .A(n3714), .B(n3662), .C(n2461), .Y(n1728) );
  OAI21X1 U1332 ( .A(n3715), .B(n3662), .C(n2648), .Y(n1729) );
  OAI21X1 U1334 ( .A(n3716), .B(n3662), .C(n2870), .Y(n1730) );
  OAI21X1 U1336 ( .A(n3717), .B(n3662), .C(n2166), .Y(n1731) );
  OAI21X1 U1338 ( .A(n3718), .B(n3662), .C(n1998), .Y(n1732) );
  OAI21X1 U1340 ( .A(n3719), .B(n3662), .C(n1997), .Y(n1733) );
  OAI21X1 U1342 ( .A(n3720), .B(n3662), .C(n2249), .Y(n1734) );
  OAI21X1 U1344 ( .A(n3721), .B(n3662), .C(n1996), .Y(n1735) );
  OAI21X1 U1346 ( .A(n3722), .B(n3662), .C(n2140), .Y(n1736) );
  OAI21X1 U1348 ( .A(n3723), .B(n3662), .C(n2192), .Y(n1737) );
  OAI21X1 U1350 ( .A(n3724), .B(n3662), .C(n2396), .Y(n1738) );
  OAI21X1 U1352 ( .A(n3725), .B(n3662), .C(n2220), .Y(n1739) );
  OAI21X1 U1354 ( .A(n3726), .B(n3662), .C(n2430), .Y(n1740) );
  OAI21X1 U1356 ( .A(n3727), .B(n3662), .C(n2250), .Y(n1741) );
  OAI21X1 U1358 ( .A(n3728), .B(n3662), .C(n2275), .Y(n1742) );
  OAI21X1 U1360 ( .A(n3729), .B(n3662), .C(n1995), .Y(n1743) );
  OAI21X1 U1362 ( .A(n3730), .B(n3662), .C(n2141), .Y(n1744) );
  OAI21X1 U1364 ( .A(n3731), .B(n3662), .C(n2301), .Y(n1745) );
  OAI21X1 U1366 ( .A(n3732), .B(n3662), .C(n2193), .Y(n1746) );
  OAI21X1 U1368 ( .A(n3733), .B(n3662), .C(n2397), .Y(n1747) );
  OAI21X1 U1370 ( .A(n3734), .B(n3662), .C(n2332), .Y(n1748) );
  OAI21X1 U1372 ( .A(n3735), .B(n3662), .C(n2431), .Y(n1749) );
  OAI21X1 U1374 ( .A(n3736), .B(n3662), .C(n2363), .Y(n1750) );
  OAI21X1 U1376 ( .A(n3737), .B(n3662), .C(n2462), .Y(n1751) );
  OAI21X1 U1378 ( .A(n3738), .B(n3662), .C(n2649), .Y(n1752) );
  OAI21X1 U1380 ( .A(n3739), .B(n3662), .C(n2871), .Y(n1753) );
  OAI21X1 U1382 ( .A(n3740), .B(n3662), .C(n2276), .Y(n1754) );
  OAI21X1 U1384 ( .A(n3741), .B(n3662), .C(n2302), .Y(n1755) );
  OAI21X1 U1386 ( .A(n3742), .B(n3662), .C(n2333), .Y(n1756) );
  OAI21X1 U1388 ( .A(n3743), .B(n3662), .C(n2364), .Y(n1757) );
  OAI21X1 U1391 ( .A(n3712), .B(n3661), .C(n1994), .Y(n1758) );
  OAI21X1 U1393 ( .A(n3713), .B(n3661), .C(n2340), .Y(n1759) );
  OAI21X1 U1395 ( .A(n3714), .B(n3661), .C(n2309), .Y(n1760) );
  OAI21X1 U1397 ( .A(n3715), .B(n3661), .C(n2404), .Y(n1761) );
  OAI21X1 U1399 ( .A(n3716), .B(n3661), .C(n2372), .Y(n1762) );
  OAI21X1 U1401 ( .A(n3717), .B(n3661), .C(n1993), .Y(n1763) );
  OAI21X1 U1403 ( .A(n3718), .B(n3661), .C(n2124), .Y(n1764) );
  OAI21X1 U1405 ( .A(n3719), .B(n3661), .C(n1992), .Y(n1765) );
  OAI21X1 U1407 ( .A(n3720), .B(n3661), .C(n2147), .Y(n1766) );
  OAI21X1 U1409 ( .A(n3721), .B(n3661), .C(n2228), .Y(n1767) );
  OAI21X1 U1411 ( .A(n3722), .B(n3661), .C(n2197), .Y(n1768) );
  OAI21X1 U1413 ( .A(n3723), .B(n3661), .C(n2283), .Y(n1769) );
  OAI21X1 U1415 ( .A(n3724), .B(n3661), .C(n2258), .Y(n1770) );
  OAI21X1 U1417 ( .A(n3725), .B(n3661), .C(n2171), .Y(n1771) );
  OAI21X1 U1419 ( .A(n3726), .B(n3661), .C(n2341), .Y(n1772) );
  OAI21X1 U1421 ( .A(n3727), .B(n3661), .C(n2148), .Y(n1773) );
  OAI21X1 U1423 ( .A(n3728), .B(n3661), .C(n2468), .Y(n1774) );
  OAI21X1 U1425 ( .A(n3729), .B(n3661), .C(n2229), .Y(n1775) );
  OAI21X1 U1427 ( .A(n3730), .B(n3661), .C(n2198), .Y(n1776) );
  OAI21X1 U1429 ( .A(n3731), .B(n3661), .C(n2438), .Y(n1777) );
  OAI21X1 U1431 ( .A(n3732), .B(n3661), .C(n2284), .Y(n1778) );
  OAI21X1 U1433 ( .A(n3733), .B(n3661), .C(n2259), .Y(n1779) );
  OAI21X1 U1435 ( .A(n3734), .B(n3661), .C(n2654), .Y(n1780) );
  OAI21X1 U1437 ( .A(n3735), .B(n3661), .C(n2342), .Y(n1781) );
  OAI21X1 U1439 ( .A(n3736), .B(n3661), .C(n2565), .Y(n1782) );
  OAI21X1 U1441 ( .A(n3737), .B(n3661), .C(n2310), .Y(n1783) );
  OAI21X1 U1443 ( .A(n3738), .B(n3661), .C(n2405), .Y(n1784) );
  OAI21X1 U1445 ( .A(n3739), .B(n3661), .C(n2373), .Y(n1785) );
  OAI21X1 U1447 ( .A(n3740), .B(n3661), .C(n2469), .Y(n1786) );
  OAI21X1 U1449 ( .A(n3741), .B(n3661), .C(n2439), .Y(n1787) );
  OAI21X1 U1451 ( .A(n3742), .B(n3661), .C(n2655), .Y(n1788) );
  OAI21X1 U1453 ( .A(n3743), .B(n3661), .C(n2566), .Y(n1789) );
  OAI21X1 U1456 ( .A(n3712), .B(n3660), .C(n2463), .Y(n1790) );
  OAI21X1 U1458 ( .A(n3713), .B(n3660), .C(n2251), .Y(n1791) );
  OAI21X1 U1460 ( .A(n3714), .B(n3660), .C(n2221), .Y(n1792) );
  OAI21X1 U1462 ( .A(n3715), .B(n3660), .C(n2277), .Y(n1793) );
  OAI21X1 U1464 ( .A(n3716), .B(n3660), .C(n2560), .Y(n1794) );
  OAI21X1 U1466 ( .A(n3717), .B(n3660), .C(n2142), .Y(n1795) );
  OAI21X1 U1468 ( .A(n3718), .B(n3660), .C(n2194), .Y(n1796) );
  OAI21X1 U1470 ( .A(n3719), .B(n3660), .C(n2167), .Y(n1797) );
  OAI21X1 U1472 ( .A(n3720), .B(n3660), .C(n1991), .Y(n1798) );
  OAI21X1 U1474 ( .A(n3721), .B(n3660), .C(n2119), .Y(n1799) );
  OAI21X1 U1476 ( .A(n3722), .B(n3660), .C(n2303), .Y(n1800) );
  OAI21X1 U1478 ( .A(n3723), .B(n3660), .C(n2365), .Y(n1801) );
  OAI21X1 U1480 ( .A(n3724), .B(n3660), .C(n2334), .Y(n1802) );
  OAI21X1 U1482 ( .A(n3725), .B(n3660), .C(n1990), .Y(n1803) );
  OAI21X1 U1484 ( .A(n3726), .B(n3660), .C(n2252), .Y(n1804) );
  OAI21X1 U1486 ( .A(n3727), .B(n3660), .C(n1989), .Y(n1805) );
  OAI21X1 U1488 ( .A(n3728), .B(n3660), .C(n2872), .Y(n1806) );
  OAI21X1 U1490 ( .A(n3729), .B(n3660), .C(n2120), .Y(n1807) );
  OAI21X1 U1492 ( .A(n3730), .B(n3660), .C(n2304), .Y(n1808) );
  OAI21X1 U1494 ( .A(n3731), .B(n3660), .C(n2650), .Y(n1809) );
  OAI21X1 U1496 ( .A(n3732), .B(n3660), .C(n2366), .Y(n1810) );
  OAI21X1 U1498 ( .A(n3733), .B(n3660), .C(n2335), .Y(n1811) );
  OAI21X1 U1500 ( .A(n3734), .B(n3660), .C(n2432), .Y(n1812) );
  OAI21X1 U1502 ( .A(n3735), .B(n3660), .C(n2253), .Y(n1813) );
  OAI21X1 U1504 ( .A(n3736), .B(n3660), .C(n2398), .Y(n1814) );
  OAI21X1 U1506 ( .A(n3737), .B(n3660), .C(n2222), .Y(n1815) );
  OAI21X1 U1508 ( .A(n3738), .B(n3660), .C(n2278), .Y(n1816) );
  OAI21X1 U1510 ( .A(n3739), .B(n3660), .C(n2561), .Y(n1817) );
  OAI21X1 U1512 ( .A(n3740), .B(n3660), .C(n2873), .Y(n1818) );
  OAI21X1 U1514 ( .A(n3741), .B(n3660), .C(n2651), .Y(n1819) );
  OAI21X1 U1516 ( .A(n3742), .B(n3660), .C(n2433), .Y(n1820) );
  OAI21X1 U1518 ( .A(n3743), .B(n3660), .C(n2399), .Y(n1821) );
  OAI21X1 U1521 ( .A(n3712), .B(n3659), .C(n2656), .Y(n1822) );
  OAI21X1 U1523 ( .A(n3713), .B(n3659), .C(n2285), .Y(n1823) );
  OAI21X1 U1525 ( .A(n3714), .B(n3659), .C(n2374), .Y(n1824) );
  OAI21X1 U1527 ( .A(n3715), .B(n3659), .C(n2343), .Y(n1825) );
  OAI21X1 U1529 ( .A(n3716), .B(n3659), .C(n2440), .Y(n1826) );
  OAI21X1 U1531 ( .A(n3717), .B(n3659), .C(n1988), .Y(n1827) );
  OAI21X1 U1533 ( .A(n3718), .B(n3659), .C(n1987), .Y(n1828) );
  OAI21X1 U1535 ( .A(n3719), .B(n3659), .C(n2149), .Y(n1829) );
  OAI21X1 U1537 ( .A(n3720), .B(n3659), .C(n2199), .Y(n1830) );
  OAI21X1 U1539 ( .A(n3721), .B(n3659), .C(n2172), .Y(n1831) );
  OAI21X1 U1541 ( .A(n3722), .B(n3659), .C(n2260), .Y(n1832) );
  OAI21X1 U1543 ( .A(n3723), .B(n3659), .C(n2230), .Y(n1833) );
  OAI21X1 U1545 ( .A(n3724), .B(n3659), .C(n2311), .Y(n1834) );
  OAI21X1 U1547 ( .A(n3725), .B(n3659), .C(n2125), .Y(n1835) );
  OAI21X1 U1549 ( .A(n3726), .B(n3659), .C(n2286), .Y(n1836) );
  OAI21X1 U1551 ( .A(n3727), .B(n3659), .C(n2200), .Y(n1837) );
  OAI21X1 U1553 ( .A(n3728), .B(n3659), .C(n2406), .Y(n1838) );
  OAI21X1 U1555 ( .A(n3729), .B(n3659), .C(n2173), .Y(n1839) );
  OAI21X1 U1557 ( .A(n3730), .B(n3659), .C(n2261), .Y(n1840) );
  OAI21X1 U1559 ( .A(n3731), .B(n3659), .C(n2567), .Y(n1841) );
  OAI21X1 U1561 ( .A(n3732), .B(n3659), .C(n2231), .Y(n1842) );
  OAI21X1 U1563 ( .A(n3733), .B(n3659), .C(n2312), .Y(n1843) );
  OAI21X1 U1565 ( .A(n3734), .B(n3659), .C(n2470), .Y(n1844) );
  OAI21X1 U1567 ( .A(n3735), .B(n3659), .C(n2287), .Y(n1845) );
  OAI21X1 U1569 ( .A(n3736), .B(n3659), .C(n2878), .Y(n1846) );
  OAI21X1 U1571 ( .A(n3737), .B(n3659), .C(n2375), .Y(n1847) );
  OAI21X1 U1573 ( .A(n3738), .B(n3659), .C(n2344), .Y(n1848) );
  OAI21X1 U1575 ( .A(n3739), .B(n3659), .C(n2441), .Y(n1849) );
  OAI21X1 U1577 ( .A(n3740), .B(n3659), .C(n2407), .Y(n1850) );
  OAI21X1 U1579 ( .A(n3741), .B(n3659), .C(n2568), .Y(n1851) );
  OAI21X1 U1581 ( .A(n3742), .B(n3659), .C(n2471), .Y(n1852) );
  OAI21X1 U1583 ( .A(n3743), .B(n3659), .C(n2879), .Y(n1853) );
  OAI21X1 U1586 ( .A(n3712), .B(n3658), .C(n2562), .Y(n1854) );
  OAI21X1 U1588 ( .A(n3713), .B(n3658), .C(n2223), .Y(n1855) );
  OAI21X1 U1590 ( .A(n3714), .B(n3658), .C(n2254), .Y(n1856) );
  OAI21X1 U1592 ( .A(n3715), .B(n3658), .C(n2305), .Y(n1857) );
  OAI21X1 U1594 ( .A(n3716), .B(n3658), .C(n2464), .Y(n1858) );
  OAI21X1 U1596 ( .A(n3717), .B(n3658), .C(n2121), .Y(n1859) );
  OAI21X1 U1598 ( .A(n3718), .B(n3658), .C(n2168), .Y(n1860) );
  OAI21X1 U1600 ( .A(n3719), .B(n3658), .C(n2195), .Y(n1861) );
  OAI21X1 U1602 ( .A(n3720), .B(n3658), .C(n1986), .Y(n1862) );
  OAI21X1 U1604 ( .A(n3721), .B(n3658), .C(n2143), .Y(n1863) );
  OAI21X1 U1606 ( .A(n3722), .B(n3658), .C(n2279), .Y(n1864) );
  OAI21X1 U1608 ( .A(n3723), .B(n3658), .C(n2336), .Y(n1865) );
  OAI21X1 U1610 ( .A(n3724), .B(n3658), .C(n2367), .Y(n1866) );
  OAI21X1 U1612 ( .A(n3725), .B(n3658), .C(n1985), .Y(n1867) );
  OAI21X1 U1614 ( .A(n3726), .B(n3658), .C(n2224), .Y(n1868) );
  OAI21X1 U1616 ( .A(n3727), .B(n3658), .C(n1984), .Y(n1869) );
  OAI21X1 U1618 ( .A(n3728), .B(n3658), .C(n2652), .Y(n1870) );
  OAI21X1 U1620 ( .A(n3729), .B(n3658), .C(n2144), .Y(n1871) );
  OAI21X1 U1622 ( .A(n3730), .B(n3658), .C(n2280), .Y(n1872) );
  OAI21X1 U1624 ( .A(n3731), .B(n3658), .C(n2874), .Y(n1873) );
  OAI21X1 U1626 ( .A(n3732), .B(n3658), .C(n2337), .Y(n1874) );
  OAI21X1 U1628 ( .A(n3733), .B(n3658), .C(n2368), .Y(n1875) );
  OAI21X1 U1630 ( .A(n3734), .B(n3658), .C(n2400), .Y(n1876) );
  OAI21X1 U1632 ( .A(n3735), .B(n3658), .C(n2225), .Y(n1877) );
  OAI21X1 U1634 ( .A(n3736), .B(n3658), .C(n2434), .Y(n1878) );
  OAI21X1 U1636 ( .A(n3737), .B(n3658), .C(n2255), .Y(n1879) );
  OAI21X1 U1638 ( .A(n3738), .B(n3658), .C(n2306), .Y(n1880) );
  OAI21X1 U1640 ( .A(n3739), .B(n3658), .C(n2465), .Y(n1881) );
  OAI21X1 U1642 ( .A(n3740), .B(n3658), .C(n2653), .Y(n1882) );
  OAI21X1 U1644 ( .A(n3741), .B(n3658), .C(n2875), .Y(n1883) );
  OAI21X1 U1646 ( .A(n3742), .B(n3658), .C(n2401), .Y(n1884) );
  OAI21X1 U1648 ( .A(n3743), .B(n3658), .C(n2435), .Y(n1885) );
  OAI21X1 U1651 ( .A(n3712), .B(n3657), .C(n2126), .Y(n1886) );
  OAI21X1 U1653 ( .A(n3713), .B(n3657), .C(n2313), .Y(n1887) );
  OAI21X1 U1655 ( .A(n3714), .B(n3657), .C(n2345), .Y(n1888) );
  OAI21X1 U1657 ( .A(n3715), .B(n3657), .C(n2376), .Y(n1889) );
  OAI21X1 U1659 ( .A(n3716), .B(n3657), .C(n2408), .Y(n1890) );
  OAI21X1 U1661 ( .A(n3717), .B(n3657), .C(n1983), .Y(n1891) );
  OAI21X1 U1663 ( .A(n3718), .B(n3657), .C(n1982), .Y(n1892) );
  OAI21X1 U1665 ( .A(n3719), .B(n3657), .C(n2127), .Y(n1893) );
  OAI21X1 U1667 ( .A(n3720), .B(n3657), .C(n2174), .Y(n1894) );
  OAI21X1 U1669 ( .A(n3721), .B(n3657), .C(n2201), .Y(n1895) );
  OAI21X1 U1671 ( .A(n3722), .B(n3657), .C(n2232), .Y(n1896) );
  OAI21X1 U1673 ( .A(n3723), .B(n3657), .C(n2262), .Y(n1897) );
  OAI21X1 U1675 ( .A(n3724), .B(n3657), .C(n2288), .Y(n1898) );
  OAI21X1 U1677 ( .A(n3725), .B(n3657), .C(n2150), .Y(n1899) );
  OAI21X1 U1679 ( .A(n3726), .B(n3657), .C(n2314), .Y(n1900) );
  OAI21X1 U1681 ( .A(n3727), .B(n3657), .C(n2175), .Y(n1901) );
  OAI21X1 U1683 ( .A(n3728), .B(n3657), .C(n2442), .Y(n1902) );
  OAI21X1 U1685 ( .A(n3729), .B(n3657), .C(n2202), .Y(n1903) );
  OAI21X1 U1687 ( .A(n3730), .B(n3657), .C(n2233), .Y(n1904) );
  OAI21X1 U1689 ( .A(n3731), .B(n3657), .C(n2472), .Y(n1905) );
  OAI21X1 U1691 ( .A(n3732), .B(n3657), .C(n2263), .Y(n1906) );
  OAI21X1 U1693 ( .A(n3733), .B(n3657), .C(n2289), .Y(n1907) );
  OAI21X1 U1695 ( .A(n3734), .B(n3657), .C(n2569), .Y(n1908) );
  OAI21X1 U1697 ( .A(n3735), .B(n3657), .C(n2315), .Y(n1909) );
  OAI21X1 U1699 ( .A(n3736), .B(n3657), .C(n2657), .Y(n1910) );
  OAI21X1 U1701 ( .A(n3737), .B(n3657), .C(n2346), .Y(n1911) );
  OAI21X1 U1703 ( .A(n3738), .B(n3657), .C(n2377), .Y(n1912) );
  OAI21X1 U1705 ( .A(n3739), .B(n3657), .C(n2409), .Y(n1913) );
  OAI21X1 U1707 ( .A(n3740), .B(n3657), .C(n2443), .Y(n1914) );
  OAI21X1 U1709 ( .A(n3741), .B(n3657), .C(n2473), .Y(n1915) );
  OAI21X1 U1711 ( .A(n3742), .B(n3657), .C(n2570), .Y(n1916) );
  OAI21X1 U1713 ( .A(n3743), .B(n3657), .C(n2658), .Y(n1917) );
  OAI21X1 U1717 ( .A(n1084), .B(n3749), .C(n2541), .Y(n1918) );
  OAI21X1 U1719 ( .A(n1084), .B(n3748), .C(n2412), .Y(n1919) );
  OAI21X1 U1721 ( .A(n1084), .B(n3747), .C(n2411), .Y(n1920) );
  OAI21X1 U1723 ( .A(n1084), .B(n3746), .C(n2659), .Y(n1921) );
  OAI21X1 U1725 ( .A(n1084), .B(n3745), .C(n2378), .Y(n1922) );
  OAI21X1 U1727 ( .A(n1364), .B(n3673), .C(n2858), .Y(n1923) );
  OAI21X1 U1729 ( .A(n1364), .B(n3674), .C(n2636), .Y(n1924) );
  OAI21X1 U1731 ( .A(n1364), .B(n3675), .C(n2540), .Y(n1925) );
  OAI21X1 U1733 ( .A(n1364), .B(n3744), .C(n2410), .Y(n1926) );
  AOI22X1 U1735 ( .A(data_out[31]), .B(n3656), .C(n75), .D(n1364), .Y(n1363)
         );
  AOI22X1 U1736 ( .A(data_out[30]), .B(n3656), .C(n76), .D(n1364), .Y(n1365)
         );
  AOI22X1 U1737 ( .A(data_out[29]), .B(n3656), .C(n77), .D(n1364), .Y(n1366)
         );
  AOI22X1 U1738 ( .A(data_out[28]), .B(n3656), .C(n78), .D(n1364), .Y(n1367)
         );
  AOI22X1 U1739 ( .A(data_out[27]), .B(n3656), .C(n79), .D(n1364), .Y(n1368)
         );
  AOI22X1 U1740 ( .A(data_out[26]), .B(n3656), .C(n80), .D(n1364), .Y(n1369)
         );
  AOI22X1 U1741 ( .A(data_out[25]), .B(n3656), .C(n81), .D(n1364), .Y(n1370)
         );
  AOI22X1 U1742 ( .A(data_out[24]), .B(n3656), .C(n82), .D(n1364), .Y(n1371)
         );
  AOI22X1 U1743 ( .A(data_out[23]), .B(n3656), .C(n83), .D(n1364), .Y(n1372)
         );
  AOI22X1 U1744 ( .A(data_out[22]), .B(n3656), .C(n84), .D(n1364), .Y(n1373)
         );
  AOI22X1 U1745 ( .A(data_out[21]), .B(n3656), .C(n85), .D(n1364), .Y(n1374)
         );
  AOI22X1 U1746 ( .A(data_out[20]), .B(n3656), .C(n86), .D(n1364), .Y(n1375)
         );
  AOI22X1 U1747 ( .A(data_out[19]), .B(n3656), .C(n87), .D(n1364), .Y(n1376)
         );
  AOI22X1 U1748 ( .A(data_out[18]), .B(n3656), .C(n88), .D(n1364), .Y(n1377)
         );
  AOI22X1 U1749 ( .A(data_out[17]), .B(n3656), .C(n89), .D(n1364), .Y(n1378)
         );
  AOI22X1 U1750 ( .A(data_out[16]), .B(n3656), .C(n90), .D(n1364), .Y(n1379)
         );
  AOI22X1 U1751 ( .A(data_out[15]), .B(n3656), .C(n91), .D(n1364), .Y(n1380)
         );
  AOI22X1 U1752 ( .A(data_out[14]), .B(n3656), .C(n92), .D(n1364), .Y(n1381)
         );
  AOI22X1 U1753 ( .A(data_out[13]), .B(n3656), .C(n93), .D(n1364), .Y(n1382)
         );
  AOI22X1 U1754 ( .A(data_out[12]), .B(n3656), .C(n94), .D(n1364), .Y(n1383)
         );
  AOI22X1 U1755 ( .A(data_out[11]), .B(n3656), .C(n95), .D(n3655), .Y(n1384)
         );
  AOI22X1 U1756 ( .A(data_out[10]), .B(n3656), .C(n96), .D(n3655), .Y(n1385)
         );
  AOI22X1 U1757 ( .A(data_out[9]), .B(n3656), .C(n97), .D(n3655), .Y(n1386) );
  AOI22X1 U1758 ( .A(data_out[8]), .B(n3656), .C(n98), .D(n3655), .Y(n1387) );
  AOI22X1 U1759 ( .A(data_out[7]), .B(n3656), .C(n99), .D(n3655), .Y(n1388) );
  AOI22X1 U1760 ( .A(data_out[6]), .B(n3656), .C(n100), .D(n3655), .Y(n1389)
         );
  AOI22X1 U1761 ( .A(data_out[5]), .B(n3656), .C(n101), .D(n3655), .Y(n1390)
         );
  AOI22X1 U1762 ( .A(data_out[4]), .B(n3656), .C(n102), .D(n3655), .Y(n1391)
         );
  AOI22X1 U1763 ( .A(data_out[3]), .B(n3656), .C(n103), .D(n3655), .Y(n1392)
         );
  AOI22X1 U1764 ( .A(data_out[2]), .B(n3656), .C(n104), .D(n3655), .Y(n1393)
         );
  AOI22X1 U1765 ( .A(data_out[1]), .B(n3656), .C(n105), .D(n3655), .Y(n1394)
         );
  AOI22X1 U1766 ( .A(data_out[0]), .B(n3656), .C(n106), .D(n3655), .Y(n1395)
         );
  OAI21X1 U1767 ( .A(n1364), .B(n3564), .C(n2444), .Y(n1927) );
  XOR2X1 U1770 ( .A(n2856), .B(n3112), .Y(n26) );
  XOR2X1 U1771 ( .A(n3112), .B(n2857), .Y(n25) );
  XOR2X1 U1775 ( .A(n2635), .B(n3111), .Y(n23) );
  XOR2X1 U1776 ( .A(n3109), .B(n1932), .Y(n22) );
  XOR2X1 U1777 ( .A(n1932), .B(n1931), .Y(n21) );
  XOR2X1 U1778 ( .A(n1931), .B(n1930), .Y(n20) );
  XOR2X1 U1779 ( .A(n1930), .B(n3676), .Y(n19) );
  NAND3X1 U1780 ( .A(full_check[4]), .B(n1928), .C(n1397), .Y(n3751) );
  NOR3X1 U1781 ( .A(full_check[1]), .B(full_check[3]), .C(full_check[2]), .Y(
        n1397) );
  NAND3X1 U1782 ( .A(n3744), .B(n1399), .C(n1400), .Y(n3750) );
  NOR3X1 U1783 ( .A(n1401), .B(n1402), .C(n1403), .Y(n1400) );
  FAX1 U1784 ( .A(n2855), .B(n1931), .C(n3110), .YC(), .YS(n1403) );
  XOR2X1 U1785 ( .A(n1932), .B(n3110), .Y(n1402) );
  FAX1 U1786 ( .A(n3107), .B(n3676), .C(n1405), .YC(), .YS(n1401) );
  XOR2X1 U1787 ( .A(n1405), .B(n3675), .Y(n1399) );
  FAX1 U1788 ( .A(n2633), .B(n3110), .C(n2855), .YC(), .YS(n1405) );
  HAX1 add_169_U1_1_1 ( .A(n1930), .B(n3676), .YC(add_169_carry[2]), .YS(n108)
         );
  HAX1 add_169_U1_1_2 ( .A(n1931), .B(add_169_carry[2]), .YC(add_169_carry[3]), 
        .YS(n109) );
  HAX1 add_169_U1_1_3 ( .A(n1932), .B(add_169_carry[3]), .YC(add_169_carry[4]), 
        .YS(n110) );
  HAX1 add_148_U1_1_1 ( .A(n2635), .B(n3111), .YC(add_148_carry[2]), .YS(n36)
         );
  HAX1 add_148_U1_1_2 ( .A(n2857), .B(add_148_carry[2]), .YC(add_148_carry[3]), 
        .YS(n37) );
  HAX1 add_148_U1_1_3 ( .A(n3112), .B(add_148_carry[3]), .YC(add_148_carry[4]), 
        .YS(n38) );
  FAX1 sub_125_U2_1 ( .A(n2635), .B(n3678), .C(sub_125_carry[1]), .YC(
        sub_125_carry[2]), .YS(full_check[1]) );
  FAX1 sub_125_U2_2 ( .A(n2857), .B(n3113), .C(sub_125_carry[2]), .YC(
        sub_125_carry[3]), .YS(full_check[2]) );
  FAX1 sub_125_U2_3 ( .A(n3112), .B(n3677), .C(sub_125_carry[3]), .YC(
        sub_125_carry[4]), .YS(full_check[3]) );
  DFFSR wr_ptr_gray_ss_reg_3_ ( .D(n1969), .CLK(rclk), .R(n3595), .S(1'b1), 
        .Q(wr_ptr_gray_ss[3]) );
  DFFSR wr_ptr_gray_ss_reg_2_ ( .D(n1971), .CLK(rclk), .R(n3595), .S(1'b1), 
        .Q(wr_ptr_gray_ss[2]) );
  DFFSR wr_ptr_gray_ss_reg_1_ ( .D(n1973), .CLK(rclk), .R(n3595), .S(1'b1), 
        .Q(wr_ptr_gray_ss[1]) );
  DFFSR wr_ptr_gray_ss_reg_0_ ( .D(n1975), .CLK(rclk), .R(n3595), .S(1'b1), 
        .Q(wr_ptr_gray_ss[0]) );
  DFFSR rd_ptr_gray_reg_3_ ( .D(n22), .CLK(rclk), .R(n3595), .S(1'b1), .Q(
        rd_ptr_gray[3]) );
  DFFSR rd_ptr_gray_reg_0_ ( .D(n19), .CLK(rclk), .R(n3595), .S(1'b1), .Q(
        rd_ptr_gray[0]) );
  DFFSR rd_ptr_gray_reg_1_ ( .D(n20), .CLK(rclk), .R(n3595), .S(1'b1), .Q(
        rd_ptr_gray[1]) );
  DFFSR rd_ptr_gray_reg_2_ ( .D(n21), .CLK(rclk), .R(n3595), .S(1'b1), .Q(
        rd_ptr_gray[2]) );
  DFFSR rd_ptr_bin_reg_4_ ( .D(n1926), .CLK(rclk), .R(n3595), .S(1'b1), .Q(
        rd_ptr_bin_4_) );
  DFFSR rd_ptr_bin_reg_3_ ( .D(n1923), .CLK(rclk), .R(n3595), .S(1'b1), .Q(n17) );
  DFFSR rd_ptr_bin_reg_2_ ( .D(n1924), .CLK(rclk), .R(n3595), .S(1'b1), .Q(n16) );
  DFFSR rd_ptr_bin_reg_1_ ( .D(n1925), .CLK(rclk), .R(n3595), .S(1'b1), .Q(n15) );
  DFFSR rd_ptr_bin_reg_0_ ( .D(n1927), .CLK(rclk), .R(n3595), .S(1'b1), .Q(n14) );
  DFFSR data_out_reg_23_ ( .D(n3703), .CLK(rclk), .R(n3595), .S(1'b1), .Q(
        n3760) );
  DFFSR data_out_reg_22_ ( .D(n3702), .CLK(rclk), .R(n3595), .S(1'b1), .Q(
        n3761) );
  DFFSR data_out_reg_21_ ( .D(n3701), .CLK(rclk), .R(n3595), .S(1'b1), .Q(
        n3762) );
  DFFSR data_out_reg_20_ ( .D(n3700), .CLK(rclk), .R(n3595), .S(1'b1), .Q(
        n3763) );
  DFFSR data_out_reg_19_ ( .D(n3699), .CLK(rclk), .R(n3595), .S(1'b1), .Q(
        n3764) );
  DFFSR data_out_reg_18_ ( .D(n3698), .CLK(rclk), .R(n3595), .S(1'b1), .Q(
        n3765) );
  DFFSR data_out_reg_17_ ( .D(n3697), .CLK(rclk), .R(n3595), .S(1'b1), .Q(
        n3766) );
  DFFSR data_out_reg_16_ ( .D(n3696), .CLK(rclk), .R(n3595), .S(1'b1), .Q(
        n3767) );
  DFFSR data_out_reg_15_ ( .D(n3695), .CLK(rclk), .R(n3595), .S(1'b1), .Q(
        n3768) );
  DFFSR data_out_reg_14_ ( .D(n3694), .CLK(rclk), .R(n3595), .S(1'b1), .Q(
        n3769) );
  DFFSR data_out_reg_13_ ( .D(n3693), .CLK(rclk), .R(n3595), .S(1'b1), .Q(
        n3770) );
  DFFSR data_out_reg_12_ ( .D(n3692), .CLK(rclk), .R(n3595), .S(1'b1), .Q(
        n3771) );
  DFFSR data_out_reg_30_ ( .D(n3710), .CLK(rclk), .R(n3595), .S(1'b1), .Q(
        n3753) );
  DFFSR data_out_reg_29_ ( .D(n3709), .CLK(rclk), .R(n3595), .S(1'b1), .Q(
        n3754) );
  DFFSR data_out_reg_28_ ( .D(n3708), .CLK(rclk), .R(n3595), .S(1'b1), .Q(
        n3755) );
  DFFSR data_out_reg_27_ ( .D(n3707), .CLK(rclk), .R(n3595), .S(1'b1), .Q(
        n3756) );
  DFFSR data_out_reg_26_ ( .D(n3706), .CLK(rclk), .R(n3595), .S(1'b1), .Q(
        n3757) );
  DFFSR data_out_reg_25_ ( .D(n3705), .CLK(rclk), .R(n3595), .S(1'b1), .Q(
        n3758) );
  DFFSR data_out_reg_24_ ( .D(n3704), .CLK(rclk), .R(n3595), .S(1'b1), .Q(
        n3759) );
  DFFSR data_out_reg_31_ ( .D(n3711), .CLK(rclk), .R(n3595), .S(1'b1), .Q(
        n3752) );
  DFFSR data_out_reg_11_ ( .D(n3691), .CLK(rclk), .R(n3679), .S(1'b1), .Q(
        n3772) );
  DFFSR data_out_reg_10_ ( .D(n3690), .CLK(rclk), .R(n3679), .S(1'b1), .Q(
        n3773) );
  DFFSR data_out_reg_9_ ( .D(n3689), .CLK(rclk), .R(n3679), .S(1'b1), .Q(n3774) );
  DFFSR data_out_reg_8_ ( .D(n3688), .CLK(rclk), .R(n3679), .S(1'b1), .Q(n3775) );
  DFFSR data_out_reg_7_ ( .D(n3687), .CLK(rclk), .R(n3679), .S(1'b1), .Q(n3776) );
  DFFSR data_out_reg_6_ ( .D(n3686), .CLK(rclk), .R(n3679), .S(1'b1), .Q(n3777) );
  DFFSR data_out_reg_5_ ( .D(n3685), .CLK(rclk), .R(n3679), .S(1'b1), .Q(n3778) );
  DFFSR data_out_reg_4_ ( .D(n3684), .CLK(rclk), .R(n3679), .S(1'b1), .Q(n3779) );
  DFFSR data_out_reg_3_ ( .D(n3683), .CLK(rclk), .R(n3679), .S(1'b1), .Q(n3780) );
  DFFSR data_out_reg_2_ ( .D(n3682), .CLK(rclk), .R(n3679), .S(1'b1), .Q(n3781) );
  DFFSR data_out_reg_1_ ( .D(n3681), .CLK(rclk), .R(n3679), .S(1'b1), .Q(n3782) );
  DFFSR data_out_reg_0_ ( .D(n3680), .CLK(rclk), .R(n3679), .S(1'b1), .Q(n3783) );
  AND2X1 U1791 ( .A(n3112), .B(n1084), .Y(n1320) );
  OR2X1 U1792 ( .A(n3114), .B(n3111), .Y(sub_125_carry[1]) );
  AND2X1 U1793 ( .A(n2491), .B(n3659), .Y(n1285) );
  AND2X1 U1794 ( .A(n2490), .B(n3659), .Y(n1278) );
  AND2X1 U1795 ( .A(n2489), .B(n3663), .Y(n1150) );
  AND2X1 U1796 ( .A(n2488), .B(n3663), .Y(n1142) );
  AND2X1 U1797 ( .A(n2578), .B(n3658), .Y(n1317) );
  AND2X1 U1798 ( .A(n2577), .B(n3658), .Y(n1316) );
  AND2X1 U1799 ( .A(n2576), .B(n3658), .Y(n1307) );
  AND2X1 U1800 ( .A(n2575), .B(n3658), .Y(n1304) );
  AND2X1 U1801 ( .A(n2487), .B(n3660), .Y(n1250) );
  AND2X1 U1802 ( .A(n2486), .B(n3660), .Y(n1249) );
  AND2X1 U1803 ( .A(n2485), .B(n3660), .Y(n1248) );
  AND2X1 U1804 ( .A(n2484), .B(n3660), .Y(n1240) );
  AND2X1 U1805 ( .A(n2483), .B(n3660), .Y(n1237) );
  AND2X1 U1806 ( .A(n2482), .B(n3660), .Y(n1225) );
  AND2X1 U1807 ( .A(n2574), .B(n3662), .Y(n1181) );
  AND2X1 U1808 ( .A(n2573), .B(n3662), .Y(n1180) );
  AND2X1 U1809 ( .A(n2572), .B(n3662), .Y(n1158) );
  AND2X1 U1810 ( .A(n2571), .B(n3662), .Y(n1157) );
  AND2X1 U1811 ( .A(n2481), .B(n3664), .Y(n1113) );
  AND2X1 U1812 ( .A(n2480), .B(n3664), .Y(n1112) );
  AND2X1 U1813 ( .A(n2479), .B(n3664), .Y(n1111) );
  AND2X1 U1814 ( .A(n2478), .B(n3664), .Y(n1090) );
  AND2X1 U1815 ( .A(n2477), .B(n3664), .Y(n1089) );
  AND2X1 U1816 ( .A(n2476), .B(n3664), .Y(n1088) );
  AND2X1 U1817 ( .A(n2666), .B(n3666), .Y(n1042) );
  AND2X1 U1818 ( .A(n2665), .B(n3666), .Y(n1019) );
  AND2X1 U1819 ( .A(n2664), .B(n3668), .Y(n974) );
  AND2X1 U1820 ( .A(n2663), .B(n3668), .Y(n965) );
  AND2X1 U1821 ( .A(n2662), .B(n3668), .Y(n952) );
  AND2X1 U1822 ( .A(n2668), .B(n3670), .Y(n906) );
  AND2X1 U1823 ( .A(n2667), .B(n3670), .Y(n897) );
  AND2X1 U1824 ( .A(n2661), .B(n3672), .Y(n836) );
  AND2X1 U1825 ( .A(n2660), .B(n3672), .Y(n827) );
  XOR2X1 U1826 ( .A(n3111), .B(n3114), .Y(n1928) );
  BUFX2 U1827 ( .A(n14), .Y(n1929) );
  BUFX2 U1828 ( .A(n15), .Y(n1930) );
  BUFX2 U1829 ( .A(n16), .Y(n1931) );
  BUFX2 U1830 ( .A(n17), .Y(n1932) );
  BUFX2 U1831 ( .A(n1395), .Y(n1933) );
  BUFX2 U1832 ( .A(n1394), .Y(n1934) );
  BUFX2 U1833 ( .A(n1393), .Y(n1935) );
  BUFX2 U1834 ( .A(n1392), .Y(n1936) );
  BUFX2 U1835 ( .A(n1391), .Y(n1937) );
  BUFX2 U1836 ( .A(n1390), .Y(n1938) );
  BUFX2 U1837 ( .A(n1389), .Y(n1939) );
  BUFX2 U1838 ( .A(n1388), .Y(n1940) );
  BUFX2 U1839 ( .A(n1387), .Y(n1941) );
  BUFX2 U1840 ( .A(n1386), .Y(n1942) );
  BUFX2 U1841 ( .A(n1385), .Y(n1943) );
  BUFX2 U1842 ( .A(n1384), .Y(n1944) );
  BUFX2 U1843 ( .A(n1383), .Y(n1945) );
  BUFX2 U1844 ( .A(n1382), .Y(n1946) );
  BUFX2 U1845 ( .A(n1381), .Y(n1947) );
  BUFX2 U1846 ( .A(n1380), .Y(n1948) );
  BUFX2 U1847 ( .A(n1379), .Y(n1949) );
  BUFX2 U1848 ( .A(n1378), .Y(n1950) );
  BUFX2 U1849 ( .A(n1377), .Y(n1951) );
  BUFX2 U1850 ( .A(n1376), .Y(n1952) );
  BUFX2 U1851 ( .A(n1375), .Y(n1953) );
  BUFX2 U1852 ( .A(n1374), .Y(n1954) );
  BUFX2 U1853 ( .A(n1373), .Y(n1955) );
  BUFX2 U1854 ( .A(n1372), .Y(n1956) );
  BUFX2 U1855 ( .A(n1371), .Y(n1957) );
  BUFX2 U1856 ( .A(n1370), .Y(n1958) );
  BUFX2 U1857 ( .A(n1369), .Y(n1959) );
  BUFX2 U1858 ( .A(n1368), .Y(n1960) );
  BUFX2 U1859 ( .A(n1367), .Y(n1961) );
  BUFX2 U1860 ( .A(n1366), .Y(n1962) );
  BUFX2 U1861 ( .A(n1365), .Y(n1963) );
  BUFX2 U1862 ( .A(n1363), .Y(n1964) );
  AND2X1 U1863 ( .A(n1152), .B(n2539), .Y(n1321) );
  AND2X1 U1864 ( .A(n1118), .B(n2539), .Y(n1287) );
  AND2X1 U1865 ( .A(n1152), .B(n1286), .Y(n1253) );
  AND2X1 U1866 ( .A(n1118), .B(n1286), .Y(n1220) );
  AND2X1 U1867 ( .A(n1152), .B(n1219), .Y(n1186) );
  AND2X1 U1868 ( .A(n1152), .B(n2538), .Y(n1119) );
  AND2X1 U1869 ( .A(n1320), .B(n3111), .Y(n1152) );
  AND2X1 U1870 ( .A(n2539), .B(n849), .Y(n1016) );
  AND2X1 U1871 ( .A(n883), .B(n2538), .Y(n850) );
  BUFX2 U1872 ( .A(rd_ptr_gray[2]), .Y(n1965) );
  BUFX2 U1873 ( .A(rd_ptr_gray[1]), .Y(n1966) );
  BUFX2 U1874 ( .A(rd_ptr_gray[0]), .Y(n1967) );
  BUFX2 U1875 ( .A(rd_ptr_gray[3]), .Y(n1968) );
  BUFX2 U1876 ( .A(wr_ptr_gray_s[3]), .Y(n1969) );
  BUFX2 U1877 ( .A(wr_ptr_gray[3]), .Y(n1970) );
  BUFX2 U1878 ( .A(wr_ptr_gray_s[2]), .Y(n1971) );
  BUFX2 U1879 ( .A(wr_ptr_gray[2]), .Y(n1972) );
  BUFX2 U1880 ( .A(wr_ptr_gray_s[1]), .Y(n1973) );
  BUFX2 U1881 ( .A(wr_ptr_gray[1]), .Y(n1974) );
  BUFX2 U1882 ( .A(wr_ptr_gray_s[0]), .Y(n1975) );
  BUFX2 U1883 ( .A(wr_ptr_gray[0]), .Y(n1976) );
  BUFX2 U1884 ( .A(rd_ptr_gray_s[3]), .Y(n1977) );
  BUFX2 U1885 ( .A(rd_ptr_gray_s[2]), .Y(n1978) );
  BUFX2 U1886 ( .A(rd_ptr_gray_s[1]), .Y(n1979) );
  BUFX2 U1887 ( .A(rd_ptr_gray_s[0]), .Y(n1980) );
  AND2X1 U1888 ( .A(n2060), .B(n2059), .Y(n24) );
  INVX1 U1889 ( .A(n24), .Y(n1981) );
  AND2X1 U1890 ( .A(n3048), .B(n3657), .Y(n1328) );
  INVX1 U1891 ( .A(n1328), .Y(n1982) );
  AND2X1 U1892 ( .A(n3047), .B(n3657), .Y(n1327) );
  INVX1 U1893 ( .A(n1327), .Y(n1983) );
  AND2X1 U1894 ( .A(n2622), .B(n3658), .Y(n1303) );
  INVX1 U1895 ( .A(n1303), .Y(n1984) );
  AND2X1 U1896 ( .A(n2620), .B(n3658), .Y(n1301) );
  INVX1 U1897 ( .A(n1301), .Y(n1985) );
  AND2X1 U1898 ( .A(n2615), .B(n3658), .Y(n1296) );
  INVX1 U1899 ( .A(n1296), .Y(n1986) );
  AND2X1 U1900 ( .A(n2830), .B(n3659), .Y(n1260) );
  INVX1 U1901 ( .A(n1260), .Y(n1987) );
  AND2X1 U1902 ( .A(n2829), .B(n3659), .Y(n1259) );
  INVX1 U1903 ( .A(n1259), .Y(n1988) );
  AND2X1 U1904 ( .A(n2528), .B(n3660), .Y(n1236) );
  INVX1 U1905 ( .A(n1236), .Y(n1989) );
  AND2X1 U1906 ( .A(n2526), .B(n3660), .Y(n1234) );
  INVX1 U1907 ( .A(n1234), .Y(n1990) );
  AND2X1 U1908 ( .A(n2521), .B(n3660), .Y(n1229) );
  INVX1 U1909 ( .A(n1229), .Y(n1991) );
  AND2X1 U1910 ( .A(n3018), .B(n3661), .Y(n1194) );
  INVX1 U1911 ( .A(n1194), .Y(n1992) );
  AND2X1 U1912 ( .A(n3016), .B(n3661), .Y(n1192) );
  INVX1 U1913 ( .A(n1192), .Y(n1993) );
  AND2X1 U1914 ( .A(n3106), .B(n3661), .Y(n1187) );
  INVX1 U1915 ( .A(n1187), .Y(n1994) );
  AND2X1 U1916 ( .A(n2595), .B(n3662), .Y(n1171) );
  INVX1 U1917 ( .A(n1171), .Y(n1995) );
  AND2X1 U1918 ( .A(n2587), .B(n3662), .Y(n1163) );
  INVX1 U1919 ( .A(n1163), .Y(n1996) );
  AND2X1 U1920 ( .A(n2585), .B(n3662), .Y(n1161) );
  INVX1 U1921 ( .A(n1161), .Y(n1997) );
  AND2X1 U1922 ( .A(n2584), .B(n3662), .Y(n1160) );
  INVX1 U1923 ( .A(n1160), .Y(n1998) );
  AND2X1 U1924 ( .A(n2802), .B(n3663), .Y(n1127) );
  INVX1 U1925 ( .A(n1127), .Y(n1999) );
  AND2X1 U1926 ( .A(n2800), .B(n3663), .Y(n1125) );
  INVX1 U1927 ( .A(n1125), .Y(n2000) );
  AND2X1 U1928 ( .A(n2505), .B(n3664), .Y(n1103) );
  INVX1 U1929 ( .A(n1103), .Y(n2001) );
  AND2X1 U1930 ( .A(n2497), .B(n3664), .Y(n1095) );
  INVX1 U1931 ( .A(n1095), .Y(n2002) );
  AND2X1 U1932 ( .A(n2495), .B(n3664), .Y(n1093) );
  INVX1 U1933 ( .A(n1093), .Y(n2003) );
  AND2X1 U1934 ( .A(n2494), .B(n3664), .Y(n1092) );
  INVX1 U1935 ( .A(n1092), .Y(n2004) );
  AND2X1 U1936 ( .A(n2994), .B(n3665), .Y(n1069) );
  INVX1 U1937 ( .A(n1069), .Y(n2005) );
  AND2X1 U1938 ( .A(n2992), .B(n3665), .Y(n1067) );
  INVX1 U1939 ( .A(n1067), .Y(n2006) );
  AND2X1 U1940 ( .A(n2990), .B(n3665), .Y(n1065) );
  INVX1 U1941 ( .A(n1065), .Y(n2007) );
  AND2X1 U1942 ( .A(n2986), .B(n3665), .Y(n1061) );
  INVX1 U1943 ( .A(n1061), .Y(n2008) );
  AND2X1 U1944 ( .A(n2985), .B(n3665), .Y(n1060) );
  INVX1 U1945 ( .A(n1060), .Y(n2009) );
  AND2X1 U1946 ( .A(n2983), .B(n3665), .Y(n1058) );
  INVX1 U1947 ( .A(n1058), .Y(n2010) );
  AND2X1 U1948 ( .A(n2982), .B(n3665), .Y(n1057) );
  INVX1 U1949 ( .A(n1057), .Y(n2011) );
  AND2X1 U1950 ( .A(n2752), .B(n3666), .Y(n1043) );
  INVX1 U1951 ( .A(n1043), .Y(n2012) );
  AND2X1 U1952 ( .A(n2748), .B(n3666), .Y(n1038) );
  INVX1 U1953 ( .A(n1038), .Y(n2013) );
  AND2X1 U1954 ( .A(n2739), .B(n3666), .Y(n1029) );
  INVX1 U1955 ( .A(n1029), .Y(n2014) );
  AND2X1 U1956 ( .A(n2730), .B(n3666), .Y(n1020) );
  INVX1 U1957 ( .A(n1020), .Y(n2015) );
  AND2X1 U1958 ( .A(n2963), .B(n3667), .Y(n1002) );
  INVX1 U1959 ( .A(n1002), .Y(n2016) );
  AND2X1 U1960 ( .A(n2962), .B(n3667), .Y(n1001) );
  INVX1 U1961 ( .A(n1001), .Y(n2017) );
  AND2X1 U1962 ( .A(n2960), .B(n3667), .Y(n999) );
  INVX1 U1963 ( .A(n999), .Y(n2018) );
  AND2X1 U1964 ( .A(n2958), .B(n3667), .Y(n997) );
  INVX1 U1965 ( .A(n997), .Y(n2019) );
  AND2X1 U1966 ( .A(n2955), .B(n3667), .Y(n994) );
  INVX1 U1967 ( .A(n994), .Y(n2020) );
  AND2X1 U1968 ( .A(n2954), .B(n3667), .Y(n993) );
  INVX1 U1969 ( .A(n993), .Y(n2021) );
  AND2X1 U1970 ( .A(n2953), .B(n3667), .Y(n992) );
  INVX1 U1971 ( .A(n992), .Y(n2022) );
  AND2X1 U1972 ( .A(n2951), .B(n3667), .Y(n990) );
  INVX1 U1973 ( .A(n990), .Y(n2023) );
  AND2X1 U1974 ( .A(n2950), .B(n3667), .Y(n989) );
  INVX1 U1975 ( .A(n989), .Y(n2024) );
  AND2X1 U1976 ( .A(n2722), .B(n3668), .Y(n977) );
  INVX1 U1977 ( .A(n977), .Y(n2025) );
  AND2X1 U1978 ( .A(n2721), .B(n3668), .Y(n976) );
  INVX1 U1979 ( .A(n976), .Y(n2026) );
  AND2X1 U1980 ( .A(n2717), .B(n3668), .Y(n971) );
  INVX1 U1981 ( .A(n971), .Y(n2027) );
  AND2X1 U1982 ( .A(n2709), .B(n3668), .Y(n962) );
  INVX1 U1983 ( .A(n962), .Y(n2028) );
  AND2X1 U1984 ( .A(n2701), .B(n3668), .Y(n954) );
  INVX1 U1985 ( .A(n954), .Y(n2029) );
  AND2X1 U1986 ( .A(n2700), .B(n3668), .Y(n953) );
  INVX1 U1987 ( .A(n953), .Y(n2030) );
  AND2X1 U1988 ( .A(n3081), .B(n3669), .Y(n925) );
  INVX1 U1989 ( .A(n925), .Y(n2031) );
  AND2X1 U1990 ( .A(n3080), .B(n3669), .Y(n924) );
  INVX1 U1991 ( .A(n924), .Y(n2032) );
  AND2X1 U1992 ( .A(n3079), .B(n3669), .Y(n923) );
  INVX1 U1993 ( .A(n923), .Y(n2033) );
  AND2X1 U1994 ( .A(n3074), .B(n3669), .Y(n918) );
  INVX1 U1995 ( .A(n918), .Y(n2034) );
  AND2X1 U1996 ( .A(n2792), .B(n3670), .Y(n914) );
  INVX1 U1997 ( .A(n914), .Y(n2035) );
  AND2X1 U1998 ( .A(n2791), .B(n3670), .Y(n913) );
  INVX1 U1999 ( .A(n913), .Y(n2036) );
  AND2X1 U2000 ( .A(n2786), .B(n3670), .Y(n908) );
  INVX1 U2001 ( .A(n908), .Y(n2037) );
  AND2X1 U2002 ( .A(n2784), .B(n3670), .Y(n905) );
  INVX1 U2003 ( .A(n905), .Y(n2038) );
  AND2X1 U2004 ( .A(n2783), .B(n3670), .Y(n904) );
  INVX1 U2005 ( .A(n904), .Y(n2039) );
  AND2X1 U2006 ( .A(n2780), .B(n3670), .Y(n901) );
  INVX1 U2007 ( .A(n901), .Y(n2040) );
  AND2X1 U2008 ( .A(n2778), .B(n3670), .Y(n899) );
  INVX1 U2009 ( .A(n899), .Y(n2041) );
  AND2X1 U2010 ( .A(n2776), .B(n3670), .Y(n896) );
  INVX1 U2011 ( .A(n896), .Y(n2042) );
  AND2X1 U2012 ( .A(n2766), .B(n3670), .Y(n886) );
  INVX1 U2013 ( .A(n886), .Y(n2043) );
  AND2X1 U2014 ( .A(n2936), .B(n3671), .Y(n874) );
  INVX1 U2015 ( .A(n874), .Y(n2044) );
  AND2X1 U2016 ( .A(n2927), .B(n3671), .Y(n865) );
  INVX1 U2017 ( .A(n865), .Y(n2045) );
  AND2X1 U2018 ( .A(n2918), .B(n3671), .Y(n856) );
  INVX1 U2019 ( .A(n856), .Y(n2046) );
  AND2X1 U2020 ( .A(n2914), .B(n3671), .Y(n852) );
  INVX1 U2021 ( .A(n852), .Y(n2047) );
  AND2X1 U2022 ( .A(n2696), .B(n3672), .Y(n845) );
  INVX1 U2023 ( .A(n845), .Y(n2048) );
  AND2X1 U2024 ( .A(n2695), .B(n3672), .Y(n844) );
  INVX1 U2025 ( .A(n844), .Y(n2049) );
  AND2X1 U2026 ( .A(n2690), .B(n3672), .Y(n839) );
  INVX1 U2027 ( .A(n839), .Y(n2050) );
  AND2X1 U2028 ( .A(n2688), .B(n3672), .Y(n837) );
  INVX1 U2029 ( .A(n837), .Y(n2051) );
  AND2X1 U2030 ( .A(n2687), .B(n3672), .Y(n835) );
  INVX1 U2031 ( .A(n835), .Y(n2052) );
  AND2X1 U2032 ( .A(n2686), .B(n3672), .Y(n834) );
  INVX1 U2033 ( .A(n834), .Y(n2053) );
  AND2X1 U2034 ( .A(n2684), .B(n3672), .Y(n832) );
  INVX1 U2035 ( .A(n832), .Y(n2054) );
  AND2X1 U2036 ( .A(n2682), .B(n3672), .Y(n830) );
  INVX1 U2037 ( .A(n830), .Y(n2055) );
  AND2X1 U2038 ( .A(n2680), .B(n3672), .Y(n828) );
  INVX1 U2039 ( .A(n828), .Y(n2056) );
  AND2X1 U2040 ( .A(n2679), .B(n3672), .Y(n826) );
  INVX1 U2041 ( .A(n826), .Y(n2057) );
  AND2X1 U2042 ( .A(n2670), .B(n3672), .Y(n817) );
  INVX1 U2043 ( .A(n817), .Y(n2058) );
  AND2X1 U2044 ( .A(n2635), .B(n3748), .Y(n1219) );
  INVX1 U2045 ( .A(n1219), .Y(n2059) );
  AND2X1 U2046 ( .A(n2857), .B(n3747), .Y(n1286) );
  INVX1 U2047 ( .A(n1286), .Y(n2060) );
  AND2X1 U2093 ( .A(n1219), .B(n883), .Y(n917) );
  AND2X1 U2094 ( .A(n2691), .B(n3672), .Y(n840) );
  INVX1 U2095 ( .A(n840), .Y(n2106) );
  AND2X1 U2096 ( .A(n2698), .B(n3672), .Y(n847) );
  INVX1 U2097 ( .A(n847), .Y(n2107) );
  AND2X1 U2098 ( .A(n2785), .B(n3670), .Y(n907) );
  INVX1 U2099 ( .A(n907), .Y(n2108) );
  AND2X1 U2100 ( .A(n2793), .B(n3670), .Y(n915) );
  INVX1 U2101 ( .A(n915), .Y(n2109) );
  AND2X1 U2102 ( .A(n2702), .B(n3668), .Y(n955) );
  INVX1 U2103 ( .A(n955), .Y(n2110) );
  AND2X1 U2104 ( .A(n2723), .B(n3668), .Y(n978) );
  INVX1 U2105 ( .A(n978), .Y(n2111) );
  AND2X1 U2106 ( .A(n2729), .B(n3666), .Y(n1018) );
  INVX1 U2107 ( .A(n1018), .Y(n2112) );
  AND2X1 U2108 ( .A(n2741), .B(n3666), .Y(n1031) );
  INVX1 U2109 ( .A(n1031), .Y(n2113) );
  AND2X1 U2110 ( .A(n2750), .B(n3666), .Y(n1040) );
  INVX1 U2111 ( .A(n1040), .Y(n2114) );
  AND2X1 U2112 ( .A(n2916), .B(n3671), .Y(n854) );
  INVX1 U2113 ( .A(n854), .Y(n2115) );
  AND2X1 U2114 ( .A(n2939), .B(n3671), .Y(n877) );
  INVX1 U2115 ( .A(n877), .Y(n2116) );
  AND2X1 U2116 ( .A(n2498), .B(n3664), .Y(n1096) );
  INVX1 U2117 ( .A(n1096), .Y(n2117) );
  AND2X1 U2118 ( .A(n2506), .B(n3664), .Y(n1104) );
  INVX1 U2119 ( .A(n1104), .Y(n2118) );
  AND2X1 U2120 ( .A(n2522), .B(n3660), .Y(n1230) );
  INVX1 U2121 ( .A(n1230), .Y(n2119) );
  AND2X1 U2122 ( .A(n2529), .B(n3660), .Y(n1238) );
  INVX1 U2123 ( .A(n1238), .Y(n2120) );
  AND2X1 U2124 ( .A(n2612), .B(n3658), .Y(n1293) );
  INVX1 U2125 ( .A(n1293), .Y(n2121) );
  AND2X1 U2126 ( .A(n2803), .B(n3663), .Y(n1128) );
  INVX1 U2127 ( .A(n1128), .Y(n2122) );
  AND2X1 U2128 ( .A(n2810), .B(n3663), .Y(n1135) );
  INVX1 U2129 ( .A(n1135), .Y(n2123) );
  AND2X1 U2130 ( .A(n3017), .B(n3661), .Y(n1193) );
  INVX1 U2131 ( .A(n1193), .Y(n2124) );
  AND2X1 U2132 ( .A(n2837), .B(n3659), .Y(n1267) );
  INVX1 U2133 ( .A(n1267), .Y(n2125) );
  AND2X1 U2134 ( .A(n3011), .B(n3657), .Y(n1322) );
  INVX1 U2135 ( .A(n1322), .Y(n2126) );
  AND2X1 U2136 ( .A(n3049), .B(n3657), .Y(n1329) );
  INVX1 U2137 ( .A(n1329), .Y(n2127) );
  AND2X1 U2138 ( .A(n1118), .B(n2538), .Y(n1085) );
  AND2X1 U2139 ( .A(n2689), .B(n3672), .Y(n838) );
  INVX1 U2140 ( .A(n838), .Y(n2128) );
  AND2X1 U2141 ( .A(n2697), .B(n3672), .Y(n846) );
  INVX1 U2142 ( .A(n846), .Y(n2129) );
  AND2X1 U2143 ( .A(n2787), .B(n3670), .Y(n909) );
  INVX1 U2144 ( .A(n909), .Y(n2130) );
  AND2X1 U2145 ( .A(n2794), .B(n3670), .Y(n916) );
  INVX1 U2146 ( .A(n916), .Y(n2131) );
  AND2X1 U2147 ( .A(n2710), .B(n3668), .Y(n963) );
  INVX1 U2148 ( .A(n963), .Y(n2132) );
  AND2X1 U2149 ( .A(n2718), .B(n3668), .Y(n972) );
  INVX1 U2150 ( .A(n972), .Y(n2133) );
  AND2X1 U2151 ( .A(n2731), .B(n3666), .Y(n1021) );
  INVX1 U2152 ( .A(n1021), .Y(n2134) );
  AND2X1 U2153 ( .A(n2753), .B(n3666), .Y(n1044) );
  INVX1 U2154 ( .A(n1044), .Y(n2135) );
  AND2X1 U2155 ( .A(n2915), .B(n3671), .Y(n853) );
  INVX1 U2156 ( .A(n853), .Y(n2136) );
  AND2X1 U2157 ( .A(n2938), .B(n3671), .Y(n876) );
  INVX1 U2158 ( .A(n876), .Y(n2137) );
  AND2X1 U2159 ( .A(n3077), .B(n3669), .Y(n921) );
  INVX1 U2160 ( .A(n921), .Y(n2138) );
  AND2X1 U2161 ( .A(n3100), .B(n3669), .Y(n944) );
  INVX1 U2162 ( .A(n944), .Y(n2139) );
  AND2X1 U2163 ( .A(n2588), .B(n3662), .Y(n1164) );
  INVX1 U2164 ( .A(n1164), .Y(n2140) );
  AND2X1 U2165 ( .A(n2596), .B(n3662), .Y(n1172) );
  INVX1 U2166 ( .A(n1172), .Y(n2141) );
  AND2X1 U2167 ( .A(n2518), .B(n3660), .Y(n1226) );
  INVX1 U2168 ( .A(n1226), .Y(n2142) );
  AND2X1 U2169 ( .A(n2616), .B(n3658), .Y(n1297) );
  INVX1 U2170 ( .A(n1297), .Y(n2143) );
  AND2X1 U2171 ( .A(n2623), .B(n3658), .Y(n1305) );
  INVX1 U2172 ( .A(n1305), .Y(n2144) );
  AND2X1 U2173 ( .A(n3009), .B(n3663), .Y(n1120) );
  INVX1 U2174 ( .A(n1120), .Y(n2145) );
  AND2X1 U2175 ( .A(n2801), .B(n3663), .Y(n1126) );
  INVX1 U2176 ( .A(n1126), .Y(n2146) );
  AND2X1 U2177 ( .A(n3019), .B(n3661), .Y(n1195) );
  INVX1 U2178 ( .A(n1195), .Y(n2147) );
  AND2X1 U2179 ( .A(n3026), .B(n3661), .Y(n1202) );
  INVX1 U2180 ( .A(n1202), .Y(n2148) );
  AND2X1 U2181 ( .A(n2831), .B(n3659), .Y(n1261) );
  INVX1 U2182 ( .A(n1261), .Y(n2149) );
  AND2X1 U2183 ( .A(n3055), .B(n3657), .Y(n1335) );
  INVX1 U2184 ( .A(n1335), .Y(n2150) );
  AND2X1 U2185 ( .A(n2539), .B(n883), .Y(n1051) );
  AND2X1 U2186 ( .A(n2673), .B(n3672), .Y(n820) );
  INVX1 U2187 ( .A(n820), .Y(n2151) );
  AND2X1 U2188 ( .A(n2694), .B(n3672), .Y(n843) );
  INVX1 U2189 ( .A(n843), .Y(n2152) );
  AND2X1 U2190 ( .A(n2767), .B(n3670), .Y(n887) );
  INVX1 U2191 ( .A(n887), .Y(n2153) );
  AND2X1 U2192 ( .A(n2788), .B(n3670), .Y(n910) );
  INVX1 U2193 ( .A(n910), .Y(n2154) );
  AND2X1 U2194 ( .A(n2720), .B(n3668), .Y(n975) );
  INVX1 U2195 ( .A(n975), .Y(n2155) );
  AND2X1 U2196 ( .A(n2727), .B(n3668), .Y(n982) );
  INVX1 U2197 ( .A(n982), .Y(n2156) );
  AND2X1 U2198 ( .A(n2749), .B(n3666), .Y(n1039) );
  INVX1 U2199 ( .A(n1039), .Y(n2157) );
  AND2X1 U2200 ( .A(n2756), .B(n3666), .Y(n1047) );
  INVX1 U2201 ( .A(n1047), .Y(n2158) );
  AND2X1 U2202 ( .A(n2932), .B(n3671), .Y(n870) );
  INVX1 U2203 ( .A(n870), .Y(n2159) );
  AND2X1 U2204 ( .A(n2942), .B(n3671), .Y(n880) );
  INVX1 U2205 ( .A(n880), .Y(n2160) );
  AND2X1 U2206 ( .A(n3090), .B(n3669), .Y(n934) );
  INVX1 U2207 ( .A(n934), .Y(n2161) );
  AND2X1 U2208 ( .A(n3102), .B(n3669), .Y(n946) );
  INVX1 U2209 ( .A(n946), .Y(n2162) );
  AND2X1 U2210 ( .A(n2499), .B(n3664), .Y(n1097) );
  INVX1 U2211 ( .A(n1097), .Y(n2163) );
  AND2X1 U2212 ( .A(n2508), .B(n3664), .Y(n1106) );
  INVX1 U2213 ( .A(n1106), .Y(n2164) );
  AND2X1 U2214 ( .A(n2795), .B(n3662), .Y(n1154) );
  INVX1 U2215 ( .A(n1154), .Y(n2165) );
  AND2X1 U2216 ( .A(n2583), .B(n3662), .Y(n1159) );
  INVX1 U2217 ( .A(n1159), .Y(n2166) );
  AND2X1 U2218 ( .A(n2520), .B(n3660), .Y(n1228) );
  INVX1 U2219 ( .A(n1228), .Y(n2167) );
  AND2X1 U2220 ( .A(n2613), .B(n3658), .Y(n1294) );
  INVX1 U2221 ( .A(n1294), .Y(n2168) );
  AND2X1 U2222 ( .A(n2805), .B(n3663), .Y(n1130) );
  INVX1 U2223 ( .A(n1130), .Y(n2169) );
  AND2X1 U2224 ( .A(n2813), .B(n3663), .Y(n1138) );
  INVX1 U2225 ( .A(n1138), .Y(n2170) );
  AND2X1 U2226 ( .A(n3024), .B(n3661), .Y(n1200) );
  INVX1 U2227 ( .A(n1200), .Y(n2171) );
  AND2X1 U2228 ( .A(n2833), .B(n3659), .Y(n1263) );
  INVX1 U2229 ( .A(n1263), .Y(n2172) );
  AND2X1 U2230 ( .A(n2841), .B(n3659), .Y(n1271) );
  INVX1 U2231 ( .A(n1271), .Y(n2173) );
  AND2X1 U2232 ( .A(n3050), .B(n3657), .Y(n1330) );
  INVX1 U2233 ( .A(n1330), .Y(n2174) );
  AND2X1 U2234 ( .A(n3057), .B(n3657), .Y(n1337) );
  INVX1 U2235 ( .A(n1337), .Y(n2175) );
  AND2X1 U2236 ( .A(n1286), .B(n883), .Y(n983) );
  AND2X1 U2237 ( .A(n3111), .B(n1050), .Y(n883) );
  AND2X1 U2238 ( .A(n2671), .B(n3672), .Y(n818) );
  INVX1 U2239 ( .A(n818), .Y(n2176) );
  AND2X1 U2240 ( .A(n2692), .B(n3672), .Y(n841) );
  INVX1 U2241 ( .A(n841), .Y(n2177) );
  AND2X1 U2242 ( .A(n2769), .B(n3670), .Y(n889) );
  INVX1 U2243 ( .A(n889), .Y(n2178) );
  AND2X1 U2244 ( .A(n2790), .B(n3670), .Y(n912) );
  INVX1 U2245 ( .A(n912), .Y(n2179) );
  AND2X1 U2246 ( .A(n2719), .B(n3668), .Y(n973) );
  INVX1 U2247 ( .A(n973), .Y(n2180) );
  AND2X1 U2248 ( .A(n2726), .B(n3668), .Y(n981) );
  INVX1 U2249 ( .A(n981), .Y(n2181) );
  AND2X1 U2250 ( .A(n2751), .B(n3666), .Y(n1041) );
  INVX1 U2251 ( .A(n1041), .Y(n2182) );
  AND2X1 U2252 ( .A(n2757), .B(n3666), .Y(n1048) );
  INVX1 U2253 ( .A(n1048), .Y(n2183) );
  AND2X1 U2254 ( .A(n2929), .B(n3671), .Y(n867) );
  INVX1 U2255 ( .A(n867), .Y(n2184) );
  AND2X1 U2256 ( .A(n2941), .B(n3671), .Y(n879) );
  INVX1 U2257 ( .A(n879), .Y(n2185) );
  AND2X1 U2258 ( .A(n3093), .B(n3669), .Y(n937) );
  INVX1 U2259 ( .A(n937), .Y(n2186) );
  AND2X1 U2260 ( .A(n3103), .B(n3669), .Y(n947) );
  INVX1 U2261 ( .A(n947), .Y(n2187) );
  AND2X1 U2262 ( .A(n2989), .B(n3665), .Y(n1064) );
  INVX1 U2263 ( .A(n1064), .Y(n2188) );
  AND2X1 U2264 ( .A(n2998), .B(n3665), .Y(n1073) );
  INVX1 U2265 ( .A(n1073), .Y(n2189) );
  AND2X1 U2266 ( .A(n2758), .B(n3664), .Y(n1086) );
  INVX1 U2267 ( .A(n1086), .Y(n2190) );
  AND2X1 U2268 ( .A(n2493), .B(n3664), .Y(n1091) );
  INVX1 U2269 ( .A(n1091), .Y(n2191) );
  AND2X1 U2270 ( .A(n2589), .B(n3662), .Y(n1165) );
  INVX1 U2271 ( .A(n1165), .Y(n2192) );
  AND2X1 U2272 ( .A(n2598), .B(n3662), .Y(n1174) );
  INVX1 U2273 ( .A(n1174), .Y(n2193) );
  AND2X1 U2274 ( .A(n2519), .B(n3660), .Y(n1227) );
  INVX1 U2275 ( .A(n1227), .Y(n2194) );
  AND2X1 U2276 ( .A(n2614), .B(n3658), .Y(n1295) );
  INVX1 U2277 ( .A(n1295), .Y(n2195) );
  AND2X1 U2278 ( .A(n2808), .B(n3663), .Y(n1133) );
  INVX1 U2279 ( .A(n1133), .Y(n2196) );
  AND2X1 U2280 ( .A(n3021), .B(n3661), .Y(n1197) );
  INVX1 U2281 ( .A(n1197), .Y(n2197) );
  AND2X1 U2282 ( .A(n3029), .B(n3661), .Y(n1205) );
  INVX1 U2283 ( .A(n1205), .Y(n2198) );
  AND2X1 U2284 ( .A(n2832), .B(n3659), .Y(n1262) );
  INVX1 U2285 ( .A(n1262), .Y(n2199) );
  AND2X1 U2286 ( .A(n2839), .B(n3659), .Y(n1269) );
  INVX1 U2287 ( .A(n1269), .Y(n2200) );
  AND2X1 U2288 ( .A(n3051), .B(n3657), .Y(n1331) );
  INVX1 U2289 ( .A(n1331), .Y(n2201) );
  AND2X1 U2290 ( .A(n3059), .B(n3657), .Y(n1339) );
  INVX1 U2291 ( .A(n1339), .Y(n2202) );
  AND2X1 U2292 ( .A(n2672), .B(n3672), .Y(n819) );
  INVX1 U2293 ( .A(n819), .Y(n2203) );
  AND2X1 U2294 ( .A(n2693), .B(n3672), .Y(n842) );
  INVX1 U2295 ( .A(n842), .Y(n2204) );
  AND2X1 U2296 ( .A(n2770), .B(n3670), .Y(n890) );
  INVX1 U2297 ( .A(n890), .Y(n2205) );
  AND2X1 U2298 ( .A(n2716), .B(n3668), .Y(n970) );
  INVX1 U2299 ( .A(n970), .Y(n2206) );
  AND2X1 U2300 ( .A(n2725), .B(n3668), .Y(n980) );
  INVX1 U2301 ( .A(n980), .Y(n2207) );
  AND2X1 U2302 ( .A(n2743), .B(n3666), .Y(n1033) );
  INVX1 U2303 ( .A(n1033), .Y(n2208) );
  AND2X1 U2304 ( .A(n2754), .B(n3666), .Y(n1045) );
  INVX1 U2305 ( .A(n1045), .Y(n2209) );
  AND2X1 U2306 ( .A(n2937), .B(n3671), .Y(n875) );
  INVX1 U2307 ( .A(n875), .Y(n2210) );
  AND2X1 U2308 ( .A(n2944), .B(n3671), .Y(n882) );
  INVX1 U2309 ( .A(n882), .Y(n2211) );
  AND2X1 U2310 ( .A(n3096), .B(n3669), .Y(n940) );
  INVX1 U2311 ( .A(n940), .Y(n2212) );
  AND2X1 U2312 ( .A(n3104), .B(n3669), .Y(n948) );
  INVX1 U2313 ( .A(n948), .Y(n2213) );
  AND2X1 U2314 ( .A(n2949), .B(n3667), .Y(n988) );
  INVX1 U2315 ( .A(n988), .Y(n2214) );
  AND2X1 U2316 ( .A(n2972), .B(n3667), .Y(n1011) );
  INVX1 U2317 ( .A(n1011), .Y(n2215) );
  AND2X1 U2318 ( .A(n2977), .B(n3665), .Y(n1052) );
  INVX1 U2319 ( .A(n1052), .Y(n2216) );
  AND2X1 U2320 ( .A(n2984), .B(n3665), .Y(n1059) );
  INVX1 U2321 ( .A(n1059), .Y(n2217) );
  AND2X1 U2322 ( .A(n2496), .B(n3664), .Y(n1094) );
  INVX1 U2323 ( .A(n1094), .Y(n2218) );
  AND2X1 U2324 ( .A(n2503), .B(n3664), .Y(n1101) );
  INVX1 U2325 ( .A(n1101), .Y(n2219) );
  AND2X1 U2326 ( .A(n2591), .B(n3662), .Y(n1167) );
  INVX1 U2327 ( .A(n1167), .Y(n2220) );
  AND2X1 U2328 ( .A(n2516), .B(n3660), .Y(n1223) );
  INVX1 U2329 ( .A(n1223), .Y(n2221) );
  AND2X1 U2330 ( .A(n2535), .B(n3660), .Y(n1246) );
  INVX1 U2331 ( .A(n1246), .Y(n2222) );
  AND2X1 U2332 ( .A(n2608), .B(n3658), .Y(n1289) );
  INVX1 U2333 ( .A(n1289), .Y(n2223) );
  AND2X1 U2334 ( .A(n2621), .B(n3658), .Y(n1302) );
  INVX1 U2335 ( .A(n1302), .Y(n2224) );
  AND2X1 U2336 ( .A(n2628), .B(n3658), .Y(n1311) );
  INVX1 U2337 ( .A(n1311), .Y(n2225) );
  AND2X1 U2338 ( .A(n2807), .B(n3663), .Y(n1132) );
  INVX1 U2339 ( .A(n1132), .Y(n2226) );
  AND2X1 U2340 ( .A(n2816), .B(n3663), .Y(n1141) );
  INVX1 U2341 ( .A(n1141), .Y(n2227) );
  AND2X1 U2342 ( .A(n3020), .B(n3661), .Y(n1196) );
  INVX1 U2343 ( .A(n1196), .Y(n2228) );
  AND2X1 U2344 ( .A(n3028), .B(n3661), .Y(n1204) );
  INVX1 U2345 ( .A(n1204), .Y(n2229) );
  AND2X1 U2346 ( .A(n2835), .B(n3659), .Y(n1265) );
  INVX1 U2347 ( .A(n1265), .Y(n2230) );
  AND2X1 U2348 ( .A(n2844), .B(n3659), .Y(n1274) );
  INVX1 U2349 ( .A(n1274), .Y(n2231) );
  AND2X1 U2350 ( .A(n3052), .B(n3657), .Y(n1332) );
  INVX1 U2351 ( .A(n1332), .Y(n2232) );
  AND2X1 U2352 ( .A(n3060), .B(n3657), .Y(n1340) );
  INVX1 U2353 ( .A(n1340), .Y(n2233) );
  AND2X1 U2354 ( .A(n2768), .B(n3670), .Y(n888) );
  INVX1 U2355 ( .A(n888), .Y(n2234) );
  AND2X1 U2356 ( .A(n2789), .B(n3670), .Y(n911) );
  INVX1 U2357 ( .A(n911), .Y(n2235) );
  AND2X1 U2358 ( .A(n2713), .B(n3668), .Y(n967) );
  INVX1 U2359 ( .A(n967), .Y(n2236) );
  AND2X1 U2360 ( .A(n2724), .B(n3668), .Y(n979) );
  INVX1 U2361 ( .A(n979), .Y(n2237) );
  AND2X1 U2362 ( .A(n2746), .B(n3666), .Y(n1036) );
  INVX1 U2363 ( .A(n1036), .Y(n2238) );
  AND2X1 U2364 ( .A(n2755), .B(n3666), .Y(n1046) );
  INVX1 U2365 ( .A(n1046), .Y(n2239) );
  AND2X1 U2366 ( .A(n2935), .B(n3671), .Y(n873) );
  INVX1 U2367 ( .A(n873), .Y(n2240) );
  AND2X1 U2368 ( .A(n2943), .B(n3671), .Y(n881) );
  INVX1 U2369 ( .A(n881), .Y(n2241) );
  AND2X1 U2370 ( .A(n3098), .B(n3669), .Y(n942) );
  INVX1 U2371 ( .A(n942), .Y(n2242) );
  AND2X1 U2372 ( .A(n3105), .B(n3669), .Y(n949) );
  INVX1 U2373 ( .A(n949), .Y(n2243) );
  AND2X1 U2374 ( .A(n2945), .B(n3667), .Y(n984) );
  INVX1 U2375 ( .A(n984), .Y(n2244) );
  AND2X1 U2376 ( .A(n2952), .B(n3667), .Y(n991) );
  INVX1 U2377 ( .A(n991), .Y(n2245) );
  AND2X1 U2378 ( .A(n2981), .B(n3665), .Y(n1056) );
  INVX1 U2379 ( .A(n1056), .Y(n2246) );
  AND2X1 U2380 ( .A(n3004), .B(n3665), .Y(n1079) );
  INVX1 U2381 ( .A(n1079), .Y(n2247) );
  AND2X1 U2382 ( .A(n2501), .B(n3664), .Y(n1099) );
  INVX1 U2383 ( .A(n1099), .Y(n2248) );
  AND2X1 U2384 ( .A(n2586), .B(n3662), .Y(n1162) );
  INVX1 U2385 ( .A(n1162), .Y(n2249) );
  AND2X1 U2386 ( .A(n2593), .B(n3662), .Y(n1169) );
  INVX1 U2387 ( .A(n1169), .Y(n2250) );
  AND2X1 U2388 ( .A(n2515), .B(n3660), .Y(n1222) );
  INVX1 U2389 ( .A(n1222), .Y(n2251) );
  AND2X1 U2390 ( .A(n2527), .B(n3660), .Y(n1235) );
  INVX1 U2391 ( .A(n1235), .Y(n2252) );
  AND2X1 U2392 ( .A(n2534), .B(n3660), .Y(n1244) );
  INVX1 U2393 ( .A(n1244), .Y(n2253) );
  AND2X1 U2394 ( .A(n2609), .B(n3658), .Y(n1290) );
  INVX1 U2395 ( .A(n1290), .Y(n2254) );
  AND2X1 U2396 ( .A(n2629), .B(n3658), .Y(n1313) );
  INVX1 U2397 ( .A(n1313), .Y(n2255) );
  AND2X1 U2398 ( .A(n2804), .B(n3663), .Y(n1129) );
  INVX1 U2399 ( .A(n1129), .Y(n2256) );
  AND2X1 U2400 ( .A(n2812), .B(n3663), .Y(n1137) );
  INVX1 U2401 ( .A(n1137), .Y(n2257) );
  AND2X1 U2402 ( .A(n3023), .B(n3661), .Y(n1199) );
  INVX1 U2403 ( .A(n1199), .Y(n2258) );
  AND2X1 U2404 ( .A(n3032), .B(n3661), .Y(n1208) );
  INVX1 U2405 ( .A(n1208), .Y(n2259) );
  AND2X1 U2406 ( .A(n2834), .B(n3659), .Y(n1264) );
  INVX1 U2407 ( .A(n1264), .Y(n2260) );
  AND2X1 U2408 ( .A(n2842), .B(n3659), .Y(n1272) );
  INVX1 U2409 ( .A(n1272), .Y(n2261) );
  AND2X1 U2410 ( .A(n3053), .B(n3657), .Y(n1333) );
  INVX1 U2411 ( .A(n1333), .Y(n2262) );
  AND2X1 U2412 ( .A(n3062), .B(n3657), .Y(n1342) );
  INVX1 U2413 ( .A(n1342), .Y(n2263) );
  AND2X1 U2414 ( .A(n2538), .B(n849), .Y(n815) );
  AND2X1 U2415 ( .A(n2703), .B(n3668), .Y(n956) );
  INVX1 U2416 ( .A(n956), .Y(n2264) );
  AND2X1 U2417 ( .A(n2733), .B(n3666), .Y(n1023) );
  INVX1 U2418 ( .A(n1023), .Y(n2265) );
  AND2X1 U2419 ( .A(n2917), .B(n3671), .Y(n855) );
  INVX1 U2420 ( .A(n855), .Y(n2266) );
  AND2X1 U2421 ( .A(n2940), .B(n3671), .Y(n878) );
  INVX1 U2422 ( .A(n878), .Y(n2267) );
  AND2X1 U2423 ( .A(n3087), .B(n3669), .Y(n931) );
  INVX1 U2424 ( .A(n931), .Y(n2268) );
  AND2X1 U2425 ( .A(n2969), .B(n3667), .Y(n1008) );
  INVX1 U2426 ( .A(n1008), .Y(n2269) );
  AND2X1 U2427 ( .A(n2976), .B(n3667), .Y(n1015) );
  INVX1 U2428 ( .A(n1015), .Y(n2270) );
  AND2X1 U2429 ( .A(n2999), .B(n3665), .Y(n1074) );
  INVX1 U2430 ( .A(n1074), .Y(n2271) );
  AND2X1 U2431 ( .A(n3007), .B(n3665), .Y(n1082) );
  INVX1 U2432 ( .A(n1082), .Y(n2272) );
  AND2X1 U2433 ( .A(n2507), .B(n3664), .Y(n1105) );
  INVX1 U2434 ( .A(n1105), .Y(n2273) );
  AND2X1 U2435 ( .A(n2513), .B(n3664), .Y(n1115) );
  INVX1 U2436 ( .A(n1115), .Y(n2274) );
  AND2X1 U2437 ( .A(n2594), .B(n3662), .Y(n1170) );
  INVX1 U2438 ( .A(n1170), .Y(n2275) );
  AND2X1 U2439 ( .A(n2603), .B(n3662), .Y(n1182) );
  INVX1 U2440 ( .A(n1182), .Y(n2276) );
  AND2X1 U2441 ( .A(n2517), .B(n3660), .Y(n1224) );
  INVX1 U2442 ( .A(n1224), .Y(n2277) );
  AND2X1 U2443 ( .A(n2536), .B(n3660), .Y(n1247) );
  INVX1 U2444 ( .A(n1247), .Y(n2278) );
  AND2X1 U2445 ( .A(n2617), .B(n3658), .Y(n1298) );
  INVX1 U2446 ( .A(n1298), .Y(n2279) );
  AND2X1 U2447 ( .A(n2624), .B(n3658), .Y(n1306) );
  INVX1 U2448 ( .A(n1306), .Y(n2280) );
  AND2X1 U2449 ( .A(n2797), .B(n3663), .Y(n1122) );
  INVX1 U2450 ( .A(n1122), .Y(n2281) );
  AND2X1 U2451 ( .A(n2819), .B(n3663), .Y(n1145) );
  INVX1 U2452 ( .A(n1145), .Y(n2282) );
  AND2X1 U2453 ( .A(n3022), .B(n3661), .Y(n1198) );
  INVX1 U2454 ( .A(n1198), .Y(n2283) );
  AND2X1 U2455 ( .A(n3031), .B(n3661), .Y(n1207) );
  INVX1 U2456 ( .A(n1207), .Y(n2284) );
  AND2X1 U2457 ( .A(n2825), .B(n3659), .Y(n1255) );
  INVX1 U2458 ( .A(n1255), .Y(n2285) );
  AND2X1 U2459 ( .A(n2838), .B(n3659), .Y(n1268) );
  INVX1 U2460 ( .A(n1268), .Y(n2286) );
  AND2X1 U2461 ( .A(n2847), .B(n3659), .Y(n1277) );
  INVX1 U2462 ( .A(n1277), .Y(n2287) );
  AND2X1 U2463 ( .A(n3054), .B(n3657), .Y(n1334) );
  INVX1 U2464 ( .A(n1334), .Y(n2288) );
  AND2X1 U2465 ( .A(n3063), .B(n3657), .Y(n1343) );
  INVX1 U2466 ( .A(n1343), .Y(n2289) );
  AND2X1 U2467 ( .A(n1219), .B(n849), .Y(n884) );
  AND2X1 U2468 ( .A(n2669), .B(n3672), .Y(n816) );
  INVX1 U2469 ( .A(n816), .Y(n2290) );
  AND2X1 U2470 ( .A(n2732), .B(n3666), .Y(n1022) );
  INVX1 U2471 ( .A(n1022), .Y(n2291) );
  AND2X1 U2472 ( .A(n2919), .B(n3671), .Y(n857) );
  INVX1 U2473 ( .A(n857), .Y(n2292) );
  AND2X1 U2474 ( .A(n3078), .B(n3669), .Y(n922) );
  INVX1 U2475 ( .A(n922), .Y(n2293) );
  AND2X1 U2476 ( .A(n3101), .B(n3669), .Y(n945) );
  INVX1 U2477 ( .A(n945), .Y(n2294) );
  AND2X1 U2478 ( .A(n2967), .B(n3667), .Y(n1006) );
  INVX1 U2479 ( .A(n1006), .Y(n2295) );
  AND2X1 U2480 ( .A(n2975), .B(n3667), .Y(n1014) );
  INVX1 U2481 ( .A(n1014), .Y(n2296) );
  AND2X1 U2482 ( .A(n3001), .B(n3665), .Y(n1076) );
  INVX1 U2483 ( .A(n1076), .Y(n2297) );
  AND2X1 U2484 ( .A(n3008), .B(n3665), .Y(n1083) );
  INVX1 U2485 ( .A(n1083), .Y(n2298) );
  AND2X1 U2486 ( .A(n2504), .B(n3664), .Y(n1102) );
  INVX1 U2487 ( .A(n1102), .Y(n2299) );
  AND2X1 U2488 ( .A(n2512), .B(n3664), .Y(n1114) );
  INVX1 U2489 ( .A(n1114), .Y(n2300) );
  AND2X1 U2490 ( .A(n2597), .B(n3662), .Y(n1173) );
  INVX1 U2491 ( .A(n1173), .Y(n2301) );
  AND2X1 U2492 ( .A(n2604), .B(n3662), .Y(n1183) );
  INVX1 U2493 ( .A(n1183), .Y(n2302) );
  AND2X1 U2494 ( .A(n2523), .B(n3660), .Y(n1231) );
  INVX1 U2495 ( .A(n1231), .Y(n2303) );
  AND2X1 U2496 ( .A(n2530), .B(n3660), .Y(n1239) );
  INVX1 U2497 ( .A(n1239), .Y(n2304) );
  AND2X1 U2498 ( .A(n2610), .B(n3658), .Y(n1291) );
  INVX1 U2499 ( .A(n1291), .Y(n2305) );
  AND2X1 U2500 ( .A(n2630), .B(n3658), .Y(n1314) );
  INVX1 U2501 ( .A(n1314), .Y(n2306) );
  AND2X1 U2502 ( .A(n2806), .B(n3663), .Y(n1131) );
  INVX1 U2503 ( .A(n1131), .Y(n2307) );
  AND2X1 U2504 ( .A(n2815), .B(n3663), .Y(n1140) );
  INVX1 U2505 ( .A(n1140), .Y(n2308) );
  AND2X1 U2506 ( .A(n3013), .B(n3661), .Y(n1189) );
  INVX1 U2507 ( .A(n1189), .Y(n2309) );
  AND2X1 U2508 ( .A(n3036), .B(n3661), .Y(n1212) );
  INVX1 U2509 ( .A(n1212), .Y(n2310) );
  AND2X1 U2510 ( .A(n2836), .B(n3659), .Y(n1266) );
  INVX1 U2511 ( .A(n1266), .Y(n2311) );
  AND2X1 U2512 ( .A(n2845), .B(n3659), .Y(n1275) );
  INVX1 U2513 ( .A(n1275), .Y(n2312) );
  AND2X1 U2514 ( .A(n3043), .B(n3657), .Y(n1323) );
  INVX1 U2515 ( .A(n1323), .Y(n2313) );
  AND2X1 U2516 ( .A(n3056), .B(n3657), .Y(n1336) );
  INVX1 U2517 ( .A(n1336), .Y(n2314) );
  AND2X1 U2518 ( .A(n3065), .B(n3657), .Y(n1345) );
  INVX1 U2519 ( .A(n1345), .Y(n2315) );
  AND2X1 U2520 ( .A(n2678), .B(n3672), .Y(n825) );
  INVX1 U2521 ( .A(n825), .Y(n2316) );
  AND2X1 U2522 ( .A(n2685), .B(n3672), .Y(n833) );
  INVX1 U2523 ( .A(n833), .Y(n2317) );
  AND2X1 U2524 ( .A(n2775), .B(n3670), .Y(n895) );
  INVX1 U2525 ( .A(n895), .Y(n2318) );
  AND2X1 U2526 ( .A(n2782), .B(n3670), .Y(n903) );
  INVX1 U2527 ( .A(n903), .Y(n2319) );
  AND2X1 U2528 ( .A(n2704), .B(n3668), .Y(n957) );
  INVX1 U2529 ( .A(n957), .Y(n2320) );
  AND2X1 U2530 ( .A(n2740), .B(n3666), .Y(n1030) );
  INVX1 U2531 ( .A(n1030), .Y(n2321) );
  AND2X1 U2532 ( .A(n2913), .B(n3671), .Y(n851) );
  INVX1 U2533 ( .A(n851), .Y(n2322) );
  AND2X1 U2534 ( .A(n2920), .B(n3671), .Y(n858) );
  INVX1 U2535 ( .A(n858), .Y(n2323) );
  AND2X1 U2536 ( .A(n3082), .B(n3669), .Y(n926) );
  INVX1 U2537 ( .A(n926), .Y(n2324) );
  AND2X1 U2538 ( .A(n3089), .B(n3669), .Y(n933) );
  INVX1 U2539 ( .A(n933), .Y(n2325) );
  AND2X1 U2540 ( .A(n2964), .B(n3667), .Y(n1003) );
  INVX1 U2541 ( .A(n1003), .Y(n2326) );
  AND2X1 U2542 ( .A(n2974), .B(n3667), .Y(n1013) );
  INVX1 U2543 ( .A(n1013), .Y(n2327) );
  AND2X1 U2544 ( .A(n2993), .B(n3665), .Y(n1068) );
  INVX1 U2545 ( .A(n1068), .Y(n2328) );
  AND2X1 U2546 ( .A(n3005), .B(n3665), .Y(n1080) );
  INVX1 U2547 ( .A(n1080), .Y(n2329) );
  AND2X1 U2548 ( .A(n2511), .B(n3664), .Y(n1110) );
  INVX1 U2549 ( .A(n1110), .Y(n2330) );
  AND2X1 U2550 ( .A(n2514), .B(n3664), .Y(n1117) );
  INVX1 U2551 ( .A(n1117), .Y(n2331) );
  AND2X1 U2552 ( .A(n2761), .B(n3662), .Y(n1176) );
  INVX1 U2553 ( .A(n1176), .Y(n2332) );
  AND2X1 U2554 ( .A(n2762), .B(n3662), .Y(n1184) );
  INVX1 U2555 ( .A(n1184), .Y(n2333) );
  AND2X1 U2556 ( .A(n2525), .B(n3660), .Y(n1233) );
  INVX1 U2557 ( .A(n1233), .Y(n2334) );
  AND2X1 U2558 ( .A(n2532), .B(n3660), .Y(n1242) );
  INVX1 U2559 ( .A(n1242), .Y(n2335) );
  AND2X1 U2560 ( .A(n2618), .B(n3658), .Y(n1299) );
  INVX1 U2561 ( .A(n1299), .Y(n2336) );
  AND2X1 U2562 ( .A(n2625), .B(n3658), .Y(n1308) );
  INVX1 U2563 ( .A(n1308), .Y(n2337) );
  AND2X1 U2564 ( .A(n2799), .B(n3663), .Y(n1124) );
  INVX1 U2565 ( .A(n1124), .Y(n2338) );
  AND2X1 U2566 ( .A(n2821), .B(n3663), .Y(n1147) );
  INVX1 U2567 ( .A(n1147), .Y(n2339) );
  AND2X1 U2568 ( .A(n3012), .B(n3661), .Y(n1188) );
  INVX1 U2569 ( .A(n1188), .Y(n2340) );
  AND2X1 U2570 ( .A(n3025), .B(n3661), .Y(n1201) );
  INVX1 U2571 ( .A(n1201), .Y(n2341) );
  AND2X1 U2572 ( .A(n3034), .B(n3661), .Y(n1210) );
  INVX1 U2573 ( .A(n1210), .Y(n2342) );
  AND2X1 U2574 ( .A(n2827), .B(n3659), .Y(n1257) );
  INVX1 U2575 ( .A(n1257), .Y(n2343) );
  AND2X1 U2576 ( .A(n2849), .B(n3659), .Y(n1280) );
  INVX1 U2577 ( .A(n1280), .Y(n2344) );
  AND2X1 U2578 ( .A(n3044), .B(n3657), .Y(n1324) );
  INVX1 U2579 ( .A(n1324), .Y(n2345) );
  AND2X1 U2580 ( .A(n3067), .B(n3657), .Y(n1347) );
  INVX1 U2581 ( .A(n1347), .Y(n2346) );
  AND2X1 U2582 ( .A(n2677), .B(n3672), .Y(n824) );
  INVX1 U2583 ( .A(n824), .Y(n2347) );
  AND2X1 U2584 ( .A(n2683), .B(n3672), .Y(n831) );
  INVX1 U2585 ( .A(n831), .Y(n2348) );
  AND2X1 U2586 ( .A(n2771), .B(n3670), .Y(n891) );
  INVX1 U2587 ( .A(n891), .Y(n2349) );
  AND2X1 U2588 ( .A(n2708), .B(n3668), .Y(n961) );
  INVX1 U2589 ( .A(n961), .Y(n2350) );
  AND2X1 U2590 ( .A(n2715), .B(n3668), .Y(n969) );
  INVX1 U2591 ( .A(n969), .Y(n2351) );
  AND2X1 U2592 ( .A(n2728), .B(n3666), .Y(n1017) );
  INVX1 U2593 ( .A(n1017), .Y(n2352) );
  AND2X1 U2594 ( .A(n2734), .B(n3666), .Y(n1024) );
  INVX1 U2595 ( .A(n1024), .Y(n2353) );
  AND2X1 U2596 ( .A(n2926), .B(n3671), .Y(n864) );
  INVX1 U2597 ( .A(n864), .Y(n2354) );
  AND2X1 U2598 ( .A(n3083), .B(n3669), .Y(n927) );
  INVX1 U2599 ( .A(n927), .Y(n2355) );
  AND2X1 U2600 ( .A(n3091), .B(n3669), .Y(n935) );
  INVX1 U2601 ( .A(n935), .Y(n2356) );
  AND2X1 U2602 ( .A(n2961), .B(n3667), .Y(n1000) );
  INVX1 U2603 ( .A(n1000), .Y(n2357) );
  AND2X1 U2604 ( .A(n2973), .B(n3667), .Y(n1012) );
  INVX1 U2605 ( .A(n1012), .Y(n2358) );
  AND2X1 U2606 ( .A(n2996), .B(n3665), .Y(n1071) );
  INVX1 U2607 ( .A(n1071), .Y(n2359) );
  AND2X1 U2608 ( .A(n3006), .B(n3665), .Y(n1081) );
  INVX1 U2609 ( .A(n1081), .Y(n2360) );
  AND2X1 U2610 ( .A(n2579), .B(n3664), .Y(n1108) );
  INVX1 U2611 ( .A(n1108), .Y(n2361) );
  AND2X1 U2612 ( .A(n2580), .B(n3664), .Y(n1116) );
  INVX1 U2613 ( .A(n1116), .Y(n2362) );
  AND2X1 U2614 ( .A(n2601), .B(n3662), .Y(n1178) );
  INVX1 U2615 ( .A(n1178), .Y(n2363) );
  AND2X1 U2616 ( .A(n2605), .B(n3662), .Y(n1185) );
  INVX1 U2617 ( .A(n1185), .Y(n2364) );
  AND2X1 U2618 ( .A(n2524), .B(n3660), .Y(n1232) );
  INVX1 U2619 ( .A(n1232), .Y(n2365) );
  AND2X1 U2620 ( .A(n2531), .B(n3660), .Y(n1241) );
  INVX1 U2621 ( .A(n1241), .Y(n2366) );
  AND2X1 U2622 ( .A(n2619), .B(n3658), .Y(n1300) );
  INVX1 U2623 ( .A(n1300), .Y(n2367) );
  AND2X1 U2624 ( .A(n2626), .B(n3658), .Y(n1309) );
  INVX1 U2625 ( .A(n1309), .Y(n2368) );
  AND2X1 U2626 ( .A(n2796), .B(n3663), .Y(n1121) );
  INVX1 U2627 ( .A(n1121), .Y(n2369) );
  AND2X1 U2628 ( .A(n2809), .B(n3663), .Y(n1134) );
  INVX1 U2629 ( .A(n1134), .Y(n2370) );
  AND2X1 U2630 ( .A(n2817), .B(n3663), .Y(n1143) );
  INVX1 U2631 ( .A(n1143), .Y(n2371) );
  AND2X1 U2632 ( .A(n3015), .B(n3661), .Y(n1191) );
  INVX1 U2633 ( .A(n1191), .Y(n2372) );
  AND2X1 U2634 ( .A(n3038), .B(n3661), .Y(n1214) );
  INVX1 U2635 ( .A(n1214), .Y(n2373) );
  AND2X1 U2636 ( .A(n2826), .B(n3659), .Y(n1256) );
  INVX1 U2637 ( .A(n1256), .Y(n2374) );
  AND2X1 U2638 ( .A(n2848), .B(n3659), .Y(n1279) );
  INVX1 U2639 ( .A(n1279), .Y(n2375) );
  AND2X1 U2640 ( .A(n3045), .B(n3657), .Y(n1325) );
  INVX1 U2641 ( .A(n1325), .Y(n2376) );
  AND2X1 U2642 ( .A(n3068), .B(n3657), .Y(n1348) );
  INVX1 U2643 ( .A(n1348), .Y(n2377) );
  AND2X1 U2644 ( .A(re), .B(empty_bar), .Y(n1364) );
  AND2X1 U2645 ( .A(n39), .B(n1084), .Y(n1358) );
  INVX1 U2646 ( .A(n1358), .Y(n2378) );
  AND2X1 U2647 ( .A(n2674), .B(n3672), .Y(n821) );
  INVX1 U2648 ( .A(n821), .Y(n2379) );
  AND2X1 U2649 ( .A(n2777), .B(n3670), .Y(n898) );
  INVX1 U2650 ( .A(n898), .Y(n2380) );
  AND2X1 U2651 ( .A(n2699), .B(n3668), .Y(n951) );
  INVX1 U2652 ( .A(n951), .Y(n2381) );
  AND2X1 U2653 ( .A(n2705), .B(n3668), .Y(n958) );
  INVX1 U2654 ( .A(n958), .Y(n2382) );
  AND2X1 U2655 ( .A(n2736), .B(n3666), .Y(n1026) );
  INVX1 U2656 ( .A(n1026), .Y(n2383) );
  AND2X1 U2657 ( .A(n2744), .B(n3666), .Y(n1034) );
  INVX1 U2658 ( .A(n1034), .Y(n2384) );
  AND2X1 U2659 ( .A(n2921), .B(n3671), .Y(n859) );
  INVX1 U2660 ( .A(n859), .Y(n2385) );
  AND2X1 U2661 ( .A(n2928), .B(n3671), .Y(n866) );
  INVX1 U2662 ( .A(n866), .Y(n2386) );
  AND2X1 U2663 ( .A(n3076), .B(n3669), .Y(n920) );
  INVX1 U2664 ( .A(n920), .Y(n2387) );
  AND2X1 U2665 ( .A(n3099), .B(n3669), .Y(n943) );
  INVX1 U2666 ( .A(n943), .Y(n2388) );
  AND2X1 U2667 ( .A(n2956), .B(n3667), .Y(n995) );
  INVX1 U2668 ( .A(n995), .Y(n2389) );
  AND2X1 U2669 ( .A(n2965), .B(n3667), .Y(n1004) );
  INVX1 U2670 ( .A(n1004), .Y(n2390) );
  AND2X1 U2671 ( .A(n2987), .B(n3665), .Y(n1062) );
  INVX1 U2672 ( .A(n1062), .Y(n2391) );
  AND2X1 U2673 ( .A(n2995), .B(n3665), .Y(n1070) );
  INVX1 U2674 ( .A(n1070), .Y(n2392) );
  AND2X1 U2675 ( .A(n2492), .B(n3664), .Y(n1087) );
  INVX1 U2676 ( .A(n1087), .Y(n2393) );
  AND2X1 U2677 ( .A(n2502), .B(n3664), .Y(n1100) );
  INVX1 U2678 ( .A(n1100), .Y(n2394) );
  AND2X1 U2679 ( .A(n2510), .B(n3664), .Y(n1109) );
  INVX1 U2680 ( .A(n1109), .Y(n2395) );
  AND2X1 U2681 ( .A(n2590), .B(n3662), .Y(n1166) );
  INVX1 U2682 ( .A(n1166), .Y(n2396) );
  AND2X1 U2683 ( .A(n2599), .B(n3662), .Y(n1175) );
  INVX1 U2684 ( .A(n1175), .Y(n2397) );
  AND2X1 U2685 ( .A(n2606), .B(n3660), .Y(n1245) );
  INVX1 U2686 ( .A(n1245), .Y(n2398) );
  AND2X1 U2687 ( .A(n2607), .B(n3660), .Y(n1252) );
  INVX1 U2688 ( .A(n1252), .Y(n2399) );
  AND2X1 U2689 ( .A(n2627), .B(n3658), .Y(n1310) );
  INVX1 U2690 ( .A(n1310), .Y(n2400) );
  AND2X1 U2691 ( .A(n2632), .B(n3658), .Y(n1318) );
  INVX1 U2692 ( .A(n1318), .Y(n2401) );
  AND2X1 U2693 ( .A(n2814), .B(n3663), .Y(n1139) );
  INVX1 U2694 ( .A(n1139), .Y(n2402) );
  AND2X1 U2695 ( .A(n2823), .B(n3663), .Y(n1149) );
  INVX1 U2696 ( .A(n1149), .Y(n2403) );
  AND2X1 U2697 ( .A(n3014), .B(n3661), .Y(n1190) );
  INVX1 U2698 ( .A(n1190), .Y(n2404) );
  AND2X1 U2699 ( .A(n3037), .B(n3661), .Y(n1213) );
  INVX1 U2700 ( .A(n1213), .Y(n2405) );
  AND2X1 U2701 ( .A(n2840), .B(n3659), .Y(n1270) );
  INVX1 U2702 ( .A(n1270), .Y(n2406) );
  AND2X1 U2703 ( .A(n2851), .B(n3659), .Y(n1282) );
  INVX1 U2704 ( .A(n1282), .Y(n2407) );
  AND2X1 U2705 ( .A(n3046), .B(n3657), .Y(n1326) );
  INVX1 U2706 ( .A(n1326), .Y(n2408) );
  AND2X1 U2707 ( .A(n3069), .B(n3657), .Y(n1349) );
  INVX1 U2708 ( .A(n1349), .Y(n2409) );
  AND2X1 U2709 ( .A(n111), .B(n1364), .Y(n1362) );
  INVX1 U2710 ( .A(n1362), .Y(n2410) );
  AND2X1 U2711 ( .A(n36), .B(n1084), .Y(n1356) );
  INVX1 U2712 ( .A(n1356), .Y(n2411) );
  AND2X1 U2713 ( .A(n37), .B(n1084), .Y(n1355) );
  INVX1 U2714 ( .A(n1355), .Y(n2412) );
  AND2X1 U2715 ( .A(we), .B(full_bar), .Y(n1084) );
  AND2X1 U2716 ( .A(n2675), .B(n3672), .Y(n822) );
  INVX1 U2717 ( .A(n822), .Y(n2413) );
  AND2X1 U2718 ( .A(n2765), .B(n3670), .Y(n885) );
  INVX1 U2719 ( .A(n885), .Y(n2414) );
  AND2X1 U2720 ( .A(n2772), .B(n3670), .Y(n892) );
  INVX1 U2721 ( .A(n892), .Y(n2415) );
  AND2X1 U2722 ( .A(n2711), .B(n3668), .Y(n964) );
  INVX1 U2723 ( .A(n964), .Y(n2416) );
  AND2X1 U2724 ( .A(n2735), .B(n3666), .Y(n1025) );
  INVX1 U2725 ( .A(n1025), .Y(n2417) );
  AND2X1 U2726 ( .A(n2742), .B(n3666), .Y(n1032) );
  INVX1 U2727 ( .A(n1032), .Y(n2418) );
  AND2X1 U2728 ( .A(n2922), .B(n3671), .Y(n860) );
  INVX1 U2729 ( .A(n860), .Y(n2419) );
  AND2X1 U2730 ( .A(n2930), .B(n3671), .Y(n868) );
  INVX1 U2731 ( .A(n868), .Y(n2420) );
  AND2X1 U2732 ( .A(n3084), .B(n3669), .Y(n928) );
  INVX1 U2733 ( .A(n928), .Y(n2421) );
  AND2X1 U2734 ( .A(n3092), .B(n3669), .Y(n936) );
  INVX1 U2735 ( .A(n936), .Y(n2422) );
  AND2X1 U2736 ( .A(n2947), .B(n3667), .Y(n986) );
  INVX1 U2737 ( .A(n986), .Y(n2423) );
  AND2X1 U2738 ( .A(n2970), .B(n3667), .Y(n1009) );
  INVX1 U2739 ( .A(n1009), .Y(n2424) );
  AND2X1 U2740 ( .A(n2988), .B(n3665), .Y(n1063) );
  INVX1 U2741 ( .A(n1063), .Y(n2425) );
  AND2X1 U2742 ( .A(n2997), .B(n3665), .Y(n1072) );
  INVX1 U2743 ( .A(n1072), .Y(n2426) );
  AND2X1 U2744 ( .A(n2500), .B(n3664), .Y(n1098) );
  INVX1 U2745 ( .A(n1098), .Y(n2427) );
  AND2X1 U2746 ( .A(n2509), .B(n3664), .Y(n1107) );
  INVX1 U2747 ( .A(n1107), .Y(n2428) );
  AND2X1 U2748 ( .A(n2581), .B(n3662), .Y(n1155) );
  INVX1 U2749 ( .A(n1155), .Y(n2429) );
  AND2X1 U2750 ( .A(n2592), .B(n3662), .Y(n1168) );
  INVX1 U2751 ( .A(n1168), .Y(n2430) );
  AND2X1 U2752 ( .A(n2600), .B(n3662), .Y(n1177) );
  INVX1 U2753 ( .A(n1177), .Y(n2431) );
  AND2X1 U2754 ( .A(n2533), .B(n3660), .Y(n1243) );
  INVX1 U2755 ( .A(n1243), .Y(n2432) );
  AND2X1 U2756 ( .A(n2537), .B(n3660), .Y(n1251) );
  INVX1 U2757 ( .A(n1251), .Y(n2433) );
  AND2X1 U2758 ( .A(n2763), .B(n3658), .Y(n1312) );
  INVX1 U2759 ( .A(n1312), .Y(n2434) );
  AND2X1 U2760 ( .A(n2764), .B(n3658), .Y(n1319) );
  INVX1 U2761 ( .A(n1319), .Y(n2435) );
  AND2X1 U2762 ( .A(n2798), .B(n3663), .Y(n1123) );
  INVX1 U2763 ( .A(n1123), .Y(n2436) );
  AND2X1 U2764 ( .A(n2820), .B(n3663), .Y(n1146) );
  INVX1 U2765 ( .A(n1146), .Y(n2437) );
  AND2X1 U2766 ( .A(n3030), .B(n3661), .Y(n1206) );
  INVX1 U2767 ( .A(n1206), .Y(n2438) );
  AND2X1 U2768 ( .A(n3040), .B(n3661), .Y(n1216) );
  INVX1 U2769 ( .A(n1216), .Y(n2439) );
  AND2X1 U2770 ( .A(n2828), .B(n3659), .Y(n1258) );
  INVX1 U2771 ( .A(n1258), .Y(n2440) );
  AND2X1 U2772 ( .A(n2850), .B(n3659), .Y(n1281) );
  INVX1 U2773 ( .A(n1281), .Y(n2441) );
  AND2X1 U2774 ( .A(n3058), .B(n3657), .Y(n1338) );
  INVX1 U2775 ( .A(n1338), .Y(n2442) );
  AND2X1 U2776 ( .A(n3070), .B(n3657), .Y(n1350) );
  INVX1 U2777 ( .A(n1350), .Y(n2443) );
  AND2X1 U2778 ( .A(n3564), .B(n3655), .Y(n1396) );
  INVX1 U2779 ( .A(n1396), .Y(n2444) );
  AND2X1 U2780 ( .A(n2676), .B(n3672), .Y(n823) );
  INVX1 U2781 ( .A(n823), .Y(n2445) );
  AND2X1 U2782 ( .A(n2774), .B(n3670), .Y(n894) );
  INVX1 U2783 ( .A(n894), .Y(n2446) );
  AND2X1 U2784 ( .A(n2781), .B(n3670), .Y(n902) );
  INVX1 U2785 ( .A(n902), .Y(n2447) );
  AND2X1 U2786 ( .A(n2706), .B(n3668), .Y(n959) );
  INVX1 U2787 ( .A(n959), .Y(n2448) );
  AND2X1 U2788 ( .A(n2712), .B(n3668), .Y(n966) );
  INVX1 U2789 ( .A(n966), .Y(n2449) );
  AND2X1 U2790 ( .A(n2737), .B(n3666), .Y(n1027) );
  INVX1 U2791 ( .A(n1027), .Y(n2450) );
  AND2X1 U2792 ( .A(n2745), .B(n3666), .Y(n1035) );
  INVX1 U2793 ( .A(n1035), .Y(n2451) );
  AND2X1 U2794 ( .A(n2925), .B(n3671), .Y(n863) );
  INVX1 U2795 ( .A(n863), .Y(n2452) );
  AND2X1 U2796 ( .A(n2934), .B(n3671), .Y(n872) );
  INVX1 U2797 ( .A(n872), .Y(n2453) );
  AND2X1 U2798 ( .A(n3085), .B(n3669), .Y(n929) );
  INVX1 U2799 ( .A(n929), .Y(n2454) );
  AND2X1 U2800 ( .A(n3094), .B(n3669), .Y(n938) );
  INVX1 U2801 ( .A(n938), .Y(n2455) );
  AND2X1 U2802 ( .A(n2948), .B(n3667), .Y(n987) );
  INVX1 U2803 ( .A(n987), .Y(n2456) );
  AND2X1 U2804 ( .A(n2971), .B(n3667), .Y(n1010) );
  INVX1 U2805 ( .A(n1010), .Y(n2457) );
  AND2X1 U2806 ( .A(n2978), .B(n3665), .Y(n1053) );
  INVX1 U2807 ( .A(n1053), .Y(n2458) );
  AND2X1 U2808 ( .A(n2991), .B(n3665), .Y(n1066) );
  INVX1 U2809 ( .A(n1066), .Y(n2459) );
  AND2X1 U2810 ( .A(n3000), .B(n3665), .Y(n1075) );
  INVX1 U2811 ( .A(n1075), .Y(n2460) );
  AND2X1 U2812 ( .A(n2582), .B(n3662), .Y(n1156) );
  INVX1 U2813 ( .A(n1156), .Y(n2461) );
  AND2X1 U2814 ( .A(n2602), .B(n3662), .Y(n1179) );
  INVX1 U2815 ( .A(n1179), .Y(n2462) );
  AND2X1 U2816 ( .A(n2759), .B(n3660), .Y(n1221) );
  INVX1 U2817 ( .A(n1221), .Y(n2463) );
  AND2X1 U2818 ( .A(n2611), .B(n3658), .Y(n1292) );
  INVX1 U2819 ( .A(n1292), .Y(n2464) );
  AND2X1 U2820 ( .A(n2631), .B(n3658), .Y(n1315) );
  INVX1 U2821 ( .A(n1315), .Y(n2465) );
  AND2X1 U2822 ( .A(n2818), .B(n3663), .Y(n1144) );
  INVX1 U2823 ( .A(n1144), .Y(n2466) );
  AND2X1 U2824 ( .A(n2824), .B(n3663), .Y(n1151) );
  INVX1 U2825 ( .A(n1151), .Y(n2467) );
  AND2X1 U2826 ( .A(n3027), .B(n3661), .Y(n1203) );
  INVX1 U2827 ( .A(n1203), .Y(n2468) );
  AND2X1 U2828 ( .A(n3039), .B(n3661), .Y(n1215) );
  INVX1 U2829 ( .A(n1215), .Y(n2469) );
  AND2X1 U2830 ( .A(n2846), .B(n3659), .Y(n1276) );
  INVX1 U2831 ( .A(n1276), .Y(n2470) );
  AND2X1 U2832 ( .A(n2853), .B(n3659), .Y(n1284) );
  INVX1 U2833 ( .A(n1284), .Y(n2471) );
  AND2X1 U2834 ( .A(n3061), .B(n3657), .Y(n1341) );
  INVX1 U2835 ( .A(n1341), .Y(n2472) );
  AND2X1 U2836 ( .A(n3071), .B(n3657), .Y(n1351) );
  INVX1 U2837 ( .A(n1351), .Y(n2473) );
  BUFX2 U2838 ( .A(n3751), .Y(full_bar) );
  BUFX2 U2839 ( .A(n3750), .Y(empty_bar) );
  BUFX2 U2840 ( .A(fifo[253]), .Y(n2476) );
  BUFX2 U2841 ( .A(fifo[252]), .Y(n2477) );
  BUFX2 U2842 ( .A(fifo[251]), .Y(n2478) );
  BUFX2 U2843 ( .A(fifo[230]), .Y(n2479) );
  BUFX2 U2844 ( .A(fifo[229]), .Y(n2480) );
  BUFX2 U2845 ( .A(fifo[228]), .Y(n2481) );
  BUFX2 U2846 ( .A(fifo[123]), .Y(n2482) );
  BUFX2 U2847 ( .A(fifo[111]), .Y(n2483) );
  BUFX2 U2848 ( .A(fifo[108]), .Y(n2484) );
  BUFX2 U2849 ( .A(fifo[100]), .Y(n2485) );
  BUFX2 U2850 ( .A(fifo[99]), .Y(n2486) );
  BUFX2 U2851 ( .A(fifo[98]), .Y(n2487) );
  BUFX2 U2852 ( .A(fifo[201]), .Y(n2488) );
  BUFX2 U2853 ( .A(fifo[193]), .Y(n2489) );
  BUFX2 U2854 ( .A(fifo[71]), .Y(n2490) );
  BUFX2 U2855 ( .A(fifo[64]), .Y(n2491) );
  BUFX2 U2856 ( .A(fifo[254]), .Y(n2492) );
  BUFX2 U2857 ( .A(fifo[250]), .Y(n2493) );
  BUFX2 U2858 ( .A(fifo[249]), .Y(n2494) );
  BUFX2 U2859 ( .A(fifo[248]), .Y(n2495) );
  BUFX2 U2860 ( .A(fifo[247]), .Y(n2496) );
  BUFX2 U2861 ( .A(fifo[246]), .Y(n2497) );
  BUFX2 U2862 ( .A(fifo[245]), .Y(n2498) );
  BUFX2 U2863 ( .A(fifo[244]), .Y(n2499) );
  BUFX2 U2864 ( .A(fifo[243]), .Y(n2500) );
  BUFX2 U2865 ( .A(fifo[242]), .Y(n2501) );
  BUFX2 U2866 ( .A(fifo[241]), .Y(n2502) );
  BUFX2 U2867 ( .A(fifo[240]), .Y(n2503) );
  BUFX2 U2868 ( .A(fifo[239]), .Y(n2504) );
  BUFX2 U2869 ( .A(fifo[238]), .Y(n2505) );
  BUFX2 U2870 ( .A(fifo[237]), .Y(n2506) );
  BUFX2 U2871 ( .A(fifo[236]), .Y(n2507) );
  BUFX2 U2872 ( .A(fifo[235]), .Y(n2508) );
  BUFX2 U2873 ( .A(fifo[234]), .Y(n2509) );
  BUFX2 U2874 ( .A(fifo[232]), .Y(n2510) );
  BUFX2 U2875 ( .A(fifo[231]), .Y(n2511) );
  BUFX2 U2876 ( .A(fifo[227]), .Y(n2512) );
  BUFX2 U2877 ( .A(fifo[226]), .Y(n2513) );
  BUFX2 U2878 ( .A(fifo[224]), .Y(n2514) );
  BUFX2 U2879 ( .A(fifo[126]), .Y(n2515) );
  BUFX2 U2880 ( .A(fifo[125]), .Y(n2516) );
  BUFX2 U2881 ( .A(fifo[124]), .Y(n2517) );
  BUFX2 U2882 ( .A(fifo[122]), .Y(n2518) );
  BUFX2 U2883 ( .A(fifo[121]), .Y(n2519) );
  BUFX2 U2884 ( .A(fifo[120]), .Y(n2520) );
  BUFX2 U2885 ( .A(fifo[119]), .Y(n2521) );
  BUFX2 U2886 ( .A(fifo[118]), .Y(n2522) );
  BUFX2 U2887 ( .A(fifo[117]), .Y(n2523) );
  BUFX2 U2888 ( .A(fifo[116]), .Y(n2524) );
  BUFX2 U2889 ( .A(fifo[115]), .Y(n2525) );
  BUFX2 U2890 ( .A(fifo[114]), .Y(n2526) );
  BUFX2 U2891 ( .A(fifo[113]), .Y(n2527) );
  BUFX2 U2892 ( .A(fifo[112]), .Y(n2528) );
  BUFX2 U2893 ( .A(fifo[110]), .Y(n2529) );
  BUFX2 U2894 ( .A(fifo[109]), .Y(n2530) );
  BUFX2 U2895 ( .A(fifo[107]), .Y(n2531) );
  BUFX2 U2896 ( .A(fifo[106]), .Y(n2532) );
  BUFX2 U2897 ( .A(fifo[105]), .Y(n2533) );
  BUFX2 U2898 ( .A(fifo[104]), .Y(n2534) );
  BUFX2 U2899 ( .A(fifo[102]), .Y(n2535) );
  BUFX2 U2900 ( .A(fifo[101]), .Y(n2536) );
  BUFX2 U2901 ( .A(fifo[97]), .Y(n2537) );
  OR2X1 U2902 ( .A(n2635), .B(n2857), .Y(n848) );
  INVX1 U2903 ( .A(n848), .Y(n2538) );
  OR2X1 U2904 ( .A(n3748), .B(n3747), .Y(n1049) );
  INVX1 U2905 ( .A(n1049), .Y(n2539) );
  AND2X1 U2906 ( .A(n1118), .B(n1219), .Y(n1153) );
  AND2X1 U2907 ( .A(n108), .B(n1364), .Y(n1361) );
  INVX1 U2908 ( .A(n1361), .Y(n2540) );
  AND2X1 U2909 ( .A(n38), .B(n1084), .Y(n1354) );
  INVX1 U2910 ( .A(n1354), .Y(n2541) );
  AND2X1 U2911 ( .A(n2681), .B(n3672), .Y(n829) );
  INVX1 U2912 ( .A(n829), .Y(n2542) );
  AND2X1 U2913 ( .A(n2773), .B(n3670), .Y(n893) );
  INVX1 U2914 ( .A(n893), .Y(n2543) );
  AND2X1 U2915 ( .A(n2779), .B(n3670), .Y(n900) );
  INVX1 U2916 ( .A(n900), .Y(n2544) );
  AND2X1 U2917 ( .A(n2707), .B(n3668), .Y(n960) );
  INVX1 U2918 ( .A(n960), .Y(n2545) );
  AND2X1 U2919 ( .A(n2714), .B(n3668), .Y(n968) );
  INVX1 U2920 ( .A(n968), .Y(n2546) );
  AND2X1 U2921 ( .A(n2738), .B(n3666), .Y(n1028) );
  INVX1 U2922 ( .A(n1028), .Y(n2547) );
  AND2X1 U2923 ( .A(n2747), .B(n3666), .Y(n1037) );
  INVX1 U2924 ( .A(n1037), .Y(n2548) );
  AND2X1 U2925 ( .A(n2923), .B(n3671), .Y(n861) );
  INVX1 U2926 ( .A(n861), .Y(n2549) );
  AND2X1 U2927 ( .A(n2931), .B(n3671), .Y(n869) );
  INVX1 U2928 ( .A(n869), .Y(n2550) );
  AND2X1 U2929 ( .A(n3075), .B(n3669), .Y(n919) );
  INVX1 U2930 ( .A(n919), .Y(n2551) );
  AND2X1 U2931 ( .A(n3088), .B(n3669), .Y(n932) );
  INVX1 U2932 ( .A(n932), .Y(n2552) );
  AND2X1 U2933 ( .A(n3097), .B(n3669), .Y(n941) );
  INVX1 U2934 ( .A(n941), .Y(n2553) );
  AND2X1 U2935 ( .A(n2957), .B(n3667), .Y(n996) );
  INVX1 U2936 ( .A(n996), .Y(n2554) );
  AND2X1 U2937 ( .A(n2966), .B(n3667), .Y(n1005) );
  INVX1 U2938 ( .A(n1005), .Y(n2555) );
  AND2X1 U2939 ( .A(n2980), .B(n3665), .Y(n1055) );
  INVX1 U2940 ( .A(n1055), .Y(n2556) );
  AND2X1 U2941 ( .A(n3003), .B(n3665), .Y(n1078) );
  INVX1 U2942 ( .A(n1078), .Y(n2557) );
  INVX1 U2943 ( .A(n1088), .Y(n2558) );
  INVX1 U2944 ( .A(n1111), .Y(n2559) );
  INVX1 U2945 ( .A(n1225), .Y(n2560) );
  INVX1 U2946 ( .A(n1248), .Y(n2561) );
  AND2X1 U2947 ( .A(n2760), .B(n3658), .Y(n1288) );
  INVX1 U2948 ( .A(n1288), .Y(n2562) );
  AND2X1 U2949 ( .A(n2811), .B(n3663), .Y(n1136) );
  INVX1 U2950 ( .A(n1136), .Y(n2563) );
  AND2X1 U2951 ( .A(n2822), .B(n3663), .Y(n1148) );
  INVX1 U2952 ( .A(n1148), .Y(n2564) );
  AND2X1 U2953 ( .A(n3035), .B(n3661), .Y(n1211) );
  INVX1 U2954 ( .A(n1211), .Y(n2565) );
  AND2X1 U2955 ( .A(n3042), .B(n3661), .Y(n1218) );
  INVX1 U2956 ( .A(n1218), .Y(n2566) );
  AND2X1 U2957 ( .A(n2843), .B(n3659), .Y(n1273) );
  INVX1 U2958 ( .A(n1273), .Y(n2567) );
  AND2X1 U2959 ( .A(n2852), .B(n3659), .Y(n1283) );
  INVX1 U2960 ( .A(n1283), .Y(n2568) );
  AND2X1 U2961 ( .A(n3064), .B(n3657), .Y(n1344) );
  INVX1 U2962 ( .A(n1344), .Y(n2569) );
  AND2X1 U2963 ( .A(n3072), .B(n3657), .Y(n1352) );
  INVX1 U2964 ( .A(n1352), .Y(n2570) );
  BUFX2 U2965 ( .A(fifo[188]), .Y(n2571) );
  BUFX2 U2966 ( .A(fifo[187]), .Y(n2572) );
  BUFX2 U2967 ( .A(fifo[165]), .Y(n2573) );
  BUFX2 U2968 ( .A(fifo[164]), .Y(n2574) );
  BUFX2 U2969 ( .A(fifo[47]), .Y(n2575) );
  BUFX2 U2970 ( .A(fifo[44]), .Y(n2576) );
  BUFX2 U2971 ( .A(fifo[35]), .Y(n2577) );
  BUFX2 U2972 ( .A(fifo[34]), .Y(n2578) );
  BUFX2 U2973 ( .A(fifo[233]), .Y(n2579) );
  BUFX2 U2974 ( .A(fifo[225]), .Y(n2580) );
  BUFX2 U2975 ( .A(fifo[190]), .Y(n2581) );
  BUFX2 U2976 ( .A(fifo[189]), .Y(n2582) );
  BUFX2 U2977 ( .A(fifo[186]), .Y(n2583) );
  BUFX2 U2978 ( .A(fifo[185]), .Y(n2584) );
  BUFX2 U2979 ( .A(fifo[184]), .Y(n2585) );
  BUFX2 U2980 ( .A(fifo[183]), .Y(n2586) );
  BUFX2 U2981 ( .A(fifo[182]), .Y(n2587) );
  BUFX2 U2982 ( .A(fifo[181]), .Y(n2588) );
  BUFX2 U2983 ( .A(fifo[180]), .Y(n2589) );
  BUFX2 U2984 ( .A(fifo[179]), .Y(n2590) );
  BUFX2 U2985 ( .A(fifo[178]), .Y(n2591) );
  BUFX2 U2986 ( .A(fifo[177]), .Y(n2592) );
  BUFX2 U2987 ( .A(fifo[176]), .Y(n2593) );
  BUFX2 U2988 ( .A(fifo[175]), .Y(n2594) );
  BUFX2 U2989 ( .A(fifo[174]), .Y(n2595) );
  BUFX2 U2990 ( .A(fifo[173]), .Y(n2596) );
  BUFX2 U2991 ( .A(fifo[172]), .Y(n2597) );
  BUFX2 U2992 ( .A(fifo[171]), .Y(n2598) );
  BUFX2 U2993 ( .A(fifo[170]), .Y(n2599) );
  BUFX2 U2994 ( .A(fifo[168]), .Y(n2600) );
  BUFX2 U2995 ( .A(fifo[167]), .Y(n2601) );
  BUFX2 U2996 ( .A(fifo[166]), .Y(n2602) );
  BUFX2 U2997 ( .A(fifo[163]), .Y(n2603) );
  BUFX2 U2998 ( .A(fifo[162]), .Y(n2604) );
  BUFX2 U2999 ( .A(fifo[160]), .Y(n2605) );
  BUFX2 U3000 ( .A(fifo[103]), .Y(n2606) );
  BUFX2 U3001 ( .A(fifo[96]), .Y(n2607) );
  BUFX2 U3002 ( .A(fifo[62]), .Y(n2608) );
  BUFX2 U3003 ( .A(fifo[61]), .Y(n2609) );
  BUFX2 U3004 ( .A(fifo[60]), .Y(n2610) );
  BUFX2 U3005 ( .A(fifo[59]), .Y(n2611) );
  BUFX2 U3006 ( .A(fifo[58]), .Y(n2612) );
  BUFX2 U3007 ( .A(fifo[57]), .Y(n2613) );
  BUFX2 U3008 ( .A(fifo[56]), .Y(n2614) );
  BUFX2 U3009 ( .A(fifo[55]), .Y(n2615) );
  BUFX2 U3010 ( .A(fifo[54]), .Y(n2616) );
  BUFX2 U3011 ( .A(fifo[53]), .Y(n2617) );
  BUFX2 U3012 ( .A(fifo[52]), .Y(n2618) );
  BUFX2 U3013 ( .A(fifo[51]), .Y(n2619) );
  BUFX2 U3014 ( .A(fifo[50]), .Y(n2620) );
  BUFX2 U3015 ( .A(fifo[49]), .Y(n2621) );
  BUFX2 U3016 ( .A(fifo[48]), .Y(n2622) );
  BUFX2 U3017 ( .A(fifo[46]), .Y(n2623) );
  BUFX2 U3018 ( .A(fifo[45]), .Y(n2624) );
  BUFX2 U3019 ( .A(fifo[43]), .Y(n2625) );
  BUFX2 U3020 ( .A(fifo[42]), .Y(n2626) );
  BUFX2 U3021 ( .A(fifo[41]), .Y(n2627) );
  BUFX2 U3022 ( .A(fifo[40]), .Y(n2628) );
  BUFX2 U3023 ( .A(fifo[38]), .Y(n2629) );
  BUFX2 U3024 ( .A(fifo[37]), .Y(n2630) );
  BUFX2 U3025 ( .A(fifo[36]), .Y(n2631) );
  BUFX2 U3026 ( .A(fifo[33]), .Y(n2632) );
  BUFX2 U3027 ( .A(wr_ptr_gray_ss[1]), .Y(n2633) );
  BUFX2 U3028 ( .A(rd_ptr_gray_ss[3]), .Y(n2634) );
  BUFX2 U3029 ( .A(wr_ptr_bin[1]), .Y(n2635) );
  AND2X1 U3030 ( .A(n1286), .B(n849), .Y(n950) );
  AND2X1 U3031 ( .A(n109), .B(n1364), .Y(n1360) );
  INVX1 U3032 ( .A(n1360), .Y(n2636) );
  AND2X1 U3033 ( .A(n2924), .B(n3671), .Y(n862) );
  INVX1 U3034 ( .A(n862), .Y(n2637) );
  AND2X1 U3035 ( .A(n2933), .B(n3671), .Y(n871) );
  INVX1 U3036 ( .A(n871), .Y(n2638) );
  AND2X1 U3037 ( .A(n3086), .B(n3669), .Y(n930) );
  INVX1 U3038 ( .A(n930), .Y(n2639) );
  AND2X1 U3039 ( .A(n3095), .B(n3669), .Y(n939) );
  INVX1 U3040 ( .A(n939), .Y(n2640) );
  AND2X1 U3041 ( .A(n2946), .B(n3667), .Y(n985) );
  INVX1 U3042 ( .A(n985), .Y(n2641) );
  AND2X1 U3043 ( .A(n2959), .B(n3667), .Y(n998) );
  INVX1 U3044 ( .A(n998), .Y(n2642) );
  AND2X1 U3045 ( .A(n2968), .B(n3667), .Y(n1007) );
  INVX1 U3046 ( .A(n1007), .Y(n2643) );
  AND2X1 U3047 ( .A(n2979), .B(n3665), .Y(n1054) );
  INVX1 U3048 ( .A(n1054), .Y(n2644) );
  AND2X1 U3049 ( .A(n3002), .B(n3665), .Y(n1077) );
  INVX1 U3050 ( .A(n1077), .Y(n2645) );
  INVX1 U3051 ( .A(n1090), .Y(n2646) );
  INVX1 U3052 ( .A(n1113), .Y(n2647) );
  INVX1 U3053 ( .A(n1157), .Y(n2648) );
  INVX1 U3054 ( .A(n1180), .Y(n2649) );
  INVX1 U3055 ( .A(n1240), .Y(n2650) );
  INVX1 U3056 ( .A(n1250), .Y(n2651) );
  INVX1 U3057 ( .A(n1304), .Y(n2652) );
  INVX1 U3058 ( .A(n1316), .Y(n2653) );
  AND2X1 U3059 ( .A(n3033), .B(n3661), .Y(n1209) );
  INVX1 U3060 ( .A(n1209), .Y(n2654) );
  AND2X1 U3061 ( .A(n3041), .B(n3661), .Y(n1217) );
  INVX1 U3062 ( .A(n1217), .Y(n2655) );
  AND2X1 U3063 ( .A(n3010), .B(n3659), .Y(n1254) );
  INVX1 U3064 ( .A(n1254), .Y(n2656) );
  AND2X1 U3065 ( .A(n3066), .B(n3657), .Y(n1346) );
  INVX1 U3066 ( .A(n1346), .Y(n2657) );
  AND2X1 U3067 ( .A(n3073), .B(n3657), .Y(n1353) );
  INVX1 U3068 ( .A(n1353), .Y(n2658) );
  AND2X1 U3069 ( .A(n3746), .B(n1084), .Y(n1357) );
  INVX1 U3070 ( .A(n1357), .Y(n2659) );
  BUFX2 U3071 ( .A(fifo[500]), .Y(n2660) );
  BUFX2 U3072 ( .A(fifo[491]), .Y(n2661) );
  BUFX2 U3073 ( .A(fifo[382]), .Y(n2662) );
  BUFX2 U3074 ( .A(fifo[369]), .Y(n2663) );
  BUFX2 U3075 ( .A(fifo[360]), .Y(n2664) );
  BUFX2 U3076 ( .A(fifo[317]), .Y(n2665) );
  BUFX2 U3077 ( .A(fifo[294]), .Y(n2666) );
  BUFX2 U3078 ( .A(fifo[435]), .Y(n2667) );
  BUFX2 U3079 ( .A(fifo[426]), .Y(n2668) );
  BUFX2 U3080 ( .A(fifo[511]), .Y(n2669) );
  BUFX2 U3081 ( .A(fifo[510]), .Y(n2670) );
  BUFX2 U3082 ( .A(fifo[509]), .Y(n2671) );
  BUFX2 U3083 ( .A(fifo[508]), .Y(n2672) );
  BUFX2 U3084 ( .A(fifo[507]), .Y(n2673) );
  BUFX2 U3085 ( .A(fifo[506]), .Y(n2674) );
  BUFX2 U3086 ( .A(fifo[505]), .Y(n2675) );
  BUFX2 U3087 ( .A(fifo[504]), .Y(n2676) );
  BUFX2 U3088 ( .A(fifo[503]), .Y(n2677) );
  BUFX2 U3089 ( .A(fifo[502]), .Y(n2678) );
  BUFX2 U3090 ( .A(fifo[501]), .Y(n2679) );
  BUFX2 U3091 ( .A(fifo[499]), .Y(n2680) );
  BUFX2 U3092 ( .A(fifo[498]), .Y(n2681) );
  BUFX2 U3093 ( .A(fifo[497]), .Y(n2682) );
  BUFX2 U3094 ( .A(fifo[496]), .Y(n2683) );
  BUFX2 U3095 ( .A(fifo[495]), .Y(n2684) );
  BUFX2 U3096 ( .A(fifo[494]), .Y(n2685) );
  BUFX2 U3097 ( .A(fifo[493]), .Y(n2686) );
  BUFX2 U3098 ( .A(fifo[492]), .Y(n2687) );
  BUFX2 U3099 ( .A(fifo[490]), .Y(n2688) );
  BUFX2 U3100 ( .A(fifo[489]), .Y(n2689) );
  BUFX2 U3101 ( .A(fifo[488]), .Y(n2690) );
  BUFX2 U3102 ( .A(fifo[487]), .Y(n2691) );
  BUFX2 U3103 ( .A(fifo[486]), .Y(n2692) );
  BUFX2 U3104 ( .A(fifo[485]), .Y(n2693) );
  BUFX2 U3105 ( .A(fifo[484]), .Y(n2694) );
  BUFX2 U3106 ( .A(fifo[483]), .Y(n2695) );
  BUFX2 U3107 ( .A(fifo[482]), .Y(n2696) );
  BUFX2 U3108 ( .A(fifo[481]), .Y(n2697) );
  BUFX2 U3109 ( .A(fifo[480]), .Y(n2698) );
  BUFX2 U3110 ( .A(fifo[383]), .Y(n2699) );
  BUFX2 U3111 ( .A(fifo[381]), .Y(n2700) );
  BUFX2 U3112 ( .A(fifo[380]), .Y(n2701) );
  BUFX2 U3113 ( .A(fifo[379]), .Y(n2702) );
  BUFX2 U3114 ( .A(fifo[378]), .Y(n2703) );
  BUFX2 U3115 ( .A(fifo[377]), .Y(n2704) );
  BUFX2 U3116 ( .A(fifo[376]), .Y(n2705) );
  BUFX2 U3117 ( .A(fifo[375]), .Y(n2706) );
  BUFX2 U3118 ( .A(fifo[374]), .Y(n2707) );
  BUFX2 U3119 ( .A(fifo[373]), .Y(n2708) );
  BUFX2 U3120 ( .A(fifo[372]), .Y(n2709) );
  BUFX2 U3121 ( .A(fifo[371]), .Y(n2710) );
  BUFX2 U3122 ( .A(fifo[370]), .Y(n2711) );
  BUFX2 U3123 ( .A(fifo[368]), .Y(n2712) );
  BUFX2 U3124 ( .A(fifo[367]), .Y(n2713) );
  BUFX2 U3125 ( .A(fifo[366]), .Y(n2714) );
  BUFX2 U3126 ( .A(fifo[365]), .Y(n2715) );
  BUFX2 U3127 ( .A(fifo[364]), .Y(n2716) );
  BUFX2 U3128 ( .A(fifo[363]), .Y(n2717) );
  BUFX2 U3129 ( .A(fifo[362]), .Y(n2718) );
  BUFX2 U3130 ( .A(fifo[361]), .Y(n2719) );
  BUFX2 U3131 ( .A(fifo[359]), .Y(n2720) );
  BUFX2 U3132 ( .A(fifo[358]), .Y(n2721) );
  BUFX2 U3133 ( .A(fifo[357]), .Y(n2722) );
  BUFX2 U3134 ( .A(fifo[356]), .Y(n2723) );
  BUFX2 U3135 ( .A(fifo[355]), .Y(n2724) );
  BUFX2 U3136 ( .A(fifo[354]), .Y(n2725) );
  BUFX2 U3137 ( .A(fifo[353]), .Y(n2726) );
  BUFX2 U3138 ( .A(fifo[352]), .Y(n2727) );
  BUFX2 U3139 ( .A(fifo[319]), .Y(n2728) );
  BUFX2 U3140 ( .A(fifo[318]), .Y(n2729) );
  BUFX2 U3141 ( .A(fifo[316]), .Y(n2730) );
  BUFX2 U3142 ( .A(fifo[315]), .Y(n2731) );
  BUFX2 U3143 ( .A(fifo[314]), .Y(n2732) );
  BUFX2 U3144 ( .A(fifo[313]), .Y(n2733) );
  BUFX2 U3145 ( .A(fifo[312]), .Y(n2734) );
  BUFX2 U3146 ( .A(fifo[311]), .Y(n2735) );
  BUFX2 U3147 ( .A(fifo[310]), .Y(n2736) );
  BUFX2 U3148 ( .A(fifo[309]), .Y(n2737) );
  BUFX2 U3149 ( .A(fifo[308]), .Y(n2738) );
  BUFX2 U3150 ( .A(fifo[307]), .Y(n2739) );
  BUFX2 U3151 ( .A(fifo[306]), .Y(n2740) );
  BUFX2 U3152 ( .A(fifo[305]), .Y(n2741) );
  BUFX2 U3153 ( .A(fifo[304]), .Y(n2742) );
  BUFX2 U3154 ( .A(fifo[303]), .Y(n2743) );
  BUFX2 U3155 ( .A(fifo[302]), .Y(n2744) );
  BUFX2 U3156 ( .A(fifo[301]), .Y(n2745) );
  BUFX2 U3157 ( .A(fifo[300]), .Y(n2746) );
  BUFX2 U3158 ( .A(fifo[299]), .Y(n2747) );
  BUFX2 U3159 ( .A(fifo[298]), .Y(n2748) );
  BUFX2 U3160 ( .A(fifo[297]), .Y(n2749) );
  BUFX2 U3161 ( .A(fifo[296]), .Y(n2750) );
  BUFX2 U3162 ( .A(fifo[295]), .Y(n2751) );
  BUFX2 U3163 ( .A(fifo[293]), .Y(n2752) );
  BUFX2 U3164 ( .A(fifo[292]), .Y(n2753) );
  BUFX2 U3165 ( .A(fifo[291]), .Y(n2754) );
  BUFX2 U3166 ( .A(fifo[290]), .Y(n2755) );
  BUFX2 U3167 ( .A(fifo[289]), .Y(n2756) );
  BUFX2 U3168 ( .A(fifo[288]), .Y(n2757) );
  BUFX2 U3169 ( .A(fifo[255]), .Y(n2758) );
  BUFX2 U3170 ( .A(fifo[127]), .Y(n2759) );
  BUFX2 U3171 ( .A(fifo[63]), .Y(n2760) );
  BUFX2 U3172 ( .A(fifo[169]), .Y(n2761) );
  BUFX2 U3173 ( .A(fifo[161]), .Y(n2762) );
  BUFX2 U3174 ( .A(fifo[39]), .Y(n2763) );
  BUFX2 U3175 ( .A(fifo[32]), .Y(n2764) );
  BUFX2 U3176 ( .A(fifo[447]), .Y(n2765) );
  BUFX2 U3177 ( .A(fifo[446]), .Y(n2766) );
  BUFX2 U3178 ( .A(fifo[445]), .Y(n2767) );
  BUFX2 U3179 ( .A(fifo[444]), .Y(n2768) );
  BUFX2 U3180 ( .A(fifo[443]), .Y(n2769) );
  BUFX2 U3181 ( .A(fifo[442]), .Y(n2770) );
  BUFX2 U3182 ( .A(fifo[441]), .Y(n2771) );
  BUFX2 U3183 ( .A(fifo[440]), .Y(n2772) );
  BUFX2 U3184 ( .A(fifo[439]), .Y(n2773) );
  BUFX2 U3185 ( .A(fifo[438]), .Y(n2774) );
  BUFX2 U3186 ( .A(fifo[437]), .Y(n2775) );
  BUFX2 U3187 ( .A(fifo[436]), .Y(n2776) );
  BUFX2 U3188 ( .A(fifo[434]), .Y(n2777) );
  BUFX2 U3189 ( .A(fifo[433]), .Y(n2778) );
  BUFX2 U3190 ( .A(fifo[432]), .Y(n2779) );
  BUFX2 U3191 ( .A(fifo[431]), .Y(n2780) );
  BUFX2 U3192 ( .A(fifo[430]), .Y(n2781) );
  BUFX2 U3193 ( .A(fifo[429]), .Y(n2782) );
  BUFX2 U3194 ( .A(fifo[428]), .Y(n2783) );
  BUFX2 U3195 ( .A(fifo[427]), .Y(n2784) );
  BUFX2 U3196 ( .A(fifo[425]), .Y(n2785) );
  BUFX2 U3197 ( .A(fifo[424]), .Y(n2786) );
  BUFX2 U3198 ( .A(fifo[423]), .Y(n2787) );
  BUFX2 U3199 ( .A(fifo[422]), .Y(n2788) );
  BUFX2 U3200 ( .A(fifo[421]), .Y(n2789) );
  BUFX2 U3201 ( .A(fifo[420]), .Y(n2790) );
  BUFX2 U3202 ( .A(fifo[419]), .Y(n2791) );
  BUFX2 U3203 ( .A(fifo[418]), .Y(n2792) );
  BUFX2 U3204 ( .A(fifo[417]), .Y(n2793) );
  BUFX2 U3205 ( .A(fifo[416]), .Y(n2794) );
  BUFX2 U3206 ( .A(fifo[191]), .Y(n2795) );
  BUFX2 U3207 ( .A(fifo[222]), .Y(n2796) );
  BUFX2 U3208 ( .A(fifo[221]), .Y(n2797) );
  BUFX2 U3209 ( .A(fifo[220]), .Y(n2798) );
  BUFX2 U3210 ( .A(fifo[219]), .Y(n2799) );
  BUFX2 U3211 ( .A(fifo[218]), .Y(n2800) );
  BUFX2 U3212 ( .A(fifo[217]), .Y(n2801) );
  BUFX2 U3213 ( .A(fifo[216]), .Y(n2802) );
  BUFX2 U3214 ( .A(fifo[215]), .Y(n2803) );
  BUFX2 U3215 ( .A(fifo[214]), .Y(n2804) );
  BUFX2 U3216 ( .A(fifo[213]), .Y(n2805) );
  BUFX2 U3217 ( .A(fifo[212]), .Y(n2806) );
  BUFX2 U3218 ( .A(fifo[211]), .Y(n2807) );
  BUFX2 U3219 ( .A(fifo[210]), .Y(n2808) );
  BUFX2 U3220 ( .A(fifo[209]), .Y(n2809) );
  BUFX2 U3221 ( .A(fifo[208]), .Y(n2810) );
  BUFX2 U3222 ( .A(fifo[207]), .Y(n2811) );
  BUFX2 U3223 ( .A(fifo[206]), .Y(n2812) );
  BUFX2 U3224 ( .A(fifo[205]), .Y(n2813) );
  BUFX2 U3225 ( .A(fifo[204]), .Y(n2814) );
  BUFX2 U3226 ( .A(fifo[203]), .Y(n2815) );
  BUFX2 U3227 ( .A(fifo[202]), .Y(n2816) );
  BUFX2 U3228 ( .A(fifo[200]), .Y(n2817) );
  BUFX2 U3229 ( .A(fifo[199]), .Y(n2818) );
  BUFX2 U3230 ( .A(fifo[198]), .Y(n2819) );
  BUFX2 U3231 ( .A(fifo[197]), .Y(n2820) );
  BUFX2 U3232 ( .A(fifo[196]), .Y(n2821) );
  BUFX2 U3233 ( .A(fifo[195]), .Y(n2822) );
  BUFX2 U3234 ( .A(fifo[194]), .Y(n2823) );
  BUFX2 U3235 ( .A(fifo[192]), .Y(n2824) );
  BUFX2 U3236 ( .A(fifo[94]), .Y(n2825) );
  BUFX2 U3237 ( .A(fifo[93]), .Y(n2826) );
  BUFX2 U3238 ( .A(fifo[92]), .Y(n2827) );
  BUFX2 U3239 ( .A(fifo[91]), .Y(n2828) );
  BUFX2 U3240 ( .A(fifo[90]), .Y(n2829) );
  BUFX2 U3241 ( .A(fifo[89]), .Y(n2830) );
  BUFX2 U3242 ( .A(fifo[88]), .Y(n2831) );
  BUFX2 U3243 ( .A(fifo[87]), .Y(n2832) );
  BUFX2 U3244 ( .A(fifo[86]), .Y(n2833) );
  BUFX2 U3245 ( .A(fifo[85]), .Y(n2834) );
  BUFX2 U3246 ( .A(fifo[84]), .Y(n2835) );
  BUFX2 U3247 ( .A(fifo[83]), .Y(n2836) );
  BUFX2 U3248 ( .A(fifo[82]), .Y(n2837) );
  BUFX2 U3249 ( .A(fifo[81]), .Y(n2838) );
  BUFX2 U3250 ( .A(fifo[80]), .Y(n2839) );
  BUFX2 U3251 ( .A(fifo[79]), .Y(n2840) );
  BUFX2 U3252 ( .A(fifo[78]), .Y(n2841) );
  BUFX2 U3253 ( .A(fifo[77]), .Y(n2842) );
  BUFX2 U3254 ( .A(fifo[76]), .Y(n2843) );
  BUFX2 U3255 ( .A(fifo[75]), .Y(n2844) );
  BUFX2 U3256 ( .A(fifo[74]), .Y(n2845) );
  BUFX2 U3257 ( .A(fifo[73]), .Y(n2846) );
  BUFX2 U3258 ( .A(fifo[72]), .Y(n2847) );
  BUFX2 U3259 ( .A(fifo[70]), .Y(n2848) );
  BUFX2 U3260 ( .A(fifo[69]), .Y(n2849) );
  BUFX2 U3261 ( .A(fifo[68]), .Y(n2850) );
  BUFX2 U3262 ( .A(fifo[67]), .Y(n2851) );
  BUFX2 U3263 ( .A(fifo[66]), .Y(n2852) );
  BUFX2 U3264 ( .A(fifo[65]), .Y(n2853) );
  BUFX2 U3265 ( .A(rd_ptr_gray_ss[1]), .Y(n2854) );
  BUFX2 U3266 ( .A(wr_ptr_gray_ss[2]), .Y(n2855) );
  BUFX2 U3267 ( .A(wr_ptr_bin[4]), .Y(n2856) );
  BUFX2 U3268 ( .A(wr_ptr_bin[2]), .Y(n2857) );
  AND2X1 U3269 ( .A(n110), .B(n1364), .Y(n1359) );
  INVX1 U3270 ( .A(n1359), .Y(n2858) );
  INVX1 U3271 ( .A(n827), .Y(n2859) );
  INVX1 U3272 ( .A(n836), .Y(n2860) );
  INVX1 U3273 ( .A(n897), .Y(n2861) );
  INVX1 U3274 ( .A(n906), .Y(n2862) );
  INVX1 U3275 ( .A(n952), .Y(n2863) );
  INVX1 U3276 ( .A(n965), .Y(n2864) );
  INVX1 U3277 ( .A(n974), .Y(n2865) );
  INVX1 U3278 ( .A(n1019), .Y(n2866) );
  INVX1 U3279 ( .A(n1042), .Y(n2867) );
  INVX1 U3280 ( .A(n1089), .Y(n2868) );
  INVX1 U3281 ( .A(n1112), .Y(n2869) );
  INVX1 U3282 ( .A(n1158), .Y(n2870) );
  INVX1 U3283 ( .A(n1181), .Y(n2871) );
  INVX1 U3284 ( .A(n1237), .Y(n2872) );
  INVX1 U3285 ( .A(n1249), .Y(n2873) );
  INVX1 U3286 ( .A(n1307), .Y(n2874) );
  INVX1 U3287 ( .A(n1317), .Y(n2875) );
  INVX1 U3288 ( .A(n1142), .Y(n2876) );
  INVX1 U3289 ( .A(n1150), .Y(n2877) );
  INVX1 U3290 ( .A(n1278), .Y(n2878) );
  INVX1 U3291 ( .A(n1285), .Y(n2879) );
  BUFX2 U3292 ( .A(rd_ptr_gray_ss[0]), .Y(n2880) );
  BUFX2 U3293 ( .A(n3783), .Y(data_out[0]) );
  BUFX2 U3294 ( .A(n3782), .Y(data_out[1]) );
  BUFX2 U3295 ( .A(n3781), .Y(data_out[2]) );
  BUFX2 U3296 ( .A(n3780), .Y(data_out[3]) );
  BUFX2 U3297 ( .A(n3779), .Y(data_out[4]) );
  BUFX2 U3298 ( .A(n3778), .Y(data_out[5]) );
  BUFX2 U3299 ( .A(n3777), .Y(data_out[6]) );
  BUFX2 U3300 ( .A(n3776), .Y(data_out[7]) );
  BUFX2 U3301 ( .A(n3775), .Y(data_out[8]) );
  BUFX2 U3302 ( .A(n3774), .Y(data_out[9]) );
  BUFX2 U3303 ( .A(n3773), .Y(data_out[10]) );
  BUFX2 U3304 ( .A(n3772), .Y(data_out[11]) );
  BUFX2 U3305 ( .A(n3771), .Y(data_out[12]) );
  BUFX2 U3306 ( .A(n3770), .Y(data_out[13]) );
  BUFX2 U3307 ( .A(n3769), .Y(data_out[14]) );
  BUFX2 U3308 ( .A(n3768), .Y(data_out[15]) );
  BUFX2 U3309 ( .A(n3767), .Y(data_out[16]) );
  BUFX2 U3310 ( .A(n3766), .Y(data_out[17]) );
  BUFX2 U3311 ( .A(n3765), .Y(data_out[18]) );
  BUFX2 U3312 ( .A(n3764), .Y(data_out[19]) );
  BUFX2 U3313 ( .A(n3763), .Y(data_out[20]) );
  BUFX2 U3314 ( .A(n3762), .Y(data_out[21]) );
  BUFX2 U3315 ( .A(n3761), .Y(data_out[22]) );
  BUFX2 U3316 ( .A(n3760), .Y(data_out[23]) );
  BUFX2 U3317 ( .A(n3759), .Y(data_out[24]) );
  BUFX2 U3318 ( .A(n3758), .Y(data_out[25]) );
  BUFX2 U3319 ( .A(n3757), .Y(data_out[26]) );
  BUFX2 U3320 ( .A(n3756), .Y(data_out[27]) );
  BUFX2 U3321 ( .A(n3755), .Y(data_out[28]) );
  BUFX2 U3322 ( .A(n3754), .Y(data_out[29]) );
  BUFX2 U3323 ( .A(n3753), .Y(data_out[30]) );
  BUFX2 U3324 ( .A(n3752), .Y(data_out[31]) );
  BUFX2 U3325 ( .A(fifo[479]), .Y(n2913) );
  BUFX2 U3326 ( .A(fifo[478]), .Y(n2914) );
  BUFX2 U3327 ( .A(fifo[477]), .Y(n2915) );
  BUFX2 U3328 ( .A(fifo[476]), .Y(n2916) );
  BUFX2 U3329 ( .A(fifo[475]), .Y(n2917) );
  BUFX2 U3330 ( .A(fifo[474]), .Y(n2918) );
  BUFX2 U3331 ( .A(fifo[473]), .Y(n2919) );
  BUFX2 U3332 ( .A(fifo[472]), .Y(n2920) );
  BUFX2 U3333 ( .A(fifo[471]), .Y(n2921) );
  BUFX2 U3334 ( .A(fifo[470]), .Y(n2922) );
  BUFX2 U3335 ( .A(fifo[469]), .Y(n2923) );
  BUFX2 U3336 ( .A(fifo[468]), .Y(n2924) );
  BUFX2 U3337 ( .A(fifo[467]), .Y(n2925) );
  BUFX2 U3338 ( .A(fifo[466]), .Y(n2926) );
  BUFX2 U3339 ( .A(fifo[465]), .Y(n2927) );
  BUFX2 U3340 ( .A(fifo[464]), .Y(n2928) );
  BUFX2 U3341 ( .A(fifo[463]), .Y(n2929) );
  BUFX2 U3342 ( .A(fifo[462]), .Y(n2930) );
  BUFX2 U3343 ( .A(fifo[461]), .Y(n2931) );
  BUFX2 U3344 ( .A(fifo[460]), .Y(n2932) );
  BUFX2 U3345 ( .A(fifo[459]), .Y(n2933) );
  BUFX2 U3346 ( .A(fifo[458]), .Y(n2934) );
  BUFX2 U3347 ( .A(fifo[457]), .Y(n2935) );
  BUFX2 U3348 ( .A(fifo[456]), .Y(n2936) );
  BUFX2 U3349 ( .A(fifo[455]), .Y(n2937) );
  BUFX2 U3350 ( .A(fifo[454]), .Y(n2938) );
  BUFX2 U3351 ( .A(fifo[453]), .Y(n2939) );
  BUFX2 U3352 ( .A(fifo[452]), .Y(n2940) );
  BUFX2 U3353 ( .A(fifo[451]), .Y(n2941) );
  BUFX2 U3354 ( .A(fifo[450]), .Y(n2942) );
  BUFX2 U3355 ( .A(fifo[449]), .Y(n2943) );
  BUFX2 U3356 ( .A(fifo[448]), .Y(n2944) );
  BUFX2 U3357 ( .A(fifo[351]), .Y(n2945) );
  BUFX2 U3358 ( .A(fifo[350]), .Y(n2946) );
  BUFX2 U3359 ( .A(fifo[349]), .Y(n2947) );
  BUFX2 U3360 ( .A(fifo[348]), .Y(n2948) );
  BUFX2 U3361 ( .A(fifo[347]), .Y(n2949) );
  BUFX2 U3362 ( .A(fifo[346]), .Y(n2950) );
  BUFX2 U3363 ( .A(fifo[345]), .Y(n2951) );
  BUFX2 U3364 ( .A(fifo[344]), .Y(n2952) );
  BUFX2 U3365 ( .A(fifo[343]), .Y(n2953) );
  BUFX2 U3366 ( .A(fifo[342]), .Y(n2954) );
  BUFX2 U3367 ( .A(fifo[341]), .Y(n2955) );
  BUFX2 U3368 ( .A(fifo[340]), .Y(n2956) );
  BUFX2 U3369 ( .A(fifo[339]), .Y(n2957) );
  BUFX2 U3370 ( .A(fifo[338]), .Y(n2958) );
  BUFX2 U3371 ( .A(fifo[337]), .Y(n2959) );
  BUFX2 U3372 ( .A(fifo[336]), .Y(n2960) );
  BUFX2 U3373 ( .A(fifo[335]), .Y(n2961) );
  BUFX2 U3374 ( .A(fifo[334]), .Y(n2962) );
  BUFX2 U3375 ( .A(fifo[333]), .Y(n2963) );
  BUFX2 U3376 ( .A(fifo[332]), .Y(n2964) );
  BUFX2 U3377 ( .A(fifo[331]), .Y(n2965) );
  BUFX2 U3378 ( .A(fifo[330]), .Y(n2966) );
  BUFX2 U3379 ( .A(fifo[329]), .Y(n2967) );
  BUFX2 U3380 ( .A(fifo[328]), .Y(n2968) );
  BUFX2 U3381 ( .A(fifo[327]), .Y(n2969) );
  BUFX2 U3382 ( .A(fifo[326]), .Y(n2970) );
  BUFX2 U3383 ( .A(fifo[325]), .Y(n2971) );
  BUFX2 U3384 ( .A(fifo[324]), .Y(n2972) );
  BUFX2 U3385 ( .A(fifo[323]), .Y(n2973) );
  BUFX2 U3386 ( .A(fifo[322]), .Y(n2974) );
  BUFX2 U3387 ( .A(fifo[321]), .Y(n2975) );
  BUFX2 U3388 ( .A(fifo[320]), .Y(n2976) );
  BUFX2 U3389 ( .A(fifo[287]), .Y(n2977) );
  BUFX2 U3390 ( .A(fifo[286]), .Y(n2978) );
  BUFX2 U3391 ( .A(fifo[285]), .Y(n2979) );
  BUFX2 U3392 ( .A(fifo[284]), .Y(n2980) );
  BUFX2 U3393 ( .A(fifo[283]), .Y(n2981) );
  BUFX2 U3394 ( .A(fifo[282]), .Y(n2982) );
  BUFX2 U3395 ( .A(fifo[281]), .Y(n2983) );
  BUFX2 U3396 ( .A(fifo[280]), .Y(n2984) );
  BUFX2 U3397 ( .A(fifo[279]), .Y(n2985) );
  BUFX2 U3398 ( .A(fifo[278]), .Y(n2986) );
  BUFX2 U3399 ( .A(fifo[277]), .Y(n2987) );
  BUFX2 U3400 ( .A(fifo[276]), .Y(n2988) );
  BUFX2 U3401 ( .A(fifo[275]), .Y(n2989) );
  BUFX2 U3402 ( .A(fifo[274]), .Y(n2990) );
  BUFX2 U3403 ( .A(fifo[273]), .Y(n2991) );
  BUFX2 U3404 ( .A(fifo[272]), .Y(n2992) );
  BUFX2 U3405 ( .A(fifo[271]), .Y(n2993) );
  BUFX2 U3406 ( .A(fifo[270]), .Y(n2994) );
  BUFX2 U3407 ( .A(fifo[269]), .Y(n2995) );
  BUFX2 U3408 ( .A(fifo[268]), .Y(n2996) );
  BUFX2 U3409 ( .A(fifo[267]), .Y(n2997) );
  BUFX2 U3410 ( .A(fifo[266]), .Y(n2998) );
  BUFX2 U3411 ( .A(fifo[265]), .Y(n2999) );
  BUFX2 U3412 ( .A(fifo[264]), .Y(n3000) );
  BUFX2 U3413 ( .A(fifo[263]), .Y(n3001) );
  BUFX2 U3414 ( .A(fifo[262]), .Y(n3002) );
  BUFX2 U3415 ( .A(fifo[261]), .Y(n3003) );
  BUFX2 U3416 ( .A(fifo[260]), .Y(n3004) );
  BUFX2 U3417 ( .A(fifo[259]), .Y(n3005) );
  BUFX2 U3418 ( .A(fifo[258]), .Y(n3006) );
  BUFX2 U3419 ( .A(fifo[257]), .Y(n3007) );
  BUFX2 U3420 ( .A(fifo[256]), .Y(n3008) );
  BUFX2 U3421 ( .A(fifo[223]), .Y(n3009) );
  BUFX2 U3422 ( .A(fifo[95]), .Y(n3010) );
  BUFX2 U3423 ( .A(fifo[31]), .Y(n3011) );
  BUFX2 U3424 ( .A(fifo[158]), .Y(n3012) );
  BUFX2 U3425 ( .A(fifo[157]), .Y(n3013) );
  BUFX2 U3426 ( .A(fifo[156]), .Y(n3014) );
  BUFX2 U3427 ( .A(fifo[155]), .Y(n3015) );
  BUFX2 U3428 ( .A(fifo[154]), .Y(n3016) );
  BUFX2 U3429 ( .A(fifo[153]), .Y(n3017) );
  BUFX2 U3430 ( .A(fifo[152]), .Y(n3018) );
  BUFX2 U3431 ( .A(fifo[151]), .Y(n3019) );
  BUFX2 U3432 ( .A(fifo[150]), .Y(n3020) );
  BUFX2 U3433 ( .A(fifo[149]), .Y(n3021) );
  BUFX2 U3434 ( .A(fifo[148]), .Y(n3022) );
  BUFX2 U3435 ( .A(fifo[147]), .Y(n3023) );
  BUFX2 U3436 ( .A(fifo[146]), .Y(n3024) );
  BUFX2 U3437 ( .A(fifo[145]), .Y(n3025) );
  BUFX2 U3438 ( .A(fifo[144]), .Y(n3026) );
  BUFX2 U3439 ( .A(fifo[143]), .Y(n3027) );
  BUFX2 U3440 ( .A(fifo[142]), .Y(n3028) );
  BUFX2 U3441 ( .A(fifo[141]), .Y(n3029) );
  BUFX2 U3442 ( .A(fifo[140]), .Y(n3030) );
  BUFX2 U3443 ( .A(fifo[139]), .Y(n3031) );
  BUFX2 U3444 ( .A(fifo[138]), .Y(n3032) );
  BUFX2 U3445 ( .A(fifo[137]), .Y(n3033) );
  BUFX2 U3446 ( .A(fifo[136]), .Y(n3034) );
  BUFX2 U3447 ( .A(fifo[135]), .Y(n3035) );
  BUFX2 U3448 ( .A(fifo[134]), .Y(n3036) );
  BUFX2 U3449 ( .A(fifo[133]), .Y(n3037) );
  BUFX2 U3450 ( .A(fifo[132]), .Y(n3038) );
  BUFX2 U3451 ( .A(fifo[131]), .Y(n3039) );
  BUFX2 U3452 ( .A(fifo[130]), .Y(n3040) );
  BUFX2 U3453 ( .A(fifo[129]), .Y(n3041) );
  BUFX2 U3454 ( .A(fifo[128]), .Y(n3042) );
  BUFX2 U3455 ( .A(fifo[30]), .Y(n3043) );
  BUFX2 U3456 ( .A(fifo[29]), .Y(n3044) );
  BUFX2 U3457 ( .A(fifo[28]), .Y(n3045) );
  BUFX2 U3458 ( .A(fifo[27]), .Y(n3046) );
  BUFX2 U3459 ( .A(fifo[26]), .Y(n3047) );
  BUFX2 U3460 ( .A(fifo[25]), .Y(n3048) );
  BUFX2 U3461 ( .A(fifo[24]), .Y(n3049) );
  BUFX2 U3462 ( .A(fifo[23]), .Y(n3050) );
  BUFX2 U3463 ( .A(fifo[22]), .Y(n3051) );
  BUFX2 U3464 ( .A(fifo[21]), .Y(n3052) );
  BUFX2 U3465 ( .A(fifo[20]), .Y(n3053) );
  BUFX2 U3466 ( .A(fifo[19]), .Y(n3054) );
  BUFX2 U3467 ( .A(fifo[18]), .Y(n3055) );
  BUFX2 U3468 ( .A(fifo[17]), .Y(n3056) );
  BUFX2 U3469 ( .A(fifo[16]), .Y(n3057) );
  BUFX2 U3470 ( .A(fifo[15]), .Y(n3058) );
  BUFX2 U3471 ( .A(fifo[14]), .Y(n3059) );
  BUFX2 U3472 ( .A(fifo[13]), .Y(n3060) );
  BUFX2 U3473 ( .A(fifo[12]), .Y(n3061) );
  BUFX2 U3474 ( .A(fifo[11]), .Y(n3062) );
  BUFX2 U3475 ( .A(fifo[10]), .Y(n3063) );
  BUFX2 U3476 ( .A(fifo[9]), .Y(n3064) );
  BUFX2 U3477 ( .A(fifo[8]), .Y(n3065) );
  BUFX2 U3478 ( .A(fifo[7]), .Y(n3066) );
  BUFX2 U3479 ( .A(fifo[6]), .Y(n3067) );
  BUFX2 U3480 ( .A(fifo[5]), .Y(n3068) );
  BUFX2 U3481 ( .A(fifo[4]), .Y(n3069) );
  BUFX2 U3482 ( .A(fifo[3]), .Y(n3070) );
  BUFX2 U3483 ( .A(fifo[2]), .Y(n3071) );
  BUFX2 U3484 ( .A(fifo[1]), .Y(n3072) );
  BUFX2 U3485 ( .A(fifo[0]), .Y(n3073) );
  BUFX2 U3486 ( .A(fifo[415]), .Y(n3074) );
  BUFX2 U3487 ( .A(fifo[414]), .Y(n3075) );
  BUFX2 U3488 ( .A(fifo[413]), .Y(n3076) );
  BUFX2 U3489 ( .A(fifo[412]), .Y(n3077) );
  BUFX2 U3490 ( .A(fifo[411]), .Y(n3078) );
  BUFX2 U3491 ( .A(fifo[410]), .Y(n3079) );
  BUFX2 U3492 ( .A(fifo[409]), .Y(n3080) );
  BUFX2 U3493 ( .A(fifo[408]), .Y(n3081) );
  BUFX2 U3494 ( .A(fifo[407]), .Y(n3082) );
  BUFX2 U3495 ( .A(fifo[406]), .Y(n3083) );
  BUFX2 U3496 ( .A(fifo[405]), .Y(n3084) );
  BUFX2 U3497 ( .A(fifo[404]), .Y(n3085) );
  BUFX2 U3498 ( .A(fifo[403]), .Y(n3086) );
  BUFX2 U3499 ( .A(fifo[402]), .Y(n3087) );
  BUFX2 U3500 ( .A(fifo[401]), .Y(n3088) );
  BUFX2 U3501 ( .A(fifo[400]), .Y(n3089) );
  BUFX2 U3502 ( .A(fifo[399]), .Y(n3090) );
  BUFX2 U3503 ( .A(fifo[398]), .Y(n3091) );
  BUFX2 U3504 ( .A(fifo[397]), .Y(n3092) );
  BUFX2 U3505 ( .A(fifo[396]), .Y(n3093) );
  BUFX2 U3506 ( .A(fifo[395]), .Y(n3094) );
  BUFX2 U3507 ( .A(fifo[394]), .Y(n3095) );
  BUFX2 U3508 ( .A(fifo[393]), .Y(n3096) );
  BUFX2 U3509 ( .A(fifo[392]), .Y(n3097) );
  BUFX2 U3510 ( .A(fifo[391]), .Y(n3098) );
  BUFX2 U3511 ( .A(fifo[390]), .Y(n3099) );
  BUFX2 U3512 ( .A(fifo[389]), .Y(n3100) );
  BUFX2 U3513 ( .A(fifo[388]), .Y(n3101) );
  BUFX2 U3514 ( .A(fifo[387]), .Y(n3102) );
  BUFX2 U3515 ( .A(fifo[386]), .Y(n3103) );
  BUFX2 U3516 ( .A(fifo[385]), .Y(n3104) );
  BUFX2 U3517 ( .A(fifo[384]), .Y(n3105) );
  BUFX2 U3518 ( .A(fifo[159]), .Y(n3106) );
  BUFX2 U3519 ( .A(wr_ptr_gray_ss[0]), .Y(n3107) );
  BUFX2 U3520 ( .A(rd_ptr_gray_ss[2]), .Y(n3108) );
  BUFX2 U3521 ( .A(rd_ptr_bin_4_), .Y(n3109) );
  BUFX2 U3522 ( .A(wr_ptr_gray_ss[3]), .Y(n3110) );
  BUFX2 U3523 ( .A(wr_ptr_bin[0]), .Y(n3111) );
  BUFX2 U3524 ( .A(wr_ptr_bin[3]), .Y(n3112) );
  INVX1 U3525 ( .A(n3564), .Y(n3583) );
  INVX1 U3526 ( .A(n3564), .Y(n3582) );
  INVX1 U3527 ( .A(n3563), .Y(n3581) );
  INVX1 U3528 ( .A(n3563), .Y(n3580) );
  INVX1 U3529 ( .A(n3563), .Y(n3579) );
  INVX1 U3530 ( .A(n3563), .Y(n3578) );
  INVX1 U3531 ( .A(n3564), .Y(n3577) );
  INVX1 U3532 ( .A(n3564), .Y(n3576) );
  INVX1 U3533 ( .A(n3564), .Y(n3575) );
  INVX1 U3534 ( .A(n3563), .Y(n3574) );
  INVX1 U3535 ( .A(n3565), .Y(n3573) );
  INVX1 U3536 ( .A(n3565), .Y(n3572) );
  INVX1 U3537 ( .A(n3565), .Y(n3571) );
  INVX1 U3538 ( .A(n3565), .Y(n3570) );
  INVX1 U3539 ( .A(n3565), .Y(n3569) );
  INVX1 U3540 ( .A(n3564), .Y(n3568) );
  INVX1 U3541 ( .A(n3564), .Y(n3567) );
  INVX1 U3542 ( .A(n3675), .Y(n3593) );
  INVX1 U3543 ( .A(n3675), .Y(n3592) );
  INVX1 U3544 ( .A(n3675), .Y(n3591) );
  INVX1 U3545 ( .A(n3675), .Y(n3590) );
  INVX1 U3546 ( .A(n3675), .Y(n3589) );
  INVX1 U3547 ( .A(n3675), .Y(n3588) );
  INVX1 U3548 ( .A(n3675), .Y(n3587) );
  INVX1 U3549 ( .A(n3563), .Y(n3586) );
  INVX1 U3550 ( .A(n3564), .Y(n3585) );
  INVX1 U3551 ( .A(n3563), .Y(n3584) );
  INVX1 U3552 ( .A(n3565), .Y(n3566) );
  INVX1 U3553 ( .A(n3675), .Y(n3594) );
  INVX1 U3554 ( .A(n1929), .Y(n3563) );
  INVX1 U3555 ( .A(n1929), .Y(n3564) );
  INVX1 U3556 ( .A(n1929), .Y(n3565) );
  INVX1 U3557 ( .A(n1220), .Y(n3660) );
  INVX1 U3558 ( .A(n1016), .Y(n3666) );
  INVX1 U3559 ( .A(n950), .Y(n3668) );
  INVX1 U3560 ( .A(n884), .Y(n3670) );
  INVX1 U3561 ( .A(n1287), .Y(n3658) );
  INVX1 U3562 ( .A(n1153), .Y(n3662) );
  INVX1 U3563 ( .A(n3653), .Y(n3602) );
  INVX1 U3564 ( .A(n3653), .Y(n3603) );
  INVX1 U3565 ( .A(n3653), .Y(n3604) );
  INVX1 U3566 ( .A(n3652), .Y(n3605) );
  INVX1 U3567 ( .A(n3652), .Y(n3606) );
  INVX1 U3568 ( .A(n3652), .Y(n3607) );
  INVX1 U3569 ( .A(n3647), .Y(n3608) );
  INVX1 U3570 ( .A(n3651), .Y(n3609) );
  INVX1 U3571 ( .A(n3650), .Y(n3610) );
  INVX1 U3572 ( .A(n3651), .Y(n3611) );
  INVX1 U3573 ( .A(n3651), .Y(n3612) );
  INVX1 U3574 ( .A(n3651), .Y(n3613) );
  INVX1 U3575 ( .A(n3650), .Y(n3614) );
  INVX1 U3576 ( .A(n3650), .Y(n3615) );
  INVX1 U3577 ( .A(n3650), .Y(n3616) );
  INVX1 U3578 ( .A(n3649), .Y(n3617) );
  INVX1 U3579 ( .A(n3649), .Y(n3618) );
  INVX1 U3580 ( .A(n3649), .Y(n3619) );
  INVX1 U3581 ( .A(n3648), .Y(n3620) );
  INVX1 U3582 ( .A(n3648), .Y(n3621) );
  INVX1 U3583 ( .A(n3648), .Y(n3622) );
  INVX1 U3584 ( .A(n3647), .Y(n3623) );
  INVX1 U3585 ( .A(n3647), .Y(n3624) );
  INVX1 U3586 ( .A(n3647), .Y(n3625) );
  INVX1 U3587 ( .A(reset), .Y(n3626) );
  INVX1 U3588 ( .A(n3646), .Y(n3627) );
  INVX1 U3589 ( .A(n3647), .Y(n3628) );
  INVX1 U3590 ( .A(n3646), .Y(n3629) );
  INVX1 U3591 ( .A(n3646), .Y(n3630) );
  INVX1 U3592 ( .A(n3646), .Y(n3631) );
  INVX1 U3593 ( .A(n3652), .Y(n3632) );
  INVX1 U3594 ( .A(n3654), .Y(n3633) );
  INVX1 U3595 ( .A(n3646), .Y(n3634) );
  INVX1 U3596 ( .A(n3649), .Y(n3635) );
  INVX1 U3597 ( .A(n3645), .Y(n3636) );
  INVX1 U3598 ( .A(n3644), .Y(n3637) );
  INVX1 U3599 ( .A(n3645), .Y(n3638) );
  INVX1 U3600 ( .A(n3645), .Y(n3639) );
  INVX1 U3601 ( .A(n3645), .Y(n3640) );
  INVX1 U3602 ( .A(n3644), .Y(n3641) );
  INVX1 U3603 ( .A(n3644), .Y(n3642) );
  INVX1 U3604 ( .A(n3644), .Y(n3643) );
  INVX1 U3605 ( .A(n3654), .Y(n3599) );
  INVX1 U3606 ( .A(n3654), .Y(n3600) );
  INVX1 U3607 ( .A(n3654), .Y(n3601) );
  INVX1 U3608 ( .A(n3656), .Y(n3655) );
  INVX1 U3609 ( .A(n1253), .Y(n3659) );
  INVX1 U3610 ( .A(n1119), .Y(n3663) );
  INVX1 U3611 ( .A(n1085), .Y(n3664) );
  INVX1 U3612 ( .A(n1321), .Y(n3657) );
  INVX1 U3613 ( .A(n1186), .Y(n3661) );
  INVX1 U3614 ( .A(n850), .Y(n3671) );
  INVX1 U3615 ( .A(n1051), .Y(n3665) );
  INVX1 U3616 ( .A(n983), .Y(n3667) );
  INVX1 U3617 ( .A(n917), .Y(n3669) );
  INVX1 U3618 ( .A(n815), .Y(n3672) );
  INVX1 U3619 ( .A(n3648), .Y(n3598) );
  INVX1 U3620 ( .A(n3597), .Y(n3653) );
  INVX1 U3621 ( .A(n3597), .Y(n3652) );
  INVX1 U3622 ( .A(n3596), .Y(n3651) );
  INVX1 U3623 ( .A(n3596), .Y(n3650) );
  INVX1 U3624 ( .A(n3596), .Y(n3649) );
  INVX1 U3625 ( .A(n3597), .Y(n3648) );
  INVX1 U3626 ( .A(n3596), .Y(n3647) );
  INVX1 U3627 ( .A(n3596), .Y(n3646) );
  INVX1 U3628 ( .A(n3595), .Y(n3645) );
  INVX1 U3629 ( .A(n3595), .Y(n3644) );
  INVX1 U3630 ( .A(n3597), .Y(n3654) );
  INVX1 U3631 ( .A(n1364), .Y(n3656) );
  INVX1 U3632 ( .A(reset), .Y(n3597) );
  INVX1 U3633 ( .A(reset), .Y(n3596) );
  INVX1 U3634 ( .A(n3653), .Y(n3595) );
  INVX1 U3635 ( .A(n3565), .Y(n3676) );
  AND2X1 U3636 ( .A(n1320), .B(n3746), .Y(n1118) );
  AND2X1 U3637 ( .A(n1050), .B(n3746), .Y(n849) );
  AND2X1 U3638 ( .A(n1084), .B(n3749), .Y(n1050) );
  INVX1 U3639 ( .A(n3109), .Y(n3744) );
  INVX1 U3640 ( .A(n1930), .Y(n3675) );
  INVX1 U3641 ( .A(n1931), .Y(n3674) );
  INVX1 U3642 ( .A(n1932), .Y(n3673) );
  INVX1 U3643 ( .A(n1964), .Y(n3711) );
  INVX1 U3644 ( .A(n1963), .Y(n3710) );
  INVX1 U3645 ( .A(n1962), .Y(n3709) );
  INVX1 U3646 ( .A(n1961), .Y(n3708) );
  INVX1 U3647 ( .A(n1960), .Y(n3707) );
  INVX1 U3648 ( .A(n1959), .Y(n3706) );
  INVX1 U3649 ( .A(n1958), .Y(n3705) );
  INVX1 U3650 ( .A(n1957), .Y(n3704) );
  INVX1 U3651 ( .A(n1956), .Y(n3703) );
  INVX1 U3652 ( .A(n1955), .Y(n3702) );
  INVX1 U3653 ( .A(n1954), .Y(n3701) );
  INVX1 U3654 ( .A(n1953), .Y(n3700) );
  INVX1 U3655 ( .A(n1952), .Y(n3699) );
  INVX1 U3656 ( .A(n1951), .Y(n3698) );
  INVX1 U3657 ( .A(n1950), .Y(n3697) );
  INVX1 U3658 ( .A(n1949), .Y(n3696) );
  INVX1 U3659 ( .A(n1948), .Y(n3695) );
  INVX1 U3660 ( .A(n1947), .Y(n3694) );
  INVX1 U3661 ( .A(n1946), .Y(n3693) );
  INVX1 U3662 ( .A(n1945), .Y(n3692) );
  INVX1 U3663 ( .A(n1944), .Y(n3691) );
  INVX1 U3664 ( .A(n1943), .Y(n3690) );
  INVX1 U3665 ( .A(n1942), .Y(n3689) );
  INVX1 U3666 ( .A(n1941), .Y(n3688) );
  INVX1 U3667 ( .A(n1940), .Y(n3687) );
  INVX1 U3668 ( .A(n1939), .Y(n3686) );
  INVX1 U3669 ( .A(n1938), .Y(n3685) );
  INVX1 U3670 ( .A(n1937), .Y(n3684) );
  INVX1 U3671 ( .A(n1936), .Y(n3683) );
  INVX1 U3672 ( .A(n1935), .Y(n3682) );
  INVX1 U3673 ( .A(n1934), .Y(n3681) );
  INVX1 U3674 ( .A(n1933), .Y(n3680) );
  XNOR2X1 U3675 ( .A(n3108), .B(n2634), .Y(n3113) );
  INVX1 U3676 ( .A(rd_ptr_bin_ss_1_), .Y(n3678) );
  INVX1 U3677 ( .A(n2856), .Y(n3745) );
  INVX1 U3678 ( .A(n2634), .Y(n3677) );
  XNOR2X1 U3679 ( .A(n2880), .B(rd_ptr_bin_ss_1_), .Y(n3114) );
  INVX1 U3680 ( .A(data_in[0]), .Y(n3743) );
  INVX1 U3681 ( .A(data_in[1]), .Y(n3742) );
  INVX1 U3682 ( .A(data_in[2]), .Y(n3741) );
  INVX1 U3683 ( .A(data_in[3]), .Y(n3740) );
  INVX1 U3684 ( .A(data_in[4]), .Y(n3739) );
  INVX1 U3685 ( .A(data_in[5]), .Y(n3738) );
  INVX1 U3686 ( .A(data_in[6]), .Y(n3737) );
  INVX1 U3687 ( .A(data_in[7]), .Y(n3736) );
  INVX1 U3688 ( .A(data_in[8]), .Y(n3735) );
  INVX1 U3689 ( .A(data_in[9]), .Y(n3734) );
  INVX1 U3690 ( .A(data_in[10]), .Y(n3733) );
  INVX1 U3691 ( .A(data_in[11]), .Y(n3732) );
  INVX1 U3692 ( .A(data_in[12]), .Y(n3731) );
  INVX1 U3693 ( .A(data_in[13]), .Y(n3730) );
  INVX1 U3694 ( .A(data_in[14]), .Y(n3729) );
  INVX1 U3695 ( .A(data_in[15]), .Y(n3728) );
  INVX1 U3696 ( .A(data_in[16]), .Y(n3727) );
  INVX1 U3697 ( .A(data_in[17]), .Y(n3726) );
  INVX1 U3698 ( .A(data_in[18]), .Y(n3725) );
  INVX1 U3699 ( .A(data_in[19]), .Y(n3724) );
  INVX1 U3700 ( .A(data_in[20]), .Y(n3723) );
  INVX1 U3701 ( .A(data_in[21]), .Y(n3722) );
  INVX1 U3702 ( .A(data_in[22]), .Y(n3721) );
  INVX1 U3703 ( .A(data_in[23]), .Y(n3720) );
  INVX1 U3704 ( .A(data_in[24]), .Y(n3719) );
  INVX1 U3705 ( .A(data_in[25]), .Y(n3718) );
  INVX1 U3706 ( .A(data_in[26]), .Y(n3717) );
  INVX1 U3707 ( .A(data_in[27]), .Y(n3716) );
  INVX1 U3708 ( .A(data_in[28]), .Y(n3715) );
  INVX1 U3709 ( .A(data_in[29]), .Y(n3714) );
  INVX1 U3710 ( .A(data_in[30]), .Y(n3713) );
  INVX1 U3711 ( .A(data_in[31]), .Y(n3712) );
  INVX1 U3712 ( .A(n3112), .Y(n3749) );
  INVX1 U3713 ( .A(n2857), .Y(n3748) );
  INVX1 U3714 ( .A(n2635), .Y(n3747) );
  INVX1 U3715 ( .A(n3111), .Y(n3746) );
  INVX1 U3716 ( .A(reset), .Y(n3679) );
  MUX2X1 U3717 ( .B(n3116), .A(n3117), .S(n3587), .Y(n3115) );
  MUX2X1 U3718 ( .B(n3119), .A(n3120), .S(n3590), .Y(n3118) );
  MUX2X1 U3719 ( .B(n3122), .A(n3123), .S(n3593), .Y(n3121) );
  MUX2X1 U3720 ( .B(n3125), .A(n3126), .S(n3592), .Y(n3124) );
  MUX2X1 U3721 ( .B(n3127), .A(n3128), .S(n1932), .Y(n106) );
  MUX2X1 U3722 ( .B(n3130), .A(n3131), .S(n3588), .Y(n3129) );
  MUX2X1 U3723 ( .B(n3133), .A(n3134), .S(n3591), .Y(n3132) );
  MUX2X1 U3724 ( .B(n3136), .A(n3137), .S(n3594), .Y(n3135) );
  MUX2X1 U3725 ( .B(n3139), .A(n3140), .S(n3588), .Y(n3138) );
  MUX2X1 U3726 ( .B(n3141), .A(n3142), .S(n1932), .Y(n105) );
  MUX2X1 U3727 ( .B(n3144), .A(n3145), .S(n3587), .Y(n3143) );
  MUX2X1 U3728 ( .B(n3147), .A(n3148), .S(n3587), .Y(n3146) );
  MUX2X1 U3729 ( .B(n3150), .A(n3151), .S(n3587), .Y(n3149) );
  MUX2X1 U3730 ( .B(n3153), .A(n3154), .S(n3587), .Y(n3152) );
  MUX2X1 U3731 ( .B(n3155), .A(n3156), .S(n1932), .Y(n104) );
  MUX2X1 U3732 ( .B(n3158), .A(n3159), .S(n3587), .Y(n3157) );
  MUX2X1 U3733 ( .B(n3161), .A(n3162), .S(n3587), .Y(n3160) );
  MUX2X1 U3734 ( .B(n3164), .A(n3165), .S(n3587), .Y(n3163) );
  MUX2X1 U3735 ( .B(n3167), .A(n3168), .S(n3587), .Y(n3166) );
  MUX2X1 U3736 ( .B(n3169), .A(n3170), .S(n1932), .Y(n103) );
  MUX2X1 U3737 ( .B(n3172), .A(n3173), .S(n3587), .Y(n3171) );
  MUX2X1 U3738 ( .B(n3175), .A(n3176), .S(n3587), .Y(n3174) );
  MUX2X1 U3739 ( .B(n3178), .A(n3179), .S(n3587), .Y(n3177) );
  MUX2X1 U3740 ( .B(n3181), .A(n3182), .S(n3587), .Y(n3180) );
  MUX2X1 U3741 ( .B(n3183), .A(n3184), .S(n1932), .Y(n102) );
  MUX2X1 U3742 ( .B(n3186), .A(n3187), .S(n3588), .Y(n3185) );
  MUX2X1 U3743 ( .B(n3189), .A(n3190), .S(n3588), .Y(n3188) );
  MUX2X1 U3744 ( .B(n3192), .A(n3193), .S(n3588), .Y(n3191) );
  MUX2X1 U3745 ( .B(n3195), .A(n3196), .S(n3588), .Y(n3194) );
  MUX2X1 U3746 ( .B(n3197), .A(n3198), .S(n1932), .Y(n101) );
  MUX2X1 U3747 ( .B(n3200), .A(n3201), .S(n3588), .Y(n3199) );
  MUX2X1 U3748 ( .B(n3203), .A(n3204), .S(n3588), .Y(n3202) );
  MUX2X1 U3749 ( .B(n3206), .A(n3207), .S(n3588), .Y(n3205) );
  MUX2X1 U3750 ( .B(n3209), .A(n3210), .S(n3588), .Y(n3208) );
  MUX2X1 U3751 ( .B(n3211), .A(n3212), .S(n1932), .Y(n100) );
  MUX2X1 U3752 ( .B(n3214), .A(n3215), .S(n3588), .Y(n3213) );
  MUX2X1 U3753 ( .B(n3217), .A(n3218), .S(n3588), .Y(n3216) );
  MUX2X1 U3754 ( .B(n3220), .A(n3221), .S(n3588), .Y(n3219) );
  MUX2X1 U3755 ( .B(n3223), .A(n3224), .S(n3588), .Y(n3222) );
  MUX2X1 U3756 ( .B(n3225), .A(n3226), .S(n1932), .Y(n99) );
  MUX2X1 U3757 ( .B(n3228), .A(n3229), .S(n3589), .Y(n3227) );
  MUX2X1 U3758 ( .B(n3231), .A(n3232), .S(n3589), .Y(n3230) );
  MUX2X1 U3759 ( .B(n3234), .A(n3235), .S(n3589), .Y(n3233) );
  MUX2X1 U3760 ( .B(n3237), .A(n3238), .S(n3589), .Y(n3236) );
  MUX2X1 U3761 ( .B(n3239), .A(n3240), .S(n1932), .Y(n98) );
  MUX2X1 U3762 ( .B(n3242), .A(n3243), .S(n3589), .Y(n3241) );
  MUX2X1 U3763 ( .B(n3245), .A(n3246), .S(n3589), .Y(n3244) );
  MUX2X1 U3764 ( .B(n3248), .A(n3249), .S(n3589), .Y(n3247) );
  MUX2X1 U3765 ( .B(n3251), .A(n3252), .S(n3589), .Y(n3250) );
  MUX2X1 U3766 ( .B(n3253), .A(n3254), .S(n1932), .Y(n97) );
  MUX2X1 U3767 ( .B(n3256), .A(n3257), .S(n3589), .Y(n3255) );
  MUX2X1 U3768 ( .B(n3259), .A(n3260), .S(n3589), .Y(n3258) );
  MUX2X1 U3769 ( .B(n3262), .A(n3263), .S(n3589), .Y(n3261) );
  MUX2X1 U3770 ( .B(n3265), .A(n3266), .S(n3589), .Y(n3264) );
  MUX2X1 U3771 ( .B(n3267), .A(n3268), .S(n1932), .Y(n96) );
  MUX2X1 U3772 ( .B(n3270), .A(n3271), .S(n3590), .Y(n3269) );
  MUX2X1 U3773 ( .B(n3273), .A(n3274), .S(n3590), .Y(n3272) );
  MUX2X1 U3774 ( .B(n3276), .A(n3277), .S(n3590), .Y(n3275) );
  MUX2X1 U3775 ( .B(n3279), .A(n3280), .S(n3590), .Y(n3278) );
  MUX2X1 U3776 ( .B(n3281), .A(n3282), .S(n1932), .Y(n95) );
  MUX2X1 U3777 ( .B(n3284), .A(n3285), .S(n3590), .Y(n3283) );
  MUX2X1 U3778 ( .B(n3287), .A(n3288), .S(n3590), .Y(n3286) );
  MUX2X1 U3779 ( .B(n3290), .A(n3291), .S(n3590), .Y(n3289) );
  MUX2X1 U3780 ( .B(n3293), .A(n3294), .S(n3590), .Y(n3292) );
  MUX2X1 U3781 ( .B(n3295), .A(n3296), .S(n1932), .Y(n94) );
  MUX2X1 U3782 ( .B(n3298), .A(n3299), .S(n3590), .Y(n3297) );
  MUX2X1 U3783 ( .B(n3301), .A(n3302), .S(n3590), .Y(n3300) );
  MUX2X1 U3784 ( .B(n3304), .A(n3305), .S(n3590), .Y(n3303) );
  MUX2X1 U3785 ( .B(n3307), .A(n3308), .S(n3590), .Y(n3306) );
  MUX2X1 U3786 ( .B(n3309), .A(n3310), .S(n1932), .Y(n93) );
  MUX2X1 U3787 ( .B(n3312), .A(n3313), .S(n3591), .Y(n3311) );
  MUX2X1 U3788 ( .B(n3315), .A(n3316), .S(n3591), .Y(n3314) );
  MUX2X1 U3789 ( .B(n3318), .A(n3319), .S(n3591), .Y(n3317) );
  MUX2X1 U3790 ( .B(n3321), .A(n3322), .S(n3591), .Y(n3320) );
  MUX2X1 U3791 ( .B(n3323), .A(n3324), .S(n1932), .Y(n92) );
  MUX2X1 U3792 ( .B(n3326), .A(n3327), .S(n3591), .Y(n3325) );
  MUX2X1 U3793 ( .B(n3329), .A(n3330), .S(n3591), .Y(n3328) );
  MUX2X1 U3794 ( .B(n3332), .A(n3333), .S(n3591), .Y(n3331) );
  MUX2X1 U3795 ( .B(n3335), .A(n3336), .S(n3591), .Y(n3334) );
  MUX2X1 U3796 ( .B(n3337), .A(n3338), .S(n1932), .Y(n91) );
  MUX2X1 U3797 ( .B(n3340), .A(n3341), .S(n3591), .Y(n3339) );
  MUX2X1 U3798 ( .B(n3343), .A(n3344), .S(n3591), .Y(n3342) );
  MUX2X1 U3799 ( .B(n3346), .A(n3347), .S(n3591), .Y(n3345) );
  MUX2X1 U3800 ( .B(n3349), .A(n3350), .S(n3591), .Y(n3348) );
  MUX2X1 U3801 ( .B(n3351), .A(n3352), .S(n1932), .Y(n90) );
  MUX2X1 U3802 ( .B(n3354), .A(n3355), .S(n3591), .Y(n3353) );
  MUX2X1 U3803 ( .B(n3357), .A(n3358), .S(n3589), .Y(n3356) );
  MUX2X1 U3804 ( .B(n3360), .A(n3361), .S(n3589), .Y(n3359) );
  MUX2X1 U3805 ( .B(n3363), .A(n3364), .S(n3587), .Y(n3362) );
  MUX2X1 U3806 ( .B(n3365), .A(n3366), .S(n1932), .Y(n89) );
  MUX2X1 U3807 ( .B(n3368), .A(n3369), .S(n3593), .Y(n3367) );
  MUX2X1 U3808 ( .B(n3371), .A(n3372), .S(n3592), .Y(n3370) );
  MUX2X1 U3809 ( .B(n3374), .A(n3375), .S(n3589), .Y(n3373) );
  MUX2X1 U3810 ( .B(n3377), .A(n3378), .S(n3588), .Y(n3376) );
  MUX2X1 U3811 ( .B(n3379), .A(n3380), .S(n1932), .Y(n88) );
  MUX2X1 U3812 ( .B(n3382), .A(n3383), .S(n3590), .Y(n3381) );
  MUX2X1 U3813 ( .B(n3385), .A(n3386), .S(n3594), .Y(n3384) );
  MUX2X1 U3814 ( .B(n3388), .A(n3389), .S(n3594), .Y(n3387) );
  MUX2X1 U3815 ( .B(n3391), .A(n3392), .S(n3591), .Y(n3390) );
  MUX2X1 U3816 ( .B(n3393), .A(n3394), .S(n1932), .Y(n87) );
  MUX2X1 U3817 ( .B(n3396), .A(n3397), .S(n3592), .Y(n3395) );
  MUX2X1 U3818 ( .B(n3399), .A(n3400), .S(n3592), .Y(n3398) );
  MUX2X1 U3819 ( .B(n3402), .A(n3403), .S(n3592), .Y(n3401) );
  MUX2X1 U3820 ( .B(n3405), .A(n3406), .S(n3592), .Y(n3404) );
  MUX2X1 U3821 ( .B(n3407), .A(n3408), .S(n1932), .Y(n86) );
  MUX2X1 U3822 ( .B(n3410), .A(n3411), .S(n3592), .Y(n3409) );
  MUX2X1 U3823 ( .B(n3413), .A(n3414), .S(n3592), .Y(n3412) );
  MUX2X1 U3824 ( .B(n3416), .A(n3417), .S(n3592), .Y(n3415) );
  MUX2X1 U3825 ( .B(n3419), .A(n3420), .S(n3592), .Y(n3418) );
  MUX2X1 U3826 ( .B(n3421), .A(n3422), .S(n1932), .Y(n85) );
  MUX2X1 U3827 ( .B(n3424), .A(n3425), .S(n3592), .Y(n3423) );
  MUX2X1 U3828 ( .B(n3427), .A(n3428), .S(n3592), .Y(n3426) );
  MUX2X1 U3829 ( .B(n3430), .A(n3431), .S(n3592), .Y(n3429) );
  MUX2X1 U3830 ( .B(n3433), .A(n3434), .S(n3592), .Y(n3432) );
  MUX2X1 U3831 ( .B(n3435), .A(n3436), .S(n1932), .Y(n84) );
  MUX2X1 U3832 ( .B(n3438), .A(n3439), .S(n3593), .Y(n3437) );
  MUX2X1 U3833 ( .B(n3441), .A(n3442), .S(n3593), .Y(n3440) );
  MUX2X1 U3834 ( .B(n3444), .A(n3445), .S(n3593), .Y(n3443) );
  MUX2X1 U3835 ( .B(n3447), .A(n3448), .S(n3593), .Y(n3446) );
  MUX2X1 U3836 ( .B(n3449), .A(n3450), .S(n1932), .Y(n83) );
  MUX2X1 U3837 ( .B(n3452), .A(n3453), .S(n3593), .Y(n3451) );
  MUX2X1 U3838 ( .B(n3455), .A(n3456), .S(n3593), .Y(n3454) );
  MUX2X1 U3839 ( .B(n3458), .A(n3459), .S(n3593), .Y(n3457) );
  MUX2X1 U3840 ( .B(n3461), .A(n3462), .S(n3593), .Y(n3460) );
  MUX2X1 U3841 ( .B(n3463), .A(n3464), .S(n1932), .Y(n82) );
  MUX2X1 U3842 ( .B(n3466), .A(n3467), .S(n3593), .Y(n3465) );
  MUX2X1 U3843 ( .B(n3469), .A(n3470), .S(n3593), .Y(n3468) );
  MUX2X1 U3844 ( .B(n3472), .A(n3473), .S(n3593), .Y(n3471) );
  MUX2X1 U3845 ( .B(n3475), .A(n3476), .S(n3593), .Y(n3474) );
  MUX2X1 U3846 ( .B(n3477), .A(n3478), .S(n1932), .Y(n81) );
  MUX2X1 U3847 ( .B(n3480), .A(n3481), .S(n3594), .Y(n3479) );
  MUX2X1 U3848 ( .B(n3483), .A(n3484), .S(n3594), .Y(n3482) );
  MUX2X1 U3849 ( .B(n3486), .A(n3487), .S(n3594), .Y(n3485) );
  MUX2X1 U3850 ( .B(n3489), .A(n3490), .S(n3594), .Y(n3488) );
  MUX2X1 U3851 ( .B(n3491), .A(n3492), .S(n1932), .Y(n80) );
  MUX2X1 U3852 ( .B(n3494), .A(n3495), .S(n3594), .Y(n3493) );
  MUX2X1 U3853 ( .B(n3497), .A(n3498), .S(n3594), .Y(n3496) );
  MUX2X1 U3854 ( .B(n3500), .A(n3501), .S(n3594), .Y(n3499) );
  MUX2X1 U3855 ( .B(n3503), .A(n3504), .S(n3594), .Y(n3502) );
  MUX2X1 U3856 ( .B(n3505), .A(n3506), .S(n1932), .Y(n79) );
  MUX2X1 U3857 ( .B(n3508), .A(n3509), .S(n3594), .Y(n3507) );
  MUX2X1 U3858 ( .B(n3511), .A(n3512), .S(n3594), .Y(n3510) );
  MUX2X1 U3859 ( .B(n3514), .A(n3515), .S(n3594), .Y(n3513) );
  MUX2X1 U3860 ( .B(n3517), .A(n3518), .S(n3594), .Y(n3516) );
  MUX2X1 U3861 ( .B(n3519), .A(n3520), .S(n1932), .Y(n78) );
  MUX2X1 U3862 ( .B(n3522), .A(n3523), .S(n3592), .Y(n3521) );
  MUX2X1 U3863 ( .B(n3525), .A(n3526), .S(n3593), .Y(n3524) );
  MUX2X1 U3864 ( .B(n3528), .A(n3529), .S(n3587), .Y(n3527) );
  MUX2X1 U3865 ( .B(n3531), .A(n3532), .S(n3590), .Y(n3530) );
  MUX2X1 U3866 ( .B(n3533), .A(n3534), .S(n1932), .Y(n77) );
  MUX2X1 U3867 ( .B(n3536), .A(n3537), .S(n3591), .Y(n3535) );
  MUX2X1 U3868 ( .B(n3539), .A(n3540), .S(n3594), .Y(n3538) );
  MUX2X1 U3869 ( .B(n3542), .A(n3543), .S(n3588), .Y(n3541) );
  MUX2X1 U3870 ( .B(n3545), .A(n3546), .S(n3593), .Y(n3544) );
  MUX2X1 U3871 ( .B(n3547), .A(n3548), .S(n1932), .Y(n76) );
  MUX2X1 U3872 ( .B(n3550), .A(n3551), .S(n3590), .Y(n3549) );
  MUX2X1 U3873 ( .B(n3553), .A(n3554), .S(n3589), .Y(n3552) );
  MUX2X1 U3874 ( .B(n3556), .A(n3557), .S(n3592), .Y(n3555) );
  MUX2X1 U3875 ( .B(n3559), .A(n3560), .S(n3587), .Y(n3558) );
  MUX2X1 U3876 ( .B(n3561), .A(n3562), .S(n1932), .Y(n75) );
  MUX2X1 U3877 ( .B(n2764), .A(n3073), .S(n3566), .Y(n3117) );
  MUX2X1 U3878 ( .B(n2607), .A(n2491), .S(n3566), .Y(n3116) );
  MUX2X1 U3879 ( .B(n2605), .A(n3042), .S(n3566), .Y(n3120) );
  MUX2X1 U3880 ( .B(n2514), .A(n2824), .S(n3566), .Y(n3119) );
  MUX2X1 U3881 ( .B(n3118), .A(n3115), .S(n1931), .Y(n3128) );
  MUX2X1 U3882 ( .B(n2757), .A(n3008), .S(n3567), .Y(n3123) );
  MUX2X1 U3883 ( .B(n2727), .A(n2976), .S(n3567), .Y(n3122) );
  MUX2X1 U3884 ( .B(n2794), .A(n3105), .S(n3567), .Y(n3126) );
  MUX2X1 U3885 ( .B(n2698), .A(n2944), .S(n3567), .Y(n3125) );
  MUX2X1 U3886 ( .B(n3124), .A(n3121), .S(n1931), .Y(n3127) );
  MUX2X1 U3887 ( .B(n2632), .A(n3072), .S(n3567), .Y(n3131) );
  MUX2X1 U3888 ( .B(n2537), .A(n2853), .S(n3567), .Y(n3130) );
  MUX2X1 U3889 ( .B(n2762), .A(n3041), .S(n3567), .Y(n3134) );
  MUX2X1 U3890 ( .B(n2580), .A(n2489), .S(n3567), .Y(n3133) );
  MUX2X1 U3891 ( .B(n3132), .A(n3129), .S(n1931), .Y(n3142) );
  MUX2X1 U3892 ( .B(n2756), .A(n3007), .S(n3567), .Y(n3137) );
  MUX2X1 U3893 ( .B(n2726), .A(n2975), .S(n3567), .Y(n3136) );
  MUX2X1 U3894 ( .B(n2793), .A(n3104), .S(n3567), .Y(n3140) );
  MUX2X1 U3895 ( .B(n2697), .A(n2943), .S(n3567), .Y(n3139) );
  MUX2X1 U3896 ( .B(n3138), .A(n3135), .S(n1931), .Y(n3141) );
  MUX2X1 U3897 ( .B(n2578), .A(n3071), .S(n3568), .Y(n3145) );
  MUX2X1 U3898 ( .B(n2487), .A(n2852), .S(n3568), .Y(n3144) );
  MUX2X1 U3899 ( .B(n2604), .A(n3040), .S(n3568), .Y(n3148) );
  MUX2X1 U3900 ( .B(n2513), .A(n2823), .S(n3568), .Y(n3147) );
  MUX2X1 U3901 ( .B(n3146), .A(n3143), .S(n1931), .Y(n3156) );
  MUX2X1 U3902 ( .B(n2755), .A(n3006), .S(n3568), .Y(n3151) );
  MUX2X1 U3903 ( .B(n2725), .A(n2974), .S(n3568), .Y(n3150) );
  MUX2X1 U3904 ( .B(n2792), .A(n3103), .S(n3568), .Y(n3154) );
  MUX2X1 U3905 ( .B(n2696), .A(n2942), .S(n3568), .Y(n3153) );
  MUX2X1 U3906 ( .B(n3152), .A(n3149), .S(n1931), .Y(n3155) );
  MUX2X1 U3907 ( .B(n2577), .A(n3070), .S(n3568), .Y(n3159) );
  MUX2X1 U3908 ( .B(n2486), .A(n2851), .S(n3568), .Y(n3158) );
  MUX2X1 U3909 ( .B(n2603), .A(n3039), .S(n3568), .Y(n3162) );
  MUX2X1 U3910 ( .B(n2512), .A(n2822), .S(n3568), .Y(n3161) );
  MUX2X1 U3911 ( .B(n3160), .A(n3157), .S(n1931), .Y(n3170) );
  MUX2X1 U3912 ( .B(n2754), .A(n3005), .S(n3569), .Y(n3165) );
  MUX2X1 U3913 ( .B(n2724), .A(n2973), .S(n3569), .Y(n3164) );
  MUX2X1 U3914 ( .B(n2791), .A(n3102), .S(n3569), .Y(n3168) );
  MUX2X1 U3915 ( .B(n2695), .A(n2941), .S(n3569), .Y(n3167) );
  MUX2X1 U3916 ( .B(n3166), .A(n3163), .S(n1931), .Y(n3169) );
  MUX2X1 U3917 ( .B(n2631), .A(n3069), .S(n3569), .Y(n3173) );
  MUX2X1 U3918 ( .B(n2485), .A(n2850), .S(n3569), .Y(n3172) );
  MUX2X1 U3919 ( .B(n2574), .A(n3038), .S(n3569), .Y(n3176) );
  MUX2X1 U3920 ( .B(n2481), .A(n2821), .S(n3569), .Y(n3175) );
  MUX2X1 U3921 ( .B(n3174), .A(n3171), .S(n1931), .Y(n3184) );
  MUX2X1 U3922 ( .B(n2753), .A(n3004), .S(n3569), .Y(n3179) );
  MUX2X1 U3923 ( .B(n2723), .A(n2972), .S(n3569), .Y(n3178) );
  MUX2X1 U3924 ( .B(n2790), .A(n3101), .S(n3569), .Y(n3182) );
  MUX2X1 U3925 ( .B(n2694), .A(n2940), .S(n3569), .Y(n3181) );
  MUX2X1 U3926 ( .B(n3180), .A(n3177), .S(n1931), .Y(n3183) );
  MUX2X1 U3927 ( .B(n2630), .A(n3068), .S(n3570), .Y(n3187) );
  MUX2X1 U3928 ( .B(n2536), .A(n2849), .S(n3570), .Y(n3186) );
  MUX2X1 U3929 ( .B(n2573), .A(n3037), .S(n3570), .Y(n3190) );
  MUX2X1 U3930 ( .B(n2480), .A(n2820), .S(n3570), .Y(n3189) );
  MUX2X1 U3931 ( .B(n3188), .A(n3185), .S(n1931), .Y(n3198) );
  MUX2X1 U3932 ( .B(n2752), .A(n3003), .S(n3570), .Y(n3193) );
  MUX2X1 U3933 ( .B(n2722), .A(n2971), .S(n3570), .Y(n3192) );
  MUX2X1 U3934 ( .B(n2789), .A(n3100), .S(n3570), .Y(n3196) );
  MUX2X1 U3935 ( .B(n2693), .A(n2939), .S(n3570), .Y(n3195) );
  MUX2X1 U3936 ( .B(n3194), .A(n3191), .S(n1931), .Y(n3197) );
  MUX2X1 U3937 ( .B(n2629), .A(n3067), .S(n3570), .Y(n3201) );
  MUX2X1 U3938 ( .B(n2535), .A(n2848), .S(n3570), .Y(n3200) );
  MUX2X1 U3939 ( .B(n2602), .A(n3036), .S(n3570), .Y(n3204) );
  MUX2X1 U3940 ( .B(n2479), .A(n2819), .S(n3570), .Y(n3203) );
  MUX2X1 U3941 ( .B(n3202), .A(n3199), .S(n1931), .Y(n3212) );
  MUX2X1 U3942 ( .B(n2666), .A(n3002), .S(n3571), .Y(n3207) );
  MUX2X1 U3943 ( .B(n2721), .A(n2970), .S(n3571), .Y(n3206) );
  MUX2X1 U3944 ( .B(n2788), .A(n3099), .S(n3571), .Y(n3210) );
  MUX2X1 U3945 ( .B(n2692), .A(n2938), .S(n3571), .Y(n3209) );
  MUX2X1 U3946 ( .B(n3208), .A(n3205), .S(n1931), .Y(n3211) );
  MUX2X1 U3947 ( .B(n2763), .A(n3066), .S(n3571), .Y(n3215) );
  MUX2X1 U3948 ( .B(n2606), .A(n2490), .S(n3571), .Y(n3214) );
  MUX2X1 U3949 ( .B(n2601), .A(n3035), .S(n3571), .Y(n3218) );
  MUX2X1 U3950 ( .B(n2511), .A(n2818), .S(n3571), .Y(n3217) );
  MUX2X1 U3951 ( .B(n3216), .A(n3213), .S(n1931), .Y(n3226) );
  MUX2X1 U3952 ( .B(n2751), .A(n3001), .S(n3571), .Y(n3221) );
  MUX2X1 U3953 ( .B(n2720), .A(n2969), .S(n3571), .Y(n3220) );
  MUX2X1 U3954 ( .B(n2787), .A(n3098), .S(n3571), .Y(n3224) );
  MUX2X1 U3955 ( .B(n2691), .A(n2937), .S(n3571), .Y(n3223) );
  MUX2X1 U3956 ( .B(n3222), .A(n3219), .S(n1931), .Y(n3225) );
  MUX2X1 U3957 ( .B(n2628), .A(n3065), .S(n3572), .Y(n3229) );
  MUX2X1 U3958 ( .B(n2534), .A(n2847), .S(n3572), .Y(n3228) );
  MUX2X1 U3959 ( .B(n2600), .A(n3034), .S(n3572), .Y(n3232) );
  MUX2X1 U3960 ( .B(n2510), .A(n2817), .S(n3572), .Y(n3231) );
  MUX2X1 U3961 ( .B(n3230), .A(n3227), .S(n1931), .Y(n3240) );
  MUX2X1 U3962 ( .B(n2750), .A(n3000), .S(n3572), .Y(n3235) );
  MUX2X1 U3963 ( .B(n2664), .A(n2968), .S(n3572), .Y(n3234) );
  MUX2X1 U3964 ( .B(n2786), .A(n3097), .S(n3572), .Y(n3238) );
  MUX2X1 U3965 ( .B(n2690), .A(n2936), .S(n3572), .Y(n3237) );
  MUX2X1 U3966 ( .B(n3236), .A(n3233), .S(n1931), .Y(n3239) );
  MUX2X1 U3967 ( .B(n2627), .A(n3064), .S(n3572), .Y(n3243) );
  MUX2X1 U3968 ( .B(n2533), .A(n2846), .S(n3572), .Y(n3242) );
  MUX2X1 U3969 ( .B(n2761), .A(n3033), .S(n3572), .Y(n3246) );
  MUX2X1 U3970 ( .B(n2579), .A(n2488), .S(n3572), .Y(n3245) );
  MUX2X1 U3971 ( .B(n3244), .A(n3241), .S(n1931), .Y(n3254) );
  MUX2X1 U3972 ( .B(n2749), .A(n2999), .S(n3573), .Y(n3249) );
  MUX2X1 U3973 ( .B(n2719), .A(n2967), .S(n3573), .Y(n3248) );
  MUX2X1 U3974 ( .B(n2785), .A(n3096), .S(n3573), .Y(n3252) );
  MUX2X1 U3975 ( .B(n2689), .A(n2935), .S(n3573), .Y(n3251) );
  MUX2X1 U3976 ( .B(n3250), .A(n3247), .S(n1931), .Y(n3253) );
  MUX2X1 U3977 ( .B(n2626), .A(n3063), .S(n3573), .Y(n3257) );
  MUX2X1 U3978 ( .B(n2532), .A(n2845), .S(n3573), .Y(n3256) );
  MUX2X1 U3979 ( .B(n2599), .A(n3032), .S(n3573), .Y(n3260) );
  MUX2X1 U3980 ( .B(n2509), .A(n2816), .S(n3573), .Y(n3259) );
  MUX2X1 U3981 ( .B(n3258), .A(n3255), .S(n1931), .Y(n3268) );
  MUX2X1 U3982 ( .B(n2748), .A(n2998), .S(n3573), .Y(n3263) );
  MUX2X1 U3983 ( .B(n2718), .A(n2966), .S(n3573), .Y(n3262) );
  MUX2X1 U3984 ( .B(n2668), .A(n3095), .S(n3573), .Y(n3266) );
  MUX2X1 U3985 ( .B(n2688), .A(n2934), .S(n3573), .Y(n3265) );
  MUX2X1 U3986 ( .B(n3264), .A(n3261), .S(n1931), .Y(n3267) );
  MUX2X1 U3987 ( .B(n2625), .A(n3062), .S(n3574), .Y(n3271) );
  MUX2X1 U3988 ( .B(n2531), .A(n2844), .S(n3574), .Y(n3270) );
  MUX2X1 U3989 ( .B(n2598), .A(n3031), .S(n3574), .Y(n3274) );
  MUX2X1 U3990 ( .B(n2508), .A(n2815), .S(n3574), .Y(n3273) );
  MUX2X1 U3991 ( .B(n3272), .A(n3269), .S(n1931), .Y(n3282) );
  MUX2X1 U3992 ( .B(n2747), .A(n2997), .S(n3574), .Y(n3277) );
  MUX2X1 U3993 ( .B(n2717), .A(n2965), .S(n3574), .Y(n3276) );
  MUX2X1 U3994 ( .B(n2784), .A(n3094), .S(n3574), .Y(n3280) );
  MUX2X1 U3995 ( .B(n2661), .A(n2933), .S(n3574), .Y(n3279) );
  MUX2X1 U3996 ( .B(n3278), .A(n3275), .S(n1931), .Y(n3281) );
  MUX2X1 U3997 ( .B(n2576), .A(n3061), .S(n3574), .Y(n3285) );
  MUX2X1 U3998 ( .B(n2484), .A(n2843), .S(n3574), .Y(n3284) );
  MUX2X1 U3999 ( .B(n2597), .A(n3030), .S(n3574), .Y(n3288) );
  MUX2X1 U4000 ( .B(n2507), .A(n2814), .S(n3574), .Y(n3287) );
  MUX2X1 U4001 ( .B(n3286), .A(n3283), .S(n1931), .Y(n3296) );
  MUX2X1 U4002 ( .B(n2746), .A(n2996), .S(n3575), .Y(n3291) );
  MUX2X1 U4003 ( .B(n2716), .A(n2964), .S(n3575), .Y(n3290) );
  MUX2X1 U4004 ( .B(n2783), .A(n3093), .S(n3575), .Y(n3294) );
  MUX2X1 U4005 ( .B(n2687), .A(n2932), .S(n3575), .Y(n3293) );
  MUX2X1 U4006 ( .B(n3292), .A(n3289), .S(n1931), .Y(n3295) );
  MUX2X1 U4007 ( .B(n2624), .A(n3060), .S(n3575), .Y(n3299) );
  MUX2X1 U4008 ( .B(n2530), .A(n2842), .S(n3575), .Y(n3298) );
  MUX2X1 U4009 ( .B(n2596), .A(n3029), .S(n3575), .Y(n3302) );
  MUX2X1 U4010 ( .B(n2506), .A(n2813), .S(n3575), .Y(n3301) );
  MUX2X1 U4011 ( .B(n3300), .A(n3297), .S(n1931), .Y(n3310) );
  MUX2X1 U4012 ( .B(n2745), .A(n2995), .S(n3575), .Y(n3305) );
  MUX2X1 U4013 ( .B(n2715), .A(n2963), .S(n3575), .Y(n3304) );
  MUX2X1 U4014 ( .B(n2782), .A(n3092), .S(n3575), .Y(n3308) );
  MUX2X1 U4015 ( .B(n2686), .A(n2931), .S(n3575), .Y(n3307) );
  MUX2X1 U4016 ( .B(n3306), .A(n3303), .S(n1931), .Y(n3309) );
  MUX2X1 U4017 ( .B(n2623), .A(n3059), .S(n3576), .Y(n3313) );
  MUX2X1 U4018 ( .B(n2529), .A(n2841), .S(n3576), .Y(n3312) );
  MUX2X1 U4019 ( .B(n2595), .A(n3028), .S(n3576), .Y(n3316) );
  MUX2X1 U4020 ( .B(n2505), .A(n2812), .S(n3576), .Y(n3315) );
  MUX2X1 U4021 ( .B(n3314), .A(n3311), .S(n1931), .Y(n3324) );
  MUX2X1 U4022 ( .B(n2744), .A(n2994), .S(n3576), .Y(n3319) );
  MUX2X1 U4023 ( .B(n2714), .A(n2962), .S(n3576), .Y(n3318) );
  MUX2X1 U4024 ( .B(n2781), .A(n3091), .S(n3576), .Y(n3322) );
  MUX2X1 U4025 ( .B(n2685), .A(n2930), .S(n3576), .Y(n3321) );
  MUX2X1 U4026 ( .B(n3320), .A(n3317), .S(n1931), .Y(n3323) );
  MUX2X1 U4027 ( .B(n2575), .A(n3058), .S(n3576), .Y(n3327) );
  MUX2X1 U4028 ( .B(n2483), .A(n2840), .S(n3576), .Y(n3326) );
  MUX2X1 U4029 ( .B(n2594), .A(n3027), .S(n3576), .Y(n3330) );
  MUX2X1 U4030 ( .B(n2504), .A(n2811), .S(n3576), .Y(n3329) );
  MUX2X1 U4031 ( .B(n3328), .A(n3325), .S(n1931), .Y(n3338) );
  MUX2X1 U4032 ( .B(n2743), .A(n2993), .S(n3577), .Y(n3333) );
  MUX2X1 U4033 ( .B(n2713), .A(n2961), .S(n3577), .Y(n3332) );
  MUX2X1 U4034 ( .B(n2780), .A(n3090), .S(n3577), .Y(n3336) );
  MUX2X1 U4035 ( .B(n2684), .A(n2929), .S(n3577), .Y(n3335) );
  MUX2X1 U4036 ( .B(n3334), .A(n3331), .S(n1931), .Y(n3337) );
  MUX2X1 U4037 ( .B(n2622), .A(n3057), .S(n3577), .Y(n3341) );
  MUX2X1 U4038 ( .B(n2528), .A(n2839), .S(n3577), .Y(n3340) );
  MUX2X1 U4039 ( .B(n2593), .A(n3026), .S(n3577), .Y(n3344) );
  MUX2X1 U4040 ( .B(n2503), .A(n2810), .S(n3577), .Y(n3343) );
  MUX2X1 U4041 ( .B(n3342), .A(n3339), .S(n1931), .Y(n3352) );
  MUX2X1 U4042 ( .B(n2742), .A(n2992), .S(n3577), .Y(n3347) );
  MUX2X1 U4043 ( .B(n2712), .A(n2960), .S(n3577), .Y(n3346) );
  MUX2X1 U4044 ( .B(n2779), .A(n3089), .S(n3577), .Y(n3350) );
  MUX2X1 U4045 ( .B(n2683), .A(n2928), .S(n3577), .Y(n3349) );
  MUX2X1 U4046 ( .B(n3348), .A(n3345), .S(n1931), .Y(n3351) );
  MUX2X1 U4047 ( .B(n2621), .A(n3056), .S(n3578), .Y(n3355) );
  MUX2X1 U4048 ( .B(n2527), .A(n2838), .S(n3578), .Y(n3354) );
  MUX2X1 U4049 ( .B(n2592), .A(n3025), .S(n3578), .Y(n3358) );
  MUX2X1 U4050 ( .B(n2502), .A(n2809), .S(n3578), .Y(n3357) );
  MUX2X1 U4051 ( .B(n3356), .A(n3353), .S(n1931), .Y(n3366) );
  MUX2X1 U4052 ( .B(n2741), .A(n2991), .S(n3578), .Y(n3361) );
  MUX2X1 U4053 ( .B(n2663), .A(n2959), .S(n3578), .Y(n3360) );
  MUX2X1 U4054 ( .B(n2778), .A(n3088), .S(n3578), .Y(n3364) );
  MUX2X1 U4055 ( .B(n2682), .A(n2927), .S(n3578), .Y(n3363) );
  MUX2X1 U4056 ( .B(n3362), .A(n3359), .S(n1931), .Y(n3365) );
  MUX2X1 U4057 ( .B(n2620), .A(n3055), .S(n3578), .Y(n3369) );
  MUX2X1 U4058 ( .B(n2526), .A(n2837), .S(n3578), .Y(n3368) );
  MUX2X1 U4059 ( .B(n2591), .A(n3024), .S(n3578), .Y(n3372) );
  MUX2X1 U4060 ( .B(n2501), .A(n2808), .S(n3578), .Y(n3371) );
  MUX2X1 U4061 ( .B(n3370), .A(n3367), .S(n1931), .Y(n3380) );
  MUX2X1 U4062 ( .B(n2740), .A(n2990), .S(n3579), .Y(n3375) );
  MUX2X1 U4063 ( .B(n2711), .A(n2958), .S(n3579), .Y(n3374) );
  MUX2X1 U4064 ( .B(n2777), .A(n3087), .S(n3579), .Y(n3378) );
  MUX2X1 U4065 ( .B(n2681), .A(n2926), .S(n3579), .Y(n3377) );
  MUX2X1 U4066 ( .B(n3376), .A(n3373), .S(n1931), .Y(n3379) );
  MUX2X1 U4067 ( .B(n2619), .A(n3054), .S(n3579), .Y(n3383) );
  MUX2X1 U4068 ( .B(n2525), .A(n2836), .S(n3579), .Y(n3382) );
  MUX2X1 U4069 ( .B(n2590), .A(n3023), .S(n3579), .Y(n3386) );
  MUX2X1 U4070 ( .B(n2500), .A(n2807), .S(n3579), .Y(n3385) );
  MUX2X1 U4071 ( .B(n3384), .A(n3381), .S(n1931), .Y(n3394) );
  MUX2X1 U4072 ( .B(n2739), .A(n2989), .S(n3579), .Y(n3389) );
  MUX2X1 U4073 ( .B(n2710), .A(n2957), .S(n3579), .Y(n3388) );
  MUX2X1 U4074 ( .B(n2667), .A(n3086), .S(n3579), .Y(n3392) );
  MUX2X1 U4075 ( .B(n2680), .A(n2925), .S(n3579), .Y(n3391) );
  MUX2X1 U4076 ( .B(n3390), .A(n3387), .S(n1931), .Y(n3393) );
  MUX2X1 U4077 ( .B(n2618), .A(n3053), .S(n3580), .Y(n3397) );
  MUX2X1 U4078 ( .B(n2524), .A(n2835), .S(n3580), .Y(n3396) );
  MUX2X1 U4079 ( .B(n2589), .A(n3022), .S(n3580), .Y(n3400) );
  MUX2X1 U4080 ( .B(n2499), .A(n2806), .S(n3580), .Y(n3399) );
  MUX2X1 U4081 ( .B(n3398), .A(n3395), .S(n1931), .Y(n3408) );
  MUX2X1 U4082 ( .B(n2738), .A(n2988), .S(n3580), .Y(n3403) );
  MUX2X1 U4083 ( .B(n2709), .A(n2956), .S(n3580), .Y(n3402) );
  MUX2X1 U4084 ( .B(n2776), .A(n3085), .S(n3580), .Y(n3406) );
  MUX2X1 U4085 ( .B(n2660), .A(n2924), .S(n3580), .Y(n3405) );
  MUX2X1 U4086 ( .B(n3404), .A(n3401), .S(n1931), .Y(n3407) );
  MUX2X1 U4087 ( .B(n2617), .A(n3052), .S(n3580), .Y(n3411) );
  MUX2X1 U4088 ( .B(n2523), .A(n2834), .S(n3580), .Y(n3410) );
  MUX2X1 U4089 ( .B(n2588), .A(n3021), .S(n3580), .Y(n3414) );
  MUX2X1 U4090 ( .B(n2498), .A(n2805), .S(n3580), .Y(n3413) );
  MUX2X1 U4091 ( .B(n3412), .A(n3409), .S(n1931), .Y(n3422) );
  MUX2X1 U4092 ( .B(n2737), .A(n2987), .S(n3581), .Y(n3417) );
  MUX2X1 U4093 ( .B(n2708), .A(n2955), .S(n3581), .Y(n3416) );
  MUX2X1 U4094 ( .B(n2775), .A(n3084), .S(n3581), .Y(n3420) );
  MUX2X1 U4095 ( .B(n2679), .A(n2923), .S(n3581), .Y(n3419) );
  MUX2X1 U4096 ( .B(n3418), .A(n3415), .S(n1931), .Y(n3421) );
  MUX2X1 U4097 ( .B(n2616), .A(n3051), .S(n3581), .Y(n3425) );
  MUX2X1 U4098 ( .B(n2522), .A(n2833), .S(n3581), .Y(n3424) );
  MUX2X1 U4099 ( .B(n2587), .A(n3020), .S(n3581), .Y(n3428) );
  MUX2X1 U4100 ( .B(n2497), .A(n2804), .S(n3581), .Y(n3427) );
  MUX2X1 U4101 ( .B(n3426), .A(n3423), .S(n1931), .Y(n3436) );
  MUX2X1 U4102 ( .B(n2736), .A(n2986), .S(n3581), .Y(n3431) );
  MUX2X1 U4103 ( .B(n2707), .A(n2954), .S(n3581), .Y(n3430) );
  MUX2X1 U4104 ( .B(n2774), .A(n3083), .S(n3581), .Y(n3434) );
  MUX2X1 U4105 ( .B(n2678), .A(n2922), .S(n3581), .Y(n3433) );
  MUX2X1 U4106 ( .B(n3432), .A(n3429), .S(n1931), .Y(n3435) );
  MUX2X1 U4107 ( .B(n2615), .A(n3050), .S(n3582), .Y(n3439) );
  MUX2X1 U4108 ( .B(n2521), .A(n2832), .S(n3582), .Y(n3438) );
  MUX2X1 U4109 ( .B(n2586), .A(n3019), .S(n3582), .Y(n3442) );
  MUX2X1 U4110 ( .B(n2496), .A(n2803), .S(n3582), .Y(n3441) );
  MUX2X1 U4111 ( .B(n3440), .A(n3437), .S(n1931), .Y(n3450) );
  MUX2X1 U4112 ( .B(n2735), .A(n2985), .S(n3582), .Y(n3445) );
  MUX2X1 U4113 ( .B(n2706), .A(n2953), .S(n3582), .Y(n3444) );
  MUX2X1 U4114 ( .B(n2773), .A(n3082), .S(n3582), .Y(n3448) );
  MUX2X1 U4115 ( .B(n2677), .A(n2921), .S(n3582), .Y(n3447) );
  MUX2X1 U4116 ( .B(n3446), .A(n3443), .S(n1931), .Y(n3449) );
  MUX2X1 U4117 ( .B(n2614), .A(n3049), .S(n3582), .Y(n3453) );
  MUX2X1 U4118 ( .B(n2520), .A(n2831), .S(n3582), .Y(n3452) );
  MUX2X1 U4119 ( .B(n2585), .A(n3018), .S(n3582), .Y(n3456) );
  MUX2X1 U4120 ( .B(n2495), .A(n2802), .S(n3582), .Y(n3455) );
  MUX2X1 U4121 ( .B(n3454), .A(n3451), .S(n1931), .Y(n3464) );
  MUX2X1 U4122 ( .B(n2734), .A(n2984), .S(n3583), .Y(n3459) );
  MUX2X1 U4123 ( .B(n2705), .A(n2952), .S(n3583), .Y(n3458) );
  MUX2X1 U4124 ( .B(n2772), .A(n3081), .S(n3583), .Y(n3462) );
  MUX2X1 U4125 ( .B(n2676), .A(n2920), .S(n3583), .Y(n3461) );
  MUX2X1 U4126 ( .B(n3460), .A(n3457), .S(n1931), .Y(n3463) );
  MUX2X1 U4127 ( .B(n2613), .A(n3048), .S(n3583), .Y(n3467) );
  MUX2X1 U4128 ( .B(n2519), .A(n2830), .S(n3583), .Y(n3466) );
  MUX2X1 U4129 ( .B(n2584), .A(n3017), .S(n3583), .Y(n3470) );
  MUX2X1 U4130 ( .B(n2494), .A(n2801), .S(n3583), .Y(n3469) );
  MUX2X1 U4131 ( .B(n3468), .A(n3465), .S(n1931), .Y(n3478) );
  MUX2X1 U4132 ( .B(n2733), .A(n2983), .S(n3583), .Y(n3473) );
  MUX2X1 U4133 ( .B(n2704), .A(n2951), .S(n3583), .Y(n3472) );
  MUX2X1 U4134 ( .B(n2771), .A(n3080), .S(n3583), .Y(n3476) );
  MUX2X1 U4135 ( .B(n2675), .A(n2919), .S(n3583), .Y(n3475) );
  MUX2X1 U4136 ( .B(n3474), .A(n3471), .S(n1931), .Y(n3477) );
  MUX2X1 U4137 ( .B(n2612), .A(n3047), .S(n3584), .Y(n3481) );
  MUX2X1 U4138 ( .B(n2518), .A(n2829), .S(n3584), .Y(n3480) );
  MUX2X1 U4139 ( .B(n2583), .A(n3016), .S(n3584), .Y(n3484) );
  MUX2X1 U4140 ( .B(n2493), .A(n2800), .S(n3584), .Y(n3483) );
  MUX2X1 U4141 ( .B(n3482), .A(n3479), .S(n1931), .Y(n3492) );
  MUX2X1 U4142 ( .B(n2732), .A(n2982), .S(n3584), .Y(n3487) );
  MUX2X1 U4143 ( .B(n2703), .A(n2950), .S(n3584), .Y(n3486) );
  MUX2X1 U4144 ( .B(n2770), .A(n3079), .S(n3584), .Y(n3490) );
  MUX2X1 U4145 ( .B(n2674), .A(n2918), .S(n3584), .Y(n3489) );
  MUX2X1 U4146 ( .B(n3488), .A(n3485), .S(n1931), .Y(n3491) );
  MUX2X1 U4147 ( .B(n2611), .A(n3046), .S(n3584), .Y(n3495) );
  MUX2X1 U4148 ( .B(n2482), .A(n2828), .S(n3584), .Y(n3494) );
  MUX2X1 U4149 ( .B(n2572), .A(n3015), .S(n3584), .Y(n3498) );
  MUX2X1 U4150 ( .B(n2478), .A(n2799), .S(n3584), .Y(n3497) );
  MUX2X1 U4151 ( .B(n3496), .A(n3493), .S(n1931), .Y(n3506) );
  MUX2X1 U4152 ( .B(n2731), .A(n2981), .S(n3585), .Y(n3501) );
  MUX2X1 U4153 ( .B(n2702), .A(n2949), .S(n3585), .Y(n3500) );
  MUX2X1 U4154 ( .B(n2769), .A(n3078), .S(n3585), .Y(n3504) );
  MUX2X1 U4155 ( .B(n2673), .A(n2917), .S(n3585), .Y(n3503) );
  MUX2X1 U4156 ( .B(n3502), .A(n3499), .S(n1931), .Y(n3505) );
  MUX2X1 U4157 ( .B(n2610), .A(n3045), .S(n3585), .Y(n3509) );
  MUX2X1 U4158 ( .B(n2517), .A(n2827), .S(n3585), .Y(n3508) );
  MUX2X1 U4159 ( .B(n2571), .A(n3014), .S(n3585), .Y(n3512) );
  MUX2X1 U4160 ( .B(n2477), .A(n2798), .S(n3585), .Y(n3511) );
  MUX2X1 U4161 ( .B(n3510), .A(n3507), .S(n1931), .Y(n3520) );
  MUX2X1 U4162 ( .B(n2730), .A(n2980), .S(n3585), .Y(n3515) );
  MUX2X1 U4163 ( .B(n2701), .A(n2948), .S(n3585), .Y(n3514) );
  MUX2X1 U4164 ( .B(n2768), .A(n3077), .S(n3585), .Y(n3518) );
  MUX2X1 U4165 ( .B(n2672), .A(n2916), .S(n3585), .Y(n3517) );
  MUX2X1 U4166 ( .B(n3516), .A(n3513), .S(n1931), .Y(n3519) );
  MUX2X1 U4167 ( .B(n2609), .A(n3044), .S(n3586), .Y(n3523) );
  MUX2X1 U4168 ( .B(n2516), .A(n2826), .S(n3586), .Y(n3522) );
  MUX2X1 U4169 ( .B(n2582), .A(n3013), .S(n3586), .Y(n3526) );
  MUX2X1 U4170 ( .B(n2476), .A(n2797), .S(n3586), .Y(n3525) );
  MUX2X1 U4171 ( .B(n3524), .A(n3521), .S(n1931), .Y(n3534) );
  MUX2X1 U4172 ( .B(n2665), .A(n2979), .S(n3586), .Y(n3529) );
  MUX2X1 U4173 ( .B(n2700), .A(n2947), .S(n3586), .Y(n3528) );
  MUX2X1 U4174 ( .B(n2767), .A(n3076), .S(n3586), .Y(n3532) );
  MUX2X1 U4175 ( .B(n2671), .A(n2915), .S(n3586), .Y(n3531) );
  MUX2X1 U4176 ( .B(n3530), .A(n3527), .S(n1931), .Y(n3533) );
  MUX2X1 U4177 ( .B(n2608), .A(n3043), .S(n3586), .Y(n3537) );
  MUX2X1 U4178 ( .B(n2515), .A(n2825), .S(n3586), .Y(n3536) );
  MUX2X1 U4179 ( .B(n2581), .A(n3012), .S(n3586), .Y(n3540) );
  MUX2X1 U4180 ( .B(n2492), .A(n2796), .S(n3586), .Y(n3539) );
  MUX2X1 U4181 ( .B(n3538), .A(n3535), .S(n1931), .Y(n3548) );
  MUX2X1 U4182 ( .B(n2729), .A(n2978), .S(n3566), .Y(n3543) );
  MUX2X1 U4183 ( .B(n2662), .A(n2946), .S(n3566), .Y(n3542) );
  MUX2X1 U4184 ( .B(n2766), .A(n3075), .S(n3566), .Y(n3546) );
  MUX2X1 U4185 ( .B(n2670), .A(n2914), .S(n3566), .Y(n3545) );
  MUX2X1 U4186 ( .B(n3544), .A(n3541), .S(n1931), .Y(n3547) );
  MUX2X1 U4187 ( .B(n2760), .A(n3011), .S(n3573), .Y(n3551) );
  MUX2X1 U4188 ( .B(n2759), .A(n3010), .S(n3566), .Y(n3550) );
  MUX2X1 U4189 ( .B(n2795), .A(n3106), .S(n3572), .Y(n3554) );
  MUX2X1 U4190 ( .B(n2758), .A(n3009), .S(n3574), .Y(n3553) );
  MUX2X1 U4191 ( .B(n3552), .A(n3549), .S(n1931), .Y(n3562) );
  MUX2X1 U4192 ( .B(n2728), .A(n2977), .S(n3566), .Y(n3557) );
  MUX2X1 U4193 ( .B(n2699), .A(n2945), .S(n3566), .Y(n3556) );
  MUX2X1 U4194 ( .B(n2765), .A(n3074), .S(n3566), .Y(n3560) );
  MUX2X1 U4195 ( .B(n2669), .A(n2913), .S(n3566), .Y(n3559) );
  MUX2X1 U4196 ( .B(n3558), .A(n3555), .S(n1931), .Y(n3561) );
  XNOR2X1 U4197 ( .A(n2856), .B(sub_125_carry[4]), .Y(full_check[4]) );
  XOR2X1 U4198 ( .A(add_148_carry[4]), .B(n2856), .Y(n39) );
  XOR2X1 U4199 ( .A(add_169_carry[4]), .B(n3109), .Y(n111) );
endmodule

